LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_15_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(8)-1 DOWNTO 0));
END L8_15_WROM;

ARCHITECTURE RTL OF L8_15_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"011010010",
  1=>"110010000",
  2=>"001110110",
  3=>"111110000",
  4=>"101001101",
  5=>"001000000",
  6=>"110011001",
  7=>"000100011",
  8=>"010110101",
  9=>"110010010",
  10=>"000000000",
  11=>"000010111",
  12=>"000100000",
  13=>"011011010",
  14=>"001110101",
  15=>"010101011",
  16=>"110101001",
  17=>"011111001",
  18=>"001001101",
  19=>"001001011",
  20=>"000001110",
  21=>"101001001",
  22=>"001101100",
  23=>"000010010",
  24=>"110000111",
  25=>"000000000",
  26=>"101000000",
  27=>"011110011",
  28=>"111001101",
  29=>"110000111",
  30=>"010001000",
  31=>"101010100",
  32=>"101101101",
  33=>"001110001",
  34=>"100101110",
  35=>"011100010",
  36=>"101110111",
  37=>"010100001",
  38=>"010001111",
  39=>"100001000",
  40=>"011011011",
  41=>"010010010",
  42=>"000100001",
  43=>"000111111",
  44=>"011001000",
  45=>"001100101",
  46=>"111110101",
  47=>"110000100",
  48=>"100100110",
  49=>"001100000",
  50=>"010100011",
  51=>"011100100",
  52=>"100001110",
  53=>"000000100",
  54=>"000111000",
  55=>"000100001",
  56=>"100000010",
  57=>"011110101",
  58=>"100110010",
  59=>"111011110",
  60=>"010100001",
  61=>"010011011",
  62=>"000100000",
  63=>"000010000",
  64=>"111101100",
  65=>"011000000",
  66=>"111011010",
  67=>"100001110",
  68=>"011100011",
  69=>"101010010",
  70=>"000111101",
  71=>"011100001",
  72=>"110000011",
  73=>"010111001",
  74=>"101111110",
  75=>"010101010",
  76=>"101011001",
  77=>"110100010",
  78=>"011011010",
  79=>"010000001",
  80=>"000001110",
  81=>"101000000",
  82=>"111001010",
  83=>"111111100",
  84=>"101100100",
  85=>"010100000",
  86=>"011001011",
  87=>"110110100",
  88=>"100101111",
  89=>"100001010",
  90=>"111111110",
  91=>"100101010",
  92=>"110110011",
  93=>"111010000",
  94=>"111001100",
  95=>"001100101",
  96=>"000100101",
  97=>"101010101",
  98=>"011100110",
  99=>"110100010",
  100=>"011111001",
  101=>"101111101",
  102=>"011111011",
  103=>"111010111",
  104=>"000000110",
  105=>"101001000",
  106=>"101100000",
  107=>"111001100",
  108=>"001001010",
  109=>"101100111",
  110=>"011111010",
  111=>"011011000",
  112=>"100000110",
  113=>"011111101",
  114=>"010111001",
  115=>"001100100",
  116=>"000001011",
  117=>"010101011",
  118=>"011100100",
  119=>"111110001",
  120=>"011110010",
  121=>"111111110",
  122=>"110011011",
  123=>"110011011",
  124=>"010000000",
  125=>"000000000",
  126=>"011011000",
  127=>"001101011",
  128=>"100101011",
  129=>"010110011",
  130=>"101101100",
  131=>"010000011",
  132=>"110100110",
  133=>"000100101",
  134=>"110101001",
  135=>"001000111",
  136=>"110111110",
  137=>"000011011",
  138=>"110000011",
  139=>"100000010",
  140=>"011000000",
  141=>"001001010",
  142=>"111001011",
  143=>"001101001",
  144=>"110010110",
  145=>"110111000",
  146=>"000010101",
  147=>"111010011",
  148=>"111000000",
  149=>"010101000",
  150=>"101010000",
  151=>"110001010",
  152=>"001101001",
  153=>"101001100",
  154=>"111000011",
  155=>"011100100",
  156=>"101100000",
  157=>"011010011",
  158=>"100101000",
  159=>"110010101",
  160=>"000100101",
  161=>"001111110",
  162=>"101110111",
  163=>"010110101",
  164=>"011110000",
  165=>"001111011",
  166=>"000001010",
  167=>"011010010",
  168=>"101100101",
  169=>"101011110",
  170=>"110100111",
  171=>"101011110",
  172=>"110111000",
  173=>"011101100",
  174=>"111110010",
  175=>"110111011",
  176=>"101000101",
  177=>"110101100",
  178=>"100110100",
  179=>"100000001",
  180=>"101110001",
  181=>"001110111",
  182=>"010011011",
  183=>"101111011",
  184=>"100000001",
  185=>"000000111",
  186=>"100011000",
  187=>"001100111",
  188=>"011001110",
  189=>"101001101",
  190=>"010110111",
  191=>"110011010",
  192=>"100110100",
  193=>"111111010",
  194=>"011100110",
  195=>"111111111",
  196=>"001000000",
  197=>"101100111",
  198=>"011000101",
  199=>"100101001",
  200=>"111101101",
  201=>"011000101",
  202=>"000100011",
  203=>"010011111",
  204=>"001011111",
  205=>"110010111",
  206=>"000100011",
  207=>"111111111",
  208=>"111000010",
  209=>"101001000",
  210=>"100001110",
  211=>"110001001",
  212=>"011000011",
  213=>"001010101",
  214=>"100001001",
  215=>"110101010",
  216=>"011111101",
  217=>"000100010",
  218=>"011111001",
  219=>"010001101",
  220=>"101100101",
  221=>"001100100",
  222=>"000100111",
  223=>"111001011",
  224=>"010010100",
  225=>"010001110",
  226=>"111010001",
  227=>"101100110",
  228=>"101101111",
  229=>"101001010",
  230=>"010000001",
  231=>"111011100",
  232=>"100101101",
  233=>"100010000",
  234=>"101101001",
  235=>"101111001",
  236=>"010010110",
  237=>"000101011",
  238=>"010010010",
  239=>"000000011",
  240=>"111010100",
  241=>"110111101",
  242=>"010010001",
  243=>"110101111",
  244=>"101000011",
  245=>"001111010",
  246=>"000011110",
  247=>"000000100",
  248=>"000011000",
  249=>"111101101",
  250=>"110011011",
  251=>"010101100",
  252=>"001100101",
  253=>"101001000",
  254=>"110110010",
  255=>"111001100",
  256=>"011111111",
  257=>"010110010",
  258=>"011110011",
  259=>"101011110",
  260=>"100011101",
  261=>"111101110",
  262=>"000101100",
  263=>"000000010",
  264=>"000000100",
  265=>"000100111",
  266=>"001101010",
  267=>"100101010",
  268=>"010000111",
  269=>"010100101",
  270=>"000011001",
  271=>"010010010",
  272=>"100000100",
  273=>"010101001",
  274=>"100010100",
  275=>"101011000",
  276=>"010101000",
  277=>"100001100",
  278=>"000001100",
  279=>"111100101",
  280=>"111101101",
  281=>"100000100",
  282=>"101110101",
  283=>"101010010",
  284=>"111101100",
  285=>"000110010",
  286=>"100001100",
  287=>"000001000",
  288=>"100001001",
  289=>"100000100",
  290=>"011100101",
  291=>"101100001",
  292=>"101100101",
  293=>"011111111",
  294=>"000101110",
  295=>"111111001",
  296=>"101001101",
  297=>"110011011",
  298=>"010000011",
  299=>"101110100",
  300=>"001110010",
  301=>"100101010",
  302=>"010010000",
  303=>"011101010",
  304=>"100011010",
  305=>"000100111",
  306=>"000100110",
  307=>"000010110",
  308=>"001101100",
  309=>"010100000",
  310=>"010111100",
  311=>"100111000",
  312=>"000101000",
  313=>"100110000",
  314=>"110000010",
  315=>"100110110",
  316=>"111001100",
  317=>"111101000",
  318=>"101000011",
  319=>"111010111",
  320=>"101100000",
  321=>"010000000",
  322=>"010110011",
  323=>"111000000",
  324=>"011010000",
  325=>"100011101",
  326=>"000001101",
  327=>"000000010",
  328=>"000001001",
  329=>"001100000",
  330=>"101100111",
  331=>"010111001",
  332=>"000100101",
  333=>"000001000",
  334=>"000110000",
  335=>"111011010",
  336=>"100001110",
  337=>"110101010",
  338=>"011000110",
  339=>"000011100",
  340=>"101111010",
  341=>"011111000",
  342=>"111100111",
  343=>"000100111",
  344=>"010100011",
  345=>"101011011",
  346=>"011000010",
  347=>"000010100",
  348=>"100100110",
  349=>"011010000",
  350=>"001110111",
  351=>"011010111",
  352=>"001010100",
  353=>"000011010",
  354=>"000111111",
  355=>"010010100",
  356=>"001101001",
  357=>"010111010",
  358=>"011101011",
  359=>"001110001",
  360=>"000001000",
  361=>"100101100",
  362=>"000111001",
  363=>"111000000",
  364=>"000001100",
  365=>"010101010",
  366=>"011111101",
  367=>"011010101",
  368=>"000110100",
  369=>"010110011",
  370=>"100111101",
  371=>"101010001",
  372=>"000111101",
  373=>"010111000",
  374=>"110110000",
  375=>"010001010",
  376=>"010100001",
  377=>"100000010",
  378=>"101000110",
  379=>"100100000",
  380=>"100000101",
  381=>"110000111",
  382=>"110001001",
  383=>"110000011",
  384=>"011110010",
  385=>"000001000",
  386=>"010001010",
  387=>"110000011",
  388=>"110001001",
  389=>"010011110",
  390=>"111011001",
  391=>"010000100",
  392=>"010011000",
  393=>"000010011",
  394=>"001110011",
  395=>"001011101",
  396=>"011010101",
  397=>"101110110",
  398=>"100001010",
  399=>"001110100",
  400=>"101101111",
  401=>"101101010",
  402=>"101010101",
  403=>"001111010",
  404=>"001000100",
  405=>"000011000",
  406=>"011101011",
  407=>"101101001",
  408=>"011100011",
  409=>"111101110",
  410=>"000010101",
  411=>"011001000",
  412=>"001011010",
  413=>"000001110",
  414=>"001111001",
  415=>"000000000",
  416=>"110000111",
  417=>"011100101",
  418=>"010011100",
  419=>"000010001",
  420=>"111100000",
  421=>"000010100",
  422=>"010010000",
  423=>"010000111",
  424=>"001000111",
  425=>"000011001",
  426=>"100011111",
  427=>"111011000",
  428=>"101001110",
  429=>"000010001",
  430=>"000000110",
  431=>"110101010",
  432=>"001101011",
  433=>"101100000",
  434=>"011101001",
  435=>"010000111",
  436=>"100011101",
  437=>"011001000",
  438=>"101110110",
  439=>"000010101",
  440=>"000101110",
  441=>"010000111",
  442=>"010001001",
  443=>"011011111",
  444=>"000100011",
  445=>"111110000",
  446=>"100010000",
  447=>"101111010",
  448=>"011100000",
  449=>"100000111",
  450=>"111011101",
  451=>"100010101",
  452=>"010011001",
  453=>"011110110",
  454=>"010000011",
  455=>"101001111",
  456=>"001001010",
  457=>"101111111",
  458=>"101000011",
  459=>"001011101",
  460=>"001011001",
  461=>"100111101",
  462=>"111101001",
  463=>"001000111",
  464=>"100000110",
  465=>"011011000",
  466=>"010010101",
  467=>"111111101",
  468=>"011100001",
  469=>"010001001",
  470=>"001101011",
  471=>"011101010",
  472=>"101101101",
  473=>"111011011",
  474=>"001110111",
  475=>"110010000",
  476=>"011000110",
  477=>"000111101",
  478=>"101011111",
  479=>"111111000",
  480=>"111110010",
  481=>"001001011",
  482=>"001100000",
  483=>"011000001",
  484=>"000001011",
  485=>"000000100",
  486=>"011110010",
  487=>"011110101",
  488=>"011111110",
  489=>"110001010",
  490=>"010101000",
  491=>"111110000",
  492=>"100001000",
  493=>"010111010",
  494=>"000101010",
  495=>"011110110",
  496=>"101100101",
  497=>"111001010",
  498=>"101011000",
  499=>"000001000",
  500=>"000011111",
  501=>"101011100",
  502=>"101010000",
  503=>"000000010",
  504=>"010010110",
  505=>"111000101",
  506=>"011010111",
  507=>"101000111",
  508=>"100011111",
  509=>"110111100",
  510=>"110010101",
  511=>"110100000",
  512=>"110111101",
  513=>"010101011",
  514=>"111010000",
  515=>"001110111",
  516=>"110110111",
  517=>"001011000",
  518=>"101000111",
  519=>"011000001",
  520=>"110000100",
  521=>"000100100",
  522=>"111111100",
  523=>"110101111",
  524=>"010111010",
  525=>"001000000",
  526=>"011010001",
  527=>"111000110",
  528=>"101111111",
  529=>"000101010",
  530=>"111101110",
  531=>"111100101",
  532=>"000011000",
  533=>"010111110",
  534=>"100111110",
  535=>"110001000",
  536=>"111000010",
  537=>"011111101",
  538=>"101100000",
  539=>"111100000",
  540=>"010100011",
  541=>"010000110",
  542=>"011100101",
  543=>"100010100",
  544=>"000011011",
  545=>"110101110",
  546=>"000101111",
  547=>"110010011",
  548=>"110010110",
  549=>"101100000",
  550=>"010111100",
  551=>"000101000",
  552=>"011000000",
  553=>"011111100",
  554=>"000100000",
  555=>"111011110",
  556=>"001110100",
  557=>"010001110",
  558=>"011100101",
  559=>"101101110",
  560=>"100110000",
  561=>"000001011",
  562=>"001101110",
  563=>"101100000",
  564=>"010111001",
  565=>"101100111",
  566=>"001010010",
  567=>"011100000",
  568=>"110101100",
  569=>"011101011",
  570=>"111101111",
  571=>"110011000",
  572=>"101000100",
  573=>"101010110",
  574=>"100000101",
  575=>"110010111",
  576=>"010101111",
  577=>"011101010",
  578=>"001000101",
  579=>"111110111",
  580=>"000101001",
  581=>"011011101",
  582=>"000011101",
  583=>"010100111",
  584=>"101100010",
  585=>"111100000",
  586=>"001100110",
  587=>"010101100",
  588=>"000101100",
  589=>"100100001",
  590=>"100000111",
  591=>"010111101",
  592=>"111111100",
  593=>"011101001",
  594=>"101000000",
  595=>"010110001",
  596=>"001111011",
  597=>"110000011",
  598=>"011011100",
  599=>"111011000",
  600=>"011101101",
  601=>"101010001",
  602=>"110011100",
  603=>"111010100",
  604=>"111100010",
  605=>"010000001",
  606=>"100010111",
  607=>"010001111",
  608=>"000001010",
  609=>"101001001",
  610=>"000000101",
  611=>"001011010",
  612=>"001010000",
  613=>"101111000",
  614=>"111100001",
  615=>"001010010",
  616=>"010111000",
  617=>"000000110",
  618=>"000101100",
  619=>"011001010",
  620=>"101000101",
  621=>"101101101",
  622=>"100100100",
  623=>"101001110",
  624=>"001111010",
  625=>"011101001",
  626=>"011000001",
  627=>"000010110",
  628=>"101100011",
  629=>"001101001",
  630=>"110010000",
  631=>"111101101",
  632=>"011011100",
  633=>"101111100",
  634=>"110000100",
  635=>"101101010",
  636=>"001110001",
  637=>"010111110",
  638=>"110000011",
  639=>"000111111",
  640=>"010011101",
  641=>"101101111",
  642=>"001000111",
  643=>"000010000",
  644=>"000110100",
  645=>"010100100",
  646=>"010101001",
  647=>"001000101",
  648=>"000100100",
  649=>"111010011",
  650=>"111000111",
  651=>"110010010",
  652=>"100000100",
  653=>"011111100",
  654=>"010001001",
  655=>"111000101",
  656=>"100001001",
  657=>"101001011",
  658=>"110110101",
  659=>"110110111",
  660=>"111010000",
  661=>"111101111",
  662=>"101000010",
  663=>"111101011",
  664=>"100110101",
  665=>"101011101",
  666=>"010000010",
  667=>"000110111",
  668=>"000010010",
  669=>"101111010",
  670=>"010011111",
  671=>"100010110",
  672=>"100001011",
  673=>"101000111",
  674=>"001110111",
  675=>"011100101",
  676=>"000010111",
  677=>"001111000",
  678=>"100001001",
  679=>"010110000",
  680=>"000000101",
  681=>"010100011",
  682=>"111000010",
  683=>"001001011",
  684=>"101100101",
  685=>"000100100",
  686=>"010110001",
  687=>"101101110",
  688=>"011100000",
  689=>"001111101",
  690=>"011010100",
  691=>"100000100",
  692=>"110011011",
  693=>"110011100",
  694=>"001111110",
  695=>"111010011",
  696=>"010011011",
  697=>"110010100",
  698=>"110111011",
  699=>"100110011",
  700=>"011110111",
  701=>"000010011",
  702=>"101010001",
  703=>"100100001",
  704=>"000001111",
  705=>"111101001",
  706=>"000011110",
  707=>"011010111",
  708=>"111100010",
  709=>"111101101",
  710=>"100000101",
  711=>"111000110",
  712=>"011001000",
  713=>"100011111",
  714=>"010001110",
  715=>"110011000",
  716=>"101101001",
  717=>"101110111",
  718=>"101000000",
  719=>"100011011",
  720=>"100111010",
  721=>"011111010",
  722=>"110010100",
  723=>"100100010",
  724=>"101001100",
  725=>"101101110",
  726=>"010101100",
  727=>"000000000",
  728=>"110010101",
  729=>"100111100",
  730=>"001101010",
  731=>"110110001",
  732=>"010101000",
  733=>"001001110",
  734=>"111101111",
  735=>"001011010",
  736=>"011011000",
  737=>"000011011",
  738=>"000110011",
  739=>"000000110",
  740=>"111111100",
  741=>"001100000",
  742=>"001010100",
  743=>"001011100",
  744=>"001101000",
  745=>"111111110",
  746=>"101011011",
  747=>"111000110",
  748=>"101001000",
  749=>"001010110",
  750=>"100011001",
  751=>"010110110",
  752=>"001011010",
  753=>"110100000",
  754=>"100110101",
  755=>"111101010",
  756=>"100011011",
  757=>"110011010",
  758=>"001001111",
  759=>"001101100",
  760=>"110110110",
  761=>"101110110",
  762=>"000111101",
  763=>"000010100",
  764=>"000011000",
  765=>"011110011",
  766=>"100101011",
  767=>"111110010",
  768=>"111100011",
  769=>"000010111",
  770=>"010111100",
  771=>"101000011",
  772=>"000110001",
  773=>"010100011",
  774=>"110011101",
  775=>"101000101",
  776=>"000111011",
  777=>"111011110",
  778=>"010000011",
  779=>"001010011",
  780=>"011000010",
  781=>"100010111",
  782=>"110100000",
  783=>"111111001",
  784=>"101000001",
  785=>"010111100",
  786=>"110000110",
  787=>"001011111",
  788=>"101100110",
  789=>"100100000",
  790=>"101111010",
  791=>"100110111",
  792=>"110001000",
  793=>"000100011",
  794=>"110011001",
  795=>"110011111",
  796=>"001010010",
  797=>"111011111",
  798=>"000010011",
  799=>"111000101",
  800=>"100000011",
  801=>"000110110",
  802=>"000100111",
  803=>"101001111",
  804=>"100010100",
  805=>"001001000",
  806=>"111010000",
  807=>"111101110",
  808=>"000111010",
  809=>"110100100",
  810=>"110011000",
  811=>"111110011",
  812=>"011011100",
  813=>"101110101",
  814=>"101010010",
  815=>"011000010",
  816=>"100110010",
  817=>"000001101",
  818=>"000010100",
  819=>"000011111",
  820=>"000111010",
  821=>"010111010",
  822=>"111001000",
  823=>"100011010",
  824=>"001000010",
  825=>"000111000",
  826=>"001100010",
  827=>"101001100",
  828=>"011001011",
  829=>"001010100",
  830=>"000000000",
  831=>"011011010",
  832=>"100100001",
  833=>"001100110",
  834=>"001000011",
  835=>"011001001",
  836=>"100011110",
  837=>"011010000",
  838=>"011010011",
  839=>"101110111",
  840=>"011110100",
  841=>"100110101",
  842=>"101101010",
  843=>"011100010",
  844=>"100100010",
  845=>"010011101",
  846=>"011000101",
  847=>"011000000",
  848=>"111100000",
  849=>"101101111",
  850=>"010011000",
  851=>"011100001",
  852=>"000100100",
  853=>"011100100",
  854=>"101110011",
  855=>"110101000",
  856=>"111101111",
  857=>"010100110",
  858=>"101101101",
  859=>"101001011",
  860=>"101110100",
  861=>"010001000",
  862=>"100000001",
  863=>"010011100",
  864=>"100010111",
  865=>"011010000",
  866=>"001111110",
  867=>"011011111",
  868=>"100010000",
  869=>"101101100",
  870=>"110101010",
  871=>"001110101",
  872=>"010000000",
  873=>"101101111",
  874=>"100101111",
  875=>"111111001",
  876=>"010100101",
  877=>"100111001",
  878=>"101000010",
  879=>"111100100",
  880=>"000110000",
  881=>"000011101",
  882=>"001000111",
  883=>"111110001",
  884=>"100100000",
  885=>"100000010",
  886=>"100001000",
  887=>"001000010",
  888=>"101101010",
  889=>"011100010",
  890=>"110001010",
  891=>"110111001",
  892=>"000100000",
  893=>"101001101",
  894=>"111100100",
  895=>"011000101",
  896=>"011011011",
  897=>"100110001",
  898=>"101011111",
  899=>"001100011",
  900=>"110101000",
  901=>"101000001",
  902=>"110000001",
  903=>"111110001",
  904=>"111100110",
  905=>"110010100",
  906=>"011011100",
  907=>"100010011",
  908=>"010110100",
  909=>"111000001",
  910=>"110110000",
  911=>"110010100",
  912=>"101101001",
  913=>"101111110",
  914=>"000110010",
  915=>"000101101",
  916=>"011100100",
  917=>"000110011",
  918=>"010111011",
  919=>"101000001",
  920=>"110100111",
  921=>"001100010",
  922=>"001101110",
  923=>"000010010",
  924=>"110110000",
  925=>"000010011",
  926=>"000010100",
  927=>"011010001",
  928=>"100011000",
  929=>"100011101",
  930=>"101001110",
  931=>"101111111",
  932=>"101000000",
  933=>"101100101",
  934=>"010010010",
  935=>"110111111",
  936=>"000001011",
  937=>"000100010",
  938=>"101001010",
  939=>"101101001",
  940=>"100111010",
  941=>"000110110",
  942=>"001000110",
  943=>"111111011",
  944=>"110110100",
  945=>"110011101",
  946=>"111011010",
  947=>"111110000",
  948=>"100100000",
  949=>"110111001",
  950=>"100101110",
  951=>"111100000",
  952=>"001000010",
  953=>"010001001",
  954=>"011110011",
  955=>"110001111",
  956=>"001110010",
  957=>"101000110",
  958=>"101011011",
  959=>"011101000",
  960=>"101010010",
  961=>"000000010",
  962=>"000000101",
  963=>"011001000",
  964=>"000101011",
  965=>"101101000",
  966=>"011100001",
  967=>"111000000",
  968=>"111101000",
  969=>"010011101",
  970=>"010110111",
  971=>"100111111",
  972=>"110111001",
  973=>"110100011",
  974=>"110100100",
  975=>"101001010",
  976=>"011110011",
  977=>"000110001",
  978=>"100010001",
  979=>"110010110",
  980=>"010110000",
  981=>"011001001",
  982=>"101001100",
  983=>"011101110",
  984=>"001010111",
  985=>"110011011",
  986=>"101011001",
  987=>"111011101",
  988=>"000110001",
  989=>"111010000",
  990=>"001000100",
  991=>"101001101",
  992=>"000010001",
  993=>"011000001",
  994=>"001100011",
  995=>"011010000",
  996=>"000000000",
  997=>"010101101",
  998=>"010101000",
  999=>"101111011",
  1000=>"000100000",
  1001=>"101100111",
  1002=>"001100100",
  1003=>"000100010",
  1004=>"101000010",
  1005=>"100011010",
  1006=>"100101100",
  1007=>"110010010",
  1008=>"011110111",
  1009=>"101011000",
  1010=>"001101110",
  1011=>"100100001",
  1012=>"101110011",
  1013=>"000010001",
  1014=>"010111111",
  1015=>"101111001",
  1016=>"011010000",
  1017=>"110110100",
  1018=>"000011110",
  1019=>"101000010",
  1020=>"001010110",
  1021=>"011011111",
  1022=>"010000100",
  1023=>"001101011",
  1024=>"000101111",
  1025=>"001010110",
  1026=>"010010101",
  1027=>"110101100",
  1028=>"111100000",
  1029=>"100100101",
  1030=>"100101111",
  1031=>"111111101",
  1032=>"000010100",
  1033=>"001000010",
  1034=>"101011000",
  1035=>"100111100",
  1036=>"100010011",
  1037=>"110100111",
  1038=>"000000110",
  1039=>"111011010",
  1040=>"101100011",
  1041=>"111111100",
  1042=>"000011110",
  1043=>"000110010",
  1044=>"111001100",
  1045=>"111010011",
  1046=>"111101111",
  1047=>"110001100",
  1048=>"100010001",
  1049=>"001110000",
  1050=>"100001111",
  1051=>"010100110",
  1052=>"010110010",
  1053=>"011100111",
  1054=>"101010001",
  1055=>"100001011",
  1056=>"010101010",
  1057=>"110101010",
  1058=>"100011111",
  1059=>"101010100",
  1060=>"101101011",
  1061=>"000101010",
  1062=>"100101011",
  1063=>"101101101",
  1064=>"001001000",
  1065=>"001100011",
  1066=>"000010110",
  1067=>"010011111",
  1068=>"101111111",
  1069=>"100110000",
  1070=>"000001100",
  1071=>"001101000",
  1072=>"110111100",
  1073=>"001001010",
  1074=>"000011000",
  1075=>"000000111",
  1076=>"001000110",
  1077=>"100101110",
  1078=>"000011101",
  1079=>"111111000",
  1080=>"101010011",
  1081=>"110101011",
  1082=>"010011101",
  1083=>"110100100",
  1084=>"111011010",
  1085=>"101011010",
  1086=>"000110011",
  1087=>"000110000",
  1088=>"001001000",
  1089=>"111110010",
  1090=>"011100010",
  1091=>"100101010",
  1092=>"010010001",
  1093=>"001010111",
  1094=>"001011001",
  1095=>"011010101",
  1096=>"110101111",
  1097=>"001101011",
  1098=>"100101011",
  1099=>"101100011",
  1100=>"100110001",
  1101=>"110010001",
  1102=>"010101001",
  1103=>"101000011",
  1104=>"100011100",
  1105=>"011010101",
  1106=>"110000110",
  1107=>"011100100",
  1108=>"101010010",
  1109=>"111100111",
  1110=>"100101101",
  1111=>"001001010",
  1112=>"110110001",
  1113=>"001110110",
  1114=>"111101011",
  1115=>"110001000",
  1116=>"101111111",
  1117=>"000000100",
  1118=>"001001100",
  1119=>"011101001",
  1120=>"110000111",
  1121=>"101000011",
  1122=>"100000111",
  1123=>"101001000",
  1124=>"101001010",
  1125=>"110101011",
  1126=>"001111101",
  1127=>"001001000",
  1128=>"111000011",
  1129=>"010100100",
  1130=>"010001110",
  1131=>"110111010",
  1132=>"010100010",
  1133=>"010100010",
  1134=>"010011101",
  1135=>"010100100",
  1136=>"101000100",
  1137=>"010111100",
  1138=>"011000001",
  1139=>"111110001",
  1140=>"010000100",
  1141=>"000000000",
  1142=>"011000000",
  1143=>"111000110",
  1144=>"111101000",
  1145=>"010011101",
  1146=>"010101110",
  1147=>"001010000",
  1148=>"010111100",
  1149=>"101010101",
  1150=>"010000001",
  1151=>"111101110",
  1152=>"011110001",
  1153=>"100000000",
  1154=>"111101001",
  1155=>"011000110",
  1156=>"000001011",
  1157=>"000100010",
  1158=>"001110110",
  1159=>"010011110",
  1160=>"000000101",
  1161=>"111011111",
  1162=>"011011111",
  1163=>"000001101",
  1164=>"010011101",
  1165=>"110111110",
  1166=>"001100111",
  1167=>"011010100",
  1168=>"010010101",
  1169=>"110110001",
  1170=>"111010010",
  1171=>"110100001",
  1172=>"000011101",
  1173=>"010110010",
  1174=>"100010000",
  1175=>"111001111",
  1176=>"100000100",
  1177=>"000100101",
  1178=>"110101110",
  1179=>"101010101",
  1180=>"010011101",
  1181=>"101000101",
  1182=>"111101111",
  1183=>"000110000",
  1184=>"000111000",
  1185=>"000010101",
  1186=>"010110011",
  1187=>"111101000",
  1188=>"110100001",
  1189=>"010110001",
  1190=>"111001101",
  1191=>"100001010",
  1192=>"110000001",
  1193=>"001001000",
  1194=>"111001111",
  1195=>"000000101",
  1196=>"101101011",
  1197=>"100011101",
  1198=>"000010100",
  1199=>"010001111",
  1200=>"010110000",
  1201=>"000101101",
  1202=>"101000011",
  1203=>"100010110",
  1204=>"010111001",
  1205=>"100000001",
  1206=>"000101011",
  1207=>"010010010",
  1208=>"010101111",
  1209=>"011111111",
  1210=>"101000110",
  1211=>"011010011",
  1212=>"111011011",
  1213=>"000000111",
  1214=>"110110110",
  1215=>"011000100",
  1216=>"110101101",
  1217=>"100111111",
  1218=>"100001101",
  1219=>"101110110",
  1220=>"001001110",
  1221=>"000000000",
  1222=>"110111011",
  1223=>"110100010",
  1224=>"000010011",
  1225=>"101101111",
  1226=>"001110011",
  1227=>"100111100",
  1228=>"010000110",
  1229=>"100010010",
  1230=>"010000111",
  1231=>"110111000",
  1232=>"010111100",
  1233=>"100011001",
  1234=>"001010110",
  1235=>"011111100",
  1236=>"011111101",
  1237=>"100100000",
  1238=>"011000010",
  1239=>"110010101",
  1240=>"000010010",
  1241=>"100101011",
  1242=>"001101000",
  1243=>"100001111",
  1244=>"010100101",
  1245=>"100011011",
  1246=>"011001000",
  1247=>"000010010",
  1248=>"000101111",
  1249=>"110110101",
  1250=>"101001000",
  1251=>"000101000",
  1252=>"010111010",
  1253=>"000111111",
  1254=>"101101010",
  1255=>"000000000",
  1256=>"111010100",
  1257=>"001110110",
  1258=>"110110001",
  1259=>"000000010",
  1260=>"001011001",
  1261=>"000011111",
  1262=>"111110101",
  1263=>"000100010",
  1264=>"011000010",
  1265=>"001110111",
  1266=>"001010011",
  1267=>"111010000",
  1268=>"001110001",
  1269=>"110010010",
  1270=>"011010110",
  1271=>"100001001",
  1272=>"011011010",
  1273=>"011001000",
  1274=>"010110101",
  1275=>"110001000",
  1276=>"010110010",
  1277=>"001000000",
  1278=>"110110110",
  1279=>"001100110",
  1280=>"000100111",
  1281=>"011101010",
  1282=>"000110101",
  1283=>"000011101",
  1284=>"111010001",
  1285=>"010001000",
  1286=>"101010111",
  1287=>"110100100",
  1288=>"111010101",
  1289=>"001101111",
  1290=>"001011001",
  1291=>"000111011",
  1292=>"101000000",
  1293=>"001100101",
  1294=>"110100111",
  1295=>"000011000",
  1296=>"001100110",
  1297=>"111100101",
  1298=>"010011101",
  1299=>"001010111",
  1300=>"000010001",
  1301=>"100001101",
  1302=>"101011111",
  1303=>"010111001",
  1304=>"000000100",
  1305=>"101111011",
  1306=>"010101011",
  1307=>"101111000",
  1308=>"101000001",
  1309=>"111001001",
  1310=>"011111010",
  1311=>"001100000",
  1312=>"000000010",
  1313=>"111110111",
  1314=>"101010110",
  1315=>"111001100",
  1316=>"111000010",
  1317=>"001001101",
  1318=>"001000101",
  1319=>"011011111",
  1320=>"100111111",
  1321=>"111010110",
  1322=>"110010011",
  1323=>"011001000",
  1324=>"100110101",
  1325=>"111101011",
  1326=>"000010010",
  1327=>"101001110",
  1328=>"100000000",
  1329=>"111000010",
  1330=>"110100111",
  1331=>"000011101",
  1332=>"010110010",
  1333=>"111110111",
  1334=>"100001010",
  1335=>"001111011",
  1336=>"111100110",
  1337=>"001010010",
  1338=>"011000001",
  1339=>"000101101",
  1340=>"100111111",
  1341=>"110110101",
  1342=>"110110001",
  1343=>"101111110",
  1344=>"001111011",
  1345=>"111000000",
  1346=>"111101000",
  1347=>"110110110",
  1348=>"011100011",
  1349=>"000001101",
  1350=>"100001010",
  1351=>"000010000",
  1352=>"001001000",
  1353=>"100110000",
  1354=>"000110001",
  1355=>"000010000",
  1356=>"011010010",
  1357=>"110011110",
  1358=>"110011100",
  1359=>"101010111",
  1360=>"111101000",
  1361=>"100101100",
  1362=>"101100101",
  1363=>"111100010",
  1364=>"000001001",
  1365=>"100011011",
  1366=>"101011001",
  1367=>"011001011",
  1368=>"010000010",
  1369=>"001100001",
  1370=>"000110100",
  1371=>"000000000",
  1372=>"011101111",
  1373=>"101110000",
  1374=>"010101100",
  1375=>"101111001",
  1376=>"000111011",
  1377=>"001000100",
  1378=>"101111100",
  1379=>"000001110",
  1380=>"101010100",
  1381=>"111101100",
  1382=>"110100000",
  1383=>"101011001",
  1384=>"110000101",
  1385=>"000000000",
  1386=>"110010100",
  1387=>"000100101",
  1388=>"001100110",
  1389=>"101011111",
  1390=>"110010010",
  1391=>"000110011",
  1392=>"101011111",
  1393=>"100001101",
  1394=>"110111011",
  1395=>"000011110",
  1396=>"011100100",
  1397=>"100111011",
  1398=>"010101010",
  1399=>"101110100",
  1400=>"000101011",
  1401=>"011101011",
  1402=>"111111000",
  1403=>"000101001",
  1404=>"001100001",
  1405=>"100110011",
  1406=>"100010101",
  1407=>"010111110",
  1408=>"100000110",
  1409=>"110000111",
  1410=>"011011011",
  1411=>"001001111",
  1412=>"101011010",
  1413=>"000101101",
  1414=>"101000100",
  1415=>"011010110",
  1416=>"011000101",
  1417=>"110000001",
  1418=>"110100101",
  1419=>"000000111",
  1420=>"111110001",
  1421=>"111101101",
  1422=>"110000101",
  1423=>"001110110",
  1424=>"110011000",
  1425=>"010010000",
  1426=>"000110011",
  1427=>"100001000",
  1428=>"001001000",
  1429=>"101100101",
  1430=>"111011000",
  1431=>"010100000",
  1432=>"011110100",
  1433=>"100110010",
  1434=>"101101011",
  1435=>"010010001",
  1436=>"001101010",
  1437=>"111101111",
  1438=>"111011100",
  1439=>"110011101",
  1440=>"001110010",
  1441=>"101111111",
  1442=>"001010111",
  1443=>"111011110",
  1444=>"000011000",
  1445=>"100100001",
  1446=>"100011010",
  1447=>"100000000",
  1448=>"000101011",
  1449=>"100010111",
  1450=>"011110111",
  1451=>"111010111",
  1452=>"010000010",
  1453=>"101111001",
  1454=>"001000000",
  1455=>"001101010",
  1456=>"111110111",
  1457=>"001101011",
  1458=>"101100101",
  1459=>"011001001",
  1460=>"100000001",
  1461=>"011001010",
  1462=>"100010110",
  1463=>"100010000",
  1464=>"111110101",
  1465=>"001110001",
  1466=>"001101011",
  1467=>"100001011",
  1468=>"001010000",
  1469=>"111110100",
  1470=>"011111100",
  1471=>"000011000",
  1472=>"010010111",
  1473=>"001011000",
  1474=>"011001011",
  1475=>"111111101",
  1476=>"110000000",
  1477=>"111001100",
  1478=>"001000100",
  1479=>"110000101",
  1480=>"101010010",
  1481=>"111111001",
  1482=>"111011111",
  1483=>"110011100",
  1484=>"100000001",
  1485=>"101001010",
  1486=>"110000001",
  1487=>"000001001",
  1488=>"010111101",
  1489=>"101001110",
  1490=>"000001011",
  1491=>"011110011",
  1492=>"111100000",
  1493=>"110001101",
  1494=>"111111110",
  1495=>"000110000",
  1496=>"000111110",
  1497=>"001011100",
  1498=>"000100001",
  1499=>"111111110",
  1500=>"001110000",
  1501=>"111000110",
  1502=>"011101011",
  1503=>"100011011",
  1504=>"111110101",
  1505=>"110000100",
  1506=>"011110000",
  1507=>"101011111",
  1508=>"011101011",
  1509=>"110100100",
  1510=>"100011101",
  1511=>"010101100",
  1512=>"010101011",
  1513=>"011111111",
  1514=>"101011011",
  1515=>"001100000",
  1516=>"100011100",
  1517=>"111110111",
  1518=>"110100011",
  1519=>"000111110",
  1520=>"110100101",
  1521=>"111100011",
  1522=>"011100100",
  1523=>"010110001",
  1524=>"100100011",
  1525=>"111101001",
  1526=>"111001000",
  1527=>"101100110",
  1528=>"101011110",
  1529=>"000110101",
  1530=>"110111110",
  1531=>"111101111",
  1532=>"100100000",
  1533=>"000111010",
  1534=>"100011010",
  1535=>"100000101",
  1536=>"101011010",
  1537=>"000110000",
  1538=>"110001010",
  1539=>"101100101",
  1540=>"011000011",
  1541=>"111110011",
  1542=>"101000111",
  1543=>"011000100",
  1544=>"100110111",
  1545=>"110111000",
  1546=>"001000100",
  1547=>"111010001",
  1548=>"011011100",
  1549=>"111101101",
  1550=>"010001011",
  1551=>"000010110",
  1552=>"111100110",
  1553=>"010110001",
  1554=>"011111110",
  1555=>"011001101",
  1556=>"111011110",
  1557=>"110011111",
  1558=>"011010010",
  1559=>"110111010",
  1560=>"100011000",
  1561=>"010111000",
  1562=>"010001100",
  1563=>"110010010",
  1564=>"000011001",
  1565=>"100011000",
  1566=>"011000110",
  1567=>"001000001",
  1568=>"110001111",
  1569=>"111011100",
  1570=>"110010000",
  1571=>"011000011",
  1572=>"010101101",
  1573=>"011011011",
  1574=>"110011111",
  1575=>"101001100",
  1576=>"101010000",
  1577=>"100101100",
  1578=>"010100011",
  1579=>"110100001",
  1580=>"111000010",
  1581=>"111001001",
  1582=>"000010010",
  1583=>"111101101",
  1584=>"101100011",
  1585=>"110100100",
  1586=>"100101011",
  1587=>"101010100",
  1588=>"001000110",
  1589=>"000101110",
  1590=>"011001010",
  1591=>"001000000",
  1592=>"111110000",
  1593=>"000011110",
  1594=>"101111100",
  1595=>"010000000",
  1596=>"000101110",
  1597=>"100100110",
  1598=>"111101000",
  1599=>"000011101",
  1600=>"100111111",
  1601=>"111100111",
  1602=>"010010101",
  1603=>"010100000",
  1604=>"001001101",
  1605=>"000011001",
  1606=>"010010000",
  1607=>"001001000",
  1608=>"101010001",
  1609=>"101111011",
  1610=>"100100001",
  1611=>"010101011",
  1612=>"001010000",
  1613=>"000000111",
  1614=>"000011010",
  1615=>"010100110",
  1616=>"101000010",
  1617=>"010111011",
  1618=>"000000000",
  1619=>"010010010",
  1620=>"000101001",
  1621=>"000001101",
  1622=>"001100000",
  1623=>"100000001",
  1624=>"000000000",
  1625=>"010101100",
  1626=>"000110011",
  1627=>"001010010",
  1628=>"111101000",
  1629=>"010000001",
  1630=>"001110100",
  1631=>"000001010",
  1632=>"100100011",
  1633=>"001001001",
  1634=>"111110000",
  1635=>"110101001",
  1636=>"010111100",
  1637=>"010000001",
  1638=>"011011010",
  1639=>"110011111",
  1640=>"001100001",
  1641=>"101010110",
  1642=>"101101111",
  1643=>"010101101",
  1644=>"010101100",
  1645=>"100010100",
  1646=>"001100011",
  1647=>"101100000",
  1648=>"110011010",
  1649=>"111111110",
  1650=>"110011010",
  1651=>"010010111",
  1652=>"011001010",
  1653=>"100001111",
  1654=>"111110100",
  1655=>"010101110",
  1656=>"011110111",
  1657=>"110100010",
  1658=>"111110110",
  1659=>"111110101",
  1660=>"000100010",
  1661=>"110001101",
  1662=>"000111011",
  1663=>"100110011",
  1664=>"101110101",
  1665=>"110100110",
  1666=>"101110101",
  1667=>"111110000",
  1668=>"111010001",
  1669=>"100100110",
  1670=>"111111010",
  1671=>"100000110",
  1672=>"000011011",
  1673=>"101100110",
  1674=>"101111000",
  1675=>"010000110",
  1676=>"000000001",
  1677=>"011001000",
  1678=>"111011101",
  1679=>"010101110",
  1680=>"010100011",
  1681=>"010110010",
  1682=>"010110010",
  1683=>"010011000",
  1684=>"110100111",
  1685=>"001100001",
  1686=>"010111101",
  1687=>"011001011",
  1688=>"001010100",
  1689=>"101010111",
  1690=>"101000111",
  1691=>"010001100",
  1692=>"111010101",
  1693=>"100000000",
  1694=>"101111101",
  1695=>"101101101",
  1696=>"111111101",
  1697=>"111001100",
  1698=>"010000000",
  1699=>"101111100",
  1700=>"010111011",
  1701=>"111000011",
  1702=>"110010010",
  1703=>"110000100",
  1704=>"111001110",
  1705=>"111001110",
  1706=>"111011010",
  1707=>"000001000",
  1708=>"000000001",
  1709=>"110000001",
  1710=>"111100010",
  1711=>"010010001",
  1712=>"111001110",
  1713=>"010011110",
  1714=>"001101010",
  1715=>"011100111",
  1716=>"111111010",
  1717=>"010010000",
  1718=>"111111111",
  1719=>"110011110",
  1720=>"000101000",
  1721=>"101110111",
  1722=>"010101011",
  1723=>"110000011",
  1724=>"011100011",
  1725=>"010010111",
  1726=>"111011101",
  1727=>"111001011",
  1728=>"111001101",
  1729=>"000000000",
  1730=>"000000000",
  1731=>"110111011",
  1732=>"001110111",
  1733=>"101000010",
  1734=>"111111101",
  1735=>"110110100",
  1736=>"001100000",
  1737=>"100001000",
  1738=>"000110010",
  1739=>"101101111",
  1740=>"101000011",
  1741=>"111001101",
  1742=>"101011111",
  1743=>"001000000",
  1744=>"100000011",
  1745=>"001001101",
  1746=>"011001110",
  1747=>"100001100",
  1748=>"111000101",
  1749=>"110011110",
  1750=>"111110001",
  1751=>"110010010",
  1752=>"000011101",
  1753=>"011000000",
  1754=>"000100111",
  1755=>"111101111",
  1756=>"000101010",
  1757=>"111100111",
  1758=>"011001100",
  1759=>"101111110",
  1760=>"101001011",
  1761=>"001110001",
  1762=>"000001011",
  1763=>"110010111",
  1764=>"010001111",
  1765=>"101000010",
  1766=>"010110011",
  1767=>"001001001",
  1768=>"100011101",
  1769=>"100000001",
  1770=>"000000100",
  1771=>"011101011",
  1772=>"101101000",
  1773=>"101010110",
  1774=>"101001100",
  1775=>"000001110",
  1776=>"111111000",
  1777=>"011110010",
  1778=>"111111110",
  1779=>"000100110",
  1780=>"010100110",
  1781=>"000111010",
  1782=>"000000000",
  1783=>"111101000",
  1784=>"101100110",
  1785=>"101000011",
  1786=>"101010111",
  1787=>"101110110",
  1788=>"110111111",
  1789=>"100000100",
  1790=>"110110100",
  1791=>"000000111",
  1792=>"011111101",
  1793=>"001001000",
  1794=>"001001011",
  1795=>"001010000",
  1796=>"110010000",
  1797=>"010011000",
  1798=>"011000101",
  1799=>"111001110",
  1800=>"001000111",
  1801=>"010011011",
  1802=>"110011110",
  1803=>"101100000",
  1804=>"011000110",
  1805=>"000111010",
  1806=>"001010011",
  1807=>"001111100",
  1808=>"110010001",
  1809=>"001100110",
  1810=>"111101111",
  1811=>"101111100",
  1812=>"000011101",
  1813=>"010010110",
  1814=>"101001001",
  1815=>"101010111",
  1816=>"011101000",
  1817=>"001010001",
  1818=>"011111110",
  1819=>"101100001",
  1820=>"010011010",
  1821=>"001000111",
  1822=>"011101000",
  1823=>"001000111",
  1824=>"011101101",
  1825=>"111011111",
  1826=>"010101000",
  1827=>"001001101",
  1828=>"100000001",
  1829=>"110111101",
  1830=>"110100001",
  1831=>"111101010",
  1832=>"000011001",
  1833=>"000101100",
  1834=>"001100100",
  1835=>"100000111",
  1836=>"010011010",
  1837=>"010001010",
  1838=>"111010100",
  1839=>"111101101",
  1840=>"000110110",
  1841=>"110111001",
  1842=>"001101010",
  1843=>"001110000",
  1844=>"000000001",
  1845=>"001011111",
  1846=>"100001111",
  1847=>"010101000",
  1848=>"000101110",
  1849=>"011100000",
  1850=>"100110010",
  1851=>"000001000",
  1852=>"000101101",
  1853=>"000000111",
  1854=>"100111000",
  1855=>"011101110",
  1856=>"110110000",
  1857=>"110011110",
  1858=>"110000110",
  1859=>"101001111",
  1860=>"111000000",
  1861=>"001111001",
  1862=>"111111101",
  1863=>"000100001",
  1864=>"101111111",
  1865=>"011011001",
  1866=>"010000010",
  1867=>"110010101",
  1868=>"100001011",
  1869=>"110100000",
  1870=>"111101111",
  1871=>"010100011",
  1872=>"010100100",
  1873=>"010001010",
  1874=>"011010011",
  1875=>"000100010",
  1876=>"111010000",
  1877=>"100001101",
  1878=>"010110010",
  1879=>"110101000",
  1880=>"101001000",
  1881=>"000100001",
  1882=>"111010011",
  1883=>"001110110",
  1884=>"001100001",
  1885=>"000110010",
  1886=>"111101100",
  1887=>"110010110",
  1888=>"010111100",
  1889=>"000110000",
  1890=>"000111111",
  1891=>"111010101",
  1892=>"000101000",
  1893=>"001001001",
  1894=>"011011101",
  1895=>"100110110",
  1896=>"010010011",
  1897=>"110111111",
  1898=>"111000101",
  1899=>"110111001",
  1900=>"000010100",
  1901=>"000001000",
  1902=>"001110111",
  1903=>"110100010",
  1904=>"000000100",
  1905=>"000000100",
  1906=>"000011010",
  1907=>"011000110",
  1908=>"000101010",
  1909=>"111111101",
  1910=>"101101000",
  1911=>"110000100",
  1912=>"001111001",
  1913=>"100011010",
  1914=>"010000110",
  1915=>"110101010",
  1916=>"101011101",
  1917=>"011010101",
  1918=>"100011101",
  1919=>"001100110",
  1920=>"000011100",
  1921=>"100111100",
  1922=>"111101000",
  1923=>"101111100",
  1924=>"111111111",
  1925=>"000010101",
  1926=>"100111100",
  1927=>"001011100",
  1928=>"001100110",
  1929=>"100000010",
  1930=>"011011110",
  1931=>"000110010",
  1932=>"001000011",
  1933=>"101100100",
  1934=>"111100011",
  1935=>"100111100",
  1936=>"000011110",
  1937=>"010110010",
  1938=>"110010111",
  1939=>"110100101",
  1940=>"001011100",
  1941=>"111011010",
  1942=>"111100101",
  1943=>"111100111",
  1944=>"000010011",
  1945=>"001010001",
  1946=>"010110100",
  1947=>"101100011",
  1948=>"011000110",
  1949=>"010010111",
  1950=>"100100111",
  1951=>"101110101",
  1952=>"111100011",
  1953=>"101011110",
  1954=>"110100010",
  1955=>"110010111",
  1956=>"110110000",
  1957=>"001000111",
  1958=>"010000101",
  1959=>"010100100",
  1960=>"100111101",
  1961=>"011100111",
  1962=>"000110001",
  1963=>"101110001",
  1964=>"101110001",
  1965=>"100101100",
  1966=>"100101000",
  1967=>"101000011",
  1968=>"010001110",
  1969=>"000110000",
  1970=>"001101000",
  1971=>"001001100",
  1972=>"111100011",
  1973=>"101000110",
  1974=>"101110100",
  1975=>"110010111",
  1976=>"000110111",
  1977=>"110011010",
  1978=>"010000101",
  1979=>"001100000",
  1980=>"000110111",
  1981=>"010001100",
  1982=>"111111111",
  1983=>"000001101",
  1984=>"001011111",
  1985=>"100001000",
  1986=>"010000011",
  1987=>"000010101",
  1988=>"010011100",
  1989=>"010100110",
  1990=>"010101000",
  1991=>"000100000",
  1992=>"111100110",
  1993=>"110101010",
  1994=>"001011100",
  1995=>"110001011",
  1996=>"111010000",
  1997=>"010110001",
  1998=>"010001111",
  1999=>"010100011",
  2000=>"110000010",
  2001=>"101000111",
  2002=>"000101100",
  2003=>"111101101",
  2004=>"000000111",
  2005=>"111010101",
  2006=>"110111000",
  2007=>"111100100",
  2008=>"110010000",
  2009=>"000010011",
  2010=>"001101011",
  2011=>"110101001",
  2012=>"000011111",
  2013=>"000110101",
  2014=>"000011010",
  2015=>"001110011",
  2016=>"111010001",
  2017=>"101101110",
  2018=>"110011100",
  2019=>"011100001",
  2020=>"000000101",
  2021=>"000001000",
  2022=>"100000000",
  2023=>"100000101",
  2024=>"010101001",
  2025=>"111010110",
  2026=>"111111001",
  2027=>"001001111",
  2028=>"010111110",
  2029=>"100000000",
  2030=>"001101110",
  2031=>"101011111",
  2032=>"100100111",
  2033=>"010101110",
  2034=>"010000010",
  2035=>"001010110",
  2036=>"010111011",
  2037=>"101011001",
  2038=>"111101111",
  2039=>"111011101",
  2040=>"000000000",
  2041=>"110110010",
  2042=>"100100110",
  2043=>"000101111",
  2044=>"010110011",
  2045=>"010100101",
  2046=>"101111101",
  2047=>"010100110",
  2048=>"111001100",
  2049=>"010000011",
  2050=>"111011010",
  2051=>"000100000",
  2052=>"010100111",
  2053=>"101000011",
  2054=>"000001010",
  2055=>"000100001",
  2056=>"000000111",
  2057=>"100101000",
  2058=>"001000101",
  2059=>"001111110",
  2060=>"000100000",
  2061=>"111011100",
  2062=>"101001010",
  2063=>"001010110",
  2064=>"111010011",
  2065=>"000000010",
  2066=>"101001011",
  2067=>"010100110",
  2068=>"111110101",
  2069=>"101001010",
  2070=>"110001100",
  2071=>"101101101",
  2072=>"011010010",
  2073=>"111000011",
  2074=>"100101000",
  2075=>"010111010",
  2076=>"110010011",
  2077=>"101110110",
  2078=>"011101110",
  2079=>"101010110",
  2080=>"000000000",
  2081=>"011101011",
  2082=>"011101011",
  2083=>"100011000",
  2084=>"101001111",
  2085=>"111000111",
  2086=>"100110010",
  2087=>"111101101",
  2088=>"111011011",
  2089=>"111001111",
  2090=>"100101111",
  2091=>"011101000",
  2092=>"110100000",
  2093=>"111100111",
  2094=>"110100010",
  2095=>"011111001",
  2096=>"011110000",
  2097=>"001011101",
  2098=>"110100100",
  2099=>"001100010",
  2100=>"101011000",
  2101=>"111101101",
  2102=>"001011100",
  2103=>"100000100",
  2104=>"111100100",
  2105=>"001000100",
  2106=>"101111100",
  2107=>"010100001",
  2108=>"001001110",
  2109=>"101001010",
  2110=>"011011100",
  2111=>"000101000",
  2112=>"001010110",
  2113=>"011100110",
  2114=>"001000110",
  2115=>"000100010",
  2116=>"111011011",
  2117=>"100011110",
  2118=>"001010111",
  2119=>"110101111",
  2120=>"011011111",
  2121=>"100111101",
  2122=>"110100111",
  2123=>"000111010",
  2124=>"010101010",
  2125=>"110010101",
  2126=>"111001001",
  2127=>"010111111",
  2128=>"111011110",
  2129=>"111100101",
  2130=>"101100010",
  2131=>"110111110",
  2132=>"100001111",
  2133=>"111001110",
  2134=>"001101100",
  2135=>"111101001",
  2136=>"100011011",
  2137=>"010001011",
  2138=>"101111110",
  2139=>"011100110",
  2140=>"001001101",
  2141=>"000010100",
  2142=>"011101110",
  2143=>"010000010",
  2144=>"000110111",
  2145=>"110100100",
  2146=>"010101110",
  2147=>"101000001",
  2148=>"010001100",
  2149=>"110100110",
  2150=>"110110111",
  2151=>"101111100",
  2152=>"110100101",
  2153=>"110011001",
  2154=>"100110000",
  2155=>"010111000",
  2156=>"010111000",
  2157=>"001100111",
  2158=>"000010101",
  2159=>"001101100",
  2160=>"100001100",
  2161=>"000001001",
  2162=>"110011001",
  2163=>"100010111",
  2164=>"111011110",
  2165=>"001010000",
  2166=>"000110100",
  2167=>"010010010",
  2168=>"100010110",
  2169=>"011010110",
  2170=>"010000001",
  2171=>"101100111",
  2172=>"010101000",
  2173=>"101000111",
  2174=>"100110111",
  2175=>"111101111",
  2176=>"101010100",
  2177=>"011000000",
  2178=>"110111011",
  2179=>"100000010",
  2180=>"011010011",
  2181=>"101111101",
  2182=>"110011101",
  2183=>"000101011",
  2184=>"111101101",
  2185=>"111101011",
  2186=>"111111100",
  2187=>"100110010",
  2188=>"111111100",
  2189=>"010111100",
  2190=>"101100111",
  2191=>"011111100",
  2192=>"010000001",
  2193=>"110001011",
  2194=>"010110011",
  2195=>"100000111",
  2196=>"011010000",
  2197=>"100101101",
  2198=>"000011000",
  2199=>"011101001",
  2200=>"000100001",
  2201=>"111011111",
  2202=>"000110010",
  2203=>"000111110",
  2204=>"010000111",
  2205=>"111110100",
  2206=>"111111011",
  2207=>"110000001",
  2208=>"000011011",
  2209=>"010011001",
  2210=>"011111011",
  2211=>"010110010",
  2212=>"011100111",
  2213=>"110110111",
  2214=>"010001111",
  2215=>"111101111",
  2216=>"010110010",
  2217=>"101011001",
  2218=>"111010000",
  2219=>"110100111",
  2220=>"000110010",
  2221=>"001110000",
  2222=>"101111011",
  2223=>"001011011",
  2224=>"101000001",
  2225=>"001011111",
  2226=>"010100000",
  2227=>"011011010",
  2228=>"000000000",
  2229=>"010100100",
  2230=>"111010101",
  2231=>"101100110",
  2232=>"010000100",
  2233=>"100001111",
  2234=>"100100111",
  2235=>"011101111",
  2236=>"010100101",
  2237=>"110010011",
  2238=>"110110010",
  2239=>"111011101",
  2240=>"010100110",
  2241=>"011111000",
  2242=>"000101101",
  2243=>"001100111",
  2244=>"011011110",
  2245=>"100111111",
  2246=>"000000101",
  2247=>"000000110",
  2248=>"110111100",
  2249=>"011000001",
  2250=>"101010111",
  2251=>"011000110",
  2252=>"010100010",
  2253=>"111110111",
  2254=>"110010000",
  2255=>"110110100",
  2256=>"011011010",
  2257=>"000101011",
  2258=>"100100110",
  2259=>"110011001",
  2260=>"111000001",
  2261=>"011101110",
  2262=>"101001001",
  2263=>"011001101",
  2264=>"001100001",
  2265=>"001000000",
  2266=>"111000001",
  2267=>"100001000",
  2268=>"010011001",
  2269=>"000000000",
  2270=>"101010001",
  2271=>"001000010",
  2272=>"111110101",
  2273=>"100011001",
  2274=>"010101101",
  2275=>"000011100",
  2276=>"001000100",
  2277=>"100100100",
  2278=>"010011101",
  2279=>"100000111",
  2280=>"001001100",
  2281=>"001111001",
  2282=>"011100011",
  2283=>"100011110",
  2284=>"110010100",
  2285=>"000001100",
  2286=>"000001100",
  2287=>"000101101",
  2288=>"001011011",
  2289=>"000001001",
  2290=>"000000011",
  2291=>"001100011",
  2292=>"111100011",
  2293=>"111110001",
  2294=>"110011110",
  2295=>"111011110",
  2296=>"101001001",
  2297=>"001011001",
  2298=>"111000101",
  2299=>"100101010",
  2300=>"010100100",
  2301=>"010011111",
  2302=>"110101010",
  2303=>"001010100",
  2304=>"100010101",
  2305=>"010001101",
  2306=>"001001010",
  2307=>"101100000",
  2308=>"010000011",
  2309=>"001111100",
  2310=>"000001001",
  2311=>"011001101",
  2312=>"100011001",
  2313=>"101100011",
  2314=>"100101101",
  2315=>"011100101",
  2316=>"101100000",
  2317=>"000010001",
  2318=>"111111110",
  2319=>"100101100",
  2320=>"011000001",
  2321=>"001000011",
  2322=>"110111001",
  2323=>"011011111",
  2324=>"101010110",
  2325=>"100011110",
  2326=>"111100111",
  2327=>"001111110",
  2328=>"111101010",
  2329=>"011101010",
  2330=>"010011111",
  2331=>"101010011",
  2332=>"100010100",
  2333=>"000001101",
  2334=>"101111011",
  2335=>"000001110",
  2336=>"000111000",
  2337=>"101110001",
  2338=>"001110001",
  2339=>"011000101",
  2340=>"001001011",
  2341=>"000000000",
  2342=>"011101110",
  2343=>"000100110",
  2344=>"000001011",
  2345=>"111010111",
  2346=>"111111110",
  2347=>"000010101",
  2348=>"010011111",
  2349=>"001010110",
  2350=>"000110000",
  2351=>"001010011",
  2352=>"100111101",
  2353=>"110001001",
  2354=>"100011110",
  2355=>"010110011",
  2356=>"001111000",
  2357=>"100011100",
  2358=>"110110010",
  2359=>"111101011",
  2360=>"001000000",
  2361=>"100111001",
  2362=>"110100100",
  2363=>"010000000",
  2364=>"011101101",
  2365=>"000011010",
  2366=>"101111011",
  2367=>"101100111",
  2368=>"100011011",
  2369=>"000010110",
  2370=>"110110111",
  2371=>"100111010",
  2372=>"000101001",
  2373=>"111101010",
  2374=>"010111100",
  2375=>"100100011",
  2376=>"101011110",
  2377=>"000110010",
  2378=>"010101001",
  2379=>"000010000",
  2380=>"001000000",
  2381=>"001100100",
  2382=>"001111011",
  2383=>"000000001",
  2384=>"000101011",
  2385=>"111101011",
  2386=>"011001011",
  2387=>"000100110",
  2388=>"000001010",
  2389=>"101000001",
  2390=>"011110000",
  2391=>"110100011",
  2392=>"001011000",
  2393=>"001010010",
  2394=>"111101110",
  2395=>"001000101",
  2396=>"100011110",
  2397=>"101001011",
  2398=>"111101001",
  2399=>"110101111",
  2400=>"101110100",
  2401=>"001110010",
  2402=>"101001010",
  2403=>"001101011",
  2404=>"001011011",
  2405=>"011010110",
  2406=>"101101101",
  2407=>"010100010",
  2408=>"001000111",
  2409=>"100001000",
  2410=>"000011101",
  2411=>"010100101",
  2412=>"000001101",
  2413=>"101111100",
  2414=>"000010110",
  2415=>"111100000",
  2416=>"100011111",
  2417=>"110000110",
  2418=>"100101111",
  2419=>"010110000",
  2420=>"001001101",
  2421=>"110001001",
  2422=>"001011010",
  2423=>"101111101",
  2424=>"000011110",
  2425=>"000101101",
  2426=>"000101101",
  2427=>"111100100",
  2428=>"000110001",
  2429=>"000101001",
  2430=>"101011011",
  2431=>"111110001",
  2432=>"000100111",
  2433=>"000000010",
  2434=>"011110110",
  2435=>"000010010",
  2436=>"100010100",
  2437=>"111010010",
  2438=>"011110111",
  2439=>"100100100",
  2440=>"100000111",
  2441=>"000000111",
  2442=>"001100101",
  2443=>"010110101",
  2444=>"011111000",
  2445=>"000001010",
  2446=>"011101111",
  2447=>"010110100",
  2448=>"100111111",
  2449=>"010010101",
  2450=>"000001111",
  2451=>"001011110",
  2452=>"010101011",
  2453=>"110001100",
  2454=>"111000110",
  2455=>"100011000",
  2456=>"001110000",
  2457=>"100000010",
  2458=>"110110110",
  2459=>"101111111",
  2460=>"111011111",
  2461=>"111100111",
  2462=>"011100000",
  2463=>"111010111",
  2464=>"111011110",
  2465=>"110101100",
  2466=>"010001100",
  2467=>"000001101",
  2468=>"111111100",
  2469=>"001000000",
  2470=>"001100001",
  2471=>"000100100",
  2472=>"011110101",
  2473=>"101011000",
  2474=>"100000101",
  2475=>"000101100",
  2476=>"000111001",
  2477=>"000100100",
  2478=>"000010011",
  2479=>"111111110",
  2480=>"110000000",
  2481=>"111111000",
  2482=>"100101010",
  2483=>"101101101",
  2484=>"111101111",
  2485=>"111010000",
  2486=>"100001001",
  2487=>"101010110",
  2488=>"000011111",
  2489=>"101000001",
  2490=>"001100011",
  2491=>"000111110",
  2492=>"110000010",
  2493=>"111011010",
  2494=>"011100000",
  2495=>"010110111",
  2496=>"001100111",
  2497=>"110110110",
  2498=>"000100111",
  2499=>"111101000",
  2500=>"001010000",
  2501=>"100100001",
  2502=>"010010101",
  2503=>"111110100",
  2504=>"000001110",
  2505=>"011101000",
  2506=>"101000000",
  2507=>"111100110",
  2508=>"101011100",
  2509=>"010000011",
  2510=>"100000100",
  2511=>"110011010",
  2512=>"100100010",
  2513=>"010001010",
  2514=>"000100101",
  2515=>"000001111",
  2516=>"101010010",
  2517=>"001001100",
  2518=>"010111001",
  2519=>"011011110",
  2520=>"011001110",
  2521=>"100100000",
  2522=>"111111011",
  2523=>"110111111",
  2524=>"110001110",
  2525=>"000110100",
  2526=>"000001010",
  2527=>"011010110",
  2528=>"010110100",
  2529=>"000111101",
  2530=>"111111100",
  2531=>"110000011",
  2532=>"110101010",
  2533=>"111110110",
  2534=>"000010111",
  2535=>"111100100",
  2536=>"000111000",
  2537=>"100000101",
  2538=>"011111100",
  2539=>"010101111",
  2540=>"101111110",
  2541=>"010110011",
  2542=>"001011001",
  2543=>"011111111",
  2544=>"110110101",
  2545=>"101110011",
  2546=>"011111000",
  2547=>"011000011",
  2548=>"100110001",
  2549=>"101101000",
  2550=>"001100101",
  2551=>"000111001",
  2552=>"110000001",
  2553=>"110000101",
  2554=>"011011010",
  2555=>"011000001",
  2556=>"100101001",
  2557=>"101101101",
  2558=>"010000100",
  2559=>"011010000",
  2560=>"111101111",
  2561=>"010110010",
  2562=>"001110001",
  2563=>"110001101",
  2564=>"011000100",
  2565=>"100111000",
  2566=>"111001000",
  2567=>"000000110",
  2568=>"000001111",
  2569=>"100001010",
  2570=>"100011011",
  2571=>"000010000",
  2572=>"000111101",
  2573=>"000100001",
  2574=>"111000011",
  2575=>"010110101",
  2576=>"000111010",
  2577=>"111000110",
  2578=>"100101111",
  2579=>"110111100",
  2580=>"101110011",
  2581=>"100000011",
  2582=>"011110101",
  2583=>"100111111",
  2584=>"010001000",
  2585=>"110111100",
  2586=>"101111111",
  2587=>"101011110",
  2588=>"101100110",
  2589=>"001001110",
  2590=>"111010110",
  2591=>"101111010",
  2592=>"100001101",
  2593=>"011101100",
  2594=>"000011111",
  2595=>"100101100",
  2596=>"001001001",
  2597=>"110010010",
  2598=>"100000111",
  2599=>"110000101",
  2600=>"011000010",
  2601=>"100011001",
  2602=>"101001111",
  2603=>"000111010",
  2604=>"100110010",
  2605=>"010001000",
  2606=>"111100011",
  2607=>"111011010",
  2608=>"110100011",
  2609=>"111001100",
  2610=>"001001100",
  2611=>"100011000",
  2612=>"010010011",
  2613=>"010010111",
  2614=>"110100101",
  2615=>"000110101",
  2616=>"000001011",
  2617=>"111010110",
  2618=>"000101011",
  2619=>"011110001",
  2620=>"000111001",
  2621=>"011010100",
  2622=>"000011001",
  2623=>"001110000",
  2624=>"111110001",
  2625=>"010101010",
  2626=>"100110011",
  2627=>"110111010",
  2628=>"111110101",
  2629=>"001111010",
  2630=>"001001011",
  2631=>"100000001",
  2632=>"111100111",
  2633=>"000001001",
  2634=>"111111110",
  2635=>"001110111",
  2636=>"000110011",
  2637=>"101100010",
  2638=>"111010100",
  2639=>"001000101",
  2640=>"011000100",
  2641=>"001001010",
  2642=>"001110001",
  2643=>"101100001",
  2644=>"011101101",
  2645=>"000110101",
  2646=>"101001010",
  2647=>"101011110",
  2648=>"101110001",
  2649=>"110011001",
  2650=>"001000110",
  2651=>"000001100",
  2652=>"010111100",
  2653=>"100101110",
  2654=>"100000000",
  2655=>"100001111",
  2656=>"011000111",
  2657=>"000101001",
  2658=>"010000000",
  2659=>"000100111",
  2660=>"001111000",
  2661=>"000000010",
  2662=>"010100001",
  2663=>"000100000",
  2664=>"000101000",
  2665=>"001011011",
  2666=>"011111010",
  2667=>"110010001",
  2668=>"110000101",
  2669=>"100110010",
  2670=>"001011110",
  2671=>"001101001",
  2672=>"100011101",
  2673=>"010001011",
  2674=>"101001101",
  2675=>"000000011",
  2676=>"010111001",
  2677=>"111000001",
  2678=>"100100110",
  2679=>"100101110",
  2680=>"101110001",
  2681=>"100100111",
  2682=>"001101101",
  2683=>"001111011",
  2684=>"100000000",
  2685=>"000101000",
  2686=>"110000110",
  2687=>"101100110",
  2688=>"001001101",
  2689=>"111101101",
  2690=>"101100110",
  2691=>"001000110",
  2692=>"011000010",
  2693=>"111100110",
  2694=>"111000011",
  2695=>"000110000",
  2696=>"010001000",
  2697=>"100011010",
  2698=>"001110001",
  2699=>"010000011",
  2700=>"010000000",
  2701=>"011111011",
  2702=>"110001110",
  2703=>"101111101",
  2704=>"110001100",
  2705=>"011001000",
  2706=>"011011101",
  2707=>"001000000",
  2708=>"101001011",
  2709=>"110111011",
  2710=>"010100010",
  2711=>"100000000",
  2712=>"101111110",
  2713=>"100101000",
  2714=>"110100000",
  2715=>"110011001",
  2716=>"100000011",
  2717=>"000001000",
  2718=>"010101110",
  2719=>"111001011",
  2720=>"011011001",
  2721=>"110000011",
  2722=>"010101000",
  2723=>"001010100",
  2724=>"100100100",
  2725=>"010000000",
  2726=>"001010000",
  2727=>"010101000",
  2728=>"011111110",
  2729=>"100000011",
  2730=>"100011110",
  2731=>"110001101",
  2732=>"100011000",
  2733=>"111110101",
  2734=>"001110111",
  2735=>"111111011",
  2736=>"000011000",
  2737=>"011000110",
  2738=>"010111100",
  2739=>"110011110",
  2740=>"001001111",
  2741=>"001011000",
  2742=>"001100010",
  2743=>"101000111",
  2744=>"000001010",
  2745=>"111000110",
  2746=>"011010000",
  2747=>"001110000",
  2748=>"111101101",
  2749=>"001100111",
  2750=>"100111111",
  2751=>"111010000",
  2752=>"111101110",
  2753=>"011010110",
  2754=>"000100101",
  2755=>"100001100",
  2756=>"010110000",
  2757=>"110101101",
  2758=>"011100101",
  2759=>"101111101",
  2760=>"000100110",
  2761=>"011010101",
  2762=>"000101100",
  2763=>"000000000",
  2764=>"000011111",
  2765=>"000110010",
  2766=>"000101010",
  2767=>"001111111",
  2768=>"010010100",
  2769=>"001010111",
  2770=>"110101010",
  2771=>"000111000",
  2772=>"101001001",
  2773=>"000000101",
  2774=>"000100100",
  2775=>"000010101",
  2776=>"000100010",
  2777=>"111110101",
  2778=>"000101010",
  2779=>"111001101",
  2780=>"000110101",
  2781=>"000111001",
  2782=>"100011110",
  2783=>"011110011",
  2784=>"001001100",
  2785=>"011001110",
  2786=>"000101100",
  2787=>"010100111",
  2788=>"000101000",
  2789=>"011001000",
  2790=>"010111100",
  2791=>"111000000",
  2792=>"000010100",
  2793=>"011000101",
  2794=>"000010011",
  2795=>"011000100",
  2796=>"000000101",
  2797=>"000010101",
  2798=>"100010000",
  2799=>"110110010",
  2800=>"110010101",
  2801=>"110001110",
  2802=>"010001100",
  2803=>"011100110",
  2804=>"100101000",
  2805=>"100000001",
  2806=>"111011001",
  2807=>"111110110",
  2808=>"110010001",
  2809=>"000011101",
  2810=>"111001110",
  2811=>"111001011",
  2812=>"001111011",
  2813=>"011101011",
  2814=>"101000000",
  2815=>"110100010",
  2816=>"000001010",
  2817=>"111010111",
  2818=>"010010100",
  2819=>"110010000",
  2820=>"100111111",
  2821=>"100010100",
  2822=>"000110110",
  2823=>"010010010",
  2824=>"001101000",
  2825=>"011111000",
  2826=>"000001111",
  2827=>"111111000",
  2828=>"101010000",
  2829=>"110011001",
  2830=>"011000101",
  2831=>"110111000",
  2832=>"001100010",
  2833=>"000100010",
  2834=>"011101010",
  2835=>"001110111",
  2836=>"111011010",
  2837=>"111110100",
  2838=>"010100011",
  2839=>"000000100",
  2840=>"110000000",
  2841=>"010001101",
  2842=>"011100011",
  2843=>"101011101",
  2844=>"100001110",
  2845=>"110110110",
  2846=>"110011101",
  2847=>"010111010",
  2848=>"100001011",
  2849=>"000101100",
  2850=>"111100000",
  2851=>"001100101",
  2852=>"010000000",
  2853=>"001111011",
  2854=>"001001001",
  2855=>"100001100",
  2856=>"110010101",
  2857=>"101101000",
  2858=>"100101101",
  2859=>"110110111",
  2860=>"010001101",
  2861=>"000111001",
  2862=>"100110101",
  2863=>"001001111",
  2864=>"011000000",
  2865=>"011010011",
  2866=>"011001110",
  2867=>"000100111",
  2868=>"011101100",
  2869=>"101011010",
  2870=>"001000000",
  2871=>"000111100",
  2872=>"010111010",
  2873=>"110011101",
  2874=>"000110111",
  2875=>"110111000",
  2876=>"100110010",
  2877=>"111110000",
  2878=>"111000000",
  2879=>"001110111",
  2880=>"011010110",
  2881=>"111011111",
  2882=>"000000100",
  2883=>"110101001",
  2884=>"111111111",
  2885=>"011011011",
  2886=>"101101110",
  2887=>"111100010",
  2888=>"110111001",
  2889=>"001110100",
  2890=>"101101011",
  2891=>"101100000",
  2892=>"010111110",
  2893=>"111100100",
  2894=>"110000101",
  2895=>"001000101",
  2896=>"010101011",
  2897=>"101100011",
  2898=>"101001110",
  2899=>"111100111",
  2900=>"010010011",
  2901=>"110001010",
  2902=>"010001100",
  2903=>"011100010",
  2904=>"011101010",
  2905=>"110110001",
  2906=>"001001101",
  2907=>"000000100",
  2908=>"110000001",
  2909=>"110110111",
  2910=>"000001110",
  2911=>"101000000",
  2912=>"111111101",
  2913=>"100111110",
  2914=>"000100011",
  2915=>"000010101",
  2916=>"110010011",
  2917=>"101010010",
  2918=>"100111110",
  2919=>"110100110",
  2920=>"000110010",
  2921=>"000010001",
  2922=>"110010000",
  2923=>"001111101",
  2924=>"011111110",
  2925=>"110010011",
  2926=>"000001010",
  2927=>"011010001",
  2928=>"110100000",
  2929=>"001000011",
  2930=>"000001110",
  2931=>"010111111",
  2932=>"111111100",
  2933=>"111011110",
  2934=>"000010111",
  2935=>"100000100",
  2936=>"100011010",
  2937=>"010010101",
  2938=>"001111101",
  2939=>"000010001",
  2940=>"101000000",
  2941=>"111111000",
  2942=>"100000111",
  2943=>"111111111",
  2944=>"100001111",
  2945=>"001110110",
  2946=>"000000111",
  2947=>"000001101",
  2948=>"100001010",
  2949=>"010111011",
  2950=>"010100010",
  2951=>"101000100",
  2952=>"110101110",
  2953=>"010100110",
  2954=>"000010000",
  2955=>"011100000",
  2956=>"111001011",
  2957=>"011111010",
  2958=>"000110010",
  2959=>"111111111",
  2960=>"000001100",
  2961=>"110100100",
  2962=>"100000111",
  2963=>"001111010",
  2964=>"110001010",
  2965=>"100011001",
  2966=>"110010110",
  2967=>"011110010",
  2968=>"000010010",
  2969=>"111000100",
  2970=>"101001000",
  2971=>"000000100",
  2972=>"011101011",
  2973=>"010000001",
  2974=>"011001110",
  2975=>"000001111",
  2976=>"110101100",
  2977=>"100000100",
  2978=>"100010011",
  2979=>"000100010",
  2980=>"110100100",
  2981=>"001000101",
  2982=>"111110000",
  2983=>"110010000",
  2984=>"011010100",
  2985=>"101100010",
  2986=>"011100101",
  2987=>"101001111",
  2988=>"000000010",
  2989=>"100001110",
  2990=>"010111111",
  2991=>"111010110",
  2992=>"010010111",
  2993=>"011010111",
  2994=>"111001110",
  2995=>"101001011",
  2996=>"111110001",
  2997=>"010101010",
  2998=>"111010011",
  2999=>"111111110",
  3000=>"110000101",
  3001=>"011111111",
  3002=>"000001000",
  3003=>"010110000",
  3004=>"010101000",
  3005=>"010100000",
  3006=>"000010101",
  3007=>"101111010",
  3008=>"110000110",
  3009=>"000001011",
  3010=>"101110110",
  3011=>"111111100",
  3012=>"110100001",
  3013=>"100010100",
  3014=>"010000111",
  3015=>"001111011",
  3016=>"000011101",
  3017=>"101001011",
  3018=>"011011011",
  3019=>"100110100",
  3020=>"011111111",
  3021=>"000000110",
  3022=>"001100000",
  3023=>"100110001",
  3024=>"001111111",
  3025=>"110110111",
  3026=>"111011011",
  3027=>"111011110",
  3028=>"000101011",
  3029=>"100000101",
  3030=>"110000010",
  3031=>"000011111",
  3032=>"000001101",
  3033=>"110111110",
  3034=>"011010000",
  3035=>"010100000",
  3036=>"111101110",
  3037=>"111011100",
  3038=>"010010010",
  3039=>"110011000",
  3040=>"000101001",
  3041=>"110101001",
  3042=>"000000111",
  3043=>"011100100",
  3044=>"111000010",
  3045=>"101000111",
  3046=>"111001010",
  3047=>"101110000",
  3048=>"000010111",
  3049=>"001000100",
  3050=>"101010100",
  3051=>"110001101",
  3052=>"100100000",
  3053=>"101100101",
  3054=>"100101000",
  3055=>"110010101",
  3056=>"101110100",
  3057=>"111011110",
  3058=>"011100111",
  3059=>"011100001",
  3060=>"010101010",
  3061=>"000101110",
  3062=>"010111000",
  3063=>"011001100",
  3064=>"010111001",
  3065=>"000000011",
  3066=>"000011000",
  3067=>"100011011",
  3068=>"110010100",
  3069=>"110011100",
  3070=>"100001001",
  3071=>"000000000",
  3072=>"000111111",
  3073=>"001111010",
  3074=>"100011011",
  3075=>"110100100",
  3076=>"110001001",
  3077=>"000011101",
  3078=>"010100111",
  3079=>"000000011",
  3080=>"010110011",
  3081=>"000101001",
  3082=>"000000110",
  3083=>"000011101",
  3084=>"111110100",
  3085=>"001010111",
  3086=>"010101010",
  3087=>"000110001",
  3088=>"001100111",
  3089=>"010111010",
  3090=>"100001000",
  3091=>"101001001",
  3092=>"000101010",
  3093=>"001010011",
  3094=>"100001000",
  3095=>"000010111",
  3096=>"001100110",
  3097=>"010111111",
  3098=>"110001111",
  3099=>"000110011",
  3100=>"000011110",
  3101=>"110000100",
  3102=>"101010110",
  3103=>"010101001",
  3104=>"000011100",
  3105=>"111111110",
  3106=>"101001001",
  3107=>"000100110",
  3108=>"101111000",
  3109=>"011010111",
  3110=>"100000111",
  3111=>"110011110",
  3112=>"001001000",
  3113=>"100111101",
  3114=>"110100010",
  3115=>"101000010",
  3116=>"110000100",
  3117=>"011110001",
  3118=>"110010000",
  3119=>"010001110",
  3120=>"000110110",
  3121=>"101101000",
  3122=>"001100010",
  3123=>"110001101",
  3124=>"111001001",
  3125=>"100011110",
  3126=>"000001100",
  3127=>"000011100",
  3128=>"000110010",
  3129=>"111110011",
  3130=>"110000000",
  3131=>"110000100",
  3132=>"000001100",
  3133=>"110100100",
  3134=>"111101111",
  3135=>"000101100",
  3136=>"100011110",
  3137=>"001111001",
  3138=>"010100111",
  3139=>"000110000",
  3140=>"111101100",
  3141=>"111010010",
  3142=>"100110010",
  3143=>"010110100",
  3144=>"001110000",
  3145=>"110011010",
  3146=>"110101010",
  3147=>"001101011",
  3148=>"111001001",
  3149=>"100010000",
  3150=>"001011001",
  3151=>"000100101",
  3152=>"110000010",
  3153=>"000011000",
  3154=>"001000101",
  3155=>"011001000",
  3156=>"111110000",
  3157=>"000011001",
  3158=>"100001010",
  3159=>"010100001",
  3160=>"111100010",
  3161=>"100101100",
  3162=>"111101010",
  3163=>"101100110",
  3164=>"000011111",
  3165=>"110101001",
  3166=>"011110010",
  3167=>"000100000",
  3168=>"100111010",
  3169=>"100100101",
  3170=>"110000010",
  3171=>"000101110",
  3172=>"001011111",
  3173=>"101110110",
  3174=>"000100000",
  3175=>"111101000",
  3176=>"001001111",
  3177=>"111101010",
  3178=>"101011011",
  3179=>"000001001",
  3180=>"011001101",
  3181=>"100001101",
  3182=>"010010100",
  3183=>"111010011",
  3184=>"101100010",
  3185=>"001110000",
  3186=>"101010101",
  3187=>"101100110",
  3188=>"100011001",
  3189=>"001101101",
  3190=>"111100001",
  3191=>"010100101",
  3192=>"000010111",
  3193=>"111111001",
  3194=>"011100000",
  3195=>"101111011",
  3196=>"000001010",
  3197=>"111000000",
  3198=>"110010011",
  3199=>"000000011",
  3200=>"101011110",
  3201=>"110100001",
  3202=>"011001011",
  3203=>"011011111",
  3204=>"000101110",
  3205=>"001001111",
  3206=>"010100100",
  3207=>"100011101",
  3208=>"101001100",
  3209=>"000000101",
  3210=>"011100111",
  3211=>"010100001",
  3212=>"000000100",
  3213=>"001111101",
  3214=>"111110111",
  3215=>"000100100",
  3216=>"001100001",
  3217=>"100110010",
  3218=>"111000000",
  3219=>"101000010",
  3220=>"001011111",
  3221=>"101010011",
  3222=>"001111101",
  3223=>"001011101",
  3224=>"111011110",
  3225=>"010100000",
  3226=>"000010110",
  3227=>"111000000",
  3228=>"100000000",
  3229=>"001010011",
  3230=>"111100010",
  3231=>"001111000",
  3232=>"000010000",
  3233=>"111100011",
  3234=>"111101101",
  3235=>"001110001",
  3236=>"010011001",
  3237=>"000010011",
  3238=>"010111100",
  3239=>"000110110",
  3240=>"101111001",
  3241=>"101100101",
  3242=>"010101010",
  3243=>"010010100",
  3244=>"110110001",
  3245=>"001011011",
  3246=>"011111110",
  3247=>"001010101",
  3248=>"100011010",
  3249=>"100100010",
  3250=>"011000100",
  3251=>"010111101",
  3252=>"001101111",
  3253=>"001100110",
  3254=>"011011100",
  3255=>"010010000",
  3256=>"011001000",
  3257=>"111011101",
  3258=>"111100000",
  3259=>"010100010",
  3260=>"111100000",
  3261=>"100011110",
  3262=>"000100010",
  3263=>"001100010",
  3264=>"000010100",
  3265=>"111101011",
  3266=>"001001000",
  3267=>"000110100",
  3268=>"110100010",
  3269=>"110100011",
  3270=>"110011000",
  3271=>"001110000",
  3272=>"000100000",
  3273=>"001001001",
  3274=>"110001011",
  3275=>"011100000",
  3276=>"001100110",
  3277=>"011110000",
  3278=>"100010000",
  3279=>"101111000",
  3280=>"101001101",
  3281=>"001100011",
  3282=>"010001010",
  3283=>"001101100",
  3284=>"000100100",
  3285=>"101110111",
  3286=>"001110100",
  3287=>"111001111",
  3288=>"100000111",
  3289=>"000101011",
  3290=>"011111111",
  3291=>"011000001",
  3292=>"000001101",
  3293=>"101001000",
  3294=>"001110101",
  3295=>"011111100",
  3296=>"100101111",
  3297=>"010111111",
  3298=>"010011111",
  3299=>"001000000",
  3300=>"001111011",
  3301=>"001100100",
  3302=>"011100000",
  3303=>"011011011",
  3304=>"000000101",
  3305=>"010101000",
  3306=>"101100111",
  3307=>"010000000",
  3308=>"110000011",
  3309=>"001110010",
  3310=>"000111111",
  3311=>"111011000",
  3312=>"011100111",
  3313=>"110001110",
  3314=>"011001100",
  3315=>"111111111",
  3316=>"111010111",
  3317=>"000010010",
  3318=>"011110000",
  3319=>"000110101",
  3320=>"000001000",
  3321=>"000111110",
  3322=>"011111111",
  3323=>"001100001",
  3324=>"101010111",
  3325=>"101010101",
  3326=>"101101110",
  3327=>"100000001",
  3328=>"000011010",
  3329=>"011011111",
  3330=>"111011001",
  3331=>"100110000",
  3332=>"100011011",
  3333=>"110001001",
  3334=>"000111110",
  3335=>"011000101",
  3336=>"011101000",
  3337=>"000000010",
  3338=>"111100111",
  3339=>"000010010",
  3340=>"110100100",
  3341=>"000010111",
  3342=>"010100010",
  3343=>"000110100",
  3344=>"001001100",
  3345=>"001111010",
  3346=>"010101010",
  3347=>"111011101",
  3348=>"000101111",
  3349=>"110000110",
  3350=>"101011100",
  3351=>"011001001",
  3352=>"101101001",
  3353=>"011010111",
  3354=>"111001100",
  3355=>"011101111",
  3356=>"110101101",
  3357=>"111100110",
  3358=>"101110000",
  3359=>"010010011",
  3360=>"011100001",
  3361=>"101111010",
  3362=>"001101100",
  3363=>"111000111",
  3364=>"001110011",
  3365=>"000111101",
  3366=>"000100000",
  3367=>"100001000",
  3368=>"011110011",
  3369=>"100111111",
  3370=>"111011110",
  3371=>"110011011",
  3372=>"001010001",
  3373=>"100000000",
  3374=>"001000010",
  3375=>"010000000",
  3376=>"000111101",
  3377=>"100001010",
  3378=>"100111111",
  3379=>"010011110",
  3380=>"000000000",
  3381=>"010111000",
  3382=>"000001011",
  3383=>"100111000",
  3384=>"111101111",
  3385=>"100100101",
  3386=>"000011001",
  3387=>"111010100",
  3388=>"101010010",
  3389=>"111111010",
  3390=>"111111010",
  3391=>"010100011",
  3392=>"010011000",
  3393=>"111010000",
  3394=>"100111010",
  3395=>"101011000",
  3396=>"010011111",
  3397=>"110001001",
  3398=>"001000010",
  3399=>"101010001",
  3400=>"011010111",
  3401=>"110001000",
  3402=>"111101011",
  3403=>"101101111",
  3404=>"110100010",
  3405=>"111000010",
  3406=>"100000000",
  3407=>"010111100",
  3408=>"101100000",
  3409=>"110111000",
  3410=>"000101011",
  3411=>"111101001",
  3412=>"111000001",
  3413=>"001110101",
  3414=>"111000001",
  3415=>"010011110",
  3416=>"000111000",
  3417=>"111010011",
  3418=>"001001000",
  3419=>"000100100",
  3420=>"010000011",
  3421=>"110001000",
  3422=>"111011000",
  3423=>"000001110",
  3424=>"101110110",
  3425=>"101100000",
  3426=>"111101111",
  3427=>"000101000",
  3428=>"110011100",
  3429=>"011111011",
  3430=>"011101100",
  3431=>"010110011",
  3432=>"110001011",
  3433=>"110001000",
  3434=>"111100111",
  3435=>"101011001",
  3436=>"000000110",
  3437=>"101110000",
  3438=>"110011000",
  3439=>"111000011",
  3440=>"101100001",
  3441=>"110100011",
  3442=>"011111011",
  3443=>"101000011",
  3444=>"001010001",
  3445=>"110001110",
  3446=>"000010101",
  3447=>"100000010",
  3448=>"011000000",
  3449=>"100000011",
  3450=>"101001000",
  3451=>"001011101",
  3452=>"001001000",
  3453=>"111000000",
  3454=>"100001101",
  3455=>"001000110",
  3456=>"101100101",
  3457=>"100001111",
  3458=>"000010011",
  3459=>"011100100",
  3460=>"001110011",
  3461=>"100010111",
  3462=>"101000100",
  3463=>"010001000",
  3464=>"101101111",
  3465=>"000011101",
  3466=>"100000110",
  3467=>"010110011",
  3468=>"110000101",
  3469=>"010000110",
  3470=>"001100001",
  3471=>"100010000",
  3472=>"101111110",
  3473=>"001100101",
  3474=>"000111000",
  3475=>"111000101",
  3476=>"011010100",
  3477=>"111111110",
  3478=>"010100000",
  3479=>"101000110",
  3480=>"100000011",
  3481=>"100010001",
  3482=>"100010101",
  3483=>"100000000",
  3484=>"010001100",
  3485=>"001110011",
  3486=>"110010000",
  3487=>"001000011",
  3488=>"101011001",
  3489=>"011011111",
  3490=>"010001111",
  3491=>"101101000",
  3492=>"001000101",
  3493=>"011000000",
  3494=>"001011100",
  3495=>"010111010",
  3496=>"010010111",
  3497=>"101001001",
  3498=>"000011000",
  3499=>"111110111",
  3500=>"011010100",
  3501=>"101100000",
  3502=>"111010110",
  3503=>"010011111",
  3504=>"111010000",
  3505=>"011110111",
  3506=>"010010001",
  3507=>"010110111",
  3508=>"100001110",
  3509=>"110001111",
  3510=>"101111000",
  3511=>"000100001",
  3512=>"111001001",
  3513=>"110110101",
  3514=>"100011001",
  3515=>"111011000",
  3516=>"000101000",
  3517=>"101110111",
  3518=>"111101110",
  3519=>"101100001",
  3520=>"100101010",
  3521=>"110101111",
  3522=>"100000001",
  3523=>"001001000",
  3524=>"001101011",
  3525=>"111011110",
  3526=>"010101011",
  3527=>"000001010",
  3528=>"101001100",
  3529=>"001101001",
  3530=>"100010111",
  3531=>"011100110",
  3532=>"001011111",
  3533=>"110010110",
  3534=>"001001110",
  3535=>"100110001",
  3536=>"000011000",
  3537=>"110101010",
  3538=>"000101100",
  3539=>"011000110",
  3540=>"010101000",
  3541=>"011000010",
  3542=>"101010101",
  3543=>"010111100",
  3544=>"100001111",
  3545=>"011010111",
  3546=>"110100111",
  3547=>"011010111",
  3548=>"111110001",
  3549=>"000000010",
  3550=>"000100111",
  3551=>"001111100",
  3552=>"101111011",
  3553=>"010011000",
  3554=>"001010101",
  3555=>"010110000",
  3556=>"111101100",
  3557=>"110001101",
  3558=>"000110000",
  3559=>"010000000",
  3560=>"111011110",
  3561=>"000011011",
  3562=>"010101010",
  3563=>"000000110",
  3564=>"101001000",
  3565=>"011010000",
  3566=>"000010001",
  3567=>"101100101",
  3568=>"000110001",
  3569=>"001100101",
  3570=>"000010000",
  3571=>"000011111",
  3572=>"101000010",
  3573=>"011011001",
  3574=>"000001111",
  3575=>"100011001",
  3576=>"101111110",
  3577=>"011101010",
  3578=>"101110000",
  3579=>"110110011",
  3580=>"110111111",
  3581=>"010100100",
  3582=>"001010000",
  3583=>"000001010",
  3584=>"010000101",
  3585=>"000101110",
  3586=>"011100111",
  3587=>"001111010",
  3588=>"011011010",
  3589=>"101010001",
  3590=>"000010101",
  3591=>"000111010",
  3592=>"000001111",
  3593=>"010110001",
  3594=>"100011111",
  3595=>"010011101",
  3596=>"000001001",
  3597=>"111101101",
  3598=>"000111001",
  3599=>"111101100",
  3600=>"100001011",
  3601=>"010100110",
  3602=>"100011111",
  3603=>"111101011",
  3604=>"111101001",
  3605=>"001010100",
  3606=>"111010000",
  3607=>"110110110",
  3608=>"100010000",
  3609=>"100110110",
  3610=>"100010111",
  3611=>"111101001",
  3612=>"110011111",
  3613=>"101100010",
  3614=>"110100100",
  3615=>"101101001",
  3616=>"110110011",
  3617=>"000110111",
  3618=>"001111110",
  3619=>"000010001",
  3620=>"110010110",
  3621=>"110000100",
  3622=>"110101010",
  3623=>"010011111",
  3624=>"101001101",
  3625=>"001101110",
  3626=>"001001101",
  3627=>"110110010",
  3628=>"110111111",
  3629=>"001011000",
  3630=>"000000101",
  3631=>"101100100",
  3632=>"010111101",
  3633=>"001010100",
  3634=>"110110000",
  3635=>"001101000",
  3636=>"011111100",
  3637=>"111011000",
  3638=>"111101101",
  3639=>"101010100",
  3640=>"010010011",
  3641=>"101010111",
  3642=>"111000001",
  3643=>"111101011",
  3644=>"001101110",
  3645=>"101010000",
  3646=>"000110110",
  3647=>"110101011",
  3648=>"000000010",
  3649=>"010000010",
  3650=>"001101011",
  3651=>"100101110",
  3652=>"011001111",
  3653=>"011111110",
  3654=>"110110001",
  3655=>"100011101",
  3656=>"101000010",
  3657=>"111111101",
  3658=>"010111010",
  3659=>"101101010",
  3660=>"011011011",
  3661=>"010111011",
  3662=>"111011100",
  3663=>"111111100",
  3664=>"011111010",
  3665=>"000111011",
  3666=>"100001100",
  3667=>"001011011",
  3668=>"101100010",
  3669=>"101101001",
  3670=>"111111110",
  3671=>"000110001",
  3672=>"000110111",
  3673=>"011110001",
  3674=>"101001010",
  3675=>"001101000",
  3676=>"111001011",
  3677=>"000000001",
  3678=>"010000100",
  3679=>"100000110",
  3680=>"000011100",
  3681=>"101101010",
  3682=>"111111000",
  3683=>"011101101",
  3684=>"111111100",
  3685=>"100110001",
  3686=>"111100010",
  3687=>"011010100",
  3688=>"110000010",
  3689=>"101000000",
  3690=>"110010101",
  3691=>"000001100",
  3692=>"011100111",
  3693=>"111000100",
  3694=>"001000010",
  3695=>"010000001",
  3696=>"101010101",
  3697=>"000100011",
  3698=>"011000110",
  3699=>"101111011",
  3700=>"100010101",
  3701=>"100100010",
  3702=>"010100111",
  3703=>"100000010",
  3704=>"101101111",
  3705=>"110111111",
  3706=>"111110001",
  3707=>"000101111",
  3708=>"010110010",
  3709=>"100100011",
  3710=>"001001000",
  3711=>"101110010",
  3712=>"010011101",
  3713=>"111011010",
  3714=>"001001100",
  3715=>"001011110",
  3716=>"000111111",
  3717=>"000111010",
  3718=>"100111100",
  3719=>"110110011",
  3720=>"101110000",
  3721=>"001010010",
  3722=>"010000100",
  3723=>"101100011",
  3724=>"001100101",
  3725=>"011010101",
  3726=>"011011000",
  3727=>"001010000",
  3728=>"001000101",
  3729=>"011111100",
  3730=>"100110111",
  3731=>"100111011",
  3732=>"011011011",
  3733=>"101100101",
  3734=>"011011000",
  3735=>"111000101",
  3736=>"110000011",
  3737=>"111011100",
  3738=>"110100111",
  3739=>"110101100",
  3740=>"000110101",
  3741=>"100011011",
  3742=>"111100110",
  3743=>"110110010",
  3744=>"000010000",
  3745=>"110101000",
  3746=>"101111010",
  3747=>"001000101",
  3748=>"110111011",
  3749=>"110010000",
  3750=>"110110100",
  3751=>"101111111",
  3752=>"000001000",
  3753=>"111110111",
  3754=>"000101100",
  3755=>"000011001",
  3756=>"000000000",
  3757=>"000101011",
  3758=>"101001000",
  3759=>"011000001",
  3760=>"111010010",
  3761=>"111011000",
  3762=>"011101001",
  3763=>"000001100",
  3764=>"011011000",
  3765=>"100000100",
  3766=>"001110101",
  3767=>"001101001",
  3768=>"101000001",
  3769=>"101000101",
  3770=>"110000010",
  3771=>"000101111",
  3772=>"110110000",
  3773=>"000110000",
  3774=>"000110010",
  3775=>"111100011",
  3776=>"000100010",
  3777=>"101010001",
  3778=>"100001100",
  3779=>"001010001",
  3780=>"100010110",
  3781=>"100111000",
  3782=>"000000011",
  3783=>"011110010",
  3784=>"011000000",
  3785=>"110110001",
  3786=>"110010011",
  3787=>"001010011",
  3788=>"110100000",
  3789=>"000101101",
  3790=>"111011001",
  3791=>"111000101",
  3792=>"100100000",
  3793=>"110001111",
  3794=>"110001110",
  3795=>"100001100",
  3796=>"000000000",
  3797=>"110000010",
  3798=>"001010100",
  3799=>"011101101",
  3800=>"100011101",
  3801=>"100000110",
  3802=>"001101111",
  3803=>"011110000",
  3804=>"010010111",
  3805=>"011110101",
  3806=>"100111100",
  3807=>"000100101",
  3808=>"000001110",
  3809=>"001100111",
  3810=>"100011000",
  3811=>"110000100",
  3812=>"000111111",
  3813=>"110101001",
  3814=>"110100100",
  3815=>"111000011",
  3816=>"000001101",
  3817=>"001000111",
  3818=>"111111101",
  3819=>"101110101",
  3820=>"001100100",
  3821=>"111001000",
  3822=>"000010101",
  3823=>"011101100",
  3824=>"110110101",
  3825=>"111010101",
  3826=>"101000000",
  3827=>"001010110",
  3828=>"010101111",
  3829=>"100100110",
  3830=>"011111001",
  3831=>"011100110",
  3832=>"111100110",
  3833=>"111001011",
  3834=>"001101101",
  3835=>"010001000",
  3836=>"010010000",
  3837=>"101001000",
  3838=>"110100001",
  3839=>"000010001",
  3840=>"001000010",
  3841=>"010110000",
  3842=>"111110111",
  3843=>"100111101",
  3844=>"111110010",
  3845=>"001111111",
  3846=>"001011010",
  3847=>"100001011",
  3848=>"101101010",
  3849=>"001111011",
  3850=>"100101010",
  3851=>"001000110",
  3852=>"101100011",
  3853=>"001010100",
  3854=>"100100111",
  3855=>"100010111",
  3856=>"001011111",
  3857=>"110001010",
  3858=>"111110111",
  3859=>"000101001",
  3860=>"000100010",
  3861=>"010010001",
  3862=>"010010111",
  3863=>"100011101",
  3864=>"011000100",
  3865=>"010010100",
  3866=>"111110011",
  3867=>"110110000",
  3868=>"011110110",
  3869=>"000010100",
  3870=>"100101110",
  3871=>"111100111",
  3872=>"011111011",
  3873=>"010111001",
  3874=>"100110011",
  3875=>"001001010",
  3876=>"110100010",
  3877=>"010011010",
  3878=>"001111100",
  3879=>"011101111",
  3880=>"011010100",
  3881=>"101110110",
  3882=>"101100010",
  3883=>"110100001",
  3884=>"100010111",
  3885=>"000011110",
  3886=>"001111101",
  3887=>"100111110",
  3888=>"010001111",
  3889=>"010010011",
  3890=>"101000101",
  3891=>"101101100",
  3892=>"011100100",
  3893=>"000001000",
  3894=>"010010000",
  3895=>"011000000",
  3896=>"101110111",
  3897=>"001110101",
  3898=>"000000010",
  3899=>"011101111",
  3900=>"010111001",
  3901=>"101100100",
  3902=>"110001100",
  3903=>"110111110",
  3904=>"110111010",
  3905=>"000100000",
  3906=>"000010101",
  3907=>"001101110",
  3908=>"101110010",
  3909=>"011001101",
  3910=>"110100111",
  3911=>"110000100",
  3912=>"101001011",
  3913=>"000110100",
  3914=>"011000011",
  3915=>"010010010",
  3916=>"110111110",
  3917=>"101001000",
  3918=>"110111100",
  3919=>"100100110",
  3920=>"101000001",
  3921=>"100011001",
  3922=>"110010000",
  3923=>"000100110",
  3924=>"011010010",
  3925=>"011010000",
  3926=>"001000010",
  3927=>"111011010",
  3928=>"000100000",
  3929=>"100011011",
  3930=>"001010000",
  3931=>"001111110",
  3932=>"000111101",
  3933=>"100110010",
  3934=>"000111001",
  3935=>"000000010",
  3936=>"111010000",
  3937=>"010111101",
  3938=>"110010111",
  3939=>"100011101",
  3940=>"100001110",
  3941=>"011000001",
  3942=>"010011011",
  3943=>"011111000",
  3944=>"011101111",
  3945=>"100110111",
  3946=>"001100110",
  3947=>"010100110",
  3948=>"110110011",
  3949=>"011110110",
  3950=>"001011111",
  3951=>"100001011",
  3952=>"010011011",
  3953=>"011111111",
  3954=>"001110011",
  3955=>"001010010",
  3956=>"010110001",
  3957=>"101111111",
  3958=>"100100001",
  3959=>"100000001",
  3960=>"110110010",
  3961=>"101001000",
  3962=>"111101000",
  3963=>"011000000",
  3964=>"100000001",
  3965=>"111011110",
  3966=>"100010001",
  3967=>"100000000",
  3968=>"111001010",
  3969=>"110111011",
  3970=>"011011000",
  3971=>"111100101",
  3972=>"100001000",
  3973=>"010000001",
  3974=>"000111110",
  3975=>"101000111",
  3976=>"101001111",
  3977=>"111000111",
  3978=>"111100010",
  3979=>"101001000",
  3980=>"001011001",
  3981=>"011001100",
  3982=>"000001110",
  3983=>"001110001",
  3984=>"010110100",
  3985=>"011110001",
  3986=>"011010000",
  3987=>"000011011",
  3988=>"101111111",
  3989=>"101101100",
  3990=>"100000011",
  3991=>"011101011",
  3992=>"101000000",
  3993=>"010001010",
  3994=>"010111010",
  3995=>"000000011",
  3996=>"000101010",
  3997=>"101111011",
  3998=>"010001010",
  3999=>"000010010",
  4000=>"001000011",
  4001=>"011111111",
  4002=>"101000111",
  4003=>"111110101",
  4004=>"100101100",
  4005=>"100110001",
  4006=>"010010111",
  4007=>"111000001",
  4008=>"011011001",
  4009=>"101111111",
  4010=>"010101100",
  4011=>"011100100",
  4012=>"000001010",
  4013=>"110011111",
  4014=>"000000000",
  4015=>"100111000",
  4016=>"101001010",
  4017=>"101110101",
  4018=>"000000000",
  4019=>"001000000",
  4020=>"100000010",
  4021=>"000000100",
  4022=>"111010100",
  4023=>"101000010",
  4024=>"111010101",
  4025=>"111011111",
  4026=>"100001010",
  4027=>"001101100",
  4028=>"111001001",
  4029=>"101000000",
  4030=>"111111111",
  4031=>"100100000",
  4032=>"110110000",
  4033=>"111000011",
  4034=>"111100100",
  4035=>"111001011",
  4036=>"101111011",
  4037=>"101100010",
  4038=>"010011001",
  4039=>"111001001",
  4040=>"101111001",
  4041=>"001111000",
  4042=>"011111101",
  4043=>"101000110",
  4044=>"000010000",
  4045=>"100011010",
  4046=>"111111110",
  4047=>"001000001",
  4048=>"010111111",
  4049=>"110000110",
  4050=>"010000000",
  4051=>"110111101",
  4052=>"010010111",
  4053=>"111001010",
  4054=>"000101000",
  4055=>"011110010",
  4056=>"110101100",
  4057=>"010111011",
  4058=>"101100100",
  4059=>"101001010",
  4060=>"110011011",
  4061=>"111101000",
  4062=>"110111111",
  4063=>"011110110",
  4064=>"001000011",
  4065=>"000011111",
  4066=>"000010101",
  4067=>"001010100",
  4068=>"000001010",
  4069=>"000011111",
  4070=>"000110111",
  4071=>"111000101",
  4072=>"011001001",
  4073=>"010110111",
  4074=>"001000010",
  4075=>"001111011",
  4076=>"100101100",
  4077=>"000101111",
  4078=>"101010101",
  4079=>"011011000",
  4080=>"000100100",
  4081=>"110101000",
  4082=>"001011111",
  4083=>"101111100",
  4084=>"000100111",
  4085=>"100110111",
  4086=>"101010110",
  4087=>"001110110",
  4088=>"001111110",
  4089=>"011011011",
  4090=>"000111010",
  4091=>"001000000",
  4092=>"001010010",
  4093=>"101110101",
  4094=>"111111100",
  4095=>"111111010",
  4096=>"110110111",
  4097=>"100001111",
  4098=>"101110011",
  4099=>"101011010",
  4100=>"010001011",
  4101=>"001111111",
  4102=>"010111010",
  4103=>"000101010",
  4104=>"001100101",
  4105=>"101001100",
  4106=>"011101010",
  4107=>"001001000",
  4108=>"011001111",
  4109=>"010001101",
  4110=>"011111000",
  4111=>"000100001",
  4112=>"101110111",
  4113=>"111010000",
  4114=>"110101010",
  4115=>"011010111",
  4116=>"011110110",
  4117=>"110110010",
  4118=>"000010110",
  4119=>"011101110",
  4120=>"100101000",
  4121=>"010110011",
  4122=>"011011011",
  4123=>"101000011",
  4124=>"101110110",
  4125=>"010110100",
  4126=>"101010010",
  4127=>"000100110",
  4128=>"010000101",
  4129=>"101111101",
  4130=>"001011110",
  4131=>"101010101",
  4132=>"110111011",
  4133=>"011010111",
  4134=>"100101110",
  4135=>"101011100",
  4136=>"010111010",
  4137=>"010011110",
  4138=>"101010101",
  4139=>"011100111",
  4140=>"011000010",
  4141=>"011001011",
  4142=>"010010100",
  4143=>"001111010",
  4144=>"101101110",
  4145=>"101010110",
  4146=>"111111110",
  4147=>"001100010",
  4148=>"111111111",
  4149=>"100000011",
  4150=>"010001011",
  4151=>"001001111",
  4152=>"000101001",
  4153=>"011010101",
  4154=>"001000100",
  4155=>"100000100",
  4156=>"100110000",
  4157=>"010100010",
  4158=>"100000000",
  4159=>"010101000",
  4160=>"110010111",
  4161=>"101010010",
  4162=>"100111100",
  4163=>"010110010",
  4164=>"101001100",
  4165=>"001001010",
  4166=>"111110010",
  4167=>"100110000",
  4168=>"101000010",
  4169=>"100011101",
  4170=>"010101000",
  4171=>"101100111",
  4172=>"111011011",
  4173=>"110001101",
  4174=>"001101100",
  4175=>"010111010",
  4176=>"100001100",
  4177=>"110010111",
  4178=>"111111001",
  4179=>"101101111",
  4180=>"111101101",
  4181=>"101110111",
  4182=>"110011001",
  4183=>"101110011",
  4184=>"011111001",
  4185=>"010101111",
  4186=>"001001001",
  4187=>"110011010",
  4188=>"000111010",
  4189=>"011100111",
  4190=>"010001111",
  4191=>"110111010",
  4192=>"010001111",
  4193=>"010100000",
  4194=>"110001101",
  4195=>"000001001",
  4196=>"001010110",
  4197=>"111011000",
  4198=>"010011101",
  4199=>"010001101",
  4200=>"010101010",
  4201=>"001100100",
  4202=>"000000110",
  4203=>"010110110",
  4204=>"100000110",
  4205=>"011001100",
  4206=>"110001100",
  4207=>"110010010",
  4208=>"011110000",
  4209=>"101101101",
  4210=>"111001000",
  4211=>"110011101",
  4212=>"000110000",
  4213=>"100000100",
  4214=>"111100010",
  4215=>"000101100",
  4216=>"001011001",
  4217=>"100111110",
  4218=>"111111011",
  4219=>"110110010",
  4220=>"000010110",
  4221=>"101100100",
  4222=>"010011010",
  4223=>"010001100",
  4224=>"001000101",
  4225=>"001101100",
  4226=>"011101111",
  4227=>"000101100",
  4228=>"001111100",
  4229=>"110101000",
  4230=>"011100000",
  4231=>"111111110",
  4232=>"010000010",
  4233=>"000000101",
  4234=>"110011011",
  4235=>"011011111",
  4236=>"001001110",
  4237=>"011010010",
  4238=>"011100001",
  4239=>"101000110",
  4240=>"110111000",
  4241=>"100100000",
  4242=>"111111010",
  4243=>"011000000",
  4244=>"100000001",
  4245=>"011000011",
  4246=>"101110111",
  4247=>"011000101",
  4248=>"011111001",
  4249=>"110000001",
  4250=>"100000011",
  4251=>"100001111",
  4252=>"100011110",
  4253=>"000100011",
  4254=>"000100101",
  4255=>"101010011",
  4256=>"011010100",
  4257=>"111100110",
  4258=>"110001000",
  4259=>"000001010",
  4260=>"001100110",
  4261=>"110000110",
  4262=>"010100010",
  4263=>"110000100",
  4264=>"111011101",
  4265=>"110000001",
  4266=>"000100101",
  4267=>"111011100",
  4268=>"010000001",
  4269=>"100011111",
  4270=>"110111111",
  4271=>"001111011",
  4272=>"000011111",
  4273=>"011101111",
  4274=>"001010000",
  4275=>"011001001",
  4276=>"011111010",
  4277=>"010111111",
  4278=>"101110111",
  4279=>"011001011",
  4280=>"001100111",
  4281=>"101000011",
  4282=>"000010100",
  4283=>"100101111",
  4284=>"110001011",
  4285=>"110001101",
  4286=>"101011011",
  4287=>"100011110",
  4288=>"011100010",
  4289=>"000100100",
  4290=>"010100110",
  4291=>"111111010",
  4292=>"000100100",
  4293=>"011100011",
  4294=>"111100100",
  4295=>"110010000",
  4296=>"000100100",
  4297=>"000101111",
  4298=>"011111110",
  4299=>"010001100",
  4300=>"010111110",
  4301=>"101011001",
  4302=>"000100000",
  4303=>"001000000",
  4304=>"111000001",
  4305=>"000100000",
  4306=>"000111010",
  4307=>"100111100",
  4308=>"111110110",
  4309=>"110101001",
  4310=>"000000001",
  4311=>"011000000",
  4312=>"011001100",
  4313=>"111011010",
  4314=>"000001010",
  4315=>"111100101",
  4316=>"100011100",
  4317=>"000110100",
  4318=>"111101001",
  4319=>"111111111",
  4320=>"001110100",
  4321=>"001100001",
  4322=>"101101110",
  4323=>"110000010",
  4324=>"110101111",
  4325=>"001111111",
  4326=>"000110000",
  4327=>"100110110",
  4328=>"010010010",
  4329=>"001111011",
  4330=>"011110100",
  4331=>"110101001",
  4332=>"000111011",
  4333=>"100110001",
  4334=>"100101110",
  4335=>"111001111",
  4336=>"011111001",
  4337=>"110000010",
  4338=>"000100000",
  4339=>"000101000",
  4340=>"111000010",
  4341=>"000111100",
  4342=>"010011110",
  4343=>"000000100",
  4344=>"010000010",
  4345=>"010011101",
  4346=>"010000111",
  4347=>"010110100",
  4348=>"000010101",
  4349=>"100100110",
  4350=>"011111010",
  4351=>"100010000",
  4352=>"101001110",
  4353=>"101001101",
  4354=>"011011111",
  4355=>"010110000",
  4356=>"011010011",
  4357=>"010101000",
  4358=>"010101001",
  4359=>"001101110",
  4360=>"110111110",
  4361=>"110000100",
  4362=>"100011001",
  4363=>"110010101",
  4364=>"001010101",
  4365=>"001111100",
  4366=>"000011001",
  4367=>"001010100",
  4368=>"000101000",
  4369=>"001001001",
  4370=>"010100101",
  4371=>"100110001",
  4372=>"101000011",
  4373=>"110001011",
  4374=>"010000001",
  4375=>"110110001",
  4376=>"000110000",
  4377=>"100101110",
  4378=>"111110001",
  4379=>"001111111",
  4380=>"111010000",
  4381=>"011111010",
  4382=>"000111011",
  4383=>"111011110",
  4384=>"100000010",
  4385=>"111000100",
  4386=>"110101100",
  4387=>"000100010",
  4388=>"110010000",
  4389=>"110010000",
  4390=>"011000010",
  4391=>"100011001",
  4392=>"001001100",
  4393=>"111010100",
  4394=>"110000000",
  4395=>"010101010",
  4396=>"011001100",
  4397=>"000000000",
  4398=>"100101000",
  4399=>"010011011",
  4400=>"110011101",
  4401=>"101110110",
  4402=>"101101100",
  4403=>"010001101",
  4404=>"000100110",
  4405=>"000100001",
  4406=>"001111000",
  4407=>"111101111",
  4408=>"000001100",
  4409=>"100010011",
  4410=>"101101101",
  4411=>"001101000",
  4412=>"010001111",
  4413=>"110101100",
  4414=>"011000101",
  4415=>"011010001",
  4416=>"010000001",
  4417=>"000010000",
  4418=>"010111101",
  4419=>"010111010",
  4420=>"000101011",
  4421=>"001001101",
  4422=>"111110110",
  4423=>"011000100",
  4424=>"000000011",
  4425=>"101001011",
  4426=>"111111101",
  4427=>"111101110",
  4428=>"110111110",
  4429=>"001001110",
  4430=>"011011110",
  4431=>"111010001",
  4432=>"110101111",
  4433=>"101110111",
  4434=>"010010001",
  4435=>"000000100",
  4436=>"001010101",
  4437=>"101011100",
  4438=>"000011001",
  4439=>"110100000",
  4440=>"001010111",
  4441=>"011110111",
  4442=>"100111100",
  4443=>"011101001",
  4444=>"000000000",
  4445=>"010000000",
  4446=>"001100000",
  4447=>"101011000",
  4448=>"100100101",
  4449=>"011011110",
  4450=>"000001011",
  4451=>"101111110",
  4452=>"101000010",
  4453=>"100001001",
  4454=>"101011110",
  4455=>"111011000",
  4456=>"100001000",
  4457=>"100100010",
  4458=>"110101011",
  4459=>"011100100",
  4460=>"001000010",
  4461=>"110001000",
  4462=>"010000100",
  4463=>"001000010",
  4464=>"000000011",
  4465=>"100110110",
  4466=>"111011000",
  4467=>"001110101",
  4468=>"100000000",
  4469=>"010101010",
  4470=>"001001011",
  4471=>"011110000",
  4472=>"100000001",
  4473=>"011111101",
  4474=>"101011010",
  4475=>"000111000",
  4476=>"110011101",
  4477=>"001010011",
  4478=>"011011101",
  4479=>"111100101",
  4480=>"111010001",
  4481=>"010010101",
  4482=>"010111100",
  4483=>"101110100",
  4484=>"101010110",
  4485=>"000110111",
  4486=>"110110100",
  4487=>"100100001",
  4488=>"101000101",
  4489=>"100101110",
  4490=>"110111101",
  4491=>"010001100",
  4492=>"110111001",
  4493=>"010010101",
  4494=>"000011111",
  4495=>"011001100",
  4496=>"101011100",
  4497=>"001001011",
  4498=>"000111000",
  4499=>"110011111",
  4500=>"010100001",
  4501=>"010111100",
  4502=>"000100000",
  4503=>"101001010",
  4504=>"110011110",
  4505=>"000111010",
  4506=>"101100110",
  4507=>"100010100",
  4508=>"011101001",
  4509=>"100001100",
  4510=>"010111101",
  4511=>"111111101",
  4512=>"000001000",
  4513=>"100000011",
  4514=>"011111000",
  4515=>"000001001",
  4516=>"010010111",
  4517=>"101011010",
  4518=>"101111111",
  4519=>"110111000",
  4520=>"101101111",
  4521=>"010111010",
  4522=>"011110110",
  4523=>"100010011",
  4524=>"111110100",
  4525=>"111101011",
  4526=>"010001111",
  4527=>"001111001",
  4528=>"000111000",
  4529=>"000111010",
  4530=>"100011100",
  4531=>"111101111",
  4532=>"100100101",
  4533=>"101000111",
  4534=>"101001111",
  4535=>"101100110",
  4536=>"110001001",
  4537=>"010111010",
  4538=>"011010110",
  4539=>"111110101",
  4540=>"001000000",
  4541=>"010010010",
  4542=>"001011111",
  4543=>"011000001",
  4544=>"001011000",
  4545=>"000010001",
  4546=>"111010100",
  4547=>"011100110",
  4548=>"100010110",
  4549=>"100110100",
  4550=>"101001001",
  4551=>"000111010",
  4552=>"110010100",
  4553=>"110110101",
  4554=>"001011000",
  4555=>"010100100",
  4556=>"011001001",
  4557=>"001100111",
  4558=>"001110011",
  4559=>"000100111",
  4560=>"011001101",
  4561=>"110101000",
  4562=>"110111111",
  4563=>"000010000",
  4564=>"011010101",
  4565=>"111101011",
  4566=>"001000100",
  4567=>"010111111",
  4568=>"010111010",
  4569=>"010111011",
  4570=>"010111101",
  4571=>"001000000",
  4572=>"100011101",
  4573=>"110000111",
  4574=>"001110011",
  4575=>"101100101",
  4576=>"111001111",
  4577=>"100001111",
  4578=>"101011001",
  4579=>"000000000",
  4580=>"110011100",
  4581=>"111001011",
  4582=>"010110101",
  4583=>"011101111",
  4584=>"101101010",
  4585=>"000101101",
  4586=>"000101111",
  4587=>"100001010",
  4588=>"111010010",
  4589=>"011101011",
  4590=>"011010010",
  4591=>"000011001",
  4592=>"000101000",
  4593=>"101001000",
  4594=>"000100110",
  4595=>"100010101",
  4596=>"101110101",
  4597=>"000110110",
  4598=>"110111111",
  4599=>"000000011",
  4600=>"010110101",
  4601=>"001011110",
  4602=>"000001000",
  4603=>"000011111",
  4604=>"011110101",
  4605=>"111111001",
  4606=>"100010000",
  4607=>"111110011",
  4608=>"000011001",
  4609=>"011010011",
  4610=>"011111000",
  4611=>"011000001",
  4612=>"011001101",
  4613=>"000100110",
  4614=>"000010010",
  4615=>"001111011",
  4616=>"010010011",
  4617=>"011011100",
  4618=>"000000110",
  4619=>"100000010",
  4620=>"011000110",
  4621=>"100100100",
  4622=>"000100101",
  4623=>"011001001",
  4624=>"000111110",
  4625=>"000010110",
  4626=>"000000000",
  4627=>"111000110",
  4628=>"111010000",
  4629=>"101100001",
  4630=>"000100110",
  4631=>"000001101",
  4632=>"011010100",
  4633=>"110101001",
  4634=>"000001001",
  4635=>"100100001",
  4636=>"100011110",
  4637=>"110110010",
  4638=>"001001011",
  4639=>"000000000",
  4640=>"101100110",
  4641=>"000100011",
  4642=>"110001101",
  4643=>"100100010",
  4644=>"110100111",
  4645=>"010110100",
  4646=>"111000000",
  4647=>"000110010",
  4648=>"000011001",
  4649=>"101011111",
  4650=>"001110100",
  4651=>"101010011",
  4652=>"000010111",
  4653=>"001011000",
  4654=>"011010001",
  4655=>"111101101",
  4656=>"110101101",
  4657=>"101011100",
  4658=>"101110000",
  4659=>"000100001",
  4660=>"110111010",
  4661=>"111011001",
  4662=>"010110010",
  4663=>"010110101",
  4664=>"110111000",
  4665=>"101110110",
  4666=>"101001011",
  4667=>"111001000",
  4668=>"000000110",
  4669=>"111001011",
  4670=>"101000011",
  4671=>"101000100",
  4672=>"000001000",
  4673=>"000100111",
  4674=>"000100000",
  4675=>"101100010",
  4676=>"111010010",
  4677=>"100011101",
  4678=>"100000010",
  4679=>"011111000",
  4680=>"010111010",
  4681=>"000001001",
  4682=>"101111101",
  4683=>"011101010",
  4684=>"111000010",
  4685=>"000010001",
  4686=>"100110000",
  4687=>"010010010",
  4688=>"000010101",
  4689=>"000001010",
  4690=>"100011011",
  4691=>"011101001",
  4692=>"001011110",
  4693=>"101010011",
  4694=>"000100000",
  4695=>"001111101",
  4696=>"111111111",
  4697=>"101101000",
  4698=>"010101101",
  4699=>"011001110",
  4700=>"010010100",
  4701=>"011010110",
  4702=>"000010110",
  4703=>"110101110",
  4704=>"001101001",
  4705=>"000111010",
  4706=>"010100111",
  4707=>"111111000",
  4708=>"011001111",
  4709=>"001100000",
  4710=>"100010000",
  4711=>"111000110",
  4712=>"100000101",
  4713=>"110000111",
  4714=>"110010111",
  4715=>"110010001",
  4716=>"000000011",
  4717=>"110111111",
  4718=>"100100100",
  4719=>"010110111",
  4720=>"001010001",
  4721=>"010011000",
  4722=>"001111000",
  4723=>"001000111",
  4724=>"010000101",
  4725=>"100011100",
  4726=>"111011010",
  4727=>"011001111",
  4728=>"111100001",
  4729=>"101010101",
  4730=>"111101110",
  4731=>"001100100",
  4732=>"110101100",
  4733=>"111110001",
  4734=>"011110010",
  4735=>"000100101",
  4736=>"011001110",
  4737=>"100001111",
  4738=>"010010001",
  4739=>"000101000",
  4740=>"011101100",
  4741=>"110010000",
  4742=>"011001011",
  4743=>"010101011",
  4744=>"010100111",
  4745=>"111101001",
  4746=>"101110001",
  4747=>"111111110",
  4748=>"100101101",
  4749=>"011000100",
  4750=>"000101001",
  4751=>"000001111",
  4752=>"110011010",
  4753=>"011110111",
  4754=>"111111101",
  4755=>"101110110",
  4756=>"100001111",
  4757=>"111010010",
  4758=>"000000111",
  4759=>"001001000",
  4760=>"110010100",
  4761=>"011110110",
  4762=>"010011001",
  4763=>"010000000",
  4764=>"101110001",
  4765=>"101000010",
  4766=>"110111000",
  4767=>"011011100",
  4768=>"111101010",
  4769=>"111011001",
  4770=>"001111100",
  4771=>"111010111",
  4772=>"000100101",
  4773=>"010111100",
  4774=>"001000000",
  4775=>"000000100",
  4776=>"010101101",
  4777=>"010000110",
  4778=>"011101100",
  4779=>"101100001",
  4780=>"011101111",
  4781=>"100101111",
  4782=>"010101001",
  4783=>"000100101",
  4784=>"000110011",
  4785=>"010000101",
  4786=>"000000001",
  4787=>"011100001",
  4788=>"100010110",
  4789=>"010111100",
  4790=>"011011111",
  4791=>"111100111",
  4792=>"101000000",
  4793=>"000001100",
  4794=>"000000101",
  4795=>"110111110",
  4796=>"101100101",
  4797=>"110001000",
  4798=>"100100011",
  4799=>"000011001",
  4800=>"000010000",
  4801=>"000000111",
  4802=>"110111100",
  4803=>"111000110",
  4804=>"010001111",
  4805=>"000100000",
  4806=>"111000011",
  4807=>"000000010",
  4808=>"101001100",
  4809=>"010111110",
  4810=>"011000001",
  4811=>"010111001",
  4812=>"000001110",
  4813=>"110111100",
  4814=>"101010001",
  4815=>"110000010",
  4816=>"101010010",
  4817=>"000011111",
  4818=>"011011000",
  4819=>"001000000",
  4820=>"111011000",
  4821=>"010101101",
  4822=>"101100011",
  4823=>"001010000",
  4824=>"010100100",
  4825=>"100110011",
  4826=>"101011001",
  4827=>"101001010",
  4828=>"110111001",
  4829=>"110100010",
  4830=>"010111111",
  4831=>"101111011",
  4832=>"111101000",
  4833=>"101101000",
  4834=>"100100011",
  4835=>"001100011",
  4836=>"111010101",
  4837=>"110011001",
  4838=>"101001101",
  4839=>"011101110",
  4840=>"101001101",
  4841=>"110100110",
  4842=>"011010011",
  4843=>"100111101",
  4844=>"000101111",
  4845=>"000010011",
  4846=>"010010100",
  4847=>"010001001",
  4848=>"000101010",
  4849=>"010000001",
  4850=>"100000000",
  4851=>"001101010",
  4852=>"101111101",
  4853=>"110110011",
  4854=>"000101001",
  4855=>"011011010",
  4856=>"101101100",
  4857=>"000110001",
  4858=>"111000101",
  4859=>"101100011",
  4860=>"010000000",
  4861=>"101100000",
  4862=>"101110110",
  4863=>"000000011",
  4864=>"110011001",
  4865=>"110100100",
  4866=>"110100010",
  4867=>"011111010",
  4868=>"001001110",
  4869=>"000111010",
  4870=>"001110110",
  4871=>"000001111",
  4872=>"001000110",
  4873=>"100110110",
  4874=>"000110011",
  4875=>"011101010",
  4876=>"111100000",
  4877=>"011100100",
  4878=>"001101001",
  4879=>"011100100",
  4880=>"101110111",
  4881=>"101101100",
  4882=>"110100010",
  4883=>"001100001",
  4884=>"010110001",
  4885=>"001001101",
  4886=>"110001001",
  4887=>"000011000",
  4888=>"111101011",
  4889=>"010010101",
  4890=>"100111110",
  4891=>"001111111",
  4892=>"011011010",
  4893=>"110100001",
  4894=>"101100100",
  4895=>"110111000",
  4896=>"010001100",
  4897=>"011001000",
  4898=>"010110110",
  4899=>"101111010",
  4900=>"011011110",
  4901=>"000100000",
  4902=>"000111111",
  4903=>"011011000",
  4904=>"110101000",
  4905=>"101010001",
  4906=>"100101010",
  4907=>"111010101",
  4908=>"001100101",
  4909=>"101010001",
  4910=>"111000101",
  4911=>"001010100",
  4912=>"000110100",
  4913=>"100111010",
  4914=>"001010011",
  4915=>"010000011",
  4916=>"100100001",
  4917=>"101010000",
  4918=>"000000010",
  4919=>"001001011",
  4920=>"101111100",
  4921=>"000010111",
  4922=>"110101101",
  4923=>"000001001",
  4924=>"001010101",
  4925=>"011001101",
  4926=>"001100001",
  4927=>"011100110",
  4928=>"100110010",
  4929=>"001101100",
  4930=>"101100000",
  4931=>"111110000",
  4932=>"011110100",
  4933=>"110111000",
  4934=>"000101000",
  4935=>"100101101",
  4936=>"111000010",
  4937=>"100111111",
  4938=>"101011110",
  4939=>"000000001",
  4940=>"111110101",
  4941=>"001001011",
  4942=>"100011010",
  4943=>"010001000",
  4944=>"001010110",
  4945=>"011010101",
  4946=>"001111100",
  4947=>"000100110",
  4948=>"000100000",
  4949=>"111111001",
  4950=>"110000101",
  4951=>"011010111",
  4952=>"101111100",
  4953=>"000000010",
  4954=>"001011000",
  4955=>"101001001",
  4956=>"111000001",
  4957=>"110111110",
  4958=>"010111100",
  4959=>"000000001",
  4960=>"010101101",
  4961=>"000000000",
  4962=>"010000011",
  4963=>"111110101",
  4964=>"111010101",
  4965=>"011010001",
  4966=>"100001110",
  4967=>"011100000",
  4968=>"100000010",
  4969=>"101011000",
  4970=>"001000000",
  4971=>"011010101",
  4972=>"100111001",
  4973=>"011100011",
  4974=>"101011010",
  4975=>"111011101",
  4976=>"011100100",
  4977=>"110100111",
  4978=>"001010111",
  4979=>"000000100",
  4980=>"011011000",
  4981=>"000010000",
  4982=>"110101110",
  4983=>"100010100",
  4984=>"111100101",
  4985=>"001101010",
  4986=>"101100010",
  4987=>"110101010",
  4988=>"011010110",
  4989=>"111111000",
  4990=>"001110000",
  4991=>"010010110",
  4992=>"011011000",
  4993=>"011001001",
  4994=>"000101000",
  4995=>"000000011",
  4996=>"010010101",
  4997=>"111111110",
  4998=>"111011100",
  4999=>"010000000",
  5000=>"000001111",
  5001=>"010110100",
  5002=>"110000000",
  5003=>"111110011",
  5004=>"011100000",
  5005=>"000001110",
  5006=>"000001101",
  5007=>"111011111",
  5008=>"000000010",
  5009=>"011001110",
  5010=>"000000000",
  5011=>"110100101",
  5012=>"001111001",
  5013=>"011110110",
  5014=>"010111101",
  5015=>"011000110",
  5016=>"000111000",
  5017=>"101101000",
  5018=>"110000101",
  5019=>"001000001",
  5020=>"010101101",
  5021=>"000110111",
  5022=>"110011111",
  5023=>"101101010",
  5024=>"100110110",
  5025=>"001011011",
  5026=>"111001000",
  5027=>"000011010",
  5028=>"001010110",
  5029=>"011110001",
  5030=>"001000001",
  5031=>"010101110",
  5032=>"101111110",
  5033=>"000101110",
  5034=>"111111000",
  5035=>"111000100",
  5036=>"100000011",
  5037=>"011000010",
  5038=>"100010011",
  5039=>"111101000",
  5040=>"010010001",
  5041=>"111111011",
  5042=>"011100101",
  5043=>"100110110",
  5044=>"110000011",
  5045=>"100011111",
  5046=>"001001000",
  5047=>"010101011",
  5048=>"001111111",
  5049=>"101011010",
  5050=>"010110101",
  5051=>"001001010",
  5052=>"010001000",
  5053=>"011011100",
  5054=>"010000101",
  5055=>"000111000",
  5056=>"101000110",
  5057=>"100010010",
  5058=>"101011110",
  5059=>"010111010",
  5060=>"111110011",
  5061=>"000110110",
  5062=>"011001010",
  5063=>"100110100",
  5064=>"101011100",
  5065=>"110101000",
  5066=>"001110001",
  5067=>"011010001",
  5068=>"110010110",
  5069=>"001111000",
  5070=>"100010010",
  5071=>"010001010",
  5072=>"111110111",
  5073=>"100010011",
  5074=>"101111110",
  5075=>"100001010",
  5076=>"111001000",
  5077=>"110011000",
  5078=>"100000000",
  5079=>"110111111",
  5080=>"000110001",
  5081=>"110000000",
  5082=>"111001101",
  5083=>"011001101",
  5084=>"100101101",
  5085=>"000001000",
  5086=>"010101011",
  5087=>"001100111",
  5088=>"001010101",
  5089=>"101101100",
  5090=>"001000000",
  5091=>"110000011",
  5092=>"100000011",
  5093=>"011100111",
  5094=>"110111101",
  5095=>"110111111",
  5096=>"001010100",
  5097=>"100110111",
  5098=>"101101000",
  5099=>"111100100",
  5100=>"101011111",
  5101=>"111000010",
  5102=>"100100110",
  5103=>"001001111",
  5104=>"000101110",
  5105=>"100010110",
  5106=>"000111100",
  5107=>"001000111",
  5108=>"000001111",
  5109=>"100010100",
  5110=>"110100111",
  5111=>"010001110",
  5112=>"111000111",
  5113=>"101111001",
  5114=>"010001100",
  5115=>"011111010",
  5116=>"001100111",
  5117=>"100011010",
  5118=>"000010001",
  5119=>"000010010",
  5120=>"000011011",
  5121=>"011110100",
  5122=>"101101111",
  5123=>"010101100",
  5124=>"010001010",
  5125=>"001101011",
  5126=>"010100110",
  5127=>"000010100",
  5128=>"001000000",
  5129=>"001100011",
  5130=>"010010000",
  5131=>"110001101",
  5132=>"010010010",
  5133=>"000100010",
  5134=>"100101001",
  5135=>"001001001",
  5136=>"100011111",
  5137=>"100111001",
  5138=>"111001011",
  5139=>"100011100",
  5140=>"011110101",
  5141=>"110001100",
  5142=>"101101111",
  5143=>"100000010",
  5144=>"001110000",
  5145=>"101000100",
  5146=>"001000100",
  5147=>"101000010",
  5148=>"001011010",
  5149=>"011001101",
  5150=>"010010010",
  5151=>"110010100",
  5152=>"000010111",
  5153=>"110110101",
  5154=>"010110100",
  5155=>"001000101",
  5156=>"100000100",
  5157=>"111100011",
  5158=>"000100110",
  5159=>"111100010",
  5160=>"100110010",
  5161=>"001011000",
  5162=>"001101011",
  5163=>"000110100",
  5164=>"011110100",
  5165=>"000101111",
  5166=>"000001110",
  5167=>"111101011",
  5168=>"101111000",
  5169=>"100100011",
  5170=>"101010101",
  5171=>"101010011",
  5172=>"100010000",
  5173=>"010010000",
  5174=>"101110001",
  5175=>"001101101",
  5176=>"000101101",
  5177=>"001000001",
  5178=>"011001011",
  5179=>"110111101",
  5180=>"001100101",
  5181=>"000111100",
  5182=>"101100111",
  5183=>"000010110",
  5184=>"011100111",
  5185=>"011000000",
  5186=>"111100110",
  5187=>"000000100",
  5188=>"010100111",
  5189=>"001001110",
  5190=>"011110001",
  5191=>"000101101",
  5192=>"101100000",
  5193=>"000011011",
  5194=>"001010100",
  5195=>"001001011",
  5196=>"010101110",
  5197=>"111100101",
  5198=>"100010111",
  5199=>"010000010",
  5200=>"101000100",
  5201=>"001111110",
  5202=>"001111111",
  5203=>"110110011",
  5204=>"011111011",
  5205=>"111110100",
  5206=>"001111010",
  5207=>"000100100",
  5208=>"111110010",
  5209=>"101110110",
  5210=>"011101011",
  5211=>"111100010",
  5212=>"101011010",
  5213=>"000001001",
  5214=>"001010001",
  5215=>"001001001",
  5216=>"011111100",
  5217=>"111100010",
  5218=>"101110001",
  5219=>"010010101",
  5220=>"100010101",
  5221=>"111111000",
  5222=>"111000100",
  5223=>"000001100",
  5224=>"011110101",
  5225=>"001111101",
  5226=>"010001111",
  5227=>"101111110",
  5228=>"100010010",
  5229=>"011110100",
  5230=>"001110111",
  5231=>"000010001",
  5232=>"110001001",
  5233=>"100000100",
  5234=>"110110101",
  5235=>"101101010",
  5236=>"110101111",
  5237=>"010100011",
  5238=>"000001011",
  5239=>"101101010",
  5240=>"101000010",
  5241=>"101111101",
  5242=>"001111111",
  5243=>"111101110",
  5244=>"100101010",
  5245=>"010111111",
  5246=>"000010100",
  5247=>"110000010",
  5248=>"110010110",
  5249=>"000001100",
  5250=>"101010010",
  5251=>"001111101",
  5252=>"010101010",
  5253=>"000110000",
  5254=>"100110100",
  5255=>"000010101",
  5256=>"100100110",
  5257=>"000010011",
  5258=>"100000001",
  5259=>"010000001",
  5260=>"001000101",
  5261=>"111010010",
  5262=>"101110111",
  5263=>"100000011",
  5264=>"011011110",
  5265=>"000000100",
  5266=>"010000011",
  5267=>"010000000",
  5268=>"000111101",
  5269=>"011101100",
  5270=>"010111110",
  5271=>"101000100",
  5272=>"000010001",
  5273=>"001100101",
  5274=>"000110100",
  5275=>"010000101",
  5276=>"110010000",
  5277=>"011001000",
  5278=>"001000100",
  5279=>"001011001",
  5280=>"001111000",
  5281=>"011101111",
  5282=>"000000000",
  5283=>"010101111",
  5284=>"101101101",
  5285=>"011010101",
  5286=>"010011111",
  5287=>"101001100",
  5288=>"000010100",
  5289=>"111000000",
  5290=>"011111110",
  5291=>"011011101",
  5292=>"111011111",
  5293=>"000000000",
  5294=>"110000111",
  5295=>"110001110",
  5296=>"000000011",
  5297=>"010010010",
  5298=>"000001000",
  5299=>"001001010",
  5300=>"000111111",
  5301=>"101111100",
  5302=>"001011111",
  5303=>"111011010",
  5304=>"000100010",
  5305=>"100101110",
  5306=>"001101000",
  5307=>"111010000",
  5308=>"100100101",
  5309=>"001010000",
  5310=>"111000101",
  5311=>"111000011",
  5312=>"011100100",
  5313=>"011000101",
  5314=>"001110001",
  5315=>"101011001",
  5316=>"101100011",
  5317=>"100110010",
  5318=>"100001011",
  5319=>"100010011",
  5320=>"100011010",
  5321=>"110111000",
  5322=>"101100111",
  5323=>"011001110",
  5324=>"110110011",
  5325=>"111110101",
  5326=>"100111010",
  5327=>"111111111",
  5328=>"111110101",
  5329=>"111011000",
  5330=>"001110000",
  5331=>"100001010",
  5332=>"001011100",
  5333=>"111111110",
  5334=>"100010000",
  5335=>"010101001",
  5336=>"101010100",
  5337=>"101010000",
  5338=>"000001010",
  5339=>"000100000",
  5340=>"101111110",
  5341=>"001011110",
  5342=>"100110101",
  5343=>"010000110",
  5344=>"010110001",
  5345=>"111100011",
  5346=>"110011001",
  5347=>"110100000",
  5348=>"110101011",
  5349=>"001010010",
  5350=>"100010110",
  5351=>"011000010",
  5352=>"101110111",
  5353=>"100100010",
  5354=>"001001010",
  5355=>"010010011",
  5356=>"011110000",
  5357=>"111110111",
  5358=>"000100110",
  5359=>"000001000",
  5360=>"011000000",
  5361=>"001010100",
  5362=>"000100011",
  5363=>"011000011",
  5364=>"001010011",
  5365=>"100000110",
  5366=>"101001111",
  5367=>"111101111",
  5368=>"101000000",
  5369=>"100101110",
  5370=>"001011110",
  5371=>"100000110",
  5372=>"110011111",
  5373=>"000001011",
  5374=>"110011010",
  5375=>"000111110",
  5376=>"111110001",
  5377=>"001100001",
  5378=>"101111100",
  5379=>"011010110",
  5380=>"110010101",
  5381=>"011010011",
  5382=>"101101110",
  5383=>"101011101",
  5384=>"010100101",
  5385=>"100010000",
  5386=>"110010010",
  5387=>"100000100",
  5388=>"100101101",
  5389=>"011111000",
  5390=>"001110100",
  5391=>"100000110",
  5392=>"011010110",
  5393=>"000100111",
  5394=>"100000100",
  5395=>"111101000",
  5396=>"101110000",
  5397=>"011010010",
  5398=>"101111111",
  5399=>"000010110",
  5400=>"010100001",
  5401=>"011001111",
  5402=>"000000010",
  5403=>"110110000",
  5404=>"000000000",
  5405=>"110101110",
  5406=>"001110111",
  5407=>"110001111",
  5408=>"110011000",
  5409=>"101110101",
  5410=>"100110001",
  5411=>"110000000",
  5412=>"110111110",
  5413=>"100100010",
  5414=>"111010101",
  5415=>"011001010",
  5416=>"111101001",
  5417=>"101011110",
  5418=>"111010010",
  5419=>"100111010",
  5420=>"000000000",
  5421=>"000011000",
  5422=>"100000010",
  5423=>"000110001",
  5424=>"101101101",
  5425=>"111010010",
  5426=>"000111111",
  5427=>"011100101",
  5428=>"101111110",
  5429=>"100010000",
  5430=>"000111010",
  5431=>"011111100",
  5432=>"000000001",
  5433=>"011000011",
  5434=>"010101010",
  5435=>"010001000",
  5436=>"000000010",
  5437=>"001001001",
  5438=>"000010100",
  5439=>"001110111",
  5440=>"010000101",
  5441=>"011110000",
  5442=>"110100101",
  5443=>"101001101",
  5444=>"011110110",
  5445=>"110001001",
  5446=>"011011101",
  5447=>"110011011",
  5448=>"110110110",
  5449=>"110100101",
  5450=>"000111101",
  5451=>"000101000",
  5452=>"000111101",
  5453=>"010000010",
  5454=>"000100100",
  5455=>"100010000",
  5456=>"100110110",
  5457=>"011111100",
  5458=>"111100101",
  5459=>"001000101",
  5460=>"110000110",
  5461=>"100010100",
  5462=>"101100110",
  5463=>"100000100",
  5464=>"111010100",
  5465=>"000000001",
  5466=>"100001111",
  5467=>"001001000",
  5468=>"111111111",
  5469=>"001111100",
  5470=>"010111101",
  5471=>"001001000",
  5472=>"101111111",
  5473=>"111101011",
  5474=>"101101101",
  5475=>"001101100",
  5476=>"011001001",
  5477=>"101100110",
  5478=>"000111111",
  5479=>"001111100",
  5480=>"000000110",
  5481=>"000101001",
  5482=>"010101110",
  5483=>"101111001",
  5484=>"000111011",
  5485=>"101101101",
  5486=>"010101000",
  5487=>"100110011",
  5488=>"100101101",
  5489=>"111001100",
  5490=>"011010100",
  5491=>"110101001",
  5492=>"001110011",
  5493=>"011001000",
  5494=>"001100101",
  5495=>"111011110",
  5496=>"000100110",
  5497=>"111100010",
  5498=>"011100101",
  5499=>"101001000",
  5500=>"101011101",
  5501=>"111000111",
  5502=>"100100001",
  5503=>"010010010",
  5504=>"101111111",
  5505=>"101111111",
  5506=>"100101101",
  5507=>"111000101",
  5508=>"010110000",
  5509=>"010010101",
  5510=>"011110011",
  5511=>"101000110",
  5512=>"000110101",
  5513=>"000111011",
  5514=>"100011001",
  5515=>"101100000",
  5516=>"010101110",
  5517=>"101110000",
  5518=>"000000010",
  5519=>"001011001",
  5520=>"010000000",
  5521=>"000111001",
  5522=>"001011101",
  5523=>"010010000",
  5524=>"111001011",
  5525=>"110101000",
  5526=>"010000001",
  5527=>"110011111",
  5528=>"110010111",
  5529=>"001000111",
  5530=>"100110111",
  5531=>"111101010",
  5532=>"011100111",
  5533=>"000000100",
  5534=>"101010101",
  5535=>"010010010",
  5536=>"000101001",
  5537=>"010100111",
  5538=>"010011111",
  5539=>"100000000",
  5540=>"011111001",
  5541=>"000010000",
  5542=>"011011000",
  5543=>"110011110",
  5544=>"010010100",
  5545=>"110100000",
  5546=>"000001101",
  5547=>"101100000",
  5548=>"000100010",
  5549=>"010011101",
  5550=>"110000000",
  5551=>"011110011",
  5552=>"110101111",
  5553=>"111001010",
  5554=>"011100101",
  5555=>"011010000",
  5556=>"011100110",
  5557=>"110100001",
  5558=>"101000111",
  5559=>"000100000",
  5560=>"010101000",
  5561=>"000001101",
  5562=>"001111011",
  5563=>"010001001",
  5564=>"011101001",
  5565=>"001001101",
  5566=>"000000110",
  5567=>"001110111",
  5568=>"100001110",
  5569=>"100011101",
  5570=>"110011011",
  5571=>"110100101",
  5572=>"100101001",
  5573=>"101111111",
  5574=>"100011101",
  5575=>"100111001",
  5576=>"100100110",
  5577=>"000110111",
  5578=>"100100111",
  5579=>"111011101",
  5580=>"110111101",
  5581=>"101110100",
  5582=>"101001100",
  5583=>"111111011",
  5584=>"000100110",
  5585=>"001000100",
  5586=>"001101000",
  5587=>"101110110",
  5588=>"010001111",
  5589=>"000011000",
  5590=>"011010001",
  5591=>"010000100",
  5592=>"000000111",
  5593=>"110110001",
  5594=>"110011100",
  5595=>"110001101",
  5596=>"111111011",
  5597=>"001010010",
  5598=>"100110000",
  5599=>"011010100",
  5600=>"001101000",
  5601=>"110010110",
  5602=>"001100001",
  5603=>"110110011",
  5604=>"000100101",
  5605=>"011000011",
  5606=>"011000011",
  5607=>"111110000",
  5608=>"001001011",
  5609=>"110100111",
  5610=>"100101001",
  5611=>"001110010",
  5612=>"110110110",
  5613=>"000110001",
  5614=>"111101110",
  5615=>"111111001",
  5616=>"000101111",
  5617=>"110011101",
  5618=>"110000100",
  5619=>"110111001",
  5620=>"111100111",
  5621=>"000001100",
  5622=>"001100111",
  5623=>"101001111",
  5624=>"101110101",
  5625=>"101110010",
  5626=>"011000011",
  5627=>"111110000",
  5628=>"111111100",
  5629=>"110000100",
  5630=>"001111111",
  5631=>"111111000",
  5632=>"000101101",
  5633=>"100000100",
  5634=>"110011000",
  5635=>"001001010",
  5636=>"000011001",
  5637=>"110000001",
  5638=>"010101000",
  5639=>"010011100",
  5640=>"110110100",
  5641=>"101111001",
  5642=>"011010100",
  5643=>"000100000",
  5644=>"000101010",
  5645=>"001010010",
  5646=>"111001100",
  5647=>"001011000",
  5648=>"111000100",
  5649=>"000111110",
  5650=>"111011100",
  5651=>"111100110",
  5652=>"010011000",
  5653=>"000010111",
  5654=>"011000110",
  5655=>"010111110",
  5656=>"111110001",
  5657=>"010001011",
  5658=>"000110101",
  5659=>"110000001",
  5660=>"110101011",
  5661=>"010011110",
  5662=>"111111111",
  5663=>"110110110",
  5664=>"101100100",
  5665=>"110011100",
  5666=>"001011011",
  5667=>"001000001",
  5668=>"101101101",
  5669=>"111101101",
  5670=>"110001111",
  5671=>"100011011",
  5672=>"110101000",
  5673=>"001110000",
  5674=>"100110010",
  5675=>"100101110",
  5676=>"111101011",
  5677=>"100000111",
  5678=>"011011111",
  5679=>"100100100",
  5680=>"110001111",
  5681=>"110110000",
  5682=>"010100001",
  5683=>"101101010",
  5684=>"101011100",
  5685=>"010110111",
  5686=>"001101111",
  5687=>"011001011",
  5688=>"110011100",
  5689=>"100100100",
  5690=>"011010111",
  5691=>"000001010",
  5692=>"101001000",
  5693=>"100010101",
  5694=>"001110010",
  5695=>"110010000",
  5696=>"010001111",
  5697=>"000110010",
  5698=>"011101010",
  5699=>"001110111",
  5700=>"100000101",
  5701=>"011000001",
  5702=>"101001110",
  5703=>"010101010",
  5704=>"111010101",
  5705=>"000110111",
  5706=>"111101000",
  5707=>"110001101",
  5708=>"101111111",
  5709=>"001010011",
  5710=>"110010011",
  5711=>"010101110",
  5712=>"101100000",
  5713=>"101000101",
  5714=>"001110110",
  5715=>"000100011",
  5716=>"100111101",
  5717=>"110101010",
  5718=>"010101110",
  5719=>"000110101",
  5720=>"111001000",
  5721=>"100011000",
  5722=>"001000001",
  5723=>"000000011",
  5724=>"001101000",
  5725=>"011010001",
  5726=>"001010111",
  5727=>"101001110",
  5728=>"111010000",
  5729=>"011010000",
  5730=>"010010101",
  5731=>"101110000",
  5732=>"001000100",
  5733=>"001101000",
  5734=>"000000000",
  5735=>"110111101",
  5736=>"100010111",
  5737=>"011100001",
  5738=>"111100000",
  5739=>"110110110",
  5740=>"101011001",
  5741=>"001110101",
  5742=>"110011111",
  5743=>"110011110",
  5744=>"010100110",
  5745=>"000000001",
  5746=>"010111011",
  5747=>"111100001",
  5748=>"111100010",
  5749=>"101101000",
  5750=>"100101010",
  5751=>"101010111",
  5752=>"101011101",
  5753=>"000100110",
  5754=>"000111000",
  5755=>"010010111",
  5756=>"010010001",
  5757=>"011101011",
  5758=>"111001000",
  5759=>"100000100",
  5760=>"100110010",
  5761=>"001001011",
  5762=>"101011101",
  5763=>"010011101",
  5764=>"111100110",
  5765=>"110010100",
  5766=>"101001100",
  5767=>"111111000",
  5768=>"011100110",
  5769=>"111001110",
  5770=>"010000000",
  5771=>"011011000",
  5772=>"110000000",
  5773=>"000100110",
  5774=>"010101110",
  5775=>"111110011",
  5776=>"011111001",
  5777=>"000110111",
  5778=>"110000101",
  5779=>"001000100",
  5780=>"001000100",
  5781=>"001011011",
  5782=>"011000011",
  5783=>"101010000",
  5784=>"000110110",
  5785=>"011001111",
  5786=>"000111010",
  5787=>"011000001",
  5788=>"111110100",
  5789=>"111100101",
  5790=>"011011110",
  5791=>"010010110",
  5792=>"010000010",
  5793=>"000000001",
  5794=>"000000111",
  5795=>"101110100",
  5796=>"100001101",
  5797=>"010110001",
  5798=>"010010110",
  5799=>"100001001",
  5800=>"000001001",
  5801=>"111011111",
  5802=>"100101000",
  5803=>"101001000",
  5804=>"010001110",
  5805=>"111010110",
  5806=>"011001010",
  5807=>"001010111",
  5808=>"010001011",
  5809=>"110001111",
  5810=>"010000001",
  5811=>"101000011",
  5812=>"010110110",
  5813=>"101111001",
  5814=>"111101101",
  5815=>"100000001",
  5816=>"010100111",
  5817=>"111010110",
  5818=>"001011000",
  5819=>"110000111",
  5820=>"010001011",
  5821=>"000101001",
  5822=>"011100011",
  5823=>"011010010",
  5824=>"010101111",
  5825=>"100111000",
  5826=>"100011010",
  5827=>"100100100",
  5828=>"000000110",
  5829=>"100101111",
  5830=>"101011001",
  5831=>"101100010",
  5832=>"100010110",
  5833=>"010001100",
  5834=>"010011011",
  5835=>"010011010",
  5836=>"000011110",
  5837=>"011001100",
  5838=>"111011110",
  5839=>"000101000",
  5840=>"000011000",
  5841=>"100111011",
  5842=>"000010100",
  5843=>"010101111",
  5844=>"111101000",
  5845=>"000111100",
  5846=>"110010001",
  5847=>"000100111",
  5848=>"001101000",
  5849=>"110010100",
  5850=>"011111010",
  5851=>"100110111",
  5852=>"001001111",
  5853=>"101000000",
  5854=>"100100111",
  5855=>"001100101",
  5856=>"001001000",
  5857=>"100011011",
  5858=>"111011010",
  5859=>"110001000",
  5860=>"000000110",
  5861=>"100111001",
  5862=>"001010011",
  5863=>"000001010",
  5864=>"011110000",
  5865=>"110111011",
  5866=>"100010110",
  5867=>"001001000",
  5868=>"101110001",
  5869=>"111010001",
  5870=>"000011100",
  5871=>"010110110",
  5872=>"111101110",
  5873=>"011000111",
  5874=>"111110111",
  5875=>"110001100",
  5876=>"110010100",
  5877=>"100111001",
  5878=>"000000011",
  5879=>"000001101",
  5880=>"111000001",
  5881=>"000000001",
  5882=>"111110100",
  5883=>"110010010",
  5884=>"001011011",
  5885=>"000111110",
  5886=>"000100011",
  5887=>"010100001",
  5888=>"111010110",
  5889=>"001110011",
  5890=>"011011110",
  5891=>"110111001",
  5892=>"010000010",
  5893=>"100110110",
  5894=>"111111001",
  5895=>"011111001",
  5896=>"101111011",
  5897=>"100100101",
  5898=>"100010011",
  5899=>"010101001",
  5900=>"110101111",
  5901=>"011000011",
  5902=>"000000101",
  5903=>"111001101",
  5904=>"000110101",
  5905=>"110101000",
  5906=>"001000101",
  5907=>"011010010",
  5908=>"110011100",
  5909=>"101110010",
  5910=>"110000000",
  5911=>"110101111",
  5912=>"001011100",
  5913=>"010010101",
  5914=>"011000110",
  5915=>"001001000",
  5916=>"101100000",
  5917=>"101000000",
  5918=>"101100111",
  5919=>"011101011",
  5920=>"000110101",
  5921=>"101001010",
  5922=>"010101110",
  5923=>"010000010",
  5924=>"101101100",
  5925=>"100111101",
  5926=>"100110111",
  5927=>"001011111",
  5928=>"110100100",
  5929=>"111011100",
  5930=>"000000110",
  5931=>"010001001",
  5932=>"011111011",
  5933=>"000110001",
  5934=>"000010010",
  5935=>"000110101",
  5936=>"101010101",
  5937=>"111101001",
  5938=>"001001010",
  5939=>"100001010",
  5940=>"101010100",
  5941=>"111100011",
  5942=>"110011100",
  5943=>"011111101",
  5944=>"100001110",
  5945=>"001001000",
  5946=>"010101110",
  5947=>"101010010",
  5948=>"110000001",
  5949=>"101111011",
  5950=>"111001101",
  5951=>"011011101",
  5952=>"101110111",
  5953=>"011001110",
  5954=>"101110110",
  5955=>"010111101",
  5956=>"111110011",
  5957=>"010011101",
  5958=>"111011111",
  5959=>"101000111",
  5960=>"001000001",
  5961=>"011111011",
  5962=>"001111001",
  5963=>"011001101",
  5964=>"111101000",
  5965=>"001110001",
  5966=>"011001100",
  5967=>"000010010",
  5968=>"111001000",
  5969=>"111011001",
  5970=>"010000110",
  5971=>"111000011",
  5972=>"011111110",
  5973=>"100100110",
  5974=>"101001110",
  5975=>"011011010",
  5976=>"110010001",
  5977=>"101001100",
  5978=>"100111111",
  5979=>"000110010",
  5980=>"001001000",
  5981=>"101101100",
  5982=>"110100100",
  5983=>"000001001",
  5984=>"011001000",
  5985=>"111001101",
  5986=>"011110101",
  5987=>"011001010",
  5988=>"011100011",
  5989=>"101101011",
  5990=>"111110100",
  5991=>"101100111",
  5992=>"000111000",
  5993=>"000101111",
  5994=>"111000101",
  5995=>"000001101",
  5996=>"110000010",
  5997=>"100001101",
  5998=>"100000100",
  5999=>"011100010",
  6000=>"010001001",
  6001=>"110110111",
  6002=>"100011010",
  6003=>"000110011",
  6004=>"100110101",
  6005=>"110011101",
  6006=>"000011001",
  6007=>"110000010",
  6008=>"110011101",
  6009=>"111011000",
  6010=>"101110110",
  6011=>"010110101",
  6012=>"011000100",
  6013=>"110111100",
  6014=>"100000101",
  6015=>"011101111",
  6016=>"000001101",
  6017=>"110110010",
  6018=>"010111010",
  6019=>"011100100",
  6020=>"100101101",
  6021=>"000000010",
  6022=>"000111010",
  6023=>"111111001",
  6024=>"000100010",
  6025=>"000000000",
  6026=>"101100010",
  6027=>"000000010",
  6028=>"001111100",
  6029=>"001010010",
  6030=>"100100010",
  6031=>"000011100",
  6032=>"110011000",
  6033=>"100110111",
  6034=>"101000100",
  6035=>"101110010",
  6036=>"100011011",
  6037=>"101100001",
  6038=>"101110011",
  6039=>"001110011",
  6040=>"101111001",
  6041=>"011111011",
  6042=>"110010101",
  6043=>"000101011",
  6044=>"010101010",
  6045=>"111001000",
  6046=>"010011101",
  6047=>"110010100",
  6048=>"010110000",
  6049=>"001110111",
  6050=>"000001111",
  6051=>"000100010",
  6052=>"000000001",
  6053=>"110011101",
  6054=>"110101111",
  6055=>"111010001",
  6056=>"111001111",
  6057=>"000010101",
  6058=>"110010010",
  6059=>"101010001",
  6060=>"100001011",
  6061=>"111011001",
  6062=>"100001110",
  6063=>"110110011",
  6064=>"011100110",
  6065=>"111010110",
  6066=>"001101111",
  6067=>"001000000",
  6068=>"001111011",
  6069=>"000010001",
  6070=>"000001111",
  6071=>"000100101",
  6072=>"100001010",
  6073=>"011001101",
  6074=>"111011010",
  6075=>"010000101",
  6076=>"100000000",
  6077=>"100111101",
  6078=>"111101101",
  6079=>"000010101",
  6080=>"100100110",
  6081=>"001110000",
  6082=>"101111011",
  6083=>"110010001",
  6084=>"000111001",
  6085=>"011100001",
  6086=>"001011000",
  6087=>"101011111",
  6088=>"000001010",
  6089=>"010000000",
  6090=>"111001100",
  6091=>"000011111",
  6092=>"101010111",
  6093=>"001100000",
  6094=>"100011100",
  6095=>"000000111",
  6096=>"011110110",
  6097=>"111000100",
  6098=>"010100111",
  6099=>"011000000",
  6100=>"011111110",
  6101=>"110111000",
  6102=>"001000010",
  6103=>"000110001",
  6104=>"010010011",
  6105=>"010001000",
  6106=>"111100010",
  6107=>"001001110",
  6108=>"111100001",
  6109=>"110101111",
  6110=>"101010111",
  6111=>"000100000",
  6112=>"100111111",
  6113=>"000001001",
  6114=>"010000111",
  6115=>"100000111",
  6116=>"000100010",
  6117=>"011100110",
  6118=>"101100110",
  6119=>"001101000",
  6120=>"000111010",
  6121=>"101100110",
  6122=>"110100101",
  6123=>"001000101",
  6124=>"111101110",
  6125=>"011101101",
  6126=>"111001110",
  6127=>"111101001",
  6128=>"001000011",
  6129=>"101111000",
  6130=>"010011010",
  6131=>"001101010",
  6132=>"111011001",
  6133=>"001011101",
  6134=>"010010001",
  6135=>"101110100",
  6136=>"000111000",
  6137=>"011111001",
  6138=>"101001110",
  6139=>"101110011",
  6140=>"101100100",
  6141=>"001010110",
  6142=>"000101100",
  6143=>"101101110",
  6144=>"000010000",
  6145=>"011000000",
  6146=>"011010001",
  6147=>"001000011",
  6148=>"110100110",
  6149=>"101001010",
  6150=>"001101100",
  6151=>"111101100",
  6152=>"101011100",
  6153=>"000101101",
  6154=>"000011000",
  6155=>"111111011",
  6156=>"000011110",
  6157=>"101011100",
  6158=>"001100110",
  6159=>"001000011",
  6160=>"111101111",
  6161=>"000100011",
  6162=>"101111001",
  6163=>"011010011",
  6164=>"000111000",
  6165=>"011100100",
  6166=>"011000111",
  6167=>"111111010",
  6168=>"011000100",
  6169=>"111111011",
  6170=>"111111000",
  6171=>"100001101",
  6172=>"101001001",
  6173=>"010001110",
  6174=>"000000001",
  6175=>"100100111",
  6176=>"011110000",
  6177=>"110001111",
  6178=>"110000010",
  6179=>"101011001",
  6180=>"001000110",
  6181=>"010101010",
  6182=>"000011110",
  6183=>"001001000",
  6184=>"101001101",
  6185=>"000111010",
  6186=>"110100101",
  6187=>"010110001",
  6188=>"111100001",
  6189=>"001110011",
  6190=>"010111011",
  6191=>"010111110",
  6192=>"001101011",
  6193=>"111000000",
  6194=>"101010010",
  6195=>"101100000",
  6196=>"010110111",
  6197=>"111110001",
  6198=>"111001010",
  6199=>"101100000",
  6200=>"010011001",
  6201=>"010010110",
  6202=>"100111011",
  6203=>"110001011",
  6204=>"011010000",
  6205=>"010000001",
  6206=>"110101111",
  6207=>"011111101",
  6208=>"111010011",
  6209=>"111001011",
  6210=>"010101111",
  6211=>"101000110",
  6212=>"010101110",
  6213=>"111101111",
  6214=>"101100011",
  6215=>"110011010",
  6216=>"011001011",
  6217=>"101111100",
  6218=>"110111101",
  6219=>"100111001",
  6220=>"100100010",
  6221=>"010010000",
  6222=>"110001101",
  6223=>"001001010",
  6224=>"110111000",
  6225=>"101000111",
  6226=>"010110111",
  6227=>"100111111",
  6228=>"001100001",
  6229=>"001100010",
  6230=>"110101010",
  6231=>"000010101",
  6232=>"111011011",
  6233=>"100011110",
  6234=>"111010010",
  6235=>"111001111",
  6236=>"010110011",
  6237=>"000011111",
  6238=>"000110110",
  6239=>"011001111",
  6240=>"101001100",
  6241=>"001001111",
  6242=>"111000011",
  6243=>"000000111",
  6244=>"101110111",
  6245=>"011011110",
  6246=>"011111000",
  6247=>"100011000",
  6248=>"100111011",
  6249=>"010111001",
  6250=>"000100111",
  6251=>"000100100",
  6252=>"110001011",
  6253=>"000101000",
  6254=>"010101011",
  6255=>"111101000",
  6256=>"111111110",
  6257=>"110010010",
  6258=>"010011111",
  6259=>"010001010",
  6260=>"011001100",
  6261=>"111001111",
  6262=>"011000011",
  6263=>"101011011",
  6264=>"000101110",
  6265=>"100000101",
  6266=>"000001010",
  6267=>"111001000",
  6268=>"011011110",
  6269=>"110110100",
  6270=>"111111110",
  6271=>"000000100",
  6272=>"110100001",
  6273=>"001111000",
  6274=>"111101010",
  6275=>"010100101",
  6276=>"010100100",
  6277=>"101000111",
  6278=>"000101010",
  6279=>"011001100",
  6280=>"010001001",
  6281=>"001101001",
  6282=>"001010100",
  6283=>"010010100",
  6284=>"111101011",
  6285=>"101100011",
  6286=>"000101111",
  6287=>"010001011",
  6288=>"011000010",
  6289=>"001000000",
  6290=>"000001010",
  6291=>"011000011",
  6292=>"001111010",
  6293=>"111111011",
  6294=>"000010001",
  6295=>"100001000",
  6296=>"110011010",
  6297=>"010111100",
  6298=>"110101010",
  6299=>"110011011",
  6300=>"000000000",
  6301=>"010011100",
  6302=>"101110101",
  6303=>"100011111",
  6304=>"000001100",
  6305=>"100101001",
  6306=>"101010101",
  6307=>"010101001",
  6308=>"111001110",
  6309=>"000001110",
  6310=>"001100100",
  6311=>"101000110",
  6312=>"110111001",
  6313=>"100000111",
  6314=>"100001010",
  6315=>"111101001",
  6316=>"101001101",
  6317=>"110110000",
  6318=>"110001111",
  6319=>"110010011",
  6320=>"000001111",
  6321=>"100111100",
  6322=>"010000011",
  6323=>"111001000",
  6324=>"000010100",
  6325=>"110101110",
  6326=>"011111011",
  6327=>"000110100",
  6328=>"110100011",
  6329=>"110011111",
  6330=>"001001011",
  6331=>"111110111",
  6332=>"000100100",
  6333=>"001001110",
  6334=>"100011000",
  6335=>"001110001",
  6336=>"100111100",
  6337=>"100111000",
  6338=>"001010011",
  6339=>"110110100",
  6340=>"100111011",
  6341=>"101100000",
  6342=>"111011010",
  6343=>"111100000",
  6344=>"101011011",
  6345=>"111101010",
  6346=>"001011011",
  6347=>"010010000",
  6348=>"011010101",
  6349=>"000000010",
  6350=>"101111100",
  6351=>"001000111",
  6352=>"001110011",
  6353=>"101000111",
  6354=>"111001000",
  6355=>"101000001",
  6356=>"101101111",
  6357=>"101000100",
  6358=>"111000010",
  6359=>"101010011",
  6360=>"100110000",
  6361=>"101000011",
  6362=>"010001100",
  6363=>"000100010",
  6364=>"000010101",
  6365=>"000111010",
  6366=>"011101100",
  6367=>"101001001",
  6368=>"101000000",
  6369=>"001110101",
  6370=>"011011010",
  6371=>"101000001",
  6372=>"110001100",
  6373=>"001011000",
  6374=>"000100111",
  6375=>"000000000",
  6376=>"100000111",
  6377=>"010110010",
  6378=>"010010010",
  6379=>"001101000",
  6380=>"001111011",
  6381=>"010101101",
  6382=>"001011101",
  6383=>"000001001",
  6384=>"000110001",
  6385=>"001101111",
  6386=>"001011100",
  6387=>"000110011",
  6388=>"100001001",
  6389=>"110100110",
  6390=>"000111101",
  6391=>"011011010",
  6392=>"100000110",
  6393=>"100111100",
  6394=>"111010010",
  6395=>"101000011",
  6396=>"111001110",
  6397=>"011001110",
  6398=>"011011011",
  6399=>"011101011",
  6400=>"101000011",
  6401=>"110011100",
  6402=>"100111010",
  6403=>"111111000",
  6404=>"100000011",
  6405=>"001110001",
  6406=>"100100011",
  6407=>"101101010",
  6408=>"010001000",
  6409=>"101010010",
  6410=>"000011111",
  6411=>"100011010",
  6412=>"100011110",
  6413=>"010101000",
  6414=>"101101100",
  6415=>"101001000",
  6416=>"111001010",
  6417=>"111110110",
  6418=>"010010011",
  6419=>"110010011",
  6420=>"010011000",
  6421=>"011001010",
  6422=>"110011101",
  6423=>"000101111",
  6424=>"011111111",
  6425=>"001101111",
  6426=>"100001000",
  6427=>"011000110",
  6428=>"000110001",
  6429=>"100011000",
  6430=>"010001101",
  6431=>"000010000",
  6432=>"010001000",
  6433=>"011010101",
  6434=>"011110011",
  6435=>"100111010",
  6436=>"011110000",
  6437=>"100101001",
  6438=>"001001100",
  6439=>"101111001",
  6440=>"010110101",
  6441=>"111010110",
  6442=>"010101101",
  6443=>"001011011",
  6444=>"101011011",
  6445=>"010001100",
  6446=>"110001100",
  6447=>"101001000",
  6448=>"100000010",
  6449=>"111101111",
  6450=>"111100000",
  6451=>"001001110",
  6452=>"110000010",
  6453=>"110101011",
  6454=>"100101011",
  6455=>"000100111",
  6456=>"000100110",
  6457=>"000000010",
  6458=>"011010000",
  6459=>"111011101",
  6460=>"111000000",
  6461=>"000000110",
  6462=>"011100001",
  6463=>"111110111",
  6464=>"100001101",
  6465=>"100101010",
  6466=>"100000011",
  6467=>"100100100",
  6468=>"001011110",
  6469=>"101110100",
  6470=>"101010100",
  6471=>"001101001",
  6472=>"001011111",
  6473=>"001101111",
  6474=>"110010010",
  6475=>"011000111",
  6476=>"000001111",
  6477=>"101000000",
  6478=>"011111110",
  6479=>"100111001",
  6480=>"111110100",
  6481=>"011111010",
  6482=>"010101101",
  6483=>"111001000",
  6484=>"010111001",
  6485=>"110000111",
  6486=>"011100111",
  6487=>"011110000",
  6488=>"011100011",
  6489=>"000111110",
  6490=>"001110000",
  6491=>"110110111",
  6492=>"000111110",
  6493=>"100110100",
  6494=>"111101001",
  6495=>"100000110",
  6496=>"111000000",
  6497=>"101101100",
  6498=>"010000100",
  6499=>"000001100",
  6500=>"010111000",
  6501=>"111001111",
  6502=>"001111011",
  6503=>"110010111",
  6504=>"101101111",
  6505=>"110011000",
  6506=>"111111111",
  6507=>"000010011",
  6508=>"000001110",
  6509=>"001100010",
  6510=>"011110000",
  6511=>"000101011",
  6512=>"101011111",
  6513=>"011011111",
  6514=>"111000011",
  6515=>"101111000",
  6516=>"110111101",
  6517=>"111110110",
  6518=>"100110010",
  6519=>"111111111",
  6520=>"011001000",
  6521=>"011011101",
  6522=>"000101001",
  6523=>"110000111",
  6524=>"010001110",
  6525=>"111110001",
  6526=>"011101111",
  6527=>"101100100",
  6528=>"000110000",
  6529=>"011010010",
  6530=>"111111001",
  6531=>"100010000",
  6532=>"101011101",
  6533=>"100110101",
  6534=>"010100101",
  6535=>"011010010",
  6536=>"100001000",
  6537=>"111011101",
  6538=>"110110001",
  6539=>"111101111",
  6540=>"011101110",
  6541=>"000000110",
  6542=>"010101111",
  6543=>"110001000",
  6544=>"011001110",
  6545=>"001011101",
  6546=>"001101101",
  6547=>"111111101",
  6548=>"100101011",
  6549=>"100000000",
  6550=>"101000010",
  6551=>"101001110",
  6552=>"010010001",
  6553=>"100111101",
  6554=>"011100010",
  6555=>"100101111",
  6556=>"001011111",
  6557=>"110011010",
  6558=>"001100101",
  6559=>"101001110",
  6560=>"000011000",
  6561=>"000010011",
  6562=>"000011101",
  6563=>"000010000",
  6564=>"010111000",
  6565=>"000010000",
  6566=>"111101111",
  6567=>"011000001",
  6568=>"100111001",
  6569=>"101011111",
  6570=>"100010101",
  6571=>"011001011",
  6572=>"010100000",
  6573=>"101110001",
  6574=>"000101001",
  6575=>"011010010",
  6576=>"011011011",
  6577=>"010010111",
  6578=>"100110011",
  6579=>"111001111",
  6580=>"101001011",
  6581=>"110111100",
  6582=>"111101110",
  6583=>"001110111",
  6584=>"001100011",
  6585=>"110011100",
  6586=>"100101111",
  6587=>"110110111",
  6588=>"010010011",
  6589=>"010001001",
  6590=>"001110000",
  6591=>"001100000",
  6592=>"110111010",
  6593=>"111111011",
  6594=>"101110011",
  6595=>"100001111",
  6596=>"011110101",
  6597=>"000101111",
  6598=>"001111110",
  6599=>"101111010",
  6600=>"100001000",
  6601=>"001001101",
  6602=>"101000010",
  6603=>"100010101",
  6604=>"000111001",
  6605=>"001100110",
  6606=>"000010010",
  6607=>"110001101",
  6608=>"011110110",
  6609=>"111111111",
  6610=>"010010000",
  6611=>"011111110",
  6612=>"000001001",
  6613=>"010001101",
  6614=>"111011011",
  6615=>"001110100",
  6616=>"100000010",
  6617=>"001000010",
  6618=>"010101100",
  6619=>"100111000",
  6620=>"110000101",
  6621=>"001011101",
  6622=>"001010111",
  6623=>"000011010",
  6624=>"000011100",
  6625=>"011100111",
  6626=>"111101100",
  6627=>"110101001",
  6628=>"001101100",
  6629=>"110111111",
  6630=>"000100000",
  6631=>"111011100",
  6632=>"100110100",
  6633=>"000010010",
  6634=>"111110100",
  6635=>"000011110",
  6636=>"100100000",
  6637=>"111001110",
  6638=>"000010100",
  6639=>"001110100",
  6640=>"011000000",
  6641=>"111111101",
  6642=>"010100111",
  6643=>"000000011",
  6644=>"100111011",
  6645=>"111111111",
  6646=>"000010000",
  6647=>"110010100",
  6648=>"001100110",
  6649=>"010110010",
  6650=>"100011000",
  6651=>"000010010",
  6652=>"100101101",
  6653=>"000001111",
  6654=>"111100111",
  6655=>"011101101",
  6656=>"100111000",
  6657=>"001111001",
  6658=>"000000101",
  6659=>"001000010",
  6660=>"001001001",
  6661=>"110010101",
  6662=>"000100110",
  6663=>"000000100",
  6664=>"111010101",
  6665=>"110100011",
  6666=>"111111010",
  6667=>"011101010",
  6668=>"100010100",
  6669=>"110111010",
  6670=>"100011110",
  6671=>"000010100",
  6672=>"110010001",
  6673=>"101000000",
  6674=>"001000011",
  6675=>"111111010",
  6676=>"111111010",
  6677=>"101101010",
  6678=>"000011010",
  6679=>"101111011",
  6680=>"010001110",
  6681=>"100010010",
  6682=>"011011001",
  6683=>"001101111",
  6684=>"011110111",
  6685=>"111111101",
  6686=>"110111110",
  6687=>"001011110",
  6688=>"011101000",
  6689=>"110101011",
  6690=>"111100010",
  6691=>"010011101",
  6692=>"010111101",
  6693=>"111100011",
  6694=>"100100111",
  6695=>"110001010",
  6696=>"011100000",
  6697=>"100011110",
  6698=>"101111101",
  6699=>"001110111",
  6700=>"101101011",
  6701=>"100111110",
  6702=>"110101001",
  6703=>"111100001",
  6704=>"001111111",
  6705=>"001110100",
  6706=>"100111100",
  6707=>"100111101",
  6708=>"100111001",
  6709=>"101010010",
  6710=>"001110011",
  6711=>"011010101",
  6712=>"111001011",
  6713=>"000110000",
  6714=>"011010101",
  6715=>"110101000",
  6716=>"000010111",
  6717=>"010001111",
  6718=>"001001001",
  6719=>"010111110",
  6720=>"100100110",
  6721=>"010010011",
  6722=>"101101110",
  6723=>"001110101",
  6724=>"100011011",
  6725=>"111111101",
  6726=>"010000010",
  6727=>"011111000",
  6728=>"010100000",
  6729=>"110100100",
  6730=>"000010011",
  6731=>"011110011",
  6732=>"011101111",
  6733=>"100001010",
  6734=>"111001011",
  6735=>"110101010",
  6736=>"000100101",
  6737=>"011101001",
  6738=>"110000010",
  6739=>"001100100",
  6740=>"101100010",
  6741=>"100010101",
  6742=>"111100110",
  6743=>"101001100",
  6744=>"100000100",
  6745=>"110101000",
  6746=>"101100101",
  6747=>"101100000",
  6748=>"010010001",
  6749=>"100010010",
  6750=>"111010010",
  6751=>"011000100",
  6752=>"110100111",
  6753=>"001111011",
  6754=>"011100001",
  6755=>"111010011",
  6756=>"000000100",
  6757=>"101011111",
  6758=>"010110011",
  6759=>"100111110",
  6760=>"111011011",
  6761=>"010010001",
  6762=>"000000111",
  6763=>"011110001",
  6764=>"001110011",
  6765=>"010101001",
  6766=>"011000100",
  6767=>"100111011",
  6768=>"110000000",
  6769=>"100110111",
  6770=>"011000111",
  6771=>"100010110",
  6772=>"011011011",
  6773=>"111000111",
  6774=>"111101110",
  6775=>"111001101",
  6776=>"000111010",
  6777=>"100000001",
  6778=>"000110111",
  6779=>"001111011",
  6780=>"000101110",
  6781=>"101001111",
  6782=>"101110010",
  6783=>"011100100",
  6784=>"110010111",
  6785=>"011110001",
  6786=>"010010000",
  6787=>"101100101",
  6788=>"001110000",
  6789=>"100011111",
  6790=>"111000010",
  6791=>"111011000",
  6792=>"110101011",
  6793=>"101010001",
  6794=>"011100110",
  6795=>"101110011",
  6796=>"110100001",
  6797=>"110011111",
  6798=>"110100011",
  6799=>"110001010",
  6800=>"000011001",
  6801=>"101100011",
  6802=>"100101011",
  6803=>"011111111",
  6804=>"001111010",
  6805=>"000000011",
  6806=>"100100011",
  6807=>"111011111",
  6808=>"100111011",
  6809=>"101101010",
  6810=>"011010000",
  6811=>"101111100",
  6812=>"110110110",
  6813=>"010001011",
  6814=>"111011100",
  6815=>"000110000",
  6816=>"011101111",
  6817=>"100011010",
  6818=>"010100100",
  6819=>"000110100",
  6820=>"001001101",
  6821=>"111110001",
  6822=>"101100011",
  6823=>"000111001",
  6824=>"110111001",
  6825=>"111010000",
  6826=>"110101001",
  6827=>"111111101",
  6828=>"000011000",
  6829=>"011000111",
  6830=>"110001000",
  6831=>"110100100",
  6832=>"000000110",
  6833=>"010110111",
  6834=>"011100111",
  6835=>"011000001",
  6836=>"000100101",
  6837=>"100110101",
  6838=>"010100110",
  6839=>"011111000",
  6840=>"001101010",
  6841=>"000000101",
  6842=>"110011111",
  6843=>"110011111",
  6844=>"101100111",
  6845=>"000000100",
  6846=>"001000110",
  6847=>"000010111",
  6848=>"111011100",
  6849=>"011100010",
  6850=>"011000101",
  6851=>"000001010",
  6852=>"101111100",
  6853=>"100001110",
  6854=>"110110010",
  6855=>"110001100",
  6856=>"111111110",
  6857=>"111110000",
  6858=>"110100101",
  6859=>"010100110",
  6860=>"011101000",
  6861=>"111000011",
  6862=>"110101001",
  6863=>"011000001",
  6864=>"001001101",
  6865=>"101000111",
  6866=>"011001110",
  6867=>"010111101",
  6868=>"010001111",
  6869=>"011111111",
  6870=>"110000001",
  6871=>"110101011",
  6872=>"100001001",
  6873=>"100110011",
  6874=>"001000101",
  6875=>"100110000",
  6876=>"100001100",
  6877=>"101001111",
  6878=>"000001011",
  6879=>"001110000",
  6880=>"110010100",
  6881=>"000001011",
  6882=>"010101101",
  6883=>"111000110",
  6884=>"010000011",
  6885=>"110100011",
  6886=>"111000001",
  6887=>"010111100",
  6888=>"111011101",
  6889=>"101100010",
  6890=>"101010100",
  6891=>"010111001",
  6892=>"100100010",
  6893=>"000110001",
  6894=>"110111101",
  6895=>"111000110",
  6896=>"100011101",
  6897=>"111111110",
  6898=>"110011110",
  6899=>"010100011",
  6900=>"100000110",
  6901=>"111111101",
  6902=>"011100111",
  6903=>"000010001",
  6904=>"100010001",
  6905=>"101111010",
  6906=>"000100010",
  6907=>"111011011",
  6908=>"000010010",
  6909=>"011000001",
  6910=>"000100011",
  6911=>"110001000",
  6912=>"110001101",
  6913=>"011100011",
  6914=>"010110000",
  6915=>"010111011",
  6916=>"111011011",
  6917=>"111010110",
  6918=>"100000011",
  6919=>"000010001",
  6920=>"000010100",
  6921=>"011011110",
  6922=>"101100110",
  6923=>"010010010",
  6924=>"110110001",
  6925=>"000001010",
  6926=>"000010110",
  6927=>"100011000",
  6928=>"100010110",
  6929=>"011000110",
  6930=>"011011011",
  6931=>"000110111",
  6932=>"001000011",
  6933=>"111110001",
  6934=>"011011010",
  6935=>"111110001",
  6936=>"101000100",
  6937=>"000011111",
  6938=>"000100100",
  6939=>"101001001",
  6940=>"011101100",
  6941=>"100010101",
  6942=>"111010000",
  6943=>"000110111",
  6944=>"011001000",
  6945=>"111011010",
  6946=>"001101110",
  6947=>"000011000",
  6948=>"110011001",
  6949=>"101001111",
  6950=>"100110111",
  6951=>"111110000",
  6952=>"100110001",
  6953=>"111101011",
  6954=>"011010010",
  6955=>"110010000",
  6956=>"110001110",
  6957=>"010101011",
  6958=>"110110111",
  6959=>"000010010",
  6960=>"000010011",
  6961=>"000100010",
  6962=>"011011000",
  6963=>"100001111",
  6964=>"111010110",
  6965=>"001011111",
  6966=>"101110101",
  6967=>"110111010",
  6968=>"111111110",
  6969=>"010111000",
  6970=>"101010001",
  6971=>"111000111",
  6972=>"001100011",
  6973=>"100010100",
  6974=>"001011110",
  6975=>"010000111",
  6976=>"010010010",
  6977=>"111101101",
  6978=>"100101101",
  6979=>"001101100",
  6980=>"110101101",
  6981=>"010100101",
  6982=>"111110110",
  6983=>"001100100",
  6984=>"111000111",
  6985=>"010100100",
  6986=>"101010100",
  6987=>"011110011",
  6988=>"010110001",
  6989=>"101010110",
  6990=>"011010001",
  6991=>"111110010",
  6992=>"101000000",
  6993=>"101100010",
  6994=>"111100101",
  6995=>"100011101",
  6996=>"111111110",
  6997=>"111011101",
  6998=>"001000001",
  6999=>"100011011",
  7000=>"010010011",
  7001=>"110101010",
  7002=>"011010011",
  7003=>"000100000",
  7004=>"000010000",
  7005=>"001011000",
  7006=>"110111011",
  7007=>"110101111",
  7008=>"111000010",
  7009=>"111010000",
  7010=>"011011001",
  7011=>"101101111",
  7012=>"110010110",
  7013=>"001001000",
  7014=>"100111101",
  7015=>"010010010",
  7016=>"111010001",
  7017=>"101010111",
  7018=>"100110010",
  7019=>"010111010",
  7020=>"101011110",
  7021=>"100101010",
  7022=>"100110111",
  7023=>"011101001",
  7024=>"100111001",
  7025=>"011010101",
  7026=>"110011101",
  7027=>"000000110",
  7028=>"000000010",
  7029=>"000111001",
  7030=>"101100111",
  7031=>"101101001",
  7032=>"101111000",
  7033=>"011101101",
  7034=>"000111010",
  7035=>"100101010",
  7036=>"001001010",
  7037=>"010100000",
  7038=>"110000100",
  7039=>"110101111",
  7040=>"010011110",
  7041=>"110011001",
  7042=>"110111001",
  7043=>"100011001",
  7044=>"011010010",
  7045=>"010101110",
  7046=>"101111101",
  7047=>"111111010",
  7048=>"101111011",
  7049=>"111101011",
  7050=>"001000011",
  7051=>"111000001",
  7052=>"100001001",
  7053=>"101111011",
  7054=>"001010001",
  7055=>"101100100",
  7056=>"011010001",
  7057=>"111100111",
  7058=>"111110001",
  7059=>"111001100",
  7060=>"101100110",
  7061=>"001101111",
  7062=>"111001000",
  7063=>"101011011",
  7064=>"000111100",
  7065=>"111001000",
  7066=>"111010110",
  7067=>"011101011",
  7068=>"011000000",
  7069=>"011110111",
  7070=>"000010100",
  7071=>"101001010",
  7072=>"111111011",
  7073=>"101000001",
  7074=>"000100011",
  7075=>"011010111",
  7076=>"010101111",
  7077=>"110101000",
  7078=>"101100100",
  7079=>"101001110",
  7080=>"001010011",
  7081=>"100000111",
  7082=>"011111000",
  7083=>"101011101",
  7084=>"001001001",
  7085=>"101101011",
  7086=>"000010001",
  7087=>"010100001",
  7088=>"101100111",
  7089=>"100000100",
  7090=>"110110100",
  7091=>"010111101",
  7092=>"111001010",
  7093=>"011000101",
  7094=>"110110111",
  7095=>"000000001",
  7096=>"001010101",
  7097=>"001100001",
  7098=>"000010101",
  7099=>"101001111",
  7100=>"111110111",
  7101=>"011000100",
  7102=>"010101010",
  7103=>"000001010",
  7104=>"000101001",
  7105=>"010111100",
  7106=>"110111100",
  7107=>"110000011",
  7108=>"001001000",
  7109=>"010001001",
  7110=>"000011001",
  7111=>"001010001",
  7112=>"110010001",
  7113=>"000100010",
  7114=>"101100101",
  7115=>"000001011",
  7116=>"011100111",
  7117=>"011010011",
  7118=>"011010001",
  7119=>"100010010",
  7120=>"010010010",
  7121=>"011111010",
  7122=>"011110110",
  7123=>"111000011",
  7124=>"011011111",
  7125=>"100100011",
  7126=>"011011010",
  7127=>"111101111",
  7128=>"010110001",
  7129=>"000010101",
  7130=>"000000001",
  7131=>"110000101",
  7132=>"100001100",
  7133=>"101000110",
  7134=>"100110100",
  7135=>"110101111",
  7136=>"000100001",
  7137=>"101101011",
  7138=>"001100010",
  7139=>"010010111",
  7140=>"110110111",
  7141=>"100010100",
  7142=>"100011100",
  7143=>"010111100",
  7144=>"111010111",
  7145=>"110010000",
  7146=>"110010111",
  7147=>"011100101",
  7148=>"101101101",
  7149=>"011011101",
  7150=>"010111111",
  7151=>"000011111",
  7152=>"101001100",
  7153=>"111010101",
  7154=>"011011001",
  7155=>"110000010",
  7156=>"110000100",
  7157=>"110100000",
  7158=>"110000101",
  7159=>"000101110",
  7160=>"000001001",
  7161=>"101110000",
  7162=>"001100010",
  7163=>"001101111",
  7164=>"111010010",
  7165=>"011010011",
  7166=>"100100111",
  7167=>"011101100",
  7168=>"111000000",
  7169=>"110100111",
  7170=>"110011111",
  7171=>"110101101",
  7172=>"010011101",
  7173=>"001110110",
  7174=>"110101100",
  7175=>"111111110",
  7176=>"101001100",
  7177=>"001110101",
  7178=>"110001011",
  7179=>"010000001",
  7180=>"011101011",
  7181=>"100100101",
  7182=>"101101111",
  7183=>"110001010",
  7184=>"101011000",
  7185=>"001011001",
  7186=>"101101111",
  7187=>"100100100",
  7188=>"000010101",
  7189=>"110011101",
  7190=>"000110110",
  7191=>"001010100",
  7192=>"101010111",
  7193=>"000100000",
  7194=>"110011011",
  7195=>"110101110",
  7196=>"101001100",
  7197=>"101010001",
  7198=>"100110100",
  7199=>"001011000",
  7200=>"110110010",
  7201=>"100000111",
  7202=>"101000110",
  7203=>"101110010",
  7204=>"000100110",
  7205=>"011011111",
  7206=>"011110010",
  7207=>"110001010",
  7208=>"010101101",
  7209=>"000100100",
  7210=>"010111110",
  7211=>"100111111",
  7212=>"101001100",
  7213=>"010010001",
  7214=>"001111100",
  7215=>"100100111",
  7216=>"010110000",
  7217=>"000011100",
  7218=>"101110101",
  7219=>"010011111",
  7220=>"110001000",
  7221=>"001101111",
  7222=>"101110100",
  7223=>"110101010",
  7224=>"100111100",
  7225=>"011110000",
  7226=>"100000100",
  7227=>"000011110",
  7228=>"000010010",
  7229=>"001001100",
  7230=>"110000100",
  7231=>"010011001",
  7232=>"100011111",
  7233=>"000100000",
  7234=>"111010001",
  7235=>"011111000",
  7236=>"100010011",
  7237=>"101111011",
  7238=>"001011111",
  7239=>"111101111",
  7240=>"001111100",
  7241=>"110110101",
  7242=>"010001000",
  7243=>"011101000",
  7244=>"110011001",
  7245=>"001011011",
  7246=>"100101101",
  7247=>"100100101",
  7248=>"001011110",
  7249=>"011110111",
  7250=>"101110100",
  7251=>"110101100",
  7252=>"101110100",
  7253=>"001111100",
  7254=>"100011001",
  7255=>"000010111",
  7256=>"011011110",
  7257=>"101000111",
  7258=>"100000100",
  7259=>"111100011",
  7260=>"100001011",
  7261=>"001111101",
  7262=>"001001010",
  7263=>"111100010",
  7264=>"110110011",
  7265=>"101000000",
  7266=>"100111010",
  7267=>"110111101",
  7268=>"011110101",
  7269=>"001110111",
  7270=>"011001000",
  7271=>"111111011",
  7272=>"000100111",
  7273=>"111100101",
  7274=>"001101010",
  7275=>"110101101",
  7276=>"111100000",
  7277=>"101011101",
  7278=>"001100111",
  7279=>"001000111",
  7280=>"001000011",
  7281=>"110111011",
  7282=>"000110111",
  7283=>"111111100",
  7284=>"010001001",
  7285=>"100011011",
  7286=>"101000111",
  7287=>"011011110",
  7288=>"101111011",
  7289=>"100010101",
  7290=>"011000010",
  7291=>"001100011",
  7292=>"011011001",
  7293=>"001001001",
  7294=>"010010010",
  7295=>"000000111",
  7296=>"100110100",
  7297=>"001010110",
  7298=>"001001010",
  7299=>"010010010",
  7300=>"000010001",
  7301=>"011011010",
  7302=>"001111111",
  7303=>"110101111",
  7304=>"101100110",
  7305=>"010010101",
  7306=>"001111111",
  7307=>"101001101",
  7308=>"000010011",
  7309=>"110101011",
  7310=>"110100001",
  7311=>"101101110",
  7312=>"000011011",
  7313=>"001100111",
  7314=>"100000110",
  7315=>"000010110",
  7316=>"111000100",
  7317=>"110010110",
  7318=>"010111101",
  7319=>"111101110",
  7320=>"100110101",
  7321=>"000101111",
  7322=>"000011110",
  7323=>"101110110",
  7324=>"000100001",
  7325=>"110101101",
  7326=>"100010110",
  7327=>"001110000",
  7328=>"100100100",
  7329=>"001001000",
  7330=>"111011010",
  7331=>"110111000",
  7332=>"010100001",
  7333=>"101001000",
  7334=>"011000101",
  7335=>"100110010",
  7336=>"010111100",
  7337=>"001011000",
  7338=>"001001101",
  7339=>"111100000",
  7340=>"011101010",
  7341=>"001000110",
  7342=>"100011100",
  7343=>"011111111",
  7344=>"001101010",
  7345=>"100110100",
  7346=>"101110101",
  7347=>"011000010",
  7348=>"101010000",
  7349=>"101111110",
  7350=>"100110010",
  7351=>"111111101",
  7352=>"001001001",
  7353=>"110011101",
  7354=>"010001100",
  7355=>"101101000",
  7356=>"110010011",
  7357=>"111111101",
  7358=>"000100000",
  7359=>"111100000",
  7360=>"011101110",
  7361=>"001011010",
  7362=>"001101101",
  7363=>"101111101",
  7364=>"101011001",
  7365=>"111001011",
  7366=>"111000000",
  7367=>"001000111",
  7368=>"111111001",
  7369=>"100111011",
  7370=>"100010101",
  7371=>"000110100",
  7372=>"011001001",
  7373=>"011101000",
  7374=>"000100000",
  7375=>"101010111",
  7376=>"001000100",
  7377=>"001001100",
  7378=>"000001100",
  7379=>"111001000",
  7380=>"010101111",
  7381=>"011010110",
  7382=>"011010111",
  7383=>"111101011",
  7384=>"100101100",
  7385=>"010001000",
  7386=>"000001100",
  7387=>"001001100",
  7388=>"011010000",
  7389=>"001110100",
  7390=>"010111010",
  7391=>"110111101",
  7392=>"010100000",
  7393=>"010100011",
  7394=>"001010111",
  7395=>"000011011",
  7396=>"000110011",
  7397=>"111000000",
  7398=>"010011011",
  7399=>"110100000",
  7400=>"001111101",
  7401=>"101111010",
  7402=>"010100101",
  7403=>"001011111",
  7404=>"000011010",
  7405=>"110011000",
  7406=>"001001010",
  7407=>"000100000",
  7408=>"001100100",
  7409=>"000111000",
  7410=>"000010011",
  7411=>"110101111",
  7412=>"001010110",
  7413=>"101000011",
  7414=>"111000000",
  7415=>"010110100",
  7416=>"011001000",
  7417=>"011000111",
  7418=>"001100100",
  7419=>"010010111",
  7420=>"100101000",
  7421=>"101100000",
  7422=>"110000100",
  7423=>"001110011",
  7424=>"001011000",
  7425=>"010110000",
  7426=>"111111111",
  7427=>"000001111",
  7428=>"010111010",
  7429=>"010100010",
  7430=>"000100011",
  7431=>"000101001",
  7432=>"100010101",
  7433=>"010110111",
  7434=>"000110101",
  7435=>"001000011",
  7436=>"100111101",
  7437=>"100101111",
  7438=>"110101001",
  7439=>"000101110",
  7440=>"001101011",
  7441=>"111111101",
  7442=>"001000011",
  7443=>"000110010",
  7444=>"001000001",
  7445=>"011100000",
  7446=>"101011001",
  7447=>"001111000",
  7448=>"100000010",
  7449=>"011100111",
  7450=>"110001101",
  7451=>"111100011",
  7452=>"011110100",
  7453=>"010100010",
  7454=>"101000011",
  7455=>"100010111",
  7456=>"011110111",
  7457=>"010000000",
  7458=>"010101100",
  7459=>"011101001",
  7460=>"101100111",
  7461=>"010101011",
  7462=>"110111101",
  7463=>"111110100",
  7464=>"001101010",
  7465=>"101111111",
  7466=>"110100111",
  7467=>"111110110",
  7468=>"100100110",
  7469=>"110011100",
  7470=>"111001101",
  7471=>"101111101",
  7472=>"011000000",
  7473=>"000000001",
  7474=>"101110001",
  7475=>"101011100",
  7476=>"111100100",
  7477=>"101001101",
  7478=>"001000001",
  7479=>"100011100",
  7480=>"100001110",
  7481=>"101011011",
  7482=>"000001110",
  7483=>"101110000",
  7484=>"111101110",
  7485=>"101000111",
  7486=>"000111110",
  7487=>"111110100",
  7488=>"001010000",
  7489=>"101000100",
  7490=>"111101110",
  7491=>"111101010",
  7492=>"101111100",
  7493=>"101011101",
  7494=>"011100011",
  7495=>"000010000",
  7496=>"101001100",
  7497=>"000010010",
  7498=>"100000111",
  7499=>"010000100",
  7500=>"000010100",
  7501=>"001101110",
  7502=>"101000010",
  7503=>"001110101",
  7504=>"001000000",
  7505=>"000010101",
  7506=>"010101111",
  7507=>"111001011",
  7508=>"011011001",
  7509=>"001001101",
  7510=>"011101111",
  7511=>"010101001",
  7512=>"001111000",
  7513=>"010001000",
  7514=>"111011011",
  7515=>"000101111",
  7516=>"101011001",
  7517=>"001110100",
  7518=>"001011010",
  7519=>"001100100",
  7520=>"110011111",
  7521=>"000100011",
  7522=>"000010010",
  7523=>"000110011",
  7524=>"100011110",
  7525=>"101100011",
  7526=>"101111010",
  7527=>"011000110",
  7528=>"001011110",
  7529=>"011100001",
  7530=>"100100101",
  7531=>"110110000",
  7532=>"000000010",
  7533=>"000111011",
  7534=>"000011011",
  7535=>"101001000",
  7536=>"000010100",
  7537=>"111000011",
  7538=>"010011011",
  7539=>"011000010",
  7540=>"111101001",
  7541=>"110101000",
  7542=>"110011011",
  7543=>"101110000",
  7544=>"111011101",
  7545=>"101010011",
  7546=>"011001101",
  7547=>"100000101",
  7548=>"001111110",
  7549=>"100100001",
  7550=>"000100001",
  7551=>"000100001",
  7552=>"011101000",
  7553=>"111111111",
  7554=>"010110111",
  7555=>"011000100",
  7556=>"100110110",
  7557=>"101010000",
  7558=>"110110111",
  7559=>"010111111",
  7560=>"101111010",
  7561=>"101100001",
  7562=>"111010100",
  7563=>"011001000",
  7564=>"010111010",
  7565=>"000011111",
  7566=>"101011000",
  7567=>"010100010",
  7568=>"111101111",
  7569=>"100001111",
  7570=>"000011100",
  7571=>"101011010",
  7572=>"011100011",
  7573=>"011011010",
  7574=>"010001111",
  7575=>"110111110",
  7576=>"000000100",
  7577=>"001100111",
  7578=>"010111100",
  7579=>"000011101",
  7580=>"011000001",
  7581=>"101001110",
  7582=>"101010000",
  7583=>"100000011",
  7584=>"101101110",
  7585=>"010011010",
  7586=>"011111100",
  7587=>"010111101",
  7588=>"011000011",
  7589=>"111001000",
  7590=>"001000111",
  7591=>"100000010",
  7592=>"001001110",
  7593=>"110001111",
  7594=>"011100011",
  7595=>"110100111",
  7596=>"101011011",
  7597=>"001011101",
  7598=>"111000111",
  7599=>"011001001",
  7600=>"010000101",
  7601=>"111000110",
  7602=>"000100010",
  7603=>"001001100",
  7604=>"101000110",
  7605=>"000011100",
  7606=>"010000001",
  7607=>"000010101",
  7608=>"100000011",
  7609=>"010100110",
  7610=>"001100010",
  7611=>"001000000",
  7612=>"101011111",
  7613=>"110111110",
  7614=>"010101100",
  7615=>"111100110",
  7616=>"001000010",
  7617=>"101001001",
  7618=>"001011001",
  7619=>"101111110",
  7620=>"111100111",
  7621=>"000000000",
  7622=>"100100000",
  7623=>"111010111",
  7624=>"001011001",
  7625=>"111111100",
  7626=>"011001010",
  7627=>"101111011",
  7628=>"001110100",
  7629=>"001100011",
  7630=>"101111110",
  7631=>"000101110",
  7632=>"111011100",
  7633=>"100100000",
  7634=>"111001001",
  7635=>"111100110",
  7636=>"000101111",
  7637=>"101111101",
  7638=>"101100001",
  7639=>"110110111",
  7640=>"101001001",
  7641=>"111001110",
  7642=>"100011111",
  7643=>"100111001",
  7644=>"101011000",
  7645=>"111110001",
  7646=>"110011100",
  7647=>"010101111",
  7648=>"001011011",
  7649=>"011100110",
  7650=>"101101111",
  7651=>"111101101",
  7652=>"100010110",
  7653=>"110110111",
  7654=>"010011111",
  7655=>"000011101",
  7656=>"111001011",
  7657=>"000010001",
  7658=>"010101001",
  7659=>"101001000",
  7660=>"101010101",
  7661=>"001001100",
  7662=>"111001001",
  7663=>"000001101",
  7664=>"011110111",
  7665=>"010101010",
  7666=>"001100010",
  7667=>"111011100",
  7668=>"101111100",
  7669=>"101110111",
  7670=>"010101001",
  7671=>"000000011",
  7672=>"100101100",
  7673=>"011111111",
  7674=>"100001011",
  7675=>"100101100",
  7676=>"010110110",
  7677=>"010000011",
  7678=>"100010101",
  7679=>"111101100",
  7680=>"011100001",
  7681=>"001001000",
  7682=>"110001110",
  7683=>"010101111",
  7684=>"011010111",
  7685=>"011101100",
  7686=>"100011000",
  7687=>"001101110",
  7688=>"011111111",
  7689=>"110110111",
  7690=>"110110111",
  7691=>"100011001",
  7692=>"100110101",
  7693=>"101101001",
  7694=>"000011001",
  7695=>"000100011",
  7696=>"001100110",
  7697=>"100111010",
  7698=>"101101110",
  7699=>"011111101",
  7700=>"001001110",
  7701=>"010110111",
  7702=>"100100110",
  7703=>"001000010",
  7704=>"000110111",
  7705=>"110001001",
  7706=>"101110001",
  7707=>"100001011",
  7708=>"001000101",
  7709=>"110000000",
  7710=>"000110010",
  7711=>"010000110",
  7712=>"101101010",
  7713=>"001101101",
  7714=>"000110011",
  7715=>"110011000",
  7716=>"101111101",
  7717=>"101011111",
  7718=>"011100011",
  7719=>"000100000",
  7720=>"011110100",
  7721=>"111100011",
  7722=>"000001001",
  7723=>"110110111",
  7724=>"011011001",
  7725=>"101101100",
  7726=>"010000000",
  7727=>"010010110",
  7728=>"111011100",
  7729=>"111000111",
  7730=>"011101100",
  7731=>"110101000",
  7732=>"000010010",
  7733=>"101101111",
  7734=>"011000101",
  7735=>"110111100",
  7736=>"100010010",
  7737=>"101000000",
  7738=>"110101010",
  7739=>"100001010",
  7740=>"100111110",
  7741=>"010011110",
  7742=>"001110101",
  7743=>"100000000",
  7744=>"011001111",
  7745=>"100111010",
  7746=>"011010111",
  7747=>"100000001",
  7748=>"011111000",
  7749=>"110000011",
  7750=>"011110001",
  7751=>"011011111",
  7752=>"101001011",
  7753=>"110110010",
  7754=>"101100101",
  7755=>"011110110",
  7756=>"001010000",
  7757=>"010000111",
  7758=>"101101000",
  7759=>"110100101",
  7760=>"011101110",
  7761=>"101000000",
  7762=>"111011001",
  7763=>"101001111",
  7764=>"000101001",
  7765=>"000111100",
  7766=>"011011100",
  7767=>"011001010",
  7768=>"101110111",
  7769=>"101110100",
  7770=>"110100000",
  7771=>"001001110",
  7772=>"100110010",
  7773=>"000100110",
  7774=>"110011101",
  7775=>"110011111",
  7776=>"010001011",
  7777=>"111111011",
  7778=>"111101011",
  7779=>"000010111",
  7780=>"000100010",
  7781=>"101000111",
  7782=>"101000110",
  7783=>"111010100",
  7784=>"010011011",
  7785=>"000001010",
  7786=>"111100111",
  7787=>"110010001",
  7788=>"000111010",
  7789=>"110111110",
  7790=>"011100010",
  7791=>"000010000",
  7792=>"101101101",
  7793=>"101100011",
  7794=>"111100001",
  7795=>"111100110",
  7796=>"110000110",
  7797=>"000010100",
  7798=>"011101001",
  7799=>"101111000",
  7800=>"101010111",
  7801=>"000000100",
  7802=>"101111000",
  7803=>"001001000",
  7804=>"000010111",
  7805=>"110000101",
  7806=>"110011101",
  7807=>"000111000",
  7808=>"111110011",
  7809=>"010011111",
  7810=>"010001000",
  7811=>"100000000",
  7812=>"010100001",
  7813=>"011110001",
  7814=>"100100000",
  7815=>"000100000",
  7816=>"101000100",
  7817=>"001001100",
  7818=>"100110010",
  7819=>"110001110",
  7820=>"010111001",
  7821=>"111110001",
  7822=>"111010111",
  7823=>"010001001",
  7824=>"010000111",
  7825=>"110001000",
  7826=>"000001000",
  7827=>"000111111",
  7828=>"101111110",
  7829=>"111001101",
  7830=>"010101111",
  7831=>"000010100",
  7832=>"111101001",
  7833=>"111101011",
  7834=>"110010101",
  7835=>"100011000",
  7836=>"101001010",
  7837=>"110101100",
  7838=>"100010100",
  7839=>"100001001",
  7840=>"011110101",
  7841=>"000110000",
  7842=>"100001101",
  7843=>"000101001",
  7844=>"110000011",
  7845=>"100101000",
  7846=>"011110111",
  7847=>"101101111",
  7848=>"110011011",
  7849=>"100001010",
  7850=>"010010100",
  7851=>"001011110",
  7852=>"010000000",
  7853=>"010010101",
  7854=>"110000100",
  7855=>"101110001",
  7856=>"000011101",
  7857=>"111111010",
  7858=>"011101100",
  7859=>"101100111",
  7860=>"010101100",
  7861=>"000111000",
  7862=>"111111001",
  7863=>"011110111",
  7864=>"111000011",
  7865=>"110110001",
  7866=>"100101001",
  7867=>"101010000",
  7868=>"001101010",
  7869=>"101011110",
  7870=>"010111111",
  7871=>"101001001",
  7872=>"101000111",
  7873=>"100100011",
  7874=>"101101000",
  7875=>"110101110",
  7876=>"101110011",
  7877=>"110110000",
  7878=>"001000100",
  7879=>"110110110",
  7880=>"000110101",
  7881=>"000000011",
  7882=>"001101101",
  7883=>"011011110",
  7884=>"111011111",
  7885=>"010111111",
  7886=>"000001111",
  7887=>"101000010",
  7888=>"101100100",
  7889=>"111110110",
  7890=>"010011101",
  7891=>"001001110",
  7892=>"010111001",
  7893=>"100110000",
  7894=>"001000111",
  7895=>"101110000",
  7896=>"100101000",
  7897=>"100100101",
  7898=>"100011110",
  7899=>"111000100",
  7900=>"000011010",
  7901=>"100011100",
  7902=>"010111110",
  7903=>"101001011",
  7904=>"111100000",
  7905=>"110111000",
  7906=>"001100100",
  7907=>"101011001",
  7908=>"011001001",
  7909=>"111000010",
  7910=>"010111010",
  7911=>"111110010",
  7912=>"001111101",
  7913=>"100100010",
  7914=>"110001111",
  7915=>"101001001",
  7916=>"001100000",
  7917=>"001101100",
  7918=>"110110001",
  7919=>"011110111",
  7920=>"111101110",
  7921=>"010010001",
  7922=>"100011000",
  7923=>"011011110",
  7924=>"101111010",
  7925=>"000001010",
  7926=>"101001010",
  7927=>"001000011",
  7928=>"101001110",
  7929=>"110110101",
  7930=>"000001010",
  7931=>"110010001",
  7932=>"110001001",
  7933=>"111101010",
  7934=>"101011001",
  7935=>"001111110",
  7936=>"000010100",
  7937=>"000100101",
  7938=>"111010011",
  7939=>"001100010",
  7940=>"000100001",
  7941=>"000010001",
  7942=>"001011111",
  7943=>"110100000",
  7944=>"100001110",
  7945=>"111111011",
  7946=>"110100000",
  7947=>"010000001",
  7948=>"110010101",
  7949=>"111110010",
  7950=>"011001110",
  7951=>"110101010",
  7952=>"001100110",
  7953=>"111011101",
  7954=>"010010111",
  7955=>"011110000",
  7956=>"110010111",
  7957=>"000100011",
  7958=>"011101000",
  7959=>"000100100",
  7960=>"101100001",
  7961=>"000000110",
  7962=>"000001000",
  7963=>"000001010",
  7964=>"000110111",
  7965=>"110110001",
  7966=>"011011101",
  7967=>"001001000",
  7968=>"110101001",
  7969=>"010110000",
  7970=>"101011110",
  7971=>"111000111",
  7972=>"110001001",
  7973=>"010101110",
  7974=>"010000100",
  7975=>"000111100",
  7976=>"100100000",
  7977=>"101000011",
  7978=>"010111110",
  7979=>"101011010",
  7980=>"010101010",
  7981=>"111001101",
  7982=>"000111000",
  7983=>"001010001",
  7984=>"010011011",
  7985=>"000010010",
  7986=>"100001110",
  7987=>"000010101",
  7988=>"011010000",
  7989=>"000100111",
  7990=>"000110010",
  7991=>"110010010",
  7992=>"100111000",
  7993=>"000010101",
  7994=>"111010110",
  7995=>"100000011",
  7996=>"000011110",
  7997=>"110001001",
  7998=>"000111111",
  7999=>"001001000",
  8000=>"100111001",
  8001=>"001001000",
  8002=>"010111111",
  8003=>"100110110",
  8004=>"100000111",
  8005=>"011000100",
  8006=>"010000000",
  8007=>"001011000",
  8008=>"111001000",
  8009=>"100000001",
  8010=>"011010010",
  8011=>"000110100",
  8012=>"001001100",
  8013=>"111101100",
  8014=>"010010101",
  8015=>"010000011",
  8016=>"010010000",
  8017=>"101000100",
  8018=>"011000001",
  8019=>"011010100",
  8020=>"000101010",
  8021=>"110000100",
  8022=>"111101010",
  8023=>"101100011",
  8024=>"001001100",
  8025=>"011100111",
  8026=>"000101111",
  8027=>"101111101",
  8028=>"010000010",
  8029=>"100000001",
  8030=>"011011110",
  8031=>"110110101",
  8032=>"100001010",
  8033=>"001000000",
  8034=>"011011100",
  8035=>"011110111",
  8036=>"101001111",
  8037=>"001001010",
  8038=>"101010100",
  8039=>"001110101",
  8040=>"010011110",
  8041=>"111000001",
  8042=>"111101001",
  8043=>"011111011",
  8044=>"011010100",
  8045=>"001011011",
  8046=>"001100000",
  8047=>"100001101",
  8048=>"001001111",
  8049=>"010011111",
  8050=>"010110111",
  8051=>"110010000",
  8052=>"001011011",
  8053=>"111111110",
  8054=>"011111101",
  8055=>"100011011",
  8056=>"000100111",
  8057=>"000110111",
  8058=>"011110011",
  8059=>"011001001",
  8060=>"001001111",
  8061=>"000111100",
  8062=>"100100110",
  8063=>"000011011",
  8064=>"101000101",
  8065=>"010110101",
  8066=>"001100111",
  8067=>"110001110",
  8068=>"001110010",
  8069=>"101111110",
  8070=>"110000111",
  8071=>"111001001",
  8072=>"000110000",
  8073=>"010101110",
  8074=>"101001110",
  8075=>"100111111",
  8076=>"010000011",
  8077=>"000000001",
  8078=>"001110101",
  8079=>"110110000",
  8080=>"110001111",
  8081=>"010010000",
  8082=>"010010000",
  8083=>"111001011",
  8084=>"111111101",
  8085=>"001011000",
  8086=>"001001101",
  8087=>"100001001",
  8088=>"001010101",
  8089=>"000111101",
  8090=>"010010011",
  8091=>"000011100",
  8092=>"111101011",
  8093=>"101111000",
  8094=>"000011111",
  8095=>"111111000",
  8096=>"000000011",
  8097=>"000000111",
  8098=>"010101100",
  8099=>"010001110",
  8100=>"100011000",
  8101=>"101000101",
  8102=>"000001010",
  8103=>"101111100",
  8104=>"011001011",
  8105=>"100000010",
  8106=>"110110010",
  8107=>"100010101",
  8108=>"000000011",
  8109=>"100010000",
  8110=>"111101100",
  8111=>"010100100",
  8112=>"110000110",
  8113=>"001010000",
  8114=>"101101111",
  8115=>"001000111",
  8116=>"011111000",
  8117=>"001101011",
  8118=>"010100110",
  8119=>"100111001",
  8120=>"011110010",
  8121=>"110011110",
  8122=>"001000111",
  8123=>"001100100",
  8124=>"100011001",
  8125=>"000000010",
  8126=>"111100001",
  8127=>"011101001",
  8128=>"110111111",
  8129=>"111101110",
  8130=>"001110100",
  8131=>"011001010",
  8132=>"010001101",
  8133=>"100100001",
  8134=>"010001000",
  8135=>"111010010",
  8136=>"010100000",
  8137=>"010001100",
  8138=>"010000010",
  8139=>"010010010",
  8140=>"000110010",
  8141=>"011010101",
  8142=>"000010110",
  8143=>"100011000",
  8144=>"110111111",
  8145=>"111010101",
  8146=>"101011110",
  8147=>"000010011",
  8148=>"001101100",
  8149=>"101111001",
  8150=>"101001111",
  8151=>"101101110",
  8152=>"101111101",
  8153=>"011001100",
  8154=>"101110010",
  8155=>"010000110",
  8156=>"001110101",
  8157=>"010000010",
  8158=>"101001011",
  8159=>"100010001",
  8160=>"100111100",
  8161=>"010110010",
  8162=>"100010100",
  8163=>"111101010",
  8164=>"101110101",
  8165=>"010111101",
  8166=>"010001100",
  8167=>"001000100",
  8168=>"001101011",
  8169=>"010110101",
  8170=>"100110000",
  8171=>"100001101",
  8172=>"001010010",
  8173=>"001001000",
  8174=>"101000100",
  8175=>"010001100",
  8176=>"010111111",
  8177=>"111011011",
  8178=>"011111110",
  8179=>"111000001",
  8180=>"100100001",
  8181=>"100100111",
  8182=>"011001101",
  8183=>"111101000",
  8184=>"101101000",
  8185=>"000011001",
  8186=>"100100100",
  8187=>"010100001",
  8188=>"000011101",
  8189=>"000010011",
  8190=>"100100011",
  8191=>"101100110",
  8192=>"110010010",
  8193=>"011011110",
  8194=>"010110101",
  8195=>"001000011",
  8196=>"010100010",
  8197=>"011111011",
  8198=>"001001010",
  8199=>"011101001",
  8200=>"011000011",
  8201=>"101111000",
  8202=>"001101111",
  8203=>"010001101",
  8204=>"011001100",
  8205=>"111101111",
  8206=>"101111110",
  8207=>"111010011",
  8208=>"011100001",
  8209=>"100110001",
  8210=>"101110001",
  8211=>"001101011",
  8212=>"100100111",
  8213=>"001000100",
  8214=>"000110111",
  8215=>"111001010",
  8216=>"000010111",
  8217=>"010111111",
  8218=>"000011010",
  8219=>"101100001",
  8220=>"001000001",
  8221=>"111101111",
  8222=>"011001011",
  8223=>"111001000",
  8224=>"010000111",
  8225=>"110101010",
  8226=>"010111111",
  8227=>"101110011",
  8228=>"110010100",
  8229=>"000010001",
  8230=>"101111110",
  8231=>"100010001",
  8232=>"011100101",
  8233=>"100000110",
  8234=>"000101011",
  8235=>"011110101",
  8236=>"111100111",
  8237=>"000001111",
  8238=>"010101001",
  8239=>"110011001",
  8240=>"100101001",
  8241=>"001111001",
  8242=>"010110001",
  8243=>"110010000",
  8244=>"111010011",
  8245=>"101101001",
  8246=>"001101010",
  8247=>"000100100",
  8248=>"111110011",
  8249=>"010111010",
  8250=>"010101001",
  8251=>"001000011",
  8252=>"011010011",
  8253=>"111101010",
  8254=>"110100011",
  8255=>"010000100",
  8256=>"001000100",
  8257=>"000010011",
  8258=>"110101101",
  8259=>"101000110",
  8260=>"000110000",
  8261=>"001000001",
  8262=>"100101000",
  8263=>"111111101",
  8264=>"000111010",
  8265=>"110000110",
  8266=>"000010101",
  8267=>"101000011",
  8268=>"110011110",
  8269=>"100011100",
  8270=>"100110011",
  8271=>"000010011",
  8272=>"001100111",
  8273=>"000000010",
  8274=>"000110110",
  8275=>"110101110",
  8276=>"111100100",
  8277=>"100101010",
  8278=>"111101011",
  8279=>"011000101",
  8280=>"001101011",
  8281=>"111100101",
  8282=>"010010110",
  8283=>"011111111",
  8284=>"010010111",
  8285=>"101101010",
  8286=>"010011111",
  8287=>"101101011",
  8288=>"001001010",
  8289=>"110101011",
  8290=>"000100001",
  8291=>"111101110",
  8292=>"011001101",
  8293=>"011011111",
  8294=>"100100000",
  8295=>"000011000",
  8296=>"111100001",
  8297=>"100100001",
  8298=>"011110100",
  8299=>"110111101",
  8300=>"101100111",
  8301=>"000101101",
  8302=>"100111010",
  8303=>"000000000",
  8304=>"111011000",
  8305=>"100001101",
  8306=>"000011010",
  8307=>"110001111",
  8308=>"000011100",
  8309=>"110001000",
  8310=>"111001011",
  8311=>"010101011",
  8312=>"101111011",
  8313=>"100001010",
  8314=>"110111111",
  8315=>"000011010",
  8316=>"010111001",
  8317=>"101010000",
  8318=>"010100001",
  8319=>"111001100",
  8320=>"110001011",
  8321=>"100100010",
  8322=>"001000101",
  8323=>"000111000",
  8324=>"111000000",
  8325=>"000000010",
  8326=>"011000010",
  8327=>"001010001",
  8328=>"010111110",
  8329=>"100001011",
  8330=>"011011111",
  8331=>"000011000",
  8332=>"110010001",
  8333=>"100111101",
  8334=>"100001000",
  8335=>"000100001",
  8336=>"001000000",
  8337=>"000110001",
  8338=>"011000101",
  8339=>"110101100",
  8340=>"010000010",
  8341=>"100000011",
  8342=>"100101100",
  8343=>"011001101",
  8344=>"011001111",
  8345=>"000011001",
  8346=>"100000000",
  8347=>"101000001",
  8348=>"101111010",
  8349=>"111101110",
  8350=>"111011101",
  8351=>"000100001",
  8352=>"100000111",
  8353=>"111110010",
  8354=>"100111011",
  8355=>"101110000",
  8356=>"010011100",
  8357=>"111110001",
  8358=>"100001010",
  8359=>"110110110",
  8360=>"111000001",
  8361=>"000001111",
  8362=>"010001101",
  8363=>"011000101",
  8364=>"011100000",
  8365=>"101001110",
  8366=>"010010110",
  8367=>"001111111",
  8368=>"100010101",
  8369=>"110101001",
  8370=>"000000010",
  8371=>"100101100",
  8372=>"111001111",
  8373=>"001001011",
  8374=>"001010100",
  8375=>"110011000",
  8376=>"110010000",
  8377=>"010010101",
  8378=>"110010111",
  8379=>"101110101",
  8380=>"011011010",
  8381=>"000000111",
  8382=>"101101100",
  8383=>"001100111",
  8384=>"100010001",
  8385=>"010110000",
  8386=>"000100000",
  8387=>"000100011",
  8388=>"011101000",
  8389=>"101010000",
  8390=>"000011010",
  8391=>"010100100",
  8392=>"001100101",
  8393=>"100001101",
  8394=>"100000111",
  8395=>"111010110",
  8396=>"111110110",
  8397=>"110000010",
  8398=>"101000000",
  8399=>"011111001",
  8400=>"111100111",
  8401=>"011010110",
  8402=>"100110000",
  8403=>"110000111",
  8404=>"110100101",
  8405=>"011111011",
  8406=>"100001010",
  8407=>"111010101",
  8408=>"011001101",
  8409=>"110111110",
  8410=>"101111100",
  8411=>"111010000",
  8412=>"000110001",
  8413=>"101011010",
  8414=>"100010100",
  8415=>"010010110",
  8416=>"110111111",
  8417=>"011101111",
  8418=>"000011101",
  8419=>"110110000",
  8420=>"001111100",
  8421=>"001000000",
  8422=>"011011101",
  8423=>"001011010",
  8424=>"101110111",
  8425=>"100100101",
  8426=>"011110001",
  8427=>"000111111",
  8428=>"111001011",
  8429=>"000010110",
  8430=>"110110010",
  8431=>"010111011",
  8432=>"101110010",
  8433=>"010011101",
  8434=>"100010001",
  8435=>"101100101",
  8436=>"001000011",
  8437=>"101000100",
  8438=>"000000110",
  8439=>"111101010",
  8440=>"000111101",
  8441=>"100100000",
  8442=>"000101010",
  8443=>"010100110",
  8444=>"100001101",
  8445=>"100011111",
  8446=>"010100110",
  8447=>"010000011",
  8448=>"001010101",
  8449=>"110100100",
  8450=>"100000001",
  8451=>"110010011",
  8452=>"000001110",
  8453=>"110010110",
  8454=>"100011001",
  8455=>"000011001",
  8456=>"011000011",
  8457=>"101111010",
  8458=>"011100001",
  8459=>"011111110",
  8460=>"100110010",
  8461=>"010100001",
  8462=>"001111110",
  8463=>"100000010",
  8464=>"101101111",
  8465=>"110001000",
  8466=>"101111111",
  8467=>"001010111",
  8468=>"010010010",
  8469=>"000011100",
  8470=>"101101001",
  8471=>"100011100",
  8472=>"011111000",
  8473=>"010001001",
  8474=>"100000110",
  8475=>"000000111",
  8476=>"011001100",
  8477=>"111011101",
  8478=>"011010110",
  8479=>"111110101",
  8480=>"000010100",
  8481=>"001101011",
  8482=>"001100010",
  8483=>"010000100",
  8484=>"101111001",
  8485=>"100101101",
  8486=>"101110010",
  8487=>"100010110",
  8488=>"000011001",
  8489=>"010110101",
  8490=>"110011111",
  8491=>"001011110",
  8492=>"001001000",
  8493=>"000001110",
  8494=>"000000010",
  8495=>"001111111",
  8496=>"011000011",
  8497=>"001110011",
  8498=>"011011010",
  8499=>"111100001",
  8500=>"110011110",
  8501=>"010001011",
  8502=>"011111100",
  8503=>"100011101",
  8504=>"001101001",
  8505=>"001111000",
  8506=>"111111101",
  8507=>"110100111",
  8508=>"000101100",
  8509=>"010110000",
  8510=>"001011011",
  8511=>"101101101",
  8512=>"010101011",
  8513=>"101100000",
  8514=>"111001010",
  8515=>"110111100",
  8516=>"000110010",
  8517=>"101100111",
  8518=>"011000111",
  8519=>"110111010",
  8520=>"100010100",
  8521=>"001100011",
  8522=>"001000000",
  8523=>"111001001",
  8524=>"100011001",
  8525=>"110000101",
  8526=>"011011011",
  8527=>"110111000",
  8528=>"100110111",
  8529=>"001001011",
  8530=>"111111100",
  8531=>"010001110",
  8532=>"011101000",
  8533=>"110101001",
  8534=>"110101010",
  8535=>"100000110",
  8536=>"100111010",
  8537=>"110100101",
  8538=>"100111011",
  8539=>"010001001",
  8540=>"000101010",
  8541=>"100010000",
  8542=>"110011111",
  8543=>"011111111",
  8544=>"111000001",
  8545=>"101011010",
  8546=>"100100000",
  8547=>"000110111",
  8548=>"100100000",
  8549=>"111010000",
  8550=>"101101001",
  8551=>"001110111",
  8552=>"001011000",
  8553=>"000111110",
  8554=>"111011001",
  8555=>"000101001",
  8556=>"100011100",
  8557=>"000111001",
  8558=>"000110110",
  8559=>"001100101",
  8560=>"010100101",
  8561=>"110110111",
  8562=>"011110000",
  8563=>"100010011",
  8564=>"000001011",
  8565=>"110101111",
  8566=>"101110111",
  8567=>"110101100",
  8568=>"000001100",
  8569=>"110100100",
  8570=>"010111101",
  8571=>"010001010",
  8572=>"000011110",
  8573=>"110011000",
  8574=>"010010000",
  8575=>"000001011",
  8576=>"000000011",
  8577=>"111100000",
  8578=>"010110011",
  8579=>"001110000",
  8580=>"001011101",
  8581=>"100111100",
  8582=>"110110001",
  8583=>"011111110",
  8584=>"001011100",
  8585=>"101011000",
  8586=>"010101011",
  8587=>"001011110",
  8588=>"101001101",
  8589=>"000100000",
  8590=>"001100001",
  8591=>"111001000",
  8592=>"101111001",
  8593=>"011110011",
  8594=>"101010101",
  8595=>"100101010",
  8596=>"000111101",
  8597=>"011001100",
  8598=>"001011011",
  8599=>"101000101",
  8600=>"110001111",
  8601=>"101101011",
  8602=>"110110110",
  8603=>"100010001",
  8604=>"010010100",
  8605=>"011110000",
  8606=>"000111000",
  8607=>"110000001",
  8608=>"111100101",
  8609=>"010010000",
  8610=>"110000110",
  8611=>"111110001",
  8612=>"110111100",
  8613=>"010011100",
  8614=>"000011110",
  8615=>"100011111",
  8616=>"001111111",
  8617=>"010010010",
  8618=>"111010010",
  8619=>"001001101",
  8620=>"100010011",
  8621=>"011011000",
  8622=>"001010001",
  8623=>"000110110",
  8624=>"101101011",
  8625=>"101111100",
  8626=>"000000011",
  8627=>"001001000",
  8628=>"010111100",
  8629=>"100101001",
  8630=>"101111110",
  8631=>"101001100",
  8632=>"101001100",
  8633=>"010010101",
  8634=>"101000100",
  8635=>"011010000",
  8636=>"011111110",
  8637=>"111111010",
  8638=>"101101111",
  8639=>"011011000",
  8640=>"000110011",
  8641=>"010010010",
  8642=>"000110100",
  8643=>"001011111",
  8644=>"100100001",
  8645=>"010011111",
  8646=>"001001111",
  8647=>"101101111",
  8648=>"111111011",
  8649=>"001001011",
  8650=>"110111111",
  8651=>"110111011",
  8652=>"110011100",
  8653=>"010000101",
  8654=>"001100011",
  8655=>"010100111",
  8656=>"100011010",
  8657=>"000111000",
  8658=>"110010100",
  8659=>"101110011",
  8660=>"001011010",
  8661=>"100010001",
  8662=>"101111111",
  8663=>"111011111",
  8664=>"110111011",
  8665=>"001111011",
  8666=>"000100001",
  8667=>"001000011",
  8668=>"101001000",
  8669=>"000010110",
  8670=>"100011011",
  8671=>"111011101",
  8672=>"111001000",
  8673=>"100000101",
  8674=>"010000110",
  8675=>"000000000",
  8676=>"110101011",
  8677=>"000101000",
  8678=>"000000111",
  8679=>"001000110",
  8680=>"011111010",
  8681=>"001000011",
  8682=>"010110000",
  8683=>"101011011",
  8684=>"010000001",
  8685=>"001100010",
  8686=>"101000101",
  8687=>"111101111",
  8688=>"000000100",
  8689=>"110010110",
  8690=>"011011101",
  8691=>"010100100",
  8692=>"001010001",
  8693=>"110010000",
  8694=>"011011111",
  8695=>"111110000",
  8696=>"110110110",
  8697=>"010111001",
  8698=>"111101101",
  8699=>"111010011",
  8700=>"101111001",
  8701=>"010111000",
  8702=>"010010100",
  8703=>"010010010",
  8704=>"111100110",
  8705=>"100010111",
  8706=>"010110111",
  8707=>"101111010",
  8708=>"000001111",
  8709=>"100011000",
  8710=>"101111000",
  8711=>"000111000",
  8712=>"101011100",
  8713=>"111110110",
  8714=>"010101101",
  8715=>"101101011",
  8716=>"000110110",
  8717=>"001000111",
  8718=>"011100000",
  8719=>"110110111",
  8720=>"000001111",
  8721=>"001101100",
  8722=>"010001111",
  8723=>"110111110",
  8724=>"100111110",
  8725=>"010011100",
  8726=>"011110011",
  8727=>"111110011",
  8728=>"100000011",
  8729=>"100101100",
  8730=>"000011101",
  8731=>"110110111",
  8732=>"110010001",
  8733=>"011111100",
  8734=>"101101100",
  8735=>"010100011",
  8736=>"100111100",
  8737=>"010011010",
  8738=>"000101110",
  8739=>"101111010",
  8740=>"100010011",
  8741=>"100111010",
  8742=>"111010101",
  8743=>"101110101",
  8744=>"101101011",
  8745=>"110111110",
  8746=>"100101111",
  8747=>"101000010",
  8748=>"010110111",
  8749=>"101110110",
  8750=>"001000011",
  8751=>"000001110",
  8752=>"100010010",
  8753=>"101100101",
  8754=>"011101111",
  8755=>"111011001",
  8756=>"101101110",
  8757=>"111001111",
  8758=>"011000111",
  8759=>"011010100",
  8760=>"111111010",
  8761=>"011110101",
  8762=>"110010110",
  8763=>"000000001",
  8764=>"100100100",
  8765=>"010001111",
  8766=>"111010111",
  8767=>"011011111",
  8768=>"010011000",
  8769=>"011111111",
  8770=>"111010000",
  8771=>"100101100",
  8772=>"110110101",
  8773=>"101001110",
  8774=>"000011110",
  8775=>"011110000",
  8776=>"100110000",
  8777=>"111001010",
  8778=>"000110111",
  8779=>"010001110",
  8780=>"111111111",
  8781=>"010101011",
  8782=>"001000011",
  8783=>"000001010",
  8784=>"110000000",
  8785=>"000011110",
  8786=>"100001110",
  8787=>"101101111",
  8788=>"111010111",
  8789=>"000111100",
  8790=>"111100100",
  8791=>"011001110",
  8792=>"100001010",
  8793=>"110110100",
  8794=>"111001101",
  8795=>"000001001",
  8796=>"111101100",
  8797=>"010110000",
  8798=>"001100100",
  8799=>"100111100",
  8800=>"010000100",
  8801=>"100000101",
  8802=>"101011000",
  8803=>"011000101",
  8804=>"111010111",
  8805=>"111100101",
  8806=>"010010000",
  8807=>"010010100",
  8808=>"101000000",
  8809=>"010011001",
  8810=>"100110011",
  8811=>"111111111",
  8812=>"000111011",
  8813=>"101110110",
  8814=>"111110101",
  8815=>"011011010",
  8816=>"110110111",
  8817=>"111100101",
  8818=>"011100000",
  8819=>"001001011",
  8820=>"110111011",
  8821=>"000100100",
  8822=>"111111111",
  8823=>"101110001",
  8824=>"000010111",
  8825=>"100000100",
  8826=>"010100000",
  8827=>"101100111",
  8828=>"111100110",
  8829=>"011011111",
  8830=>"000101000",
  8831=>"001010011",
  8832=>"000011011",
  8833=>"111110101",
  8834=>"101011100",
  8835=>"001000010",
  8836=>"110101100",
  8837=>"101000101",
  8838=>"010100001",
  8839=>"101101000",
  8840=>"100000110",
  8841=>"010101101",
  8842=>"011101100",
  8843=>"000001110",
  8844=>"101011101",
  8845=>"101001000",
  8846=>"000000100",
  8847=>"011010010",
  8848=>"101010011",
  8849=>"100110000",
  8850=>"011101010",
  8851=>"111000010",
  8852=>"110010010",
  8853=>"110101111",
  8854=>"011001010",
  8855=>"101010000",
  8856=>"111101101",
  8857=>"111110000",
  8858=>"101110011",
  8859=>"100011010",
  8860=>"110101010",
  8861=>"000111111",
  8862=>"111111101",
  8863=>"100101011",
  8864=>"100010100",
  8865=>"001001111",
  8866=>"001101101",
  8867=>"001000001",
  8868=>"011001000",
  8869=>"011100001",
  8870=>"001001011",
  8871=>"000100110",
  8872=>"111111111",
  8873=>"111011001",
  8874=>"000000000",
  8875=>"001011100",
  8876=>"011101011",
  8877=>"011100100",
  8878=>"101011111",
  8879=>"011101010",
  8880=>"000100100",
  8881=>"110010101",
  8882=>"001000011",
  8883=>"111111110",
  8884=>"110000011",
  8885=>"100000000",
  8886=>"101111111",
  8887=>"110110010",
  8888=>"110001111",
  8889=>"111110100",
  8890=>"001111011",
  8891=>"000100111",
  8892=>"011101100",
  8893=>"100111100",
  8894=>"001101101",
  8895=>"001100011",
  8896=>"100110011",
  8897=>"101110111",
  8898=>"101011100",
  8899=>"101111111",
  8900=>"011100101",
  8901=>"110001010",
  8902=>"111011101",
  8903=>"100000111",
  8904=>"101110001",
  8905=>"000000101",
  8906=>"110100010",
  8907=>"011010100",
  8908=>"000001011",
  8909=>"011001000",
  8910=>"001010011",
  8911=>"110101000",
  8912=>"110001011",
  8913=>"111100111",
  8914=>"001110000",
  8915=>"100100010",
  8916=>"101001000",
  8917=>"011001101",
  8918=>"100111010",
  8919=>"110111101",
  8920=>"111111101",
  8921=>"110000000",
  8922=>"111001001",
  8923=>"101011010",
  8924=>"001010001",
  8925=>"001000111",
  8926=>"000110100",
  8927=>"011010001",
  8928=>"110001100",
  8929=>"011000011",
  8930=>"000001011",
  8931=>"011000011",
  8932=>"010000000",
  8933=>"011001011",
  8934=>"100000011",
  8935=>"111011101",
  8936=>"110111100",
  8937=>"000101111",
  8938=>"100100110",
  8939=>"001000000",
  8940=>"010001101",
  8941=>"100100101",
  8942=>"010000100",
  8943=>"100000111",
  8944=>"111110101",
  8945=>"101101011",
  8946=>"001100011",
  8947=>"110010101",
  8948=>"110111011",
  8949=>"110000101",
  8950=>"000010011",
  8951=>"110001111",
  8952=>"010100101",
  8953=>"101011111",
  8954=>"101110101",
  8955=>"110101110",
  8956=>"011111000",
  8957=>"011101111",
  8958=>"111011101",
  8959=>"000101001",
  8960=>"000011011",
  8961=>"001101011",
  8962=>"101001111",
  8963=>"101000110",
  8964=>"011010100",
  8965=>"100000111",
  8966=>"001011100",
  8967=>"011001100",
  8968=>"101010011",
  8969=>"110011011",
  8970=>"010010000",
  8971=>"010110000",
  8972=>"100001111",
  8973=>"010100010",
  8974=>"010010000",
  8975=>"110111110",
  8976=>"011110011",
  8977=>"110011101",
  8978=>"000011100",
  8979=>"100101001",
  8980=>"011111111",
  8981=>"000001011",
  8982=>"010000100",
  8983=>"101101000",
  8984=>"011101111",
  8985=>"110111110",
  8986=>"100000001",
  8987=>"111111101",
  8988=>"110001001",
  8989=>"110011100",
  8990=>"110010011",
  8991=>"100101000",
  8992=>"000100001",
  8993=>"100011111",
  8994=>"000011011",
  8995=>"111110110",
  8996=>"111101011",
  8997=>"000001101",
  8998=>"010000010",
  8999=>"001100100",
  9000=>"111001100",
  9001=>"000011110",
  9002=>"011000011",
  9003=>"100111010",
  9004=>"101011100",
  9005=>"010011000",
  9006=>"101110101",
  9007=>"100001101",
  9008=>"111110100",
  9009=>"100110101",
  9010=>"100000111",
  9011=>"010100010",
  9012=>"100001011",
  9013=>"110101100",
  9014=>"011100100",
  9015=>"110010111",
  9016=>"101000110",
  9017=>"111111001",
  9018=>"100001011",
  9019=>"101000010",
  9020=>"000011100",
  9021=>"011010010",
  9022=>"000010101",
  9023=>"000000010",
  9024=>"011111100",
  9025=>"100010111",
  9026=>"011110101",
  9027=>"011011111",
  9028=>"000100000",
  9029=>"100001111",
  9030=>"111110110",
  9031=>"101111101",
  9032=>"000010011",
  9033=>"111111100",
  9034=>"000000110",
  9035=>"110111001",
  9036=>"111101000",
  9037=>"011010100",
  9038=>"001011100",
  9039=>"101100011",
  9040=>"010100000",
  9041=>"000000010",
  9042=>"111011101",
  9043=>"111011100",
  9044=>"000000011",
  9045=>"101110101",
  9046=>"110111000",
  9047=>"111101111",
  9048=>"010110010",
  9049=>"100100001",
  9050=>"011111100",
  9051=>"010110110",
  9052=>"001110100",
  9053=>"101111101",
  9054=>"110000110",
  9055=>"010000100",
  9056=>"100100111",
  9057=>"000011001",
  9058=>"101100010",
  9059=>"110110111",
  9060=>"100100111",
  9061=>"110100101",
  9062=>"100101110",
  9063=>"001101110",
  9064=>"111101001",
  9065=>"010100001",
  9066=>"011010000",
  9067=>"000100111",
  9068=>"011000001",
  9069=>"101101000",
  9070=>"110000000",
  9071=>"100011110",
  9072=>"000111010",
  9073=>"001100100",
  9074=>"011000011",
  9075=>"010111101",
  9076=>"011011011",
  9077=>"110111111",
  9078=>"100111011",
  9079=>"101011110",
  9080=>"110101111",
  9081=>"100011000",
  9082=>"001100010",
  9083=>"111100110",
  9084=>"110110011",
  9085=>"100100101",
  9086=>"000000010",
  9087=>"110111110",
  9088=>"000010011",
  9089=>"100111111",
  9090=>"111100001",
  9091=>"110000000",
  9092=>"100100111",
  9093=>"011010100",
  9094=>"101100000",
  9095=>"111001000",
  9096=>"111101100",
  9097=>"101000101",
  9098=>"000100011",
  9099=>"001001011",
  9100=>"000011000",
  9101=>"100100101",
  9102=>"011101111",
  9103=>"001101111",
  9104=>"011010001",
  9105=>"001111001",
  9106=>"101001001",
  9107=>"110000000",
  9108=>"011010100",
  9109=>"111111011",
  9110=>"101111000",
  9111=>"110001100",
  9112=>"101010101",
  9113=>"000001010",
  9114=>"001111110",
  9115=>"010101011",
  9116=>"111010001",
  9117=>"101011000",
  9118=>"000011000",
  9119=>"011000001",
  9120=>"111100011",
  9121=>"100000101",
  9122=>"000001000",
  9123=>"001000101",
  9124=>"000011001",
  9125=>"000010101",
  9126=>"001011101",
  9127=>"000110010",
  9128=>"110001110",
  9129=>"110101110",
  9130=>"110110111",
  9131=>"110010010",
  9132=>"101101011",
  9133=>"110111100",
  9134=>"001111010",
  9135=>"001011011",
  9136=>"111101110",
  9137=>"101001101",
  9138=>"101110001",
  9139=>"001001011",
  9140=>"000101100",
  9141=>"100011101",
  9142=>"001110000",
  9143=>"101001111",
  9144=>"001010101",
  9145=>"010001010",
  9146=>"011111110",
  9147=>"000111100",
  9148=>"101111111",
  9149=>"010000010",
  9150=>"011111111",
  9151=>"010110111",
  9152=>"101111111",
  9153=>"011110010",
  9154=>"000101000",
  9155=>"001100101",
  9156=>"011110111",
  9157=>"011010111",
  9158=>"011100001",
  9159=>"110010110",
  9160=>"001000110",
  9161=>"000110100",
  9162=>"010001001",
  9163=>"000000111",
  9164=>"010111000",
  9165=>"101000100",
  9166=>"100000001",
  9167=>"101010111",
  9168=>"100000100",
  9169=>"100011100",
  9170=>"001000110",
  9171=>"010101001",
  9172=>"001000001",
  9173=>"101110100",
  9174=>"100101100",
  9175=>"001111110",
  9176=>"011110110",
  9177=>"000101110",
  9178=>"111101001",
  9179=>"111111110",
  9180=>"111010110",
  9181=>"110110010",
  9182=>"000010100",
  9183=>"010001011",
  9184=>"111111111",
  9185=>"111101001",
  9186=>"011110100",
  9187=>"101110110",
  9188=>"010000100",
  9189=>"100011010",
  9190=>"101101110",
  9191=>"001111110",
  9192=>"111001111",
  9193=>"110001101",
  9194=>"011011000",
  9195=>"100101001",
  9196=>"111110110",
  9197=>"111110010",
  9198=>"101010011",
  9199=>"101111011",
  9200=>"000101010",
  9201=>"011111111",
  9202=>"101011001",
  9203=>"010101011",
  9204=>"011111000",
  9205=>"010010100",
  9206=>"011001010",
  9207=>"000100101",
  9208=>"010101111",
  9209=>"001111011",
  9210=>"111001110",
  9211=>"011010011",
  9212=>"110010010",
  9213=>"101011101",
  9214=>"101100101",
  9215=>"101100101",
  9216=>"011001010",
  9217=>"101101000",
  9218=>"000011101",
  9219=>"000111000",
  9220=>"001100111",
  9221=>"111100011",
  9222=>"000110010",
  9223=>"000001010",
  9224=>"111001100",
  9225=>"011010011",
  9226=>"111011100",
  9227=>"111000000",
  9228=>"100011110",
  9229=>"011011111",
  9230=>"001110100",
  9231=>"011111110",
  9232=>"101111100",
  9233=>"100011001",
  9234=>"000000111",
  9235=>"001100010",
  9236=>"000000011",
  9237=>"010100001",
  9238=>"001010101",
  9239=>"110101000",
  9240=>"010000111",
  9241=>"000111110",
  9242=>"001000011",
  9243=>"110010010",
  9244=>"000100101",
  9245=>"000000000",
  9246=>"010100001",
  9247=>"000011000",
  9248=>"001100000",
  9249=>"111011010",
  9250=>"110110110",
  9251=>"101001100",
  9252=>"101011010",
  9253=>"100111011",
  9254=>"001101111",
  9255=>"101110111",
  9256=>"011110100",
  9257=>"111111010",
  9258=>"011101101",
  9259=>"000000011",
  9260=>"010001010",
  9261=>"000111000",
  9262=>"000111001",
  9263=>"001000011",
  9264=>"100111100",
  9265=>"111000110",
  9266=>"001000110",
  9267=>"010110010",
  9268=>"000100110",
  9269=>"000000110",
  9270=>"110010001",
  9271=>"111111000",
  9272=>"001001100",
  9273=>"101000010",
  9274=>"101100101",
  9275=>"111100011",
  9276=>"100101110",
  9277=>"010111011",
  9278=>"011000000",
  9279=>"000001011",
  9280=>"010000011",
  9281=>"000001010",
  9282=>"110011011",
  9283=>"001100010",
  9284=>"010110111",
  9285=>"000011101",
  9286=>"110010111",
  9287=>"011100001",
  9288=>"010101100",
  9289=>"001110010",
  9290=>"101111000",
  9291=>"110110010",
  9292=>"001111010",
  9293=>"101101100",
  9294=>"101000010",
  9295=>"111000010",
  9296=>"100000001",
  9297=>"111110111",
  9298=>"000100110",
  9299=>"100000011",
  9300=>"111000000",
  9301=>"000100000",
  9302=>"000100101",
  9303=>"010100010",
  9304=>"111100101",
  9305=>"001111100",
  9306=>"001010101",
  9307=>"100010110",
  9308=>"111011010",
  9309=>"001100001",
  9310=>"101001111",
  9311=>"100011111",
  9312=>"000011001",
  9313=>"010110010",
  9314=>"011101000",
  9315=>"000010111",
  9316=>"110001110",
  9317=>"000110011",
  9318=>"011111100",
  9319=>"001101011",
  9320=>"111000110",
  9321=>"101001001",
  9322=>"101000000",
  9323=>"000100110",
  9324=>"011111010",
  9325=>"000011001",
  9326=>"000100000",
  9327=>"111111111",
  9328=>"000111011",
  9329=>"110101100",
  9330=>"000001010",
  9331=>"000110010",
  9332=>"010011110",
  9333=>"110110010",
  9334=>"001110000",
  9335=>"111101100",
  9336=>"110010011",
  9337=>"101110001",
  9338=>"100111011",
  9339=>"010100010",
  9340=>"001010001",
  9341=>"001110000",
  9342=>"111111111",
  9343=>"001001011",
  9344=>"000100110",
  9345=>"101000011",
  9346=>"100100111",
  9347=>"111001101",
  9348=>"110100111",
  9349=>"100010011",
  9350=>"000011111",
  9351=>"101001001",
  9352=>"011101101",
  9353=>"000000000",
  9354=>"001110100",
  9355=>"101100011",
  9356=>"011100000",
  9357=>"111101101",
  9358=>"100010011",
  9359=>"001110110",
  9360=>"010000010",
  9361=>"000100010",
  9362=>"111010111",
  9363=>"011111101",
  9364=>"000001110",
  9365=>"101000000",
  9366=>"010111100",
  9367=>"010110000",
  9368=>"011010000",
  9369=>"000111000",
  9370=>"110110010",
  9371=>"001010100",
  9372=>"000111110",
  9373=>"000001101",
  9374=>"001110011",
  9375=>"010101011",
  9376=>"000011010",
  9377=>"000010000",
  9378=>"001100010",
  9379=>"000101101",
  9380=>"110101000",
  9381=>"011110000",
  9382=>"110001001",
  9383=>"001010110",
  9384=>"111001010",
  9385=>"110110111",
  9386=>"111111111",
  9387=>"010111101",
  9388=>"001001110",
  9389=>"010100110",
  9390=>"011110010",
  9391=>"100110011",
  9392=>"011010111",
  9393=>"000011001",
  9394=>"000101000",
  9395=>"010110101",
  9396=>"101001111",
  9397=>"011000001",
  9398=>"100001101",
  9399=>"100110000",
  9400=>"000111110",
  9401=>"000001000",
  9402=>"011111011",
  9403=>"101010010",
  9404=>"000110110",
  9405=>"001101000",
  9406=>"110000000",
  9407=>"011011101",
  9408=>"100010101",
  9409=>"001100010",
  9410=>"111100000",
  9411=>"000111000",
  9412=>"101010011",
  9413=>"011101010",
  9414=>"011010111",
  9415=>"110001000",
  9416=>"000111100",
  9417=>"001110100",
  9418=>"101100001",
  9419=>"111000000",
  9420=>"011001100",
  9421=>"001010010",
  9422=>"011100101",
  9423=>"000110010",
  9424=>"100011110",
  9425=>"001000001",
  9426=>"110111110",
  9427=>"110011110",
  9428=>"010110100",
  9429=>"000001010",
  9430=>"011000110",
  9431=>"001010000",
  9432=>"000001000",
  9433=>"111100001",
  9434=>"100001110",
  9435=>"011101100",
  9436=>"001011001",
  9437=>"100100000",
  9438=>"001000100",
  9439=>"111000111",
  9440=>"010111001",
  9441=>"001101101",
  9442=>"101011011",
  9443=>"110010100",
  9444=>"011101110",
  9445=>"110001001",
  9446=>"100101000",
  9447=>"101100000",
  9448=>"111110010",
  9449=>"100000111",
  9450=>"000000001",
  9451=>"111001111",
  9452=>"111101001",
  9453=>"101110000",
  9454=>"100110110",
  9455=>"111001111",
  9456=>"111100101",
  9457=>"111000000",
  9458=>"000111010",
  9459=>"011010101",
  9460=>"110111010",
  9461=>"101000101",
  9462=>"101001110",
  9463=>"000110111",
  9464=>"011111000",
  9465=>"000011000",
  9466=>"101110000",
  9467=>"011001010",
  9468=>"101001101",
  9469=>"101110111",
  9470=>"111101101",
  9471=>"011111111",
  9472=>"001011001",
  9473=>"000000101",
  9474=>"111000010",
  9475=>"001100111",
  9476=>"011000101",
  9477=>"101011111",
  9478=>"010001110",
  9479=>"101111101",
  9480=>"111101000",
  9481=>"100000100",
  9482=>"000100010",
  9483=>"110100110",
  9484=>"000101111",
  9485=>"000010000",
  9486=>"111111000",
  9487=>"011100010",
  9488=>"101110110",
  9489=>"000110011",
  9490=>"001000000",
  9491=>"111000000",
  9492=>"000100101",
  9493=>"000110011",
  9494=>"001000111",
  9495=>"111001110",
  9496=>"010011010",
  9497=>"110000000",
  9498=>"000000100",
  9499=>"100000101",
  9500=>"000100011",
  9501=>"011100100",
  9502=>"101000101",
  9503=>"011011111",
  9504=>"010101101",
  9505=>"101010000",
  9506=>"010001101",
  9507=>"011100010",
  9508=>"011111101",
  9509=>"101011011",
  9510=>"001011110",
  9511=>"010110011",
  9512=>"010110111",
  9513=>"100000010",
  9514=>"100000010",
  9515=>"001001000",
  9516=>"111001010",
  9517=>"111000000",
  9518=>"000000001",
  9519=>"001011001",
  9520=>"000100010",
  9521=>"101111101",
  9522=>"001000010",
  9523=>"100111000",
  9524=>"111011101",
  9525=>"101010001",
  9526=>"101100001",
  9527=>"011000111",
  9528=>"010000011",
  9529=>"011100100",
  9530=>"110100000",
  9531=>"001011000",
  9532=>"101001011",
  9533=>"001111001",
  9534=>"000101100",
  9535=>"111111111",
  9536=>"110000010",
  9537=>"101111101",
  9538=>"000110010",
  9539=>"101101101",
  9540=>"001001110",
  9541=>"111100000",
  9542=>"101100101",
  9543=>"000001010",
  9544=>"100000010",
  9545=>"000001000",
  9546=>"110101111",
  9547=>"111001110",
  9548=>"101101010",
  9549=>"111011011",
  9550=>"110110011",
  9551=>"101010001",
  9552=>"010100111",
  9553=>"011011000",
  9554=>"000001000",
  9555=>"011010101",
  9556=>"010000001",
  9557=>"100010011",
  9558=>"110100000",
  9559=>"100001100",
  9560=>"000000000",
  9561=>"110010010",
  9562=>"001011001",
  9563=>"010001001",
  9564=>"110010001",
  9565=>"011111111",
  9566=>"001001111",
  9567=>"100100100",
  9568=>"110101011",
  9569=>"001111110",
  9570=>"000001001",
  9571=>"110110110",
  9572=>"101100001",
  9573=>"011100110",
  9574=>"000010110",
  9575=>"100010100",
  9576=>"011001101",
  9577=>"001011110",
  9578=>"011100100",
  9579=>"100010111",
  9580=>"011011100",
  9581=>"000110111",
  9582=>"100001111",
  9583=>"011100010",
  9584=>"000101110",
  9585=>"111001111",
  9586=>"000111001",
  9587=>"000101011",
  9588=>"101011101",
  9589=>"110100101",
  9590=>"100110101",
  9591=>"100100100",
  9592=>"001011111",
  9593=>"101100110",
  9594=>"000100000",
  9595=>"101001111",
  9596=>"000001001",
  9597=>"000000001",
  9598=>"010010110",
  9599=>"100111010",
  9600=>"101101111",
  9601=>"110101100",
  9602=>"000101010",
  9603=>"000110010",
  9604=>"100100101",
  9605=>"001110100",
  9606=>"001011000",
  9607=>"000001010",
  9608=>"010100011",
  9609=>"110010011",
  9610=>"101000101",
  9611=>"010000010",
  9612=>"111101100",
  9613=>"001100100",
  9614=>"011010111",
  9615=>"100010010",
  9616=>"101001000",
  9617=>"110011100",
  9618=>"000100100",
  9619=>"011100001",
  9620=>"011011000",
  9621=>"110000111",
  9622=>"010111011",
  9623=>"110000000",
  9624=>"110010010",
  9625=>"100001111",
  9626=>"100100100",
  9627=>"000000111",
  9628=>"101000010",
  9629=>"000001010",
  9630=>"111000101",
  9631=>"000011110",
  9632=>"001100000",
  9633=>"110000110",
  9634=>"011111101",
  9635=>"001001010",
  9636=>"111011010",
  9637=>"011010000",
  9638=>"001000101",
  9639=>"101110101",
  9640=>"011110001",
  9641=>"000110011",
  9642=>"011100011",
  9643=>"001011010",
  9644=>"010000001",
  9645=>"011111111",
  9646=>"111001000",
  9647=>"000110011",
  9648=>"010001001",
  9649=>"110010000",
  9650=>"110011000",
  9651=>"011011101",
  9652=>"100001100",
  9653=>"001010001",
  9654=>"011001011",
  9655=>"100101110",
  9656=>"110111100",
  9657=>"110111100",
  9658=>"100111101",
  9659=>"101110010",
  9660=>"101010110",
  9661=>"100100110",
  9662=>"110010000",
  9663=>"110100010",
  9664=>"001110010",
  9665=>"000110100",
  9666=>"011101110",
  9667=>"011100000",
  9668=>"110011111",
  9669=>"001110110",
  9670=>"000000001",
  9671=>"101101111",
  9672=>"110011111",
  9673=>"010100111",
  9674=>"011000101",
  9675=>"100101111",
  9676=>"101100101",
  9677=>"000011010",
  9678=>"101101000",
  9679=>"010110101",
  9680=>"100010011",
  9681=>"000111100",
  9682=>"110100000",
  9683=>"010111100",
  9684=>"100011111",
  9685=>"001111110",
  9686=>"010000111",
  9687=>"001000110",
  9688=>"001110111",
  9689=>"111110000",
  9690=>"110010001",
  9691=>"110101010",
  9692=>"110101011",
  9693=>"011100011",
  9694=>"110000100",
  9695=>"010111001",
  9696=>"000101011",
  9697=>"000011110",
  9698=>"000110000",
  9699=>"111010000",
  9700=>"100010101",
  9701=>"111111000",
  9702=>"101101110",
  9703=>"111000010",
  9704=>"110100101",
  9705=>"011100100",
  9706=>"111100011",
  9707=>"001000011",
  9708=>"100011010",
  9709=>"100110100",
  9710=>"000000010",
  9711=>"000010010",
  9712=>"101010011",
  9713=>"000110011",
  9714=>"010100111",
  9715=>"001101101",
  9716=>"101110111",
  9717=>"111001110",
  9718=>"010000011",
  9719=>"101100111",
  9720=>"101100010",
  9721=>"110001001",
  9722=>"011101000",
  9723=>"111000010",
  9724=>"100110111",
  9725=>"100001000",
  9726=>"010001110",
  9727=>"100000111",
  9728=>"100000001",
  9729=>"011011100",
  9730=>"110110001",
  9731=>"010001011",
  9732=>"100000011",
  9733=>"001011011",
  9734=>"011000111",
  9735=>"000010001",
  9736=>"000000010",
  9737=>"000110000",
  9738=>"101000011",
  9739=>"110001100",
  9740=>"011111111",
  9741=>"001001010",
  9742=>"011011010",
  9743=>"111011011",
  9744=>"110111001",
  9745=>"011100101",
  9746=>"011110010",
  9747=>"110111001",
  9748=>"110101011",
  9749=>"000010101",
  9750=>"011111101",
  9751=>"101111111",
  9752=>"100100000",
  9753=>"010101110",
  9754=>"010010010",
  9755=>"111001101",
  9756=>"000000010",
  9757=>"110000010",
  9758=>"101110111",
  9759=>"001011111",
  9760=>"011110011",
  9761=>"001011010",
  9762=>"000111110",
  9763=>"000111111",
  9764=>"111101011",
  9765=>"010000100",
  9766=>"110010010",
  9767=>"010010101",
  9768=>"000000111",
  9769=>"010000001",
  9770=>"111110111",
  9771=>"011100001",
  9772=>"011110001",
  9773=>"000000010",
  9774=>"110101011",
  9775=>"100111101",
  9776=>"010001000",
  9777=>"110101110",
  9778=>"100010011",
  9779=>"001001010",
  9780=>"010011000",
  9781=>"111001011",
  9782=>"000001010",
  9783=>"101101101",
  9784=>"110111100",
  9785=>"001011000",
  9786=>"000000111",
  9787=>"011010010",
  9788=>"000111011",
  9789=>"010111111",
  9790=>"011111010",
  9791=>"101001011",
  9792=>"001110101",
  9793=>"111111000",
  9794=>"110000111",
  9795=>"101001010",
  9796=>"010000011",
  9797=>"100101001",
  9798=>"100000101",
  9799=>"100111011",
  9800=>"011000000",
  9801=>"011111101",
  9802=>"000101110",
  9803=>"000110111",
  9804=>"001110000",
  9805=>"000001001",
  9806=>"011100000",
  9807=>"010011110",
  9808=>"011001100",
  9809=>"010000001",
  9810=>"110011011",
  9811=>"110010100",
  9812=>"101111100",
  9813=>"111100100",
  9814=>"000101001",
  9815=>"011101111",
  9816=>"111010011",
  9817=>"001011011",
  9818=>"010101101",
  9819=>"111011001",
  9820=>"110011001",
  9821=>"110110111",
  9822=>"101001000",
  9823=>"001100010",
  9824=>"110011110",
  9825=>"010001110",
  9826=>"000101101",
  9827=>"111100001",
  9828=>"110001010",
  9829=>"100110011",
  9830=>"101100001",
  9831=>"100010010",
  9832=>"111100100",
  9833=>"000100011",
  9834=>"101011101",
  9835=>"111100101",
  9836=>"001000100",
  9837=>"101100011",
  9838=>"001111111",
  9839=>"010010001",
  9840=>"111110001",
  9841=>"001001101",
  9842=>"001001011",
  9843=>"101011000",
  9844=>"110001100",
  9845=>"100110111",
  9846=>"000110110",
  9847=>"000000000",
  9848=>"000000001",
  9849=>"011111011",
  9850=>"110011111",
  9851=>"100011011",
  9852=>"111111111",
  9853=>"010111111",
  9854=>"001000111",
  9855=>"100100111",
  9856=>"000110101",
  9857=>"010001011",
  9858=>"011001110",
  9859=>"100101011",
  9860=>"011001100",
  9861=>"011011101",
  9862=>"101101100",
  9863=>"011111011",
  9864=>"010111101",
  9865=>"001110011",
  9866=>"011000000",
  9867=>"011101111",
  9868=>"001101001",
  9869=>"011111101",
  9870=>"000010000",
  9871=>"110010110",
  9872=>"110110010",
  9873=>"100101010",
  9874=>"011101110",
  9875=>"101100010",
  9876=>"111100001",
  9877=>"000111100",
  9878=>"011000011",
  9879=>"110100101",
  9880=>"100000010",
  9881=>"010110111",
  9882=>"101011010",
  9883=>"100001100",
  9884=>"010001110",
  9885=>"101001011",
  9886=>"001000000",
  9887=>"001000000",
  9888=>"000010101",
  9889=>"110111010",
  9890=>"011001101",
  9891=>"000001000",
  9892=>"101110111",
  9893=>"101110100",
  9894=>"011001110",
  9895=>"000010000",
  9896=>"001001100",
  9897=>"010100111",
  9898=>"000000111",
  9899=>"111001000",
  9900=>"101010100",
  9901=>"011001010",
  9902=>"111111010",
  9903=>"011011100",
  9904=>"000110111",
  9905=>"001010011",
  9906=>"011010000",
  9907=>"010101011",
  9908=>"110100110",
  9909=>"001000110",
  9910=>"010011000",
  9911=>"011010001",
  9912=>"101101000",
  9913=>"000001111",
  9914=>"100000110",
  9915=>"001000011",
  9916=>"110010001",
  9917=>"010100110",
  9918=>"101000010",
  9919=>"010011010",
  9920=>"000110001",
  9921=>"100110011",
  9922=>"101001000",
  9923=>"000010011",
  9924=>"011010001",
  9925=>"011001100",
  9926=>"011010000",
  9927=>"101111100",
  9928=>"101100111",
  9929=>"110011111",
  9930=>"010011011",
  9931=>"101001110",
  9932=>"010101101",
  9933=>"100001001",
  9934=>"010111010",
  9935=>"011110110",
  9936=>"101100000",
  9937=>"111010111",
  9938=>"011101101",
  9939=>"000010010",
  9940=>"001010001",
  9941=>"110110111",
  9942=>"001001101",
  9943=>"100100010",
  9944=>"100111101",
  9945=>"011000100",
  9946=>"100001000",
  9947=>"111101110",
  9948=>"111101110",
  9949=>"100110000",
  9950=>"101100111",
  9951=>"111110100",
  9952=>"011101101",
  9953=>"001000010",
  9954=>"110111001",
  9955=>"111001010",
  9956=>"100101011",
  9957=>"101111100",
  9958=>"110111010",
  9959=>"101110000",
  9960=>"101011001",
  9961=>"100101110",
  9962=>"111110010",
  9963=>"110111101",
  9964=>"100011111",
  9965=>"000100110",
  9966=>"011011001",
  9967=>"001110101",
  9968=>"010011100",
  9969=>"101000111",
  9970=>"000000110",
  9971=>"110100000",
  9972=>"111111010",
  9973=>"001000100",
  9974=>"000110000",
  9975=>"000100011",
  9976=>"001011011",
  9977=>"001100011",
  9978=>"011010100",
  9979=>"110110010",
  9980=>"000001101",
  9981=>"100000001",
  9982=>"100110011",
  9983=>"101001111",
  9984=>"000100101",
  9985=>"010110000",
  9986=>"010010001",
  9987=>"111001001",
  9988=>"000101001",
  9989=>"001110100",
  9990=>"000101010",
  9991=>"000001111",
  9992=>"110101010",
  9993=>"111111110",
  9994=>"111001101",
  9995=>"011010011",
  9996=>"001110010",
  9997=>"001101101",
  9998=>"110001110",
  9999=>"101111101",
  10000=>"110011001",
  10001=>"100110100",
  10002=>"100101100",
  10003=>"110111101",
  10004=>"101010110",
  10005=>"100010110",
  10006=>"001101111",
  10007=>"111001011",
  10008=>"000011111",
  10009=>"101010000",
  10010=>"100110110",
  10011=>"010010110",
  10012=>"101111100",
  10013=>"100001110",
  10014=>"100011000",
  10015=>"100010100",
  10016=>"000000001",
  10017=>"100010010",
  10018=>"011111101",
  10019=>"011000000",
  10020=>"010111001",
  10021=>"111111001",
  10022=>"001101111",
  10023=>"011101011",
  10024=>"111001011",
  10025=>"111110100",
  10026=>"111001011",
  10027=>"001110100",
  10028=>"000101111",
  10029=>"000101111",
  10030=>"011010101",
  10031=>"110000010",
  10032=>"100000110",
  10033=>"101111110",
  10034=>"111110110",
  10035=>"111110001",
  10036=>"000000000",
  10037=>"100011000",
  10038=>"111000000",
  10039=>"101011101",
  10040=>"011110110",
  10041=>"100010110",
  10042=>"111111000",
  10043=>"111010001",
  10044=>"000100000",
  10045=>"001110000",
  10046=>"010001001",
  10047=>"000010100",
  10048=>"011101101",
  10049=>"110011111",
  10050=>"111000110",
  10051=>"101010110",
  10052=>"101100110",
  10053=>"101001000",
  10054=>"111011100",
  10055=>"000110010",
  10056=>"000010001",
  10057=>"111011111",
  10058=>"101101001",
  10059=>"000010000",
  10060=>"011000110",
  10061=>"101000001",
  10062=>"000111100",
  10063=>"011101101",
  10064=>"101110100",
  10065=>"110110101",
  10066=>"000110110",
  10067=>"110111011",
  10068=>"001010110",
  10069=>"000101010",
  10070=>"001001110",
  10071=>"101011000",
  10072=>"111110010",
  10073=>"111001011",
  10074=>"001100001",
  10075=>"101001011",
  10076=>"010100010",
  10077=>"111111101",
  10078=>"001001111",
  10079=>"101000101",
  10080=>"100100100",
  10081=>"111000101",
  10082=>"100110111",
  10083=>"100010011",
  10084=>"000101001",
  10085=>"010100100",
  10086=>"011011011",
  10087=>"100110101",
  10088=>"110011000",
  10089=>"101110110",
  10090=>"101010010",
  10091=>"010101101",
  10092=>"100010010",
  10093=>"111000101",
  10094=>"001000110",
  10095=>"111011011",
  10096=>"101100101",
  10097=>"101100110",
  10098=>"101011010",
  10099=>"001010110",
  10100=>"000001000",
  10101=>"110111110",
  10102=>"100110110",
  10103=>"111010111",
  10104=>"101010010",
  10105=>"100110010",
  10106=>"011011111",
  10107=>"010110110",
  10108=>"001010011",
  10109=>"111100100",
  10110=>"001000000",
  10111=>"111101001",
  10112=>"011010000",
  10113=>"001011001",
  10114=>"011001011",
  10115=>"000110011",
  10116=>"110000110",
  10117=>"100001000",
  10118=>"011111010",
  10119=>"011101110",
  10120=>"011111100",
  10121=>"001100001",
  10122=>"000011010",
  10123=>"000011100",
  10124=>"111100000",
  10125=>"101000001",
  10126=>"000011011",
  10127=>"011101000",
  10128=>"001110101",
  10129=>"110110010",
  10130=>"011111000",
  10131=>"011001101",
  10132=>"010001000",
  10133=>"000111000",
  10134=>"100000000",
  10135=>"001100001",
  10136=>"001000111",
  10137=>"000000101",
  10138=>"101000111",
  10139=>"100001001",
  10140=>"111101111",
  10141=>"100001001",
  10142=>"101000111",
  10143=>"000010100",
  10144=>"101000110",
  10145=>"100101011",
  10146=>"100100010",
  10147=>"100011101",
  10148=>"000011101",
  10149=>"010100111",
  10150=>"000011111",
  10151=>"110010100",
  10152=>"010010110",
  10153=>"010111000",
  10154=>"110100100",
  10155=>"110000110",
  10156=>"001100000",
  10157=>"100000110",
  10158=>"101000001",
  10159=>"000010001",
  10160=>"110001000",
  10161=>"100101001",
  10162=>"000011000",
  10163=>"111100011",
  10164=>"110001001",
  10165=>"100111111",
  10166=>"001101100",
  10167=>"001010111",
  10168=>"011011010",
  10169=>"100011011",
  10170=>"111100001",
  10171=>"110001101",
  10172=>"111100000",
  10173=>"111010000",
  10174=>"010011011",
  10175=>"000111110",
  10176=>"011011111",
  10177=>"001111100",
  10178=>"001001101",
  10179=>"010110011",
  10180=>"111000010",
  10181=>"110100111",
  10182=>"101010000",
  10183=>"100111011",
  10184=>"001100001",
  10185=>"011101100",
  10186=>"111000010",
  10187=>"011000011",
  10188=>"110100000",
  10189=>"111000101",
  10190=>"100010010",
  10191=>"110010000",
  10192=>"001101110",
  10193=>"001001100",
  10194=>"100010101",
  10195=>"111000111",
  10196=>"011010101",
  10197=>"110110010",
  10198=>"001100000",
  10199=>"100011111",
  10200=>"001110101",
  10201=>"111111011",
  10202=>"101001100",
  10203=>"011101111",
  10204=>"111111101",
  10205=>"000111101",
  10206=>"011101100",
  10207=>"101000000",
  10208=>"101001001",
  10209=>"101001000",
  10210=>"100011010",
  10211=>"101110000",
  10212=>"000000001",
  10213=>"110100011",
  10214=>"011111111",
  10215=>"101001000",
  10216=>"010110100",
  10217=>"011110100",
  10218=>"101101010",
  10219=>"011001110",
  10220=>"111111111",
  10221=>"010110010",
  10222=>"001000000",
  10223=>"101001010",
  10224=>"010111000",
  10225=>"110110000",
  10226=>"100101011",
  10227=>"011100111",
  10228=>"001111000",
  10229=>"110111000",
  10230=>"101111001",
  10231=>"110101110",
  10232=>"001110010",
  10233=>"100001011",
  10234=>"101100001",
  10235=>"000100100",
  10236=>"000001111",
  10237=>"111111100",
  10238=>"011101010",
  10239=>"100101011",
  10240=>"110110101",
  10241=>"011111011",
  10242=>"010111011",
  10243=>"110100100",
  10244=>"010111111",
  10245=>"010000011",
  10246=>"000101110",
  10247=>"100111001",
  10248=>"000110010",
  10249=>"000001101",
  10250=>"001101101",
  10251=>"100100000",
  10252=>"000110000",
  10253=>"111000100",
  10254=>"101001010",
  10255=>"111000000",
  10256=>"010100011",
  10257=>"010000010",
  10258=>"000110000",
  10259=>"101111000",
  10260=>"111111100",
  10261=>"011110110",
  10262=>"010111100",
  10263=>"011000000",
  10264=>"100000110",
  10265=>"011011000",
  10266=>"101100011",
  10267=>"111100010",
  10268=>"110110010",
  10269=>"111111111",
  10270=>"101110111",
  10271=>"110001111",
  10272=>"110100001",
  10273=>"000000110",
  10274=>"101000101",
  10275=>"110011110",
  10276=>"101110010",
  10277=>"001100010",
  10278=>"100000110",
  10279=>"101101110",
  10280=>"110100100",
  10281=>"100000110",
  10282=>"000011011",
  10283=>"111001001",
  10284=>"111010001",
  10285=>"110001110",
  10286=>"011100011",
  10287=>"101001101",
  10288=>"011111011",
  10289=>"000111100",
  10290=>"110001011",
  10291=>"110001000",
  10292=>"100111000",
  10293=>"000011001",
  10294=>"111100111",
  10295=>"001101011",
  10296=>"100100110",
  10297=>"101001010",
  10298=>"000110110",
  10299=>"000001011",
  10300=>"010000100",
  10301=>"000111101",
  10302=>"000001110",
  10303=>"011100000",
  10304=>"101000000",
  10305=>"101001000",
  10306=>"011001011",
  10307=>"110000001",
  10308=>"110110001",
  10309=>"011101011",
  10310=>"011110111",
  10311=>"100100111",
  10312=>"101111001",
  10313=>"010110101",
  10314=>"101101011",
  10315=>"001100110",
  10316=>"000001111",
  10317=>"011010100",
  10318=>"101110010",
  10319=>"111100101",
  10320=>"100110111",
  10321=>"100101110",
  10322=>"111111101",
  10323=>"000100001",
  10324=>"001111011",
  10325=>"101001110",
  10326=>"010011011",
  10327=>"110001011",
  10328=>"100111111",
  10329=>"010000101",
  10330=>"011001001",
  10331=>"001001110",
  10332=>"110011111",
  10333=>"100100011",
  10334=>"101001010",
  10335=>"100001010",
  10336=>"101110101",
  10337=>"101101010",
  10338=>"001010111",
  10339=>"000010011",
  10340=>"010011100",
  10341=>"010100111",
  10342=>"101001011",
  10343=>"110100101",
  10344=>"010101111",
  10345=>"111000010",
  10346=>"100010100",
  10347=>"000110100",
  10348=>"110001010",
  10349=>"011110001",
  10350=>"000100101",
  10351=>"000011000",
  10352=>"110011011",
  10353=>"000011001",
  10354=>"100100111",
  10355=>"110111111",
  10356=>"100101100",
  10357=>"000000011",
  10358=>"011101100",
  10359=>"000000110",
  10360=>"011110110",
  10361=>"010001000",
  10362=>"110100000",
  10363=>"001100110",
  10364=>"111001110",
  10365=>"010000001",
  10366=>"000110111",
  10367=>"100001000",
  10368=>"101100011",
  10369=>"001100101",
  10370=>"111001100",
  10371=>"000111110",
  10372=>"100100001",
  10373=>"011010111",
  10374=>"100101011",
  10375=>"101000011",
  10376=>"011001110",
  10377=>"010011011",
  10378=>"111111111",
  10379=>"011101101",
  10380=>"101100101",
  10381=>"010101001",
  10382=>"000000100",
  10383=>"001011100",
  10384=>"001100101",
  10385=>"111111110",
  10386=>"110110101",
  10387=>"000100011",
  10388=>"111010100",
  10389=>"110101101",
  10390=>"000110100",
  10391=>"010100100",
  10392=>"000110101",
  10393=>"010000000",
  10394=>"000100000",
  10395=>"011011100",
  10396=>"011100100",
  10397=>"111110001",
  10398=>"101110000",
  10399=>"110110000",
  10400=>"100011100",
  10401=>"111011010",
  10402=>"111100000",
  10403=>"001100110",
  10404=>"001100010",
  10405=>"010101010",
  10406=>"111101101",
  10407=>"010001010",
  10408=>"100000010",
  10409=>"100010001",
  10410=>"011011001",
  10411=>"011100000",
  10412=>"110110111",
  10413=>"100000000",
  10414=>"110101100",
  10415=>"100011011",
  10416=>"101111110",
  10417=>"100110011",
  10418=>"001010100",
  10419=>"001001111",
  10420=>"010110000",
  10421=>"111010010",
  10422=>"100101001",
  10423=>"000111000",
  10424=>"100000111",
  10425=>"001001000",
  10426=>"111011010",
  10427=>"010011111",
  10428=>"100011110",
  10429=>"111110010",
  10430=>"111101000",
  10431=>"101111000",
  10432=>"111110100",
  10433=>"101101001",
  10434=>"001111011",
  10435=>"111101100",
  10436=>"011000111",
  10437=>"001010101",
  10438=>"111100000",
  10439=>"011110000",
  10440=>"110001000",
  10441=>"000001110",
  10442=>"100000100",
  10443=>"100000111",
  10444=>"011110000",
  10445=>"010000111",
  10446=>"011000010",
  10447=>"101000110",
  10448=>"100000001",
  10449=>"100001010",
  10450=>"001111000",
  10451=>"010110100",
  10452=>"111001100",
  10453=>"111101011",
  10454=>"010001011",
  10455=>"111110001",
  10456=>"000110010",
  10457=>"101000111",
  10458=>"001111110",
  10459=>"011100010",
  10460=>"011010111",
  10461=>"011101100",
  10462=>"011111011",
  10463=>"000110011",
  10464=>"101010110",
  10465=>"100100111",
  10466=>"001010100",
  10467=>"111111000",
  10468=>"100100001",
  10469=>"011000101",
  10470=>"000010011",
  10471=>"101011010",
  10472=>"111101110",
  10473=>"110010110",
  10474=>"100110110",
  10475=>"111001001",
  10476=>"100101011",
  10477=>"111011001",
  10478=>"000111010",
  10479=>"010111110",
  10480=>"000011100",
  10481=>"111001101",
  10482=>"000000111",
  10483=>"101101011",
  10484=>"101000101",
  10485=>"111100111",
  10486=>"000000111",
  10487=>"000010000",
  10488=>"000011101",
  10489=>"000001101",
  10490=>"101111011",
  10491=>"011101100",
  10492=>"111110010",
  10493=>"100100001",
  10494=>"011001110",
  10495=>"001000011",
  10496=>"011110110",
  10497=>"000011110",
  10498=>"101110110",
  10499=>"110100000",
  10500=>"110100000",
  10501=>"001010010",
  10502=>"000111110",
  10503=>"000110110",
  10504=>"110101100",
  10505=>"001011001",
  10506=>"001011110",
  10507=>"111001001",
  10508=>"000001000",
  10509=>"011011010",
  10510=>"010101000",
  10511=>"000101011",
  10512=>"100011111",
  10513=>"000000010",
  10514=>"001110000",
  10515=>"110100011",
  10516=>"100011111",
  10517=>"101010001",
  10518=>"000001100",
  10519=>"001000011",
  10520=>"011111100",
  10521=>"101101110",
  10522=>"110111100",
  10523=>"111111010",
  10524=>"000101011",
  10525=>"011001101",
  10526=>"111110001",
  10527=>"010011000",
  10528=>"011000110",
  10529=>"010000111",
  10530=>"000100011",
  10531=>"101000001",
  10532=>"100111111",
  10533=>"010011010",
  10534=>"011010011",
  10535=>"010001000",
  10536=>"000100011",
  10537=>"000110101",
  10538=>"101111110",
  10539=>"110110011",
  10540=>"000010000",
  10541=>"010010001",
  10542=>"110100100",
  10543=>"000010110",
  10544=>"000011000",
  10545=>"001010111",
  10546=>"100111000",
  10547=>"110111100",
  10548=>"100010110",
  10549=>"001110010",
  10550=>"110011101",
  10551=>"000010100",
  10552=>"011101001",
  10553=>"100010001",
  10554=>"001000011",
  10555=>"100110110",
  10556=>"000000100",
  10557=>"001110101",
  10558=>"111100100",
  10559=>"111001011",
  10560=>"000100000",
  10561=>"101011000",
  10562=>"100000100",
  10563=>"110011011",
  10564=>"110000101",
  10565=>"110011010",
  10566=>"010100110",
  10567=>"001011000",
  10568=>"000010110",
  10569=>"001100001",
  10570=>"100100110",
  10571=>"010001111",
  10572=>"011001111",
  10573=>"101011010",
  10574=>"111101000",
  10575=>"101100001",
  10576=>"001111111",
  10577=>"010101110",
  10578=>"000000010",
  10579=>"101011100",
  10580=>"011110100",
  10581=>"110101011",
  10582=>"101010100",
  10583=>"010011110",
  10584=>"101001100",
  10585=>"000010100",
  10586=>"110001111",
  10587=>"101000001",
  10588=>"101000000",
  10589=>"010101110",
  10590=>"111111001",
  10591=>"000000101",
  10592=>"100111110",
  10593=>"111100000",
  10594=>"000010100",
  10595=>"110001100",
  10596=>"100111010",
  10597=>"000101101",
  10598=>"001001100",
  10599=>"101111101",
  10600=>"101011101",
  10601=>"101000000",
  10602=>"011101010",
  10603=>"011011101",
  10604=>"010010111",
  10605=>"110111000",
  10606=>"110010101",
  10607=>"110001100",
  10608=>"010011000",
  10609=>"101001011",
  10610=>"000010000",
  10611=>"010100010",
  10612=>"000111110",
  10613=>"011111001",
  10614=>"011111001",
  10615=>"011110000",
  10616=>"101100111",
  10617=>"011100111",
  10618=>"111100110",
  10619=>"110111111",
  10620=>"001100110",
  10621=>"100100010",
  10622=>"100110011",
  10623=>"111010110",
  10624=>"000000100",
  10625=>"010000010",
  10626=>"010011011",
  10627=>"011110101",
  10628=>"010111111",
  10629=>"011001010",
  10630=>"010111011",
  10631=>"101010000",
  10632=>"001000111",
  10633=>"100000000",
  10634=>"001100110",
  10635=>"001000000",
  10636=>"110010111",
  10637=>"001000001",
  10638=>"110010000",
  10639=>"000110100",
  10640=>"001101010",
  10641=>"010011101",
  10642=>"001000100",
  10643=>"010011101",
  10644=>"110110110",
  10645=>"110111101",
  10646=>"110001001",
  10647=>"100100011",
  10648=>"111110000",
  10649=>"010010010",
  10650=>"001000110",
  10651=>"100110001",
  10652=>"101111001",
  10653=>"010100011",
  10654=>"111101100",
  10655=>"011101101",
  10656=>"100010101",
  10657=>"011000011",
  10658=>"011111010",
  10659=>"001111001",
  10660=>"001000101",
  10661=>"111010100",
  10662=>"111110001",
  10663=>"011110111",
  10664=>"000100010",
  10665=>"110101100",
  10666=>"010000001",
  10667=>"111101100",
  10668=>"000001111",
  10669=>"000100110",
  10670=>"010010000",
  10671=>"111010000",
  10672=>"100111001",
  10673=>"001001110",
  10674=>"000100000",
  10675=>"000000110",
  10676=>"011001110",
  10677=>"110111011",
  10678=>"001010100",
  10679=>"010001111",
  10680=>"111000111",
  10681=>"001101110",
  10682=>"011111111",
  10683=>"110111111",
  10684=>"100100001",
  10685=>"011000111",
  10686=>"000010101",
  10687=>"000001100",
  10688=>"010010101",
  10689=>"011110001",
  10690=>"000001011",
  10691=>"001010110",
  10692=>"110011011",
  10693=>"011000100",
  10694=>"010010101",
  10695=>"010010100",
  10696=>"001001011",
  10697=>"000011011",
  10698=>"110100000",
  10699=>"100111011",
  10700=>"010111000",
  10701=>"111111101",
  10702=>"010001001",
  10703=>"010110010",
  10704=>"110110100",
  10705=>"011011111",
  10706=>"001101100",
  10707=>"001011110",
  10708=>"011001010",
  10709=>"101100100",
  10710=>"000001001",
  10711=>"101100100",
  10712=>"011000011",
  10713=>"011101010",
  10714=>"111101001",
  10715=>"000010000",
  10716=>"010001010",
  10717=>"000011110",
  10718=>"111011110",
  10719=>"110010000",
  10720=>"000110110",
  10721=>"111111001",
  10722=>"110001111",
  10723=>"101100101",
  10724=>"011010100",
  10725=>"000010000",
  10726=>"010110111",
  10727=>"101101111",
  10728=>"100100000",
  10729=>"010101100",
  10730=>"111010110",
  10731=>"001010011",
  10732=>"111111000",
  10733=>"010011011",
  10734=>"000111111",
  10735=>"111001000",
  10736=>"100100011",
  10737=>"001101000",
  10738=>"111001001",
  10739=>"000101000",
  10740=>"101100001",
  10741=>"111100110",
  10742=>"011000001",
  10743=>"101100111",
  10744=>"111001101",
  10745=>"111010011",
  10746=>"000111100",
  10747=>"101000101",
  10748=>"101101011",
  10749=>"111001101",
  10750=>"110100110",
  10751=>"101100100",
  10752=>"011110110",
  10753=>"010110001",
  10754=>"000011011",
  10755=>"000001100",
  10756=>"010001110",
  10757=>"011000000",
  10758=>"100110110",
  10759=>"111010000",
  10760=>"100000111",
  10761=>"000111110",
  10762=>"010011010",
  10763=>"010111010",
  10764=>"110000010",
  10765=>"011001001",
  10766=>"100000100",
  10767=>"110111100",
  10768=>"011011100",
  10769=>"000000110",
  10770=>"111101011",
  10771=>"011010011",
  10772=>"011001111",
  10773=>"111000010",
  10774=>"001100100",
  10775=>"110110110",
  10776=>"001000110",
  10777=>"100101101",
  10778=>"110101000",
  10779=>"000101011",
  10780=>"101011111",
  10781=>"110101001",
  10782=>"001001110",
  10783=>"001011110",
  10784=>"000011000",
  10785=>"000101001",
  10786=>"011011000",
  10787=>"110100100",
  10788=>"110101010",
  10789=>"100111111",
  10790=>"011111111",
  10791=>"010000110",
  10792=>"000011010",
  10793=>"001011000",
  10794=>"100101101",
  10795=>"101001011",
  10796=>"100110111",
  10797=>"110100101",
  10798=>"011010100",
  10799=>"101010111",
  10800=>"111100111",
  10801=>"001111111",
  10802=>"101111101",
  10803=>"010101001",
  10804=>"101100011",
  10805=>"000110111",
  10806=>"110011111",
  10807=>"001101011",
  10808=>"001001101",
  10809=>"110100111",
  10810=>"101001011",
  10811=>"010101101",
  10812=>"000010101",
  10813=>"000100010",
  10814=>"011011111",
  10815=>"001011011",
  10816=>"000010111",
  10817=>"110100000",
  10818=>"111100110",
  10819=>"101010010",
  10820=>"011101001",
  10821=>"011011000",
  10822=>"111101110",
  10823=>"000001001",
  10824=>"001000010",
  10825=>"010000100",
  10826=>"000101110",
  10827=>"010000011",
  10828=>"101101100",
  10829=>"001101000",
  10830=>"001010111",
  10831=>"011000101",
  10832=>"001001010",
  10833=>"001001010",
  10834=>"001001110",
  10835=>"100000000",
  10836=>"010001011",
  10837=>"110011110",
  10838=>"111110010",
  10839=>"010110001",
  10840=>"011001110",
  10841=>"000101000",
  10842=>"100100000",
  10843=>"001010101",
  10844=>"010001011",
  10845=>"000110100",
  10846=>"011001110",
  10847=>"000110101",
  10848=>"111111111",
  10849=>"110010101",
  10850=>"010101011",
  10851=>"110001101",
  10852=>"110010111",
  10853=>"110011110",
  10854=>"111101110",
  10855=>"000010100",
  10856=>"111111101",
  10857=>"110101100",
  10858=>"011000111",
  10859=>"101101110",
  10860=>"000101001",
  10861=>"011001011",
  10862=>"000111111",
  10863=>"011001101",
  10864=>"100000110",
  10865=>"011111011",
  10866=>"011110100",
  10867=>"000001011",
  10868=>"001010000",
  10869=>"011100000",
  10870=>"111000101",
  10871=>"000011100",
  10872=>"001001001",
  10873=>"101001001",
  10874=>"011110011",
  10875=>"111010110",
  10876=>"011000010",
  10877=>"110011011",
  10878=>"011101100",
  10879=>"100010111",
  10880=>"100010101",
  10881=>"001000000",
  10882=>"101110101",
  10883=>"001101001",
  10884=>"001001110",
  10885=>"001001010",
  10886=>"011011111",
  10887=>"101010010",
  10888=>"111011101",
  10889=>"011000000",
  10890=>"100110101",
  10891=>"111000100",
  10892=>"000011101",
  10893=>"100000000",
  10894=>"011010010",
  10895=>"111101000",
  10896=>"010011010",
  10897=>"110000111",
  10898=>"101010110",
  10899=>"010111110",
  10900=>"101111000",
  10901=>"011011100",
  10902=>"110101001",
  10903=>"111011001",
  10904=>"011011111",
  10905=>"101000011",
  10906=>"011111000",
  10907=>"011111110",
  10908=>"011100100",
  10909=>"000110110",
  10910=>"100100001",
  10911=>"111100100",
  10912=>"011110010",
  10913=>"011111001",
  10914=>"010100000",
  10915=>"001101110",
  10916=>"011100110",
  10917=>"100001000",
  10918=>"000110011",
  10919=>"101011100",
  10920=>"101110000",
  10921=>"100011110",
  10922=>"000001111",
  10923=>"100100111",
  10924=>"111010100",
  10925=>"010100101",
  10926=>"100100100",
  10927=>"010010010",
  10928=>"001111001",
  10929=>"110001101",
  10930=>"001101001",
  10931=>"001110011",
  10932=>"011100001",
  10933=>"111111100",
  10934=>"010111010",
  10935=>"001100000",
  10936=>"001101111",
  10937=>"100111111",
  10938=>"000011000",
  10939=>"100001001",
  10940=>"111100111",
  10941=>"101111000",
  10942=>"101011000",
  10943=>"000011110",
  10944=>"100011000",
  10945=>"110011111",
  10946=>"101101001",
  10947=>"000001111",
  10948=>"011110001",
  10949=>"110010111",
  10950=>"111101000",
  10951=>"111011001",
  10952=>"101010100",
  10953=>"001001011",
  10954=>"001111000",
  10955=>"001101111",
  10956=>"011101101",
  10957=>"001011111",
  10958=>"011110010",
  10959=>"001110111",
  10960=>"111000011",
  10961=>"010001111",
  10962=>"011100010",
  10963=>"001000111",
  10964=>"100101000",
  10965=>"001101011",
  10966=>"000111001",
  10967=>"111011101",
  10968=>"000110101",
  10969=>"011101111",
  10970=>"101011000",
  10971=>"101010110",
  10972=>"001001100",
  10973=>"111111011",
  10974=>"101011101",
  10975=>"010101101",
  10976=>"000010001",
  10977=>"111101011",
  10978=>"001111111",
  10979=>"100000100",
  10980=>"001010111",
  10981=>"111010010",
  10982=>"111101101",
  10983=>"000001100",
  10984=>"101000000",
  10985=>"111111001",
  10986=>"000000001",
  10987=>"011110010",
  10988=>"001111100",
  10989=>"010111111",
  10990=>"000111111",
  10991=>"111001000",
  10992=>"111110010",
  10993=>"101001000",
  10994=>"110010111",
  10995=>"011100100",
  10996=>"100111100",
  10997=>"000111101",
  10998=>"110000111",
  10999=>"001101110",
  11000=>"111010101",
  11001=>"101001101",
  11002=>"101111001",
  11003=>"101000111",
  11004=>"100100101",
  11005=>"011010111",
  11006=>"001011000",
  11007=>"010001001",
  11008=>"101001010",
  11009=>"000110100",
  11010=>"100101000",
  11011=>"111101110",
  11012=>"011011101",
  11013=>"111101110",
  11014=>"010100000",
  11015=>"111111000",
  11016=>"001101110",
  11017=>"011100110",
  11018=>"000001010",
  11019=>"000011110",
  11020=>"001001001",
  11021=>"000101111",
  11022=>"001100011",
  11023=>"000011000",
  11024=>"100110100",
  11025=>"000000100",
  11026=>"111110100",
  11027=>"100101110",
  11028=>"001101100",
  11029=>"101011010",
  11030=>"100101111",
  11031=>"110111101",
  11032=>"010000110",
  11033=>"000011101",
  11034=>"000010110",
  11035=>"100000101",
  11036=>"111100001",
  11037=>"000110110",
  11038=>"101110010",
  11039=>"000000010",
  11040=>"011011110",
  11041=>"100000011",
  11042=>"001110000",
  11043=>"000011001",
  11044=>"011111110",
  11045=>"111101100",
  11046=>"000011001",
  11047=>"110111000",
  11048=>"011001000",
  11049=>"000101010",
  11050=>"101110100",
  11051=>"110111111",
  11052=>"110110011",
  11053=>"110111011",
  11054=>"101111111",
  11055=>"101001001",
  11056=>"100001110",
  11057=>"010101101",
  11058=>"000011100",
  11059=>"000010001",
  11060=>"110101010",
  11061=>"011111010",
  11062=>"010001001",
  11063=>"101011011",
  11064=>"001100000",
  11065=>"010111001",
  11066=>"000100110",
  11067=>"010000101",
  11068=>"100111001",
  11069=>"101100101",
  11070=>"000000100",
  11071=>"001100000",
  11072=>"001110111",
  11073=>"010001010",
  11074=>"111100100",
  11075=>"000001001",
  11076=>"000000100",
  11077=>"010000000",
  11078=>"110110001",
  11079=>"101101010",
  11080=>"011110011",
  11081=>"001011101",
  11082=>"011110101",
  11083=>"001010101",
  11084=>"011111101",
  11085=>"011110110",
  11086=>"100101010",
  11087=>"011011110",
  11088=>"001111111",
  11089=>"010010111",
  11090=>"110000010",
  11091=>"101010000",
  11092=>"100110100",
  11093=>"001011001",
  11094=>"101101100",
  11095=>"010100010",
  11096=>"010000000",
  11097=>"111100010",
  11098=>"101000001",
  11099=>"101111000",
  11100=>"110000101",
  11101=>"101000101",
  11102=>"010110000",
  11103=>"001000001",
  11104=>"100110011",
  11105=>"110111100",
  11106=>"011010010",
  11107=>"001101011",
  11108=>"111010001",
  11109=>"000101111",
  11110=>"101101110",
  11111=>"010101000",
  11112=>"110010011",
  11113=>"001010111",
  11114=>"100111010",
  11115=>"100110010",
  11116=>"101111100",
  11117=>"110101000",
  11118=>"001001101",
  11119=>"110101100",
  11120=>"111011101",
  11121=>"011010010",
  11122=>"001010110",
  11123=>"011100001",
  11124=>"110010001",
  11125=>"000101011",
  11126=>"010110010",
  11127=>"100110110",
  11128=>"010111011",
  11129=>"101000100",
  11130=>"111001111",
  11131=>"010010110",
  11132=>"001000111",
  11133=>"011001011",
  11134=>"001100001",
  11135=>"001001101",
  11136=>"100101000",
  11137=>"011110111",
  11138=>"100110010",
  11139=>"011011001",
  11140=>"010010010",
  11141=>"101000010",
  11142=>"000110011",
  11143=>"000001001",
  11144=>"110101101",
  11145=>"111000110",
  11146=>"111011010",
  11147=>"011000000",
  11148=>"001000000",
  11149=>"101110001",
  11150=>"001010111",
  11151=>"000110100",
  11152=>"001111001",
  11153=>"001110110",
  11154=>"010111100",
  11155=>"101001100",
  11156=>"001000111",
  11157=>"001101110",
  11158=>"010010111",
  11159=>"001111010",
  11160=>"111110010",
  11161=>"010101100",
  11162=>"111000011",
  11163=>"001100110",
  11164=>"101100001",
  11165=>"111000010",
  11166=>"000001111",
  11167=>"011001000",
  11168=>"100101000",
  11169=>"110010111",
  11170=>"011010100",
  11171=>"111110001",
  11172=>"010111001",
  11173=>"111000100",
  11174=>"100010010",
  11175=>"001110101",
  11176=>"001111010",
  11177=>"101101111",
  11178=>"010011100",
  11179=>"001011110",
  11180=>"100111001",
  11181=>"100101001",
  11182=>"100000100",
  11183=>"101011010",
  11184=>"111011101",
  11185=>"110011111",
  11186=>"010000000",
  11187=>"010111001",
  11188=>"110111100",
  11189=>"110010010",
  11190=>"101001010",
  11191=>"010111001",
  11192=>"010100101",
  11193=>"011011011",
  11194=>"101100101",
  11195=>"111011100",
  11196=>"101101110",
  11197=>"000010110",
  11198=>"111100101",
  11199=>"100110101",
  11200=>"111101011",
  11201=>"010111111",
  11202=>"101111110",
  11203=>"000000110",
  11204=>"000011010",
  11205=>"001100010",
  11206=>"111101111",
  11207=>"100011110",
  11208=>"001101000",
  11209=>"101101100",
  11210=>"011010110",
  11211=>"000110001",
  11212=>"001010011",
  11213=>"000001111",
  11214=>"100010011",
  11215=>"010000110",
  11216=>"001000000",
  11217=>"000101000",
  11218=>"010000111",
  11219=>"100010101",
  11220=>"000111111",
  11221=>"010000000",
  11222=>"011110011",
  11223=>"010000110",
  11224=>"011001101",
  11225=>"101001101",
  11226=>"111111101",
  11227=>"011010010",
  11228=>"111001001",
  11229=>"001010111",
  11230=>"110101001",
  11231=>"111100000",
  11232=>"011011011",
  11233=>"111000110",
  11234=>"111001100",
  11235=>"100010100",
  11236=>"010000110",
  11237=>"010100000",
  11238=>"110010011",
  11239=>"110001010",
  11240=>"110011001",
  11241=>"011111010",
  11242=>"110001010",
  11243=>"000011111",
  11244=>"100001111",
  11245=>"000101111",
  11246=>"110001010",
  11247=>"011101000",
  11248=>"110000111",
  11249=>"010110010",
  11250=>"000000000",
  11251=>"000100100",
  11252=>"110001000",
  11253=>"000010001",
  11254=>"110100111",
  11255=>"100010000",
  11256=>"011101001",
  11257=>"111000011",
  11258=>"110101110",
  11259=>"100001100",
  11260=>"100111110",
  11261=>"000101000",
  11262=>"110110001",
  11263=>"111101000",
  11264=>"010000011",
  11265=>"011101101",
  11266=>"001100001",
  11267=>"100000010",
  11268=>"100000001",
  11269=>"001101011",
  11270=>"011100001",
  11271=>"110000101",
  11272=>"111100010",
  11273=>"001011010",
  11274=>"001100111",
  11275=>"101010011",
  11276=>"011111111",
  11277=>"010101111",
  11278=>"010000110",
  11279=>"011101010",
  11280=>"000100100",
  11281=>"000001000",
  11282=>"101011100",
  11283=>"011111110",
  11284=>"001111100",
  11285=>"101100101",
  11286=>"110101111",
  11287=>"110101011",
  11288=>"000011111",
  11289=>"000110010",
  11290=>"100111101",
  11291=>"010111011",
  11292=>"111111011",
  11293=>"011011010",
  11294=>"011111110",
  11295=>"110110010",
  11296=>"011011101",
  11297=>"011100110",
  11298=>"101001001",
  11299=>"011100100",
  11300=>"010000110",
  11301=>"101110001",
  11302=>"001111000",
  11303=>"101111001",
  11304=>"100110000",
  11305=>"110001000",
  11306=>"100001000",
  11307=>"111000011",
  11308=>"100010100",
  11309=>"000101100",
  11310=>"100001101",
  11311=>"100111101",
  11312=>"011101111",
  11313=>"110111111",
  11314=>"110100000",
  11315=>"000100111",
  11316=>"000000111",
  11317=>"000000111",
  11318=>"100010110",
  11319=>"011100011",
  11320=>"000111100",
  11321=>"010000010",
  11322=>"110110100",
  11323=>"100100000",
  11324=>"001010001",
  11325=>"011000101",
  11326=>"101011110",
  11327=>"000110000",
  11328=>"111111001",
  11329=>"111011101",
  11330=>"011110011",
  11331=>"111111011",
  11332=>"001111100",
  11333=>"000010110",
  11334=>"111111000",
  11335=>"000110110",
  11336=>"100110010",
  11337=>"000001010",
  11338=>"001111100",
  11339=>"111011101",
  11340=>"000011101",
  11341=>"111001110",
  11342=>"000100001",
  11343=>"011010000",
  11344=>"111101011",
  11345=>"000011001",
  11346=>"111011000",
  11347=>"111010101",
  11348=>"110111000",
  11349=>"100000000",
  11350=>"111001010",
  11351=>"101000100",
  11352=>"100011000",
  11353=>"011100111",
  11354=>"001110010",
  11355=>"110000100",
  11356=>"110100010",
  11357=>"100110011",
  11358=>"011010001",
  11359=>"100011011",
  11360=>"101100101",
  11361=>"100010000",
  11362=>"000000000",
  11363=>"000000111",
  11364=>"111110001",
  11365=>"001010111",
  11366=>"111011011",
  11367=>"100110001",
  11368=>"001101110",
  11369=>"010111111",
  11370=>"010110000",
  11371=>"001101000",
  11372=>"110010010",
  11373=>"001101101",
  11374=>"100001110",
  11375=>"110101101",
  11376=>"100101100",
  11377=>"010000100",
  11378=>"001111110",
  11379=>"100011110",
  11380=>"101101111",
  11381=>"110001100",
  11382=>"101101111",
  11383=>"000110001",
  11384=>"101100010",
  11385=>"101110010",
  11386=>"001111011",
  11387=>"000000001",
  11388=>"000111000",
  11389=>"001010000",
  11390=>"110110101",
  11391=>"100101100",
  11392=>"001111100",
  11393=>"101000011",
  11394=>"001000010",
  11395=>"011000101",
  11396=>"010111011",
  11397=>"100111110",
  11398=>"101001110",
  11399=>"100001100",
  11400=>"000101010",
  11401=>"100110101",
  11402=>"110110100",
  11403=>"100000101",
  11404=>"000100100",
  11405=>"000110111",
  11406=>"010100110",
  11407=>"001111100",
  11408=>"010010110",
  11409=>"110101100",
  11410=>"101101010",
  11411=>"100000110",
  11412=>"101000010",
  11413=>"001001111",
  11414=>"011110011",
  11415=>"000000001",
  11416=>"110110101",
  11417=>"110100000",
  11418=>"001110000",
  11419=>"111001101",
  11420=>"101011000",
  11421=>"010001001",
  11422=>"001111001",
  11423=>"110111000",
  11424=>"101011011",
  11425=>"001110100",
  11426=>"111110101",
  11427=>"001000001",
  11428=>"111101100",
  11429=>"111000111",
  11430=>"101110101",
  11431=>"100100010",
  11432=>"000001001",
  11433=>"011100101",
  11434=>"011110100",
  11435=>"110111101",
  11436=>"000001001",
  11437=>"001001011",
  11438=>"011110101",
  11439=>"001111110",
  11440=>"110000000",
  11441=>"011110100",
  11442=>"000100101",
  11443=>"100010000",
  11444=>"111000111",
  11445=>"000010111",
  11446=>"011001101",
  11447=>"110011000",
  11448=>"001000100",
  11449=>"011101101",
  11450=>"010000011",
  11451=>"001101000",
  11452=>"100100100",
  11453=>"111101000",
  11454=>"011011100",
  11455=>"111010100",
  11456=>"110011010",
  11457=>"111110101",
  11458=>"100010101",
  11459=>"110011101",
  11460=>"100100011",
  11461=>"110100101",
  11462=>"100001001",
  11463=>"011110000",
  11464=>"001010001",
  11465=>"011101111",
  11466=>"010100001",
  11467=>"110111101",
  11468=>"101011001",
  11469=>"111100010",
  11470=>"000011000",
  11471=>"110010011",
  11472=>"100001011",
  11473=>"101010110",
  11474=>"101011100",
  11475=>"100100010",
  11476=>"100110110",
  11477=>"011000101",
  11478=>"000111011",
  11479=>"111111011",
  11480=>"110111111",
  11481=>"110110100",
  11482=>"111011011",
  11483=>"101110110",
  11484=>"100101110",
  11485=>"100111101",
  11486=>"100001011",
  11487=>"000000100",
  11488=>"100111011",
  11489=>"100000010",
  11490=>"111000000",
  11491=>"111001011",
  11492=>"001110000",
  11493=>"110101000",
  11494=>"110110010",
  11495=>"000010100",
  11496=>"110001011",
  11497=>"000001110",
  11498=>"010001000",
  11499=>"100101001",
  11500=>"011100010",
  11501=>"110011111",
  11502=>"101100000",
  11503=>"001001001",
  11504=>"000001010",
  11505=>"010101101",
  11506=>"001010010",
  11507=>"111011100",
  11508=>"111101011",
  11509=>"111110001",
  11510=>"111000110",
  11511=>"100110100",
  11512=>"010100100",
  11513=>"110000101",
  11514=>"010010000",
  11515=>"101011010",
  11516=>"100000100",
  11517=>"001001000",
  11518=>"111110011",
  11519=>"001110010",
  11520=>"011110111",
  11521=>"111101111",
  11522=>"110011001",
  11523=>"010001110",
  11524=>"110100101",
  11525=>"010000011",
  11526=>"010111000",
  11527=>"101001001",
  11528=>"111001100",
  11529=>"011001001",
  11530=>"001001000",
  11531=>"010100101",
  11532=>"000111010",
  11533=>"100100011",
  11534=>"001001100",
  11535=>"001100010",
  11536=>"001001010",
  11537=>"100100010",
  11538=>"101010111",
  11539=>"011111010",
  11540=>"100100111",
  11541=>"010110010",
  11542=>"010000011",
  11543=>"001001101",
  11544=>"110000110",
  11545=>"000010000",
  11546=>"000000010",
  11547=>"101111001",
  11548=>"001101110",
  11549=>"111001010",
  11550=>"011110010",
  11551=>"000100001",
  11552=>"001101001",
  11553=>"001111111",
  11554=>"110111010",
  11555=>"101000101",
  11556=>"011010000",
  11557=>"101111100",
  11558=>"111100000",
  11559=>"101010100",
  11560=>"101101010",
  11561=>"101010000",
  11562=>"011100111",
  11563=>"100100110",
  11564=>"111110111",
  11565=>"010001010",
  11566=>"001000000",
  11567=>"110000000",
  11568=>"101101111",
  11569=>"000111101",
  11570=>"010111000",
  11571=>"011001010",
  11572=>"101000111",
  11573=>"000011101",
  11574=>"100011100",
  11575=>"000000001",
  11576=>"111000111",
  11577=>"010011011",
  11578=>"001011111",
  11579=>"100000110",
  11580=>"110000101",
  11581=>"010010011",
  11582=>"001011101",
  11583=>"111011101",
  11584=>"100010011",
  11585=>"011101011",
  11586=>"111101010",
  11587=>"101111110",
  11588=>"101111000",
  11589=>"011110001",
  11590=>"000011100",
  11591=>"010110100",
  11592=>"111101111",
  11593=>"000100000",
  11594=>"101011111",
  11595=>"000000000",
  11596=>"111110110",
  11597=>"111011001",
  11598=>"110001000",
  11599=>"110100110",
  11600=>"101101001",
  11601=>"000001001",
  11602=>"110111011",
  11603=>"111110100",
  11604=>"111100100",
  11605=>"101001101",
  11606=>"001000100",
  11607=>"001111111",
  11608=>"000110101",
  11609=>"001010000",
  11610=>"011101101",
  11611=>"010001011",
  11612=>"111011001",
  11613=>"000000100",
  11614=>"101001111",
  11615=>"001110001",
  11616=>"010110000",
  11617=>"010000110",
  11618=>"101111011",
  11619=>"001000000",
  11620=>"000110111",
  11621=>"000110000",
  11622=>"000101110",
  11623=>"110101110",
  11624=>"011100110",
  11625=>"000100011",
  11626=>"101110100",
  11627=>"011010001",
  11628=>"101111000",
  11629=>"100111011",
  11630=>"100011101",
  11631=>"000100101",
  11632=>"010110100",
  11633=>"010101110",
  11634=>"010011010",
  11635=>"100101111",
  11636=>"010110001",
  11637=>"111000111",
  11638=>"111111100",
  11639=>"100111110",
  11640=>"100000101",
  11641=>"110100001",
  11642=>"001010011",
  11643=>"011000111",
  11644=>"011011000",
  11645=>"010010010",
  11646=>"010111100",
  11647=>"110101110",
  11648=>"011011101",
  11649=>"000000011",
  11650=>"001001111",
  11651=>"001001110",
  11652=>"101011110",
  11653=>"001100011",
  11654=>"101101110",
  11655=>"011100011",
  11656=>"001001000",
  11657=>"011111000",
  11658=>"001110111",
  11659=>"110011001",
  11660=>"001001000",
  11661=>"110001101",
  11662=>"001001110",
  11663=>"000101101",
  11664=>"110100110",
  11665=>"010001000",
  11666=>"010110111",
  11667=>"001010101",
  11668=>"110100011",
  11669=>"001000110",
  11670=>"110001100",
  11671=>"111111000",
  11672=>"011100010",
  11673=>"000001001",
  11674=>"010010110",
  11675=>"011010010",
  11676=>"000100000",
  11677=>"011011000",
  11678=>"101100110",
  11679=>"001110110",
  11680=>"011011100",
  11681=>"001010010",
  11682=>"110010001",
  11683=>"000010010",
  11684=>"110011000",
  11685=>"000101101",
  11686=>"100010110",
  11687=>"111000010",
  11688=>"010011001",
  11689=>"011110001",
  11690=>"100100100",
  11691=>"001010111",
  11692=>"001111011",
  11693=>"011001011",
  11694=>"110010100",
  11695=>"011010001",
  11696=>"100101100",
  11697=>"011111010",
  11698=>"111111111",
  11699=>"000100000",
  11700=>"000000000",
  11701=>"110010110",
  11702=>"011011010",
  11703=>"100101011",
  11704=>"010000110",
  11705=>"111010100",
  11706=>"100010010",
  11707=>"001001110",
  11708=>"110001011",
  11709=>"101100100",
  11710=>"011000000",
  11711=>"101101101",
  11712=>"100111111",
  11713=>"110110101",
  11714=>"000100000",
  11715=>"000011100",
  11716=>"010111111",
  11717=>"001100100",
  11718=>"100001010",
  11719=>"111011000",
  11720=>"101000011",
  11721=>"111111010",
  11722=>"100011001",
  11723=>"000010110",
  11724=>"101010001",
  11725=>"010110110",
  11726=>"001001010",
  11727=>"000100111",
  11728=>"111111100",
  11729=>"010100001",
  11730=>"001010010",
  11731=>"101001111",
  11732=>"111101011",
  11733=>"110011101",
  11734=>"110001001",
  11735=>"101011011",
  11736=>"010000110",
  11737=>"000001001",
  11738=>"011001101",
  11739=>"110000101",
  11740=>"111100010",
  11741=>"101111101",
  11742=>"100011111",
  11743=>"100000011",
  11744=>"011110111",
  11745=>"101110111",
  11746=>"011100110",
  11747=>"110011011",
  11748=>"110110101",
  11749=>"111110010",
  11750=>"010101100",
  11751=>"110001000",
  11752=>"111001010",
  11753=>"001011011",
  11754=>"110000000",
  11755=>"011100111",
  11756=>"011011000",
  11757=>"111100100",
  11758=>"110010100",
  11759=>"011101100",
  11760=>"101110000",
  11761=>"001000000",
  11762=>"111001111",
  11763=>"101100000",
  11764=>"101111101",
  11765=>"011011111",
  11766=>"111000001",
  11767=>"000010110",
  11768=>"001000011",
  11769=>"011100101",
  11770=>"000100010",
  11771=>"111100000",
  11772=>"000001001",
  11773=>"000001100",
  11774=>"000001101",
  11775=>"110111110",
  11776=>"011000010",
  11777=>"011010001",
  11778=>"010011001",
  11779=>"111000111",
  11780=>"110100010",
  11781=>"110100001",
  11782=>"000100000",
  11783=>"011011101",
  11784=>"010001011",
  11785=>"001010100",
  11786=>"101010100",
  11787=>"000100110",
  11788=>"000111101",
  11789=>"011011111",
  11790=>"010011010",
  11791=>"010010110",
  11792=>"111111110",
  11793=>"110011101",
  11794=>"000100010",
  11795=>"101010111",
  11796=>"001110100",
  11797=>"111000100",
  11798=>"010111001",
  11799=>"110001010",
  11800=>"010100010",
  11801=>"001011101",
  11802=>"001101010",
  11803=>"110011110",
  11804=>"100011111",
  11805=>"101010001",
  11806=>"010011011",
  11807=>"011111110",
  11808=>"010000010",
  11809=>"101001000",
  11810=>"111000101",
  11811=>"011010011",
  11812=>"011111010",
  11813=>"100011110",
  11814=>"100011111",
  11815=>"011011100",
  11816=>"110111010",
  11817=>"010100111",
  11818=>"110111111",
  11819=>"111010011",
  11820=>"001001011",
  11821=>"111010011",
  11822=>"011101001",
  11823=>"111111100",
  11824=>"011101101",
  11825=>"111100111",
  11826=>"000000110",
  11827=>"000001010",
  11828=>"011111101",
  11829=>"111101101",
  11830=>"001001000",
  11831=>"111111010",
  11832=>"000100011",
  11833=>"010000101",
  11834=>"111001110",
  11835=>"100100010",
  11836=>"000010110",
  11837=>"110011010",
  11838=>"111001000",
  11839=>"100110001",
  11840=>"000000110",
  11841=>"111111100",
  11842=>"000111111",
  11843=>"011111111",
  11844=>"011001000",
  11845=>"110101101",
  11846=>"010100100",
  11847=>"010011100",
  11848=>"000110011",
  11849=>"111001101",
  11850=>"011101101",
  11851=>"001111101",
  11852=>"000101110",
  11853=>"110111011",
  11854=>"010100011",
  11855=>"001010111",
  11856=>"100110001",
  11857=>"011010010",
  11858=>"110011000",
  11859=>"010110010",
  11860=>"000000000",
  11861=>"111000000",
  11862=>"100011010",
  11863=>"110101001",
  11864=>"100011100",
  11865=>"101100000",
  11866=>"111101000",
  11867=>"010000000",
  11868=>"000011111",
  11869=>"011000011",
  11870=>"000001010",
  11871=>"100001011",
  11872=>"100001010",
  11873=>"010010010",
  11874=>"000000101",
  11875=>"110011111",
  11876=>"100110101",
  11877=>"011100100",
  11878=>"111101110",
  11879=>"101111111",
  11880=>"101111101",
  11881=>"100001010",
  11882=>"111111101",
  11883=>"011000101",
  11884=>"110010111",
  11885=>"010000111",
  11886=>"101010000",
  11887=>"000000011",
  11888=>"101001110",
  11889=>"100001011",
  11890=>"111101000",
  11891=>"010010001",
  11892=>"011110101",
  11893=>"100010011",
  11894=>"110010011",
  11895=>"110001000",
  11896=>"111001111",
  11897=>"011101100",
  11898=>"010000001",
  11899=>"101111010",
  11900=>"001011100",
  11901=>"001100101",
  11902=>"100101011",
  11903=>"001010111",
  11904=>"010100011",
  11905=>"110011100",
  11906=>"100100010",
  11907=>"111100011",
  11908=>"110111010",
  11909=>"111010101",
  11910=>"011010100",
  11911=>"001101001",
  11912=>"111110111",
  11913=>"110111111",
  11914=>"111001101",
  11915=>"111111110",
  11916=>"000001000",
  11917=>"110000000",
  11918=>"101001001",
  11919=>"000110110",
  11920=>"100101011",
  11921=>"010010100",
  11922=>"101110010",
  11923=>"001101001",
  11924=>"000000011",
  11925=>"110000100",
  11926=>"010001011",
  11927=>"001101000",
  11928=>"110101111",
  11929=>"000101111",
  11930=>"011111110",
  11931=>"000110100",
  11932=>"001010001",
  11933=>"100000100",
  11934=>"101000110",
  11935=>"111011000",
  11936=>"011001110",
  11937=>"010110110",
  11938=>"110111001",
  11939=>"011010011",
  11940=>"011000001",
  11941=>"111111011",
  11942=>"111110000",
  11943=>"110011000",
  11944=>"110111000",
  11945=>"101000010",
  11946=>"101011111",
  11947=>"011001000",
  11948=>"001100010",
  11949=>"100010000",
  11950=>"011101110",
  11951=>"010101111",
  11952=>"100000000",
  11953=>"110110000",
  11954=>"001101101",
  11955=>"000101001",
  11956=>"010101001",
  11957=>"011010101",
  11958=>"010001100",
  11959=>"000010000",
  11960=>"000100111",
  11961=>"110010100",
  11962=>"011101101",
  11963=>"111010100",
  11964=>"110101011",
  11965=>"001111000",
  11966=>"100001001",
  11967=>"001101011",
  11968=>"110001010",
  11969=>"001010000",
  11970=>"011000110",
  11971=>"110010101",
  11972=>"010110110",
  11973=>"101011100",
  11974=>"001101110",
  11975=>"000101010",
  11976=>"111100001",
  11977=>"000100111",
  11978=>"111000110",
  11979=>"111000001",
  11980=>"111001100",
  11981=>"100011111",
  11982=>"011111001",
  11983=>"100010100",
  11984=>"100101111",
  11985=>"110001010",
  11986=>"001011011",
  11987=>"000100000",
  11988=>"000101110",
  11989=>"110010110",
  11990=>"100111110",
  11991=>"110010010",
  11992=>"100101111",
  11993=>"101001011",
  11994=>"100101001",
  11995=>"010111011",
  11996=>"000000100",
  11997=>"110001001",
  11998=>"000011111",
  11999=>"011000001",
  12000=>"011101111",
  12001=>"011110011",
  12002=>"100110011",
  12003=>"011101111",
  12004=>"000010011",
  12005=>"001101001",
  12006=>"001111111",
  12007=>"011000101",
  12008=>"101000011",
  12009=>"010111011",
  12010=>"000110000",
  12011=>"010001010",
  12012=>"011110000",
  12013=>"110011111",
  12014=>"011010110",
  12015=>"100011101",
  12016=>"010111101",
  12017=>"110001110",
  12018=>"100111111",
  12019=>"011100011",
  12020=>"101001100",
  12021=>"011110001",
  12022=>"101110110",
  12023=>"111111100",
  12024=>"010110010",
  12025=>"100101010",
  12026=>"000110111",
  12027=>"011101010",
  12028=>"100101111",
  12029=>"010100110",
  12030=>"100110000",
  12031=>"100011101",
  12032=>"000010100",
  12033=>"000111100",
  12034=>"111011101",
  12035=>"111010110",
  12036=>"000010110",
  12037=>"110000101",
  12038=>"101001111",
  12039=>"000011000",
  12040=>"000011100",
  12041=>"001010100",
  12042=>"111000011",
  12043=>"111011001",
  12044=>"000100000",
  12045=>"000100111",
  12046=>"111011111",
  12047=>"100100111",
  12048=>"101010111",
  12049=>"100010000",
  12050=>"001110000",
  12051=>"010111110",
  12052=>"100100010",
  12053=>"110111110",
  12054=>"111000111",
  12055=>"001000010",
  12056=>"101001100",
  12057=>"000001011",
  12058=>"111010001",
  12059=>"000000001",
  12060=>"000111110",
  12061=>"100001010",
  12062=>"001100110",
  12063=>"101000101",
  12064=>"011101110",
  12065=>"010100010",
  12066=>"110111101",
  12067=>"000000001",
  12068=>"100000000",
  12069=>"010101001",
  12070=>"000100011",
  12071=>"001101001",
  12072=>"011010001",
  12073=>"101001000",
  12074=>"010111101",
  12075=>"101010101",
  12076=>"010101100",
  12077=>"000111010",
  12078=>"111000010",
  12079=>"100110110",
  12080=>"010100001",
  12081=>"001110100",
  12082=>"001100011",
  12083=>"000001110",
  12084=>"100111100",
  12085=>"001010000",
  12086=>"000010010",
  12087=>"010011100",
  12088=>"001100111",
  12089=>"110001000",
  12090=>"100001010",
  12091=>"000110111",
  12092=>"100000000",
  12093=>"001001000",
  12094=>"010100100",
  12095=>"111010100",
  12096=>"010011011",
  12097=>"001001110",
  12098=>"100000011",
  12099=>"001001110",
  12100=>"010100100",
  12101=>"101100000",
  12102=>"101010011",
  12103=>"000110000",
  12104=>"100110100",
  12105=>"011011000",
  12106=>"001010111",
  12107=>"001101000",
  12108=>"011110000",
  12109=>"111101011",
  12110=>"000110110",
  12111=>"110100010",
  12112=>"111010100",
  12113=>"011100111",
  12114=>"000110111",
  12115=>"000000100",
  12116=>"101011000",
  12117=>"000011100",
  12118=>"000100011",
  12119=>"100000101",
  12120=>"010001110",
  12121=>"101011000",
  12122=>"101100101",
  12123=>"000100011",
  12124=>"111010111",
  12125=>"001010001",
  12126=>"000100001",
  12127=>"001101100",
  12128=>"000110100",
  12129=>"000111111",
  12130=>"011100101",
  12131=>"100101000",
  12132=>"000000111",
  12133=>"000010010",
  12134=>"101010011",
  12135=>"111100010",
  12136=>"010101111",
  12137=>"010101111",
  12138=>"111011011",
  12139=>"010101111",
  12140=>"110001110",
  12141=>"111011111",
  12142=>"001010010",
  12143=>"100101111",
  12144=>"101010101",
  12145=>"101100110",
  12146=>"111010010",
  12147=>"010101000",
  12148=>"100001010",
  12149=>"011111001",
  12150=>"101000101",
  12151=>"000000100",
  12152=>"001001010",
  12153=>"101001110",
  12154=>"100001011",
  12155=>"010011010",
  12156=>"111000100",
  12157=>"111110110",
  12158=>"111100100",
  12159=>"100000100",
  12160=>"011001000",
  12161=>"000001011",
  12162=>"110111010",
  12163=>"010111000",
  12164=>"010011100",
  12165=>"010001001",
  12166=>"001011111",
  12167=>"111010100",
  12168=>"011010010",
  12169=>"000000110",
  12170=>"011101000",
  12171=>"101000000",
  12172=>"100010111",
  12173=>"001010001",
  12174=>"110110110",
  12175=>"001001101",
  12176=>"111110001",
  12177=>"110000011",
  12178=>"001001100",
  12179=>"100001111",
  12180=>"100110111",
  12181=>"100111001",
  12182=>"000010000",
  12183=>"110010111",
  12184=>"111010100",
  12185=>"010110110",
  12186=>"000110110",
  12187=>"101111000",
  12188=>"111100010",
  12189=>"010100010",
  12190=>"000100010",
  12191=>"011101011",
  12192=>"010000101",
  12193=>"000010001",
  12194=>"111011000",
  12195=>"111101001",
  12196=>"100000001",
  12197=>"100111011",
  12198=>"100101011",
  12199=>"011011111",
  12200=>"110110100",
  12201=>"101100110",
  12202=>"111101000",
  12203=>"111001100",
  12204=>"011101011",
  12205=>"011101110",
  12206=>"111101110",
  12207=>"110001110",
  12208=>"101011101",
  12209=>"000111110",
  12210=>"000001000",
  12211=>"101010001",
  12212=>"101000000",
  12213=>"011110111",
  12214=>"001001001",
  12215=>"001011110",
  12216=>"000000110",
  12217=>"101000110",
  12218=>"111111101",
  12219=>"011011100",
  12220=>"100100100",
  12221=>"001000110",
  12222=>"101110000",
  12223=>"010010010",
  12224=>"011110101",
  12225=>"000001110",
  12226=>"110000110",
  12227=>"111001000",
  12228=>"001110110",
  12229=>"011101110",
  12230=>"001010111",
  12231=>"110011111",
  12232=>"001010001",
  12233=>"110110011",
  12234=>"110101101",
  12235=>"100001111",
  12236=>"110100111",
  12237=>"001100010",
  12238=>"011101000",
  12239=>"111011001",
  12240=>"100100000",
  12241=>"101000101",
  12242=>"110100011",
  12243=>"000101010",
  12244=>"000100100",
  12245=>"001100011",
  12246=>"001000100",
  12247=>"110000010",
  12248=>"111001011",
  12249=>"111111110",
  12250=>"000011101",
  12251=>"000001110",
  12252=>"101001010",
  12253=>"000001000",
  12254=>"111111000",
  12255=>"000110101",
  12256=>"000100110",
  12257=>"111010100",
  12258=>"000110111",
  12259=>"000010101",
  12260=>"101110110",
  12261=>"011100101",
  12262=>"000001001",
  12263=>"100111011",
  12264=>"110010001",
  12265=>"000000110",
  12266=>"101111100",
  12267=>"010110011",
  12268=>"111101110",
  12269=>"000101000",
  12270=>"010101000",
  12271=>"001011100",
  12272=>"111010011",
  12273=>"111111011",
  12274=>"011110001",
  12275=>"000011111",
  12276=>"000101010",
  12277=>"001111110",
  12278=>"101111111",
  12279=>"000100001",
  12280=>"010010010",
  12281=>"101000111",
  12282=>"000011110",
  12283=>"101100110",
  12284=>"010011011",
  12285=>"101000101",
  12286=>"011001000",
  12287=>"101011000",
  12288=>"111100010",
  12289=>"111111000",
  12290=>"000011000",
  12291=>"101000111",
  12292=>"000111000",
  12293=>"111100010",
  12294=>"110010110",
  12295=>"110111101",
  12296=>"110101100",
  12297=>"111100101",
  12298=>"000100001",
  12299=>"101011011",
  12300=>"011000000",
  12301=>"001000100",
  12302=>"101011101",
  12303=>"001100110",
  12304=>"111101010",
  12305=>"001101011",
  12306=>"011010101",
  12307=>"010010001",
  12308=>"011110001",
  12309=>"000111010",
  12310=>"111011101",
  12311=>"000011100",
  12312=>"110011111",
  12313=>"101110101",
  12314=>"110001000",
  12315=>"111111110",
  12316=>"000110010",
  12317=>"110100100",
  12318=>"010111011",
  12319=>"011001010",
  12320=>"110101011",
  12321=>"010011001",
  12322=>"111110001",
  12323=>"010111010",
  12324=>"111110101",
  12325=>"110010100",
  12326=>"010100000",
  12327=>"001000101",
  12328=>"011110101",
  12329=>"100100001",
  12330=>"111111010",
  12331=>"010010011",
  12332=>"111101000",
  12333=>"110011000",
  12334=>"111010000",
  12335=>"111000000",
  12336=>"111001000",
  12337=>"010100010",
  12338=>"100111110",
  12339=>"000010100",
  12340=>"111111010",
  12341=>"101111111",
  12342=>"011011101",
  12343=>"101010001",
  12344=>"100101010",
  12345=>"010000100",
  12346=>"101000100",
  12347=>"011000100",
  12348=>"010100110",
  12349=>"000111101",
  12350=>"111100001",
  12351=>"010101110",
  12352=>"011010001",
  12353=>"110001000",
  12354=>"110110010",
  12355=>"101000010",
  12356=>"000000010",
  12357=>"001000110",
  12358=>"011110101",
  12359=>"101111111",
  12360=>"110010110",
  12361=>"100010110",
  12362=>"000101000",
  12363=>"001100101",
  12364=>"011001110",
  12365=>"100100101",
  12366=>"101110000",
  12367=>"111010100",
  12368=>"001100110",
  12369=>"010100110",
  12370=>"101000110",
  12371=>"010101111",
  12372=>"111010100",
  12373=>"010111000",
  12374=>"011011011",
  12375=>"101110010",
  12376=>"011101011",
  12377=>"101101111",
  12378=>"010010010",
  12379=>"110101101",
  12380=>"001100011",
  12381=>"010100110",
  12382=>"111001001",
  12383=>"100110010",
  12384=>"000100010",
  12385=>"001001001",
  12386=>"101100100",
  12387=>"001010010",
  12388=>"011000010",
  12389=>"100101101",
  12390=>"011000010",
  12391=>"011101110",
  12392=>"100000010",
  12393=>"010110100",
  12394=>"010000010",
  12395=>"011000110",
  12396=>"101010010",
  12397=>"100110010",
  12398=>"100101110",
  12399=>"100000100",
  12400=>"111111011",
  12401=>"000111010",
  12402=>"011100100",
  12403=>"100111001",
  12404=>"011110011",
  12405=>"101111100",
  12406=>"100011100",
  12407=>"100001001",
  12408=>"001100011",
  12409=>"011010011",
  12410=>"111101000",
  12411=>"000000001",
  12412=>"001110110",
  12413=>"111011011",
  12414=>"001000100",
  12415=>"111010111",
  12416=>"000000011",
  12417=>"111001010",
  12418=>"111101000",
  12419=>"100001010",
  12420=>"011011100",
  12421=>"101110111",
  12422=>"100010011",
  12423=>"011111010",
  12424=>"110001101",
  12425=>"000010011",
  12426=>"100001111",
  12427=>"010110010",
  12428=>"111111000",
  12429=>"101010000",
  12430=>"000111011",
  12431=>"010011101",
  12432=>"111100100",
  12433=>"111001001",
  12434=>"011100001",
  12435=>"101001010",
  12436=>"011101000",
  12437=>"010010111",
  12438=>"101101110",
  12439=>"110111011",
  12440=>"011100001",
  12441=>"111011100",
  12442=>"111011111",
  12443=>"010010111",
  12444=>"111100000",
  12445=>"000001100",
  12446=>"111111001",
  12447=>"111010101",
  12448=>"000011101",
  12449=>"100011001",
  12450=>"111101000",
  12451=>"101010101",
  12452=>"110010011",
  12453=>"111110110",
  12454=>"010101010",
  12455=>"000010110",
  12456=>"101101011",
  12457=>"000101110",
  12458=>"011110101",
  12459=>"001111111",
  12460=>"101001111",
  12461=>"111110000",
  12462=>"001011111",
  12463=>"000110111",
  12464=>"000011011",
  12465=>"000100110",
  12466=>"001101001",
  12467=>"010001011",
  12468=>"101011110",
  12469=>"001111000",
  12470=>"001101001",
  12471=>"011001111",
  12472=>"110100111",
  12473=>"000101101",
  12474=>"000010101",
  12475=>"101011011",
  12476=>"101111110",
  12477=>"010001111",
  12478=>"111101101",
  12479=>"110111011",
  12480=>"001000101",
  12481=>"011000000",
  12482=>"100010101",
  12483=>"111101000",
  12484=>"000110101",
  12485=>"110000111",
  12486=>"010100110",
  12487=>"110100110",
  12488=>"110001111",
  12489=>"111100010",
  12490=>"010101001",
  12491=>"111101010",
  12492=>"110110000",
  12493=>"000101000",
  12494=>"110100100",
  12495=>"100111010",
  12496=>"111100100",
  12497=>"100001000",
  12498=>"010101000",
  12499=>"111011110",
  12500=>"111001001",
  12501=>"011001100",
  12502=>"111100110",
  12503=>"110101010",
  12504=>"101111100",
  12505=>"100010000",
  12506=>"000001010",
  12507=>"111010101",
  12508=>"011100011",
  12509=>"010101101",
  12510=>"101100001",
  12511=>"100001010",
  12512=>"011110010",
  12513=>"101001101",
  12514=>"110110111",
  12515=>"100100100",
  12516=>"001001100",
  12517=>"011000001",
  12518=>"111111010",
  12519=>"000001011",
  12520=>"100110011",
  12521=>"010010010",
  12522=>"010011100",
  12523=>"101000111",
  12524=>"110001001",
  12525=>"111110010",
  12526=>"001000011",
  12527=>"000000010",
  12528=>"011100011",
  12529=>"001100010",
  12530=>"110100101",
  12531=>"100000000",
  12532=>"010000011",
  12533=>"000111110",
  12534=>"010111110",
  12535=>"111000000",
  12536=>"111010001",
  12537=>"010010100",
  12538=>"000001111",
  12539=>"100010110",
  12540=>"000100100",
  12541=>"001110101",
  12542=>"110010010",
  12543=>"110010010",
  12544=>"110010101",
  12545=>"011101100",
  12546=>"001001000",
  12547=>"110011000",
  12548=>"101000011",
  12549=>"001100011",
  12550=>"110000001",
  12551=>"110000110",
  12552=>"111010001",
  12553=>"111001011",
  12554=>"010010010",
  12555=>"101101110",
  12556=>"001111000",
  12557=>"011111000",
  12558=>"010101010",
  12559=>"100001100",
  12560=>"000111111",
  12561=>"100100011",
  12562=>"100010010",
  12563=>"111100001",
  12564=>"010000101",
  12565=>"111000011",
  12566=>"111111001",
  12567=>"011001010",
  12568=>"000111100",
  12569=>"101101110",
  12570=>"001101110",
  12571=>"101100100",
  12572=>"110110000",
  12573=>"101111100",
  12574=>"001000010",
  12575=>"000000111",
  12576=>"001010110",
  12577=>"101010010",
  12578=>"000100001",
  12579=>"001101100",
  12580=>"000011100",
  12581=>"000010011",
  12582=>"011101000",
  12583=>"010100100",
  12584=>"000010100",
  12585=>"111100101",
  12586=>"101101111",
  12587=>"010001110",
  12588=>"110011101",
  12589=>"100010011",
  12590=>"001011101",
  12591=>"001100001",
  12592=>"010100110",
  12593=>"001100011",
  12594=>"110100110",
  12595=>"000001011",
  12596=>"101111011",
  12597=>"001110111",
  12598=>"011111011",
  12599=>"010111011",
  12600=>"100100000",
  12601=>"100001110",
  12602=>"011001110",
  12603=>"010010110",
  12604=>"101010011",
  12605=>"011000011",
  12606=>"000110100",
  12607=>"011111001",
  12608=>"101101011",
  12609=>"101101010",
  12610=>"111111010",
  12611=>"010011100",
  12612=>"001001110",
  12613=>"010101011",
  12614=>"100001000",
  12615=>"000001010",
  12616=>"001111101",
  12617=>"000000011",
  12618=>"000100011",
  12619=>"100001010",
  12620=>"100111010",
  12621=>"101000100",
  12622=>"000110001",
  12623=>"000001110",
  12624=>"010000001",
  12625=>"001100001",
  12626=>"100000110",
  12627=>"000111000",
  12628=>"110111111",
  12629=>"101110101",
  12630=>"001111100",
  12631=>"111110000",
  12632=>"100110001",
  12633=>"000000001",
  12634=>"110110001",
  12635=>"010000101",
  12636=>"100110111",
  12637=>"011111010",
  12638=>"011100111",
  12639=>"101100011",
  12640=>"111110111",
  12641=>"011110111",
  12642=>"100001001",
  12643=>"101100010",
  12644=>"111111010",
  12645=>"000000010",
  12646=>"011000110",
  12647=>"010001011",
  12648=>"110000000",
  12649=>"100110011",
  12650=>"111110000",
  12651=>"111001001",
  12652=>"110101000",
  12653=>"110001001",
  12654=>"001110011",
  12655=>"101101100",
  12656=>"100000011",
  12657=>"001000011",
  12658=>"101001110",
  12659=>"010110011",
  12660=>"001111101",
  12661=>"001111111",
  12662=>"000000010",
  12663=>"111100011",
  12664=>"011010111",
  12665=>"000010100",
  12666=>"001001111",
  12667=>"101100100",
  12668=>"110000110",
  12669=>"111101101",
  12670=>"101001011",
  12671=>"010101110",
  12672=>"011101101",
  12673=>"100010001",
  12674=>"100101100",
  12675=>"001110001",
  12676=>"001010001",
  12677=>"101001010",
  12678=>"110101100",
  12679=>"001011010",
  12680=>"100011010",
  12681=>"100101010",
  12682=>"000001001",
  12683=>"111001101",
  12684=>"001000100",
  12685=>"010010101",
  12686=>"101101011",
  12687=>"000010110",
  12688=>"001110100",
  12689=>"010001100",
  12690=>"110111010",
  12691=>"011001010",
  12692=>"110010101",
  12693=>"001100110",
  12694=>"100100000",
  12695=>"010011111",
  12696=>"011100110",
  12697=>"000001111",
  12698=>"100010001",
  12699=>"100101000",
  12700=>"111000100",
  12701=>"010111110",
  12702=>"011111011",
  12703=>"000001111",
  12704=>"010010100",
  12705=>"100000100",
  12706=>"000001001",
  12707=>"000000011",
  12708=>"110100011",
  12709=>"001011110",
  12710=>"001010010",
  12711=>"110100010",
  12712=>"010000000",
  12713=>"100011010",
  12714=>"000001011",
  12715=>"101000011",
  12716=>"111110101",
  12717=>"001000010",
  12718=>"100010001",
  12719=>"101000010",
  12720=>"010010010",
  12721=>"011010100",
  12722=>"000011001",
  12723=>"100000010",
  12724=>"110111101",
  12725=>"001111111",
  12726=>"101001000",
  12727=>"011100110",
  12728=>"111000101",
  12729=>"000110100",
  12730=>"000101010",
  12731=>"110001101",
  12732=>"010100100",
  12733=>"110010101",
  12734=>"011000000",
  12735=>"000000100",
  12736=>"010001111",
  12737=>"100001100",
  12738=>"111000000",
  12739=>"101100010",
  12740=>"101111101",
  12741=>"011110010",
  12742=>"111011110",
  12743=>"011011101",
  12744=>"100010001",
  12745=>"001101011",
  12746=>"000000000",
  12747=>"000010001",
  12748=>"001110111",
  12749=>"001001010",
  12750=>"101001111",
  12751=>"100011010",
  12752=>"100100010",
  12753=>"000000101",
  12754=>"111100100",
  12755=>"011101110",
  12756=>"100001110",
  12757=>"111101101",
  12758=>"010000001",
  12759=>"101001110",
  12760=>"011100001",
  12761=>"001001110",
  12762=>"011011010",
  12763=>"001010001",
  12764=>"000010011",
  12765=>"001001101",
  12766=>"100000111",
  12767=>"110000110",
  12768=>"100101111",
  12769=>"010010011",
  12770=>"110000100",
  12771=>"111110101",
  12772=>"001001110",
  12773=>"100000110",
  12774=>"101011110",
  12775=>"001011011",
  12776=>"111100111",
  12777=>"001111000",
  12778=>"010000000",
  12779=>"011000110",
  12780=>"011100011",
  12781=>"000011010",
  12782=>"001000011",
  12783=>"000100100",
  12784=>"110111110",
  12785=>"111010100",
  12786=>"001110001",
  12787=>"100001111",
  12788=>"111011011",
  12789=>"011011100",
  12790=>"011101001",
  12791=>"011011110",
  12792=>"111010111",
  12793=>"110111011",
  12794=>"001001100",
  12795=>"011100000",
  12796=>"101001001",
  12797=>"011111110",
  12798=>"011110001",
  12799=>"110110101",
  12800=>"000001100",
  12801=>"100111111",
  12802=>"100110000",
  12803=>"100011011",
  12804=>"000100101",
  12805=>"111111001",
  12806=>"110100011",
  12807=>"100100111",
  12808=>"010111111",
  12809=>"111011001",
  12810=>"101101011",
  12811=>"111000000",
  12812=>"000000101",
  12813=>"111011010",
  12814=>"011011001",
  12815=>"111100100",
  12816=>"100010111",
  12817=>"111101110",
  12818=>"110010100",
  12819=>"111010111",
  12820=>"010111010",
  12821=>"111000001",
  12822=>"000101101",
  12823=>"011000110",
  12824=>"100101110",
  12825=>"110100111",
  12826=>"001011001",
  12827=>"111010011",
  12828=>"011000100",
  12829=>"010101100",
  12830=>"010010101",
  12831=>"000010011",
  12832=>"011011010",
  12833=>"111010000",
  12834=>"000000000",
  12835=>"010001001",
  12836=>"011000111",
  12837=>"010010000",
  12838=>"111000010",
  12839=>"011110001",
  12840=>"010010001",
  12841=>"100101010",
  12842=>"101011101",
  12843=>"001111000",
  12844=>"111000011",
  12845=>"000000010",
  12846=>"111010011",
  12847=>"110101000",
  12848=>"011110101",
  12849=>"100011101",
  12850=>"110101010",
  12851=>"101110100",
  12852=>"010011111",
  12853=>"111010011",
  12854=>"111011110",
  12855=>"100111000",
  12856=>"110101000",
  12857=>"100001000",
  12858=>"010111111",
  12859=>"011110110",
  12860=>"000111101",
  12861=>"101001010",
  12862=>"111000101",
  12863=>"001111111",
  12864=>"101001000",
  12865=>"000011101",
  12866=>"000001110",
  12867=>"110001111",
  12868=>"101000000",
  12869=>"100000111",
  12870=>"001101100",
  12871=>"111000010",
  12872=>"011010111",
  12873=>"110101001",
  12874=>"100111101",
  12875=>"100111100",
  12876=>"100000110",
  12877=>"001010011",
  12878=>"110100000",
  12879=>"110011110",
  12880=>"110100110",
  12881=>"101100100",
  12882=>"011010011",
  12883=>"101000000",
  12884=>"011010000",
  12885=>"011010111",
  12886=>"000000100",
  12887=>"100000011",
  12888=>"011101000",
  12889=>"100110011",
  12890=>"000100000",
  12891=>"001100101",
  12892=>"010100011",
  12893=>"001010001",
  12894=>"100000110",
  12895=>"111110011",
  12896=>"000011110",
  12897=>"001100001",
  12898=>"100011101",
  12899=>"101010001",
  12900=>"100001001",
  12901=>"011001001",
  12902=>"000001110",
  12903=>"110110011",
  12904=>"010101101",
  12905=>"110011111",
  12906=>"010000101",
  12907=>"111110111",
  12908=>"011000110",
  12909=>"000101010",
  12910=>"010111001",
  12911=>"101110011",
  12912=>"100101000",
  12913=>"000001000",
  12914=>"001001100",
  12915=>"000101010",
  12916=>"100001111",
  12917=>"101010100",
  12918=>"111010010",
  12919=>"110110001",
  12920=>"010101000",
  12921=>"101010000",
  12922=>"001111110",
  12923=>"010110000",
  12924=>"001011001",
  12925=>"101010001",
  12926=>"101010110",
  12927=>"111000111",
  12928=>"100101100",
  12929=>"111111011",
  12930=>"100001000",
  12931=>"001001011",
  12932=>"110111000",
  12933=>"010000011",
  12934=>"010111001",
  12935=>"001110010",
  12936=>"100010011",
  12937=>"110100010",
  12938=>"000000100",
  12939=>"100111101",
  12940=>"100100111",
  12941=>"010001011",
  12942=>"111000001",
  12943=>"101100010",
  12944=>"110100001",
  12945=>"111100111",
  12946=>"100110111",
  12947=>"101011111",
  12948=>"110111010",
  12949=>"001101111",
  12950=>"010010000",
  12951=>"111111110",
  12952=>"110100100",
  12953=>"111101111",
  12954=>"011010000",
  12955=>"000110110",
  12956=>"010000111",
  12957=>"000001110",
  12958=>"101111101",
  12959=>"011110001",
  12960=>"101011011",
  12961=>"000100111",
  12962=>"001111011",
  12963=>"100110000",
  12964=>"101010110",
  12965=>"010111100",
  12966=>"110111100",
  12967=>"000001110",
  12968=>"100001001",
  12969=>"100000011",
  12970=>"011110111",
  12971=>"110010110",
  12972=>"001010110",
  12973=>"101000011",
  12974=>"111001011",
  12975=>"000101000",
  12976=>"000111111",
  12977=>"111110101",
  12978=>"100001111",
  12979=>"000010110",
  12980=>"001001001",
  12981=>"111001101",
  12982=>"101011111",
  12983=>"000010011",
  12984=>"001101101",
  12985=>"000010101",
  12986=>"111011100",
  12987=>"010001001",
  12988=>"110100101",
  12989=>"001011101",
  12990=>"111001011",
  12991=>"100000110",
  12992=>"110101101",
  12993=>"110111110",
  12994=>"100101111",
  12995=>"101101001",
  12996=>"010001001",
  12997=>"001010100",
  12998=>"101010010",
  12999=>"001011101",
  13000=>"111011000",
  13001=>"011111101",
  13002=>"110011111",
  13003=>"001010100",
  13004=>"011110101",
  13005=>"010111111",
  13006=>"000110010",
  13007=>"011000111",
  13008=>"010011010",
  13009=>"100000100",
  13010=>"010111001",
  13011=>"011010010",
  13012=>"001111100",
  13013=>"010001111",
  13014=>"101111100",
  13015=>"110110110",
  13016=>"111111101",
  13017=>"101110011",
  13018=>"100011011",
  13019=>"100111001",
  13020=>"101100010",
  13021=>"001001001",
  13022=>"000100011",
  13023=>"100111111",
  13024=>"000000110",
  13025=>"101100111",
  13026=>"000011100",
  13027=>"111010011",
  13028=>"110010101",
  13029=>"011111001",
  13030=>"101000110",
  13031=>"100110010",
  13032=>"111011111",
  13033=>"101000001",
  13034=>"101101011",
  13035=>"110001111",
  13036=>"000001001",
  13037=>"000000101",
  13038=>"101001010",
  13039=>"011000110",
  13040=>"111100110",
  13041=>"101011000",
  13042=>"010011010",
  13043=>"011100110",
  13044=>"111010110",
  13045=>"100101001",
  13046=>"111100100",
  13047=>"110000010",
  13048=>"011001101",
  13049=>"000100000",
  13050=>"010111000",
  13051=>"000111001",
  13052=>"001000000",
  13053=>"101100100",
  13054=>"101000001",
  13055=>"010100101",
  13056=>"011000011",
  13057=>"111010101",
  13058=>"110110010",
  13059=>"101010100",
  13060=>"000100101",
  13061=>"111010100",
  13062=>"111010111",
  13063=>"011011110",
  13064=>"000110101",
  13065=>"110111010",
  13066=>"111111100",
  13067=>"101100100",
  13068=>"010100010",
  13069=>"101011000",
  13070=>"101111111",
  13071=>"101101000",
  13072=>"100111110",
  13073=>"001110011",
  13074=>"000001001",
  13075=>"100001110",
  13076=>"000011000",
  13077=>"011110000",
  13078=>"100101101",
  13079=>"011111111",
  13080=>"000100101",
  13081=>"000010100",
  13082=>"010010101",
  13083=>"101011000",
  13084=>"100101111",
  13085=>"111000001",
  13086=>"011001010",
  13087=>"001110111",
  13088=>"000110110",
  13089=>"100110111",
  13090=>"011111001",
  13091=>"001101001",
  13092=>"100101111",
  13093=>"000101011",
  13094=>"010000101",
  13095=>"011001111",
  13096=>"111011111",
  13097=>"101101111",
  13098=>"010101100",
  13099=>"111101011",
  13100=>"100111000",
  13101=>"001000011",
  13102=>"010001010",
  13103=>"101000010",
  13104=>"100111111",
  13105=>"011001011",
  13106=>"101010100",
  13107=>"010001110",
  13108=>"001011111",
  13109=>"010010011",
  13110=>"010011111",
  13111=>"010111110",
  13112=>"011001111",
  13113=>"100010100",
  13114=>"011001010",
  13115=>"100000010",
  13116=>"000001011",
  13117=>"010100100",
  13118=>"111010010",
  13119=>"100001011",
  13120=>"011100001",
  13121=>"000011010",
  13122=>"000110110",
  13123=>"100000101",
  13124=>"001000011",
  13125=>"010001110",
  13126=>"100010011",
  13127=>"111100000",
  13128=>"011011001",
  13129=>"010011111",
  13130=>"101101010",
  13131=>"001111110",
  13132=>"001001110",
  13133=>"100100010",
  13134=>"011000101",
  13135=>"010101000",
  13136=>"001010010",
  13137=>"111011000",
  13138=>"010101010",
  13139=>"100101111",
  13140=>"010011011",
  13141=>"110011001",
  13142=>"111101000",
  13143=>"000001100",
  13144=>"111111111",
  13145=>"011011110",
  13146=>"010111011",
  13147=>"101110101",
  13148=>"000110111",
  13149=>"011011101",
  13150=>"010001101",
  13151=>"001000011",
  13152=>"000000010",
  13153=>"110011000",
  13154=>"100010010",
  13155=>"011100111",
  13156=>"110001001",
  13157=>"010110110",
  13158=>"011011011",
  13159=>"000100001",
  13160=>"010111010",
  13161=>"001010010",
  13162=>"000000000",
  13163=>"010111111",
  13164=>"111101010",
  13165=>"110100000",
  13166=>"000100111",
  13167=>"111101011",
  13168=>"101010110",
  13169=>"001010100",
  13170=>"100111110",
  13171=>"011010001",
  13172=>"000111010",
  13173=>"111001001",
  13174=>"000010011",
  13175=>"101010110",
  13176=>"110101000",
  13177=>"000011100",
  13178=>"100010000",
  13179=>"100111001",
  13180=>"001000010",
  13181=>"000111100",
  13182=>"001110100",
  13183=>"011011010",
  13184=>"000010111",
  13185=>"001110111",
  13186=>"000111100",
  13187=>"100000010",
  13188=>"000001010",
  13189=>"001010010",
  13190=>"100000000",
  13191=>"100110011",
  13192=>"100001001",
  13193=>"010111111",
  13194=>"101000110",
  13195=>"001101001",
  13196=>"111110011",
  13197=>"101101011",
  13198=>"011011111",
  13199=>"010011101",
  13200=>"110001111",
  13201=>"111111011",
  13202=>"001110010",
  13203=>"111000110",
  13204=>"010010100",
  13205=>"000110000",
  13206=>"000001010",
  13207=>"001101100",
  13208=>"101001000",
  13209=>"111010001",
  13210=>"100110111",
  13211=>"000010101",
  13212=>"111010001",
  13213=>"111000001",
  13214=>"000111111",
  13215=>"010100001",
  13216=>"000001000",
  13217=>"011011111",
  13218=>"011110101",
  13219=>"010101001",
  13220=>"000010001",
  13221=>"001100110",
  13222=>"100110110",
  13223=>"110010001",
  13224=>"010010000",
  13225=>"001010110",
  13226=>"101011001",
  13227=>"001011100",
  13228=>"101001011",
  13229=>"100101101",
  13230=>"011111111",
  13231=>"011101000",
  13232=>"001011111",
  13233=>"000101110",
  13234=>"000011101",
  13235=>"110111101",
  13236=>"010000001",
  13237=>"111000011",
  13238=>"010101011",
  13239=>"111001101",
  13240=>"011001111",
  13241=>"110111110",
  13242=>"110011001",
  13243=>"110001001",
  13244=>"010110111",
  13245=>"001111111",
  13246=>"000000110",
  13247=>"000000101",
  13248=>"110111111",
  13249=>"111000010",
  13250=>"101111011",
  13251=>"011000000",
  13252=>"111010011",
  13253=>"001001111",
  13254=>"001000001",
  13255=>"010110011",
  13256=>"111010010",
  13257=>"010000000",
  13258=>"111010101",
  13259=>"110100010",
  13260=>"100101110",
  13261=>"000010010",
  13262=>"001000111",
  13263=>"001001111",
  13264=>"011101111",
  13265=>"000011001",
  13266=>"111110110",
  13267=>"010000110",
  13268=>"100000001",
  13269=>"110111101",
  13270=>"101011011",
  13271=>"011010101",
  13272=>"101100110",
  13273=>"101001101",
  13274=>"011010000",
  13275=>"010111111",
  13276=>"001001110",
  13277=>"101000101",
  13278=>"001011100",
  13279=>"001100000",
  13280=>"000000010",
  13281=>"011000111",
  13282=>"100110101",
  13283=>"010111110",
  13284=>"011011101",
  13285=>"110100000",
  13286=>"100010110",
  13287=>"000110100",
  13288=>"010100000",
  13289=>"100011100",
  13290=>"101111100",
  13291=>"111011010",
  13292=>"100001101",
  13293=>"010110111",
  13294=>"001011101",
  13295=>"010101011",
  13296=>"110010111",
  13297=>"100000010",
  13298=>"100010110",
  13299=>"000010111",
  13300=>"101111000",
  13301=>"101000111",
  13302=>"011110001",
  13303=>"010011100",
  13304=>"011010110",
  13305=>"010001011",
  13306=>"001001000",
  13307=>"001111100",
  13308=>"000111011",
  13309=>"111011110",
  13310=>"111011110",
  13311=>"111110110",
  13312=>"100100000",
  13313=>"000011010",
  13314=>"011101000",
  13315=>"001010100",
  13316=>"111000010",
  13317=>"110100110",
  13318=>"111101111",
  13319=>"100001000",
  13320=>"101101000",
  13321=>"011101001",
  13322=>"010111110",
  13323=>"110111101",
  13324=>"111110101",
  13325=>"011001111",
  13326=>"000010110",
  13327=>"000100001",
  13328=>"110100100",
  13329=>"010100010",
  13330=>"100010010",
  13331=>"101000110",
  13332=>"111011101",
  13333=>"111010111",
  13334=>"100010100",
  13335=>"010111100",
  13336=>"011011011",
  13337=>"110000111",
  13338=>"010110111",
  13339=>"100001010",
  13340=>"100111100",
  13341=>"011010000",
  13342=>"101001100",
  13343=>"011011100",
  13344=>"011111000",
  13345=>"111100010",
  13346=>"001000011",
  13347=>"101010100",
  13348=>"000010000",
  13349=>"110010011",
  13350=>"011001000",
  13351=>"000111101",
  13352=>"010010010",
  13353=>"111101010",
  13354=>"010101010",
  13355=>"010011001",
  13356=>"111111001",
  13357=>"010010111",
  13358=>"100000000",
  13359=>"010100011",
  13360=>"101100100",
  13361=>"100010110",
  13362=>"001111111",
  13363=>"111111001",
  13364=>"111010001",
  13365=>"111111001",
  13366=>"111010011",
  13367=>"010010010",
  13368=>"000101111",
  13369=>"100100111",
  13370=>"111100001",
  13371=>"110110111",
  13372=>"101110110",
  13373=>"100101100",
  13374=>"011100010",
  13375=>"111111001",
  13376=>"010111111",
  13377=>"100100100",
  13378=>"100100111",
  13379=>"111001111",
  13380=>"111110111",
  13381=>"001010110",
  13382=>"111001011",
  13383=>"000110101",
  13384=>"010110100",
  13385=>"100101010",
  13386=>"101000100",
  13387=>"000100000",
  13388=>"011000100",
  13389=>"110010111",
  13390=>"010010111",
  13391=>"010000010",
  13392=>"111110011",
  13393=>"001010000",
  13394=>"010100010",
  13395=>"100101010",
  13396=>"101000100",
  13397=>"110100010",
  13398=>"010011000",
  13399=>"011010011",
  13400=>"110001100",
  13401=>"001110000",
  13402=>"011010001",
  13403=>"001100111",
  13404=>"100101101",
  13405=>"101110111",
  13406=>"111101000",
  13407=>"111110011",
  13408=>"101001001",
  13409=>"010100110",
  13410=>"100110010",
  13411=>"110011100",
  13412=>"101000101",
  13413=>"000101001",
  13414=>"110100000",
  13415=>"001000110",
  13416=>"101111001",
  13417=>"111100101",
  13418=>"100101110",
  13419=>"101001110",
  13420=>"101000011",
  13421=>"111000101",
  13422=>"010011010",
  13423=>"110010000",
  13424=>"111001001",
  13425=>"000101010",
  13426=>"000011001",
  13427=>"001110110",
  13428=>"011001000",
  13429=>"011111111",
  13430=>"100011100",
  13431=>"000000011",
  13432=>"111100110",
  13433=>"110000101",
  13434=>"000100011",
  13435=>"010110010",
  13436=>"111101100",
  13437=>"001011100",
  13438=>"010010110",
  13439=>"011110110",
  13440=>"111111110",
  13441=>"001100100",
  13442=>"001000110",
  13443=>"001000110",
  13444=>"001100011",
  13445=>"111011110",
  13446=>"011010000",
  13447=>"101111000",
  13448=>"101010001",
  13449=>"001000110",
  13450=>"101111101",
  13451=>"111010111",
  13452=>"010010111",
  13453=>"011101101",
  13454=>"100001100",
  13455=>"000101011",
  13456=>"000110100",
  13457=>"110000011",
  13458=>"001100100",
  13459=>"001010011",
  13460=>"110010000",
  13461=>"101010011",
  13462=>"100111100",
  13463=>"110111101",
  13464=>"111010001",
  13465=>"110001001",
  13466=>"111000010",
  13467=>"110011011",
  13468=>"101111111",
  13469=>"001011111",
  13470=>"111110101",
  13471=>"100010000",
  13472=>"110110010",
  13473=>"110100011",
  13474=>"011111011",
  13475=>"101111110",
  13476=>"000000110",
  13477=>"101100101",
  13478=>"101011011",
  13479=>"100100010",
  13480=>"000000111",
  13481=>"011101010",
  13482=>"111100101",
  13483=>"010111100",
  13484=>"111100111",
  13485=>"111100101",
  13486=>"100000111",
  13487=>"110000010",
  13488=>"111000100",
  13489=>"110111111",
  13490=>"100111110",
  13491=>"110100101",
  13492=>"101011001",
  13493=>"100101101",
  13494=>"000110010",
  13495=>"011011111",
  13496=>"100100111",
  13497=>"001001101",
  13498=>"001010111",
  13499=>"110011001",
  13500=>"100101011",
  13501=>"101100010",
  13502=>"111001110",
  13503=>"000100011",
  13504=>"100011011",
  13505=>"110100111",
  13506=>"010011011",
  13507=>"111001011",
  13508=>"000010100",
  13509=>"011110000",
  13510=>"111100010",
  13511=>"001101111",
  13512=>"111111111",
  13513=>"010011101",
  13514=>"110010011",
  13515=>"101000000",
  13516=>"111011100",
  13517=>"001100000",
  13518=>"111101111",
  13519=>"001111101",
  13520=>"011110100",
  13521=>"101011100",
  13522=>"100000010",
  13523=>"010110100",
  13524=>"111010101",
  13525=>"110001010",
  13526=>"101101010",
  13527=>"011101111",
  13528=>"101101001",
  13529=>"100110111",
  13530=>"010110111",
  13531=>"001001001",
  13532=>"011100001",
  13533=>"000111000",
  13534=>"000011111",
  13535=>"000000001",
  13536=>"111011010",
  13537=>"110001000",
  13538=>"000110011",
  13539=>"000011111",
  13540=>"010100111",
  13541=>"010100011",
  13542=>"001010100",
  13543=>"011101101",
  13544=>"011101100",
  13545=>"100110100",
  13546=>"000100101",
  13547=>"001101011",
  13548=>"111000001",
  13549=>"100000011",
  13550=>"101000000",
  13551=>"100101100",
  13552=>"110010110",
  13553=>"100111101",
  13554=>"101110000",
  13555=>"100111000",
  13556=>"110110001",
  13557=>"111011111",
  13558=>"111110100",
  13559=>"111101100",
  13560=>"000101111",
  13561=>"100010011",
  13562=>"110001101",
  13563=>"110100101",
  13564=>"110111101",
  13565=>"110101101",
  13566=>"101101100",
  13567=>"100011100",
  13568=>"000111000",
  13569=>"101111100",
  13570=>"111111001",
  13571=>"110000110",
  13572=>"100100100",
  13573=>"000110011",
  13574=>"011010111",
  13575=>"111101001",
  13576=>"111101111",
  13577=>"011110100",
  13578=>"100001010",
  13579=>"110101110",
  13580=>"011010010",
  13581=>"000101111",
  13582=>"111110001",
  13583=>"101011110",
  13584=>"010110101",
  13585=>"010001101",
  13586=>"000100101",
  13587=>"001101110",
  13588=>"010000100",
  13589=>"111001101",
  13590=>"110000011",
  13591=>"110110000",
  13592=>"010100010",
  13593=>"000010000",
  13594=>"011001100",
  13595=>"100110000",
  13596=>"110100000",
  13597=>"110111111",
  13598=>"000101110",
  13599=>"101011011",
  13600=>"100111110",
  13601=>"010011111",
  13602=>"001001011",
  13603=>"101111111",
  13604=>"011100110",
  13605=>"001000101",
  13606=>"111111001",
  13607=>"001000110",
  13608=>"011001011",
  13609=>"100010101",
  13610=>"111110000",
  13611=>"110010110",
  13612=>"101110001",
  13613=>"011110110",
  13614=>"100010010",
  13615=>"010101000",
  13616=>"101001110",
  13617=>"110100101",
  13618=>"011001011",
  13619=>"001100000",
  13620=>"110011110",
  13621=>"110000000",
  13622=>"101101110",
  13623=>"100010010",
  13624=>"111101011",
  13625=>"101001111",
  13626=>"111111010",
  13627=>"001110011",
  13628=>"100110011",
  13629=>"100110011",
  13630=>"101011001",
  13631=>"000010101",
  13632=>"001101111",
  13633=>"010011111",
  13634=>"010000100",
  13635=>"001000110",
  13636=>"110000101",
  13637=>"100110111",
  13638=>"010110010",
  13639=>"100110000",
  13640=>"000100010",
  13641=>"010111100",
  13642=>"010000100",
  13643=>"001000100",
  13644=>"001010011",
  13645=>"100010001",
  13646=>"001110111",
  13647=>"101110111",
  13648=>"110000010",
  13649=>"011100101",
  13650=>"011110011",
  13651=>"000010000",
  13652=>"010010110",
  13653=>"101000001",
  13654=>"000110000",
  13655=>"001011000",
  13656=>"011110011",
  13657=>"000011000",
  13658=>"111100001",
  13659=>"011101111",
  13660=>"110100101",
  13661=>"010110110",
  13662=>"001000010",
  13663=>"000101000",
  13664=>"000010011",
  13665=>"010110011",
  13666=>"011010111",
  13667=>"101100011",
  13668=>"001000001",
  13669=>"001010100",
  13670=>"000110110",
  13671=>"111011101",
  13672=>"111110000",
  13673=>"101001000",
  13674=>"100111111",
  13675=>"111010000",
  13676=>"111111011",
  13677=>"000101010",
  13678=>"111101101",
  13679=>"110000111",
  13680=>"001010010",
  13681=>"111110101",
  13682=>"110011011",
  13683=>"111100000",
  13684=>"101100001",
  13685=>"000111111",
  13686=>"110000010",
  13687=>"100111110",
  13688=>"101100100",
  13689=>"110011100",
  13690=>"111000000",
  13691=>"011110011",
  13692=>"101001000",
  13693=>"001000001",
  13694=>"111001110",
  13695=>"001100000",
  13696=>"111000111",
  13697=>"111010011",
  13698=>"001110100",
  13699=>"111010011",
  13700=>"100011110",
  13701=>"101001010",
  13702=>"011100011",
  13703=>"101111110",
  13704=>"010100101",
  13705=>"100011000",
  13706=>"110110111",
  13707=>"101100010",
  13708=>"101000100",
  13709=>"111110001",
  13710=>"101011111",
  13711=>"011000010",
  13712=>"001101001",
  13713=>"101011000",
  13714=>"111110011",
  13715=>"000111110",
  13716=>"100010101",
  13717=>"010110001",
  13718=>"111000110",
  13719=>"110110110",
  13720=>"101110111",
  13721=>"010001011",
  13722=>"001111100",
  13723=>"011010100",
  13724=>"000011010",
  13725=>"000011000",
  13726=>"100100110",
  13727=>"011011000",
  13728=>"000100111",
  13729=>"001111110",
  13730=>"100101011",
  13731=>"011110111",
  13732=>"111011011",
  13733=>"011101010",
  13734=>"000101111",
  13735=>"100111100",
  13736=>"001000010",
  13737=>"000100101",
  13738=>"110010000",
  13739=>"011000111",
  13740=>"010000011",
  13741=>"110000111",
  13742=>"010110100",
  13743=>"001101100",
  13744=>"100101100",
  13745=>"111010110",
  13746=>"111111111",
  13747=>"101111101",
  13748=>"111101111",
  13749=>"100011110",
  13750=>"011101101",
  13751=>"000011100",
  13752=>"111001011",
  13753=>"010111110",
  13754=>"111001000",
  13755=>"101010111",
  13756=>"101010110",
  13757=>"101000011",
  13758=>"011001110",
  13759=>"000001111",
  13760=>"100001110",
  13761=>"001100001",
  13762=>"101000100",
  13763=>"100111000",
  13764=>"110100111",
  13765=>"001000111",
  13766=>"101011111",
  13767=>"011111111",
  13768=>"010101110",
  13769=>"101011011",
  13770=>"100111000",
  13771=>"000110100",
  13772=>"111110001",
  13773=>"000101010",
  13774=>"001110111",
  13775=>"011001001",
  13776=>"001111001",
  13777=>"010111000",
  13778=>"100000011",
  13779=>"010111010",
  13780=>"001000000",
  13781=>"111000000",
  13782=>"111111111",
  13783=>"100111100",
  13784=>"101000100",
  13785=>"110010010",
  13786=>"101001111",
  13787=>"101101111",
  13788=>"001001000",
  13789=>"111100011",
  13790=>"010111111",
  13791=>"001111110",
  13792=>"011000011",
  13793=>"100101001",
  13794=>"101101001",
  13795=>"010011001",
  13796=>"110000101",
  13797=>"111000101",
  13798=>"111111111",
  13799=>"111101011",
  13800=>"101110000",
  13801=>"100010011",
  13802=>"111001010",
  13803=>"101010010",
  13804=>"001110001",
  13805=>"010011111",
  13806=>"011001011",
  13807=>"110110010",
  13808=>"110000000",
  13809=>"010011101",
  13810=>"110101111",
  13811=>"001010100",
  13812=>"111010010",
  13813=>"010110100",
  13814=>"100100110",
  13815=>"000011110",
  13816=>"110011001",
  13817=>"111101001",
  13818=>"001110110",
  13819=>"010111110",
  13820=>"101010000",
  13821=>"011010111",
  13822=>"100110101",
  13823=>"001111011",
  13824=>"000011111",
  13825=>"100010111",
  13826=>"101111101",
  13827=>"100001010",
  13828=>"010110110",
  13829=>"011110000",
  13830=>"010111000",
  13831=>"111010010",
  13832=>"110011011",
  13833=>"010110111",
  13834=>"100111101",
  13835=>"111110111",
  13836=>"010110011",
  13837=>"111101101",
  13838=>"110001100",
  13839=>"011000100",
  13840=>"001011001",
  13841=>"011001010",
  13842=>"111011111",
  13843=>"101001011",
  13844=>"101010011",
  13845=>"011010111",
  13846=>"001000101",
  13847=>"111001000",
  13848=>"111011100",
  13849=>"110101100",
  13850=>"101100110",
  13851=>"011111110",
  13852=>"110110010",
  13853=>"111100100",
  13854=>"101011110",
  13855=>"000011110",
  13856=>"110011010",
  13857=>"000100100",
  13858=>"101101111",
  13859=>"011101010",
  13860=>"011000100",
  13861=>"111100111",
  13862=>"101010111",
  13863=>"010111100",
  13864=>"110010010",
  13865=>"101110001",
  13866=>"000100110",
  13867=>"100100000",
  13868=>"011010000",
  13869=>"000011101",
  13870=>"111110000",
  13871=>"100000011",
  13872=>"000001110",
  13873=>"001011110",
  13874=>"110001000",
  13875=>"100000011",
  13876=>"010101001",
  13877=>"010011110",
  13878=>"101111000",
  13879=>"000011101",
  13880=>"000111011",
  13881=>"010101100",
  13882=>"100111011",
  13883=>"101100011",
  13884=>"001100011",
  13885=>"110100011",
  13886=>"111011111",
  13887=>"011111011",
  13888=>"010000000",
  13889=>"100001011",
  13890=>"011111111",
  13891=>"010000110",
  13892=>"101010010",
  13893=>"000101010",
  13894=>"001100011",
  13895=>"010100100",
  13896=>"110010010",
  13897=>"100001100",
  13898=>"001111011",
  13899=>"100011001",
  13900=>"001100100",
  13901=>"101101110",
  13902=>"111111011",
  13903=>"101000001",
  13904=>"000110000",
  13905=>"010010001",
  13906=>"100111111",
  13907=>"000110111",
  13908=>"111011100",
  13909=>"001001010",
  13910=>"100110001",
  13911=>"110011001",
  13912=>"101110010",
  13913=>"101100101",
  13914=>"101101110",
  13915=>"111110011",
  13916=>"010111001",
  13917=>"111011011",
  13918=>"000100011",
  13919=>"100000101",
  13920=>"001001110",
  13921=>"111010111",
  13922=>"100010001",
  13923=>"101000110",
  13924=>"001100000",
  13925=>"100011100",
  13926=>"111101110",
  13927=>"101010010",
  13928=>"101111101",
  13929=>"010110111",
  13930=>"001000010",
  13931=>"011001011",
  13932=>"010000000",
  13933=>"011110011",
  13934=>"110001110",
  13935=>"000101110",
  13936=>"110111101",
  13937=>"011111011",
  13938=>"100011011",
  13939=>"001010110",
  13940=>"110110000",
  13941=>"110010010",
  13942=>"111111001",
  13943=>"111111111",
  13944=>"111011000",
  13945=>"101010100",
  13946=>"111101000",
  13947=>"011110111",
  13948=>"000010101",
  13949=>"011010111",
  13950=>"000100011",
  13951=>"100111111",
  13952=>"110110000",
  13953=>"101001010",
  13954=>"100011100",
  13955=>"011111110",
  13956=>"110100101",
  13957=>"001011010",
  13958=>"101000100",
  13959=>"001110010",
  13960=>"100111001",
  13961=>"011110011",
  13962=>"001110001",
  13963=>"011000111",
  13964=>"000101111",
  13965=>"110001111",
  13966=>"100101110",
  13967=>"100100100",
  13968=>"011000111",
  13969=>"000001001",
  13970=>"011111110",
  13971=>"100000110",
  13972=>"011100000",
  13973=>"010000111",
  13974=>"000101000",
  13975=>"010001101",
  13976=>"110011111",
  13977=>"000100110",
  13978=>"000100111",
  13979=>"001101111",
  13980=>"100110000",
  13981=>"110110111",
  13982=>"000111111",
  13983=>"000100100",
  13984=>"011010010",
  13985=>"111110111",
  13986=>"101101110",
  13987=>"010111111",
  13988=>"100011101",
  13989=>"010010000",
  13990=>"011000100",
  13991=>"011101011",
  13992=>"101011010",
  13993=>"000100010",
  13994=>"011110010",
  13995=>"011101110",
  13996=>"001011110",
  13997=>"100001110",
  13998=>"101000101",
  13999=>"010101110",
  14000=>"111100100",
  14001=>"110110111",
  14002=>"000111000",
  14003=>"101010000",
  14004=>"000100011",
  14005=>"110111110",
  14006=>"011011001",
  14007=>"001010010",
  14008=>"110011101",
  14009=>"110100100",
  14010=>"010111100",
  14011=>"010001011",
  14012=>"111001111",
  14013=>"001000000",
  14014=>"001000011",
  14015=>"000010110",
  14016=>"001110111",
  14017=>"000111111",
  14018=>"100010111",
  14019=>"010000001",
  14020=>"011001000",
  14021=>"100110100",
  14022=>"101101011",
  14023=>"001111010",
  14024=>"001101111",
  14025=>"100100111",
  14026=>"000101100",
  14027=>"111111111",
  14028=>"000111010",
  14029=>"010010111",
  14030=>"001101001",
  14031=>"110100000",
  14032=>"000111111",
  14033=>"100101001",
  14034=>"001001111",
  14035=>"001101110",
  14036=>"000110110",
  14037=>"101001011",
  14038=>"111111001",
  14039=>"001111100",
  14040=>"100111111",
  14041=>"010110001",
  14042=>"110001010",
  14043=>"110001110",
  14044=>"101111101",
  14045=>"111111111",
  14046=>"101101000",
  14047=>"111011100",
  14048=>"101001010",
  14049=>"101001001",
  14050=>"000000011",
  14051=>"001011001",
  14052=>"001110000",
  14053=>"100100011",
  14054=>"011111111",
  14055=>"011011111",
  14056=>"110101100",
  14057=>"101001110",
  14058=>"101000000",
  14059=>"101100110",
  14060=>"111101110",
  14061=>"011110111",
  14062=>"100000110",
  14063=>"010110100",
  14064=>"110100010",
  14065=>"101000010",
  14066=>"111111010",
  14067=>"000000001",
  14068=>"111110111",
  14069=>"100000010",
  14070=>"001001111",
  14071=>"011011100",
  14072=>"100000011",
  14073=>"000000001",
  14074=>"001011010",
  14075=>"110101111",
  14076=>"000001111",
  14077=>"010011101",
  14078=>"100101010",
  14079=>"111100100",
  14080=>"111110100",
  14081=>"110001001",
  14082=>"100000101",
  14083=>"111010100",
  14084=>"000010100",
  14085=>"001000101",
  14086=>"101011100",
  14087=>"110000010",
  14088=>"000011101",
  14089=>"000100110",
  14090=>"100100000",
  14091=>"110001101",
  14092=>"001000011",
  14093=>"101101100",
  14094=>"110011011",
  14095=>"100010000",
  14096=>"110101111",
  14097=>"010000111",
  14098=>"010011001",
  14099=>"011000101",
  14100=>"010010100",
  14101=>"111011011",
  14102=>"101101010",
  14103=>"111110101",
  14104=>"111001000",
  14105=>"010010100",
  14106=>"110001010",
  14107=>"011010001",
  14108=>"101111100",
  14109=>"010100111",
  14110=>"011101000",
  14111=>"000111010",
  14112=>"110110000",
  14113=>"000001001",
  14114=>"010110111",
  14115=>"110101000",
  14116=>"001001100",
  14117=>"101101111",
  14118=>"111100001",
  14119=>"100111001",
  14120=>"010100110",
  14121=>"000101111",
  14122=>"011110100",
  14123=>"101010000",
  14124=>"000110100",
  14125=>"110011110",
  14126=>"111101000",
  14127=>"011101100",
  14128=>"011001001",
  14129=>"001100010",
  14130=>"111011010",
  14131=>"100010010",
  14132=>"101111011",
  14133=>"111110100",
  14134=>"101100001",
  14135=>"011110001",
  14136=>"111100111",
  14137=>"110000000",
  14138=>"100000011",
  14139=>"001001111",
  14140=>"000000011",
  14141=>"001000100",
  14142=>"111101101",
  14143=>"000100001",
  14144=>"101010010",
  14145=>"010111001",
  14146=>"110010110",
  14147=>"111001010",
  14148=>"100011011",
  14149=>"111111001",
  14150=>"000101000",
  14151=>"000110111",
  14152=>"110010011",
  14153=>"010100110",
  14154=>"101001101",
  14155=>"101111001",
  14156=>"000010010",
  14157=>"110100111",
  14158=>"100100111",
  14159=>"100100011",
  14160=>"010101100",
  14161=>"101000011",
  14162=>"110100101",
  14163=>"110010001",
  14164=>"101111101",
  14165=>"001000110",
  14166=>"000111000",
  14167=>"010001101",
  14168=>"111100010",
  14169=>"001001101",
  14170=>"011001010",
  14171=>"110110010",
  14172=>"111101010",
  14173=>"001101111",
  14174=>"010010101",
  14175=>"110111101",
  14176=>"110011010",
  14177=>"100110000",
  14178=>"010000001",
  14179=>"000011111",
  14180=>"010101111",
  14181=>"111001100",
  14182=>"101111111",
  14183=>"110011000",
  14184=>"101111111",
  14185=>"010111001",
  14186=>"011110100",
  14187=>"100001011",
  14188=>"100110111",
  14189=>"101001100",
  14190=>"100100000",
  14191=>"000011010",
  14192=>"101000100",
  14193=>"001000110",
  14194=>"000000010",
  14195=>"110011011",
  14196=>"111110100",
  14197=>"100100010",
  14198=>"111011100",
  14199=>"011110110",
  14200=>"100111111",
  14201=>"010010110",
  14202=>"100111001",
  14203=>"001010111",
  14204=>"100010010",
  14205=>"110100110",
  14206=>"101011000",
  14207=>"001010111",
  14208=>"101111111",
  14209=>"111101111",
  14210=>"111111100",
  14211=>"110101100",
  14212=>"011100111",
  14213=>"111101000",
  14214=>"010110001",
  14215=>"101000001",
  14216=>"110000110",
  14217=>"011110100",
  14218=>"111111011",
  14219=>"111001101",
  14220=>"100000100",
  14221=>"011010101",
  14222=>"100011111",
  14223=>"000000101",
  14224=>"000000100",
  14225=>"000110111",
  14226=>"111100000",
  14227=>"101000000",
  14228=>"101101111",
  14229=>"110110101",
  14230=>"100000011",
  14231=>"010000000",
  14232=>"010110011",
  14233=>"101101011",
  14234=>"011101000",
  14235=>"000001101",
  14236=>"100110011",
  14237=>"111101101",
  14238=>"000101110",
  14239=>"110001101",
  14240=>"110110000",
  14241=>"011101110",
  14242=>"110101111",
  14243=>"100011101",
  14244=>"100011101",
  14245=>"001110100",
  14246=>"101010001",
  14247=>"111100101",
  14248=>"110101000",
  14249=>"011101101",
  14250=>"011010010",
  14251=>"001101011",
  14252=>"000111001",
  14253=>"000010100",
  14254=>"011110111",
  14255=>"010000011",
  14256=>"100110010",
  14257=>"011010010",
  14258=>"000101001",
  14259=>"000001100",
  14260=>"000010011",
  14261=>"000011011",
  14262=>"110001110",
  14263=>"111110000",
  14264=>"001110000",
  14265=>"101111000",
  14266=>"100011111",
  14267=>"011010111",
  14268=>"000001100",
  14269=>"101000001",
  14270=>"000110010",
  14271=>"111110110",
  14272=>"011101011",
  14273=>"010011100",
  14274=>"010011001",
  14275=>"000110001",
  14276=>"011000100",
  14277=>"001101100",
  14278=>"111000001",
  14279=>"010011101",
  14280=>"010011101",
  14281=>"101110100",
  14282=>"110101111",
  14283=>"101101010",
  14284=>"111001111",
  14285=>"110101001",
  14286=>"110111000",
  14287=>"000101001",
  14288=>"101010011",
  14289=>"011111001",
  14290=>"100110100",
  14291=>"001100001",
  14292=>"100110111",
  14293=>"111000001",
  14294=>"100010000",
  14295=>"011011110",
  14296=>"101110001",
  14297=>"101001101",
  14298=>"101010010",
  14299=>"000111110",
  14300=>"110101001",
  14301=>"010111100",
  14302=>"001010111",
  14303=>"001101010",
  14304=>"000100100",
  14305=>"000101100",
  14306=>"001000100",
  14307=>"111111100",
  14308=>"001111101",
  14309=>"111101111",
  14310=>"111100001",
  14311=>"001000111",
  14312=>"110111111",
  14313=>"000110100",
  14314=>"011101111",
  14315=>"110001011",
  14316=>"000010101",
  14317=>"000100000",
  14318=>"110100110",
  14319=>"101110111",
  14320=>"100010101",
  14321=>"011111101",
  14322=>"101001000",
  14323=>"100010100",
  14324=>"101101010",
  14325=>"110110010",
  14326=>"000110100",
  14327=>"011000001",
  14328=>"010100011",
  14329=>"001000011",
  14330=>"111111010",
  14331=>"100010111",
  14332=>"111101011",
  14333=>"001010010",
  14334=>"111000110",
  14335=>"101011100",
  14336=>"011001010",
  14337=>"100001100",
  14338=>"011001111",
  14339=>"000000011",
  14340=>"011101111",
  14341=>"110110110",
  14342=>"010000111",
  14343=>"101101010",
  14344=>"010001001",
  14345=>"010100111",
  14346=>"000100010",
  14347=>"000001101",
  14348=>"010100011",
  14349=>"010110011",
  14350=>"101101000",
  14351=>"100110110",
  14352=>"110101100",
  14353=>"001001000",
  14354=>"000011111",
  14355=>"011010001",
  14356=>"011110000",
  14357=>"000011110",
  14358=>"110011100",
  14359=>"011111000",
  14360=>"010101000",
  14361=>"000011001",
  14362=>"000111101",
  14363=>"001011011",
  14364=>"010000010",
  14365=>"000001000",
  14366=>"010111000",
  14367=>"010111110",
  14368=>"001001100",
  14369=>"000111001",
  14370=>"101000010",
  14371=>"110010111",
  14372=>"100111000",
  14373=>"011101101",
  14374=>"101100101",
  14375=>"001010011",
  14376=>"111010011",
  14377=>"101110100",
  14378=>"101101001",
  14379=>"110111001",
  14380=>"111100101",
  14381=>"110011010",
  14382=>"101011111",
  14383=>"111100001",
  14384=>"111011101",
  14385=>"000101111",
  14386=>"110111101",
  14387=>"010101111",
  14388=>"000110001",
  14389=>"101000101",
  14390=>"111001110",
  14391=>"001010010",
  14392=>"000000111",
  14393=>"000010010",
  14394=>"000000000",
  14395=>"111100101",
  14396=>"000001110",
  14397=>"100000011",
  14398=>"100011111",
  14399=>"110000111",
  14400=>"111111111",
  14401=>"001001100",
  14402=>"011111001",
  14403=>"110000101",
  14404=>"000001111",
  14405=>"111111010",
  14406=>"001011000",
  14407=>"110001000",
  14408=>"111000010",
  14409=>"110110101",
  14410=>"001101011",
  14411=>"001011011",
  14412=>"001100010",
  14413=>"111010010",
  14414=>"100110010",
  14415=>"010000000",
  14416=>"100010110",
  14417=>"100010101",
  14418=>"001001010",
  14419=>"010111111",
  14420=>"000001001",
  14421=>"100100001",
  14422=>"111100011",
  14423=>"001101011",
  14424=>"000010000",
  14425=>"011110011",
  14426=>"100101010",
  14427=>"011111001",
  14428=>"110010010",
  14429=>"101010011",
  14430=>"010010111",
  14431=>"101111000",
  14432=>"101111101",
  14433=>"000000010",
  14434=>"011110001",
  14435=>"000000010",
  14436=>"101100101",
  14437=>"100100101",
  14438=>"100101010",
  14439=>"011110000",
  14440=>"010111011",
  14441=>"011011110",
  14442=>"001100110",
  14443=>"100000100",
  14444=>"111001000",
  14445=>"101110110",
  14446=>"000000001",
  14447=>"001111111",
  14448=>"010010010",
  14449=>"001100010",
  14450=>"111111110",
  14451=>"101000111",
  14452=>"110100101",
  14453=>"101001000",
  14454=>"010100111",
  14455=>"111001101",
  14456=>"000011101",
  14457=>"100010101",
  14458=>"001110101",
  14459=>"110000000",
  14460=>"110110111",
  14461=>"000110110",
  14462=>"000100010",
  14463=>"010000110",
  14464=>"011010101",
  14465=>"110010011",
  14466=>"111000111",
  14467=>"010010100",
  14468=>"111111011",
  14469=>"000000111",
  14470=>"110010111",
  14471=>"011010100",
  14472=>"111000110",
  14473=>"001101011",
  14474=>"011010110",
  14475=>"011000001",
  14476=>"001100101",
  14477=>"000110111",
  14478=>"001111010",
  14479=>"010010111",
  14480=>"101010101",
  14481=>"110011000",
  14482=>"100111001",
  14483=>"101101100",
  14484=>"000010000",
  14485=>"110011111",
  14486=>"010010110",
  14487=>"101111011",
  14488=>"101101100",
  14489=>"001001010",
  14490=>"110110000",
  14491=>"011101110",
  14492=>"011101001",
  14493=>"100010010",
  14494=>"010110011",
  14495=>"000001011",
  14496=>"000001110",
  14497=>"000011001",
  14498=>"110011110",
  14499=>"000000010",
  14500=>"111000011",
  14501=>"010000100",
  14502=>"010001000",
  14503=>"010100110",
  14504=>"101111011",
  14505=>"100111111",
  14506=>"010001101",
  14507=>"101101101",
  14508=>"000001010",
  14509=>"001000011",
  14510=>"100110110",
  14511=>"010101011",
  14512=>"001011110",
  14513=>"001010010",
  14514=>"100101000",
  14515=>"111111001",
  14516=>"110001110",
  14517=>"101011010",
  14518=>"110110100",
  14519=>"111010111",
  14520=>"011111000",
  14521=>"010110011",
  14522=>"100110001",
  14523=>"110011101",
  14524=>"101011000",
  14525=>"100001111",
  14526=>"101110000",
  14527=>"001100101",
  14528=>"010011101",
  14529=>"010111000",
  14530=>"111010100",
  14531=>"111110110",
  14532=>"000110010",
  14533=>"111111111",
  14534=>"111011101",
  14535=>"111011001",
  14536=>"110111000",
  14537=>"011110011",
  14538=>"111110111",
  14539=>"100111100",
  14540=>"010110011",
  14541=>"010111101",
  14542=>"100000011",
  14543=>"000010110",
  14544=>"101000100",
  14545=>"100000110",
  14546=>"100101010",
  14547=>"111100111",
  14548=>"000000010",
  14549=>"100000001",
  14550=>"100011010",
  14551=>"001111111",
  14552=>"000011100",
  14553=>"100000100",
  14554=>"010110111",
  14555=>"011111001",
  14556=>"000011100",
  14557=>"101010010",
  14558=>"100101011",
  14559=>"101110100",
  14560=>"010010000",
  14561=>"111101101",
  14562=>"110011001",
  14563=>"010000101",
  14564=>"110111101",
  14565=>"000001001",
  14566=>"011111110",
  14567=>"101111100",
  14568=>"001011001",
  14569=>"010111010",
  14570=>"010001101",
  14571=>"000110000",
  14572=>"100100000",
  14573=>"111010011",
  14574=>"110001111",
  14575=>"011011010",
  14576=>"000010001",
  14577=>"111001111",
  14578=>"111011111",
  14579=>"100011000",
  14580=>"011001010",
  14581=>"110111011",
  14582=>"010111001",
  14583=>"100000100",
  14584=>"110001010",
  14585=>"000100010",
  14586=>"100111001",
  14587=>"011100011",
  14588=>"100001101",
  14589=>"001011011",
  14590=>"110101101",
  14591=>"100001101",
  14592=>"000001100",
  14593=>"110110110",
  14594=>"100010010",
  14595=>"111010110",
  14596=>"110010111",
  14597=>"100111000",
  14598=>"010001001",
  14599=>"011101110",
  14600=>"000001111",
  14601=>"010000100",
  14602=>"100110001",
  14603=>"111010110",
  14604=>"100010000",
  14605=>"001100011",
  14606=>"100111000",
  14607=>"001011001",
  14608=>"001111101",
  14609=>"101111111",
  14610=>"011101000",
  14611=>"101011100",
  14612=>"111101011",
  14613=>"110100011",
  14614=>"010100000",
  14615=>"010110000",
  14616=>"101100010",
  14617=>"000001011",
  14618=>"100111000",
  14619=>"011101000",
  14620=>"100010110",
  14621=>"100101101",
  14622=>"101010101",
  14623=>"111110001",
  14624=>"010111011",
  14625=>"001100100",
  14626=>"001110110",
  14627=>"110000110",
  14628=>"101000010",
  14629=>"001101101",
  14630=>"000010100",
  14631=>"100110000",
  14632=>"000100001",
  14633=>"110000111",
  14634=>"100100000",
  14635=>"010101000",
  14636=>"100100111",
  14637=>"010100000",
  14638=>"000100101",
  14639=>"111110100",
  14640=>"001101101",
  14641=>"111111110",
  14642=>"010111010",
  14643=>"000111100",
  14644=>"000111001",
  14645=>"100011001",
  14646=>"010001110",
  14647=>"101110011",
  14648=>"100101101",
  14649=>"000100011",
  14650=>"001000010",
  14651=>"011011101",
  14652=>"010000001",
  14653=>"100101011",
  14654=>"101011101",
  14655=>"111110101",
  14656=>"011101010",
  14657=>"111100101",
  14658=>"101011011",
  14659=>"101110011",
  14660=>"111011110",
  14661=>"011101110",
  14662=>"111010001",
  14663=>"000001100",
  14664=>"100101001",
  14665=>"100110101",
  14666=>"001101001",
  14667=>"010110100",
  14668=>"111101100",
  14669=>"010111011",
  14670=>"011011010",
  14671=>"101101011",
  14672=>"111111001",
  14673=>"100110100",
  14674=>"011101000",
  14675=>"001010001",
  14676=>"100100000",
  14677=>"110101111",
  14678=>"101000000",
  14679=>"111110001",
  14680=>"000111111",
  14681=>"001010010",
  14682=>"011010000",
  14683=>"101011000",
  14684=>"000010010",
  14685=>"010001001",
  14686=>"111100010",
  14687=>"011101100",
  14688=>"101101111",
  14689=>"101010010",
  14690=>"000000111",
  14691=>"000101000",
  14692=>"011111111",
  14693=>"000100111",
  14694=>"000000100",
  14695=>"111111000",
  14696=>"000000110",
  14697=>"011111000",
  14698=>"010101010",
  14699=>"011001100",
  14700=>"111100010",
  14701=>"111000001",
  14702=>"100010100",
  14703=>"111101101",
  14704=>"010010000",
  14705=>"111011011",
  14706=>"001111011",
  14707=>"100101110",
  14708=>"111101111",
  14709=>"111001001",
  14710=>"000100111",
  14711=>"011000011",
  14712=>"111001010",
  14713=>"110101000",
  14714=>"111000011",
  14715=>"011101010",
  14716=>"011011110",
  14717=>"000010000",
  14718=>"111111101",
  14719=>"011101111",
  14720=>"000000010",
  14721=>"000000011",
  14722=>"100011001",
  14723=>"110000011",
  14724=>"111000110",
  14725=>"111101110",
  14726=>"011011001",
  14727=>"000000000",
  14728=>"000011010",
  14729=>"101001111",
  14730=>"011100011",
  14731=>"100000011",
  14732=>"000010011",
  14733=>"010110111",
  14734=>"101011000",
  14735=>"111101100",
  14736=>"011000011",
  14737=>"110010000",
  14738=>"011001011",
  14739=>"010101001",
  14740=>"111001100",
  14741=>"010100111",
  14742=>"000000000",
  14743=>"001111101",
  14744=>"000000101",
  14745=>"001100111",
  14746=>"011010010",
  14747=>"111101110",
  14748=>"011111001",
  14749=>"010001101",
  14750=>"011010100",
  14751=>"100111110",
  14752=>"010110000",
  14753=>"111101111",
  14754=>"100001110",
  14755=>"011000100",
  14756=>"100000010",
  14757=>"001100110",
  14758=>"100000100",
  14759=>"010111001",
  14760=>"001101111",
  14761=>"011101001",
  14762=>"000011101",
  14763=>"001111010",
  14764=>"101110000",
  14765=>"100111111",
  14766=>"111110001",
  14767=>"011001000",
  14768=>"111110001",
  14769=>"000110001",
  14770=>"110110011",
  14771=>"000111010",
  14772=>"101100111",
  14773=>"101010111",
  14774=>"111111111",
  14775=>"001111111",
  14776=>"111101111",
  14777=>"110101001",
  14778=>"000000101",
  14779=>"010010101",
  14780=>"110010001",
  14781=>"111111111",
  14782=>"000000100",
  14783=>"001101000",
  14784=>"111110000",
  14785=>"100011001",
  14786=>"111001101",
  14787=>"110001111",
  14788=>"100111010",
  14789=>"111111011",
  14790=>"111100001",
  14791=>"010110011",
  14792=>"110011000",
  14793=>"110011001",
  14794=>"110010011",
  14795=>"101000101",
  14796=>"100001000",
  14797=>"111100110",
  14798=>"011000100",
  14799=>"110100110",
  14800=>"110110101",
  14801=>"100101100",
  14802=>"100110111",
  14803=>"100111010",
  14804=>"001100101",
  14805=>"111011011",
  14806=>"100011011",
  14807=>"000101111",
  14808=>"111001011",
  14809=>"010101010",
  14810=>"001100000",
  14811=>"011000010",
  14812=>"101101100",
  14813=>"110110101",
  14814=>"001001111",
  14815=>"110010001",
  14816=>"001000001",
  14817=>"111010011",
  14818=>"011100011",
  14819=>"101000011",
  14820=>"001011001",
  14821=>"000011110",
  14822=>"000010000",
  14823=>"001010111",
  14824=>"100011101",
  14825=>"001001001",
  14826=>"001100101",
  14827=>"111111010",
  14828=>"000100111",
  14829=>"000110011",
  14830=>"001000000",
  14831=>"010110001",
  14832=>"111101111",
  14833=>"000111000",
  14834=>"110100111",
  14835=>"000001010",
  14836=>"011110100",
  14837=>"110100000",
  14838=>"000110100",
  14839=>"100100111",
  14840=>"010001001",
  14841=>"101010000",
  14842=>"100101111",
  14843=>"011001010",
  14844=>"000111110",
  14845=>"100101001",
  14846=>"101100101",
  14847=>"010001110",
  14848=>"110100001",
  14849=>"000000001",
  14850=>"010011111",
  14851=>"001110110",
  14852=>"010001000",
  14853=>"000011001",
  14854=>"101011001",
  14855=>"000000100",
  14856=>"111110100",
  14857=>"110001110",
  14858=>"111001110",
  14859=>"101011100",
  14860=>"001011101",
  14861=>"100010100",
  14862=>"111101000",
  14863=>"001111101",
  14864=>"111010111",
  14865=>"011001001",
  14866=>"110001101",
  14867=>"111111011",
  14868=>"001000100",
  14869=>"001001000",
  14870=>"010100001",
  14871=>"001010010",
  14872=>"001100101",
  14873=>"110111111",
  14874=>"110001000",
  14875=>"000111111",
  14876=>"111111101",
  14877=>"010011001",
  14878=>"111011011",
  14879=>"100101010",
  14880=>"000100001",
  14881=>"111111011",
  14882=>"110010000",
  14883=>"011000101",
  14884=>"000001100",
  14885=>"000100001",
  14886=>"010110100",
  14887=>"010001001",
  14888=>"001110100",
  14889=>"110110010",
  14890=>"010110010",
  14891=>"001011100",
  14892=>"111010011",
  14893=>"111100011",
  14894=>"101000111",
  14895=>"111101001",
  14896=>"010110000",
  14897=>"110011000",
  14898=>"001010000",
  14899=>"111011111",
  14900=>"100010101",
  14901=>"000000101",
  14902=>"110010011",
  14903=>"101101011",
  14904=>"011000000",
  14905=>"000010000",
  14906=>"110101010",
  14907=>"111000100",
  14908=>"011011111",
  14909=>"000011001",
  14910=>"100100110",
  14911=>"001110011",
  14912=>"011110010",
  14913=>"100000100",
  14914=>"010101011",
  14915=>"111100100",
  14916=>"001010100",
  14917=>"001000101",
  14918=>"100000010",
  14919=>"000011000",
  14920=>"001001110",
  14921=>"010011011",
  14922=>"110000111",
  14923=>"110000100",
  14924=>"111100111",
  14925=>"001011011",
  14926=>"100100110",
  14927=>"000010011",
  14928=>"111111000",
  14929=>"011111011",
  14930=>"010011111",
  14931=>"010010000",
  14932=>"100001000",
  14933=>"001110101",
  14934=>"011001000",
  14935=>"110011110",
  14936=>"111000001",
  14937=>"101001000",
  14938=>"110000111",
  14939=>"111101101",
  14940=>"101111100",
  14941=>"111110010",
  14942=>"011000101",
  14943=>"011111111",
  14944=>"000110011",
  14945=>"111001011",
  14946=>"001111000",
  14947=>"001001101",
  14948=>"110010011",
  14949=>"111000011",
  14950=>"100110100",
  14951=>"110111110",
  14952=>"110011101",
  14953=>"101000100",
  14954=>"010000000",
  14955=>"001111111",
  14956=>"000001001",
  14957=>"100101010",
  14958=>"001110101",
  14959=>"010001111",
  14960=>"010010011",
  14961=>"010011100",
  14962=>"110010110",
  14963=>"100110111",
  14964=>"000001111",
  14965=>"000100011",
  14966=>"111000011",
  14967=>"111000000",
  14968=>"011000000",
  14969=>"010001010",
  14970=>"000010010",
  14971=>"011010011",
  14972=>"000001000",
  14973=>"010100001",
  14974=>"001000110",
  14975=>"101110110",
  14976=>"111100110",
  14977=>"011110100",
  14978=>"010010101",
  14979=>"110000010",
  14980=>"100111111",
  14981=>"101001100",
  14982=>"100000111",
  14983=>"110011000",
  14984=>"111111110",
  14985=>"001011101",
  14986=>"110110111",
  14987=>"110100001",
  14988=>"011011000",
  14989=>"001111010",
  14990=>"011001000",
  14991=>"110110000",
  14992=>"010110100",
  14993=>"010101100",
  14994=>"010101111",
  14995=>"101101001",
  14996=>"100010000",
  14997=>"100001110",
  14998=>"111000001",
  14999=>"101001101",
  15000=>"101100011",
  15001=>"110101111",
  15002=>"101110000",
  15003=>"010101101",
  15004=>"101010001",
  15005=>"100011001",
  15006=>"001110001",
  15007=>"011000111",
  15008=>"111110000",
  15009=>"000101101",
  15010=>"110001111",
  15011=>"010010111",
  15012=>"001010100",
  15013=>"000101010",
  15014=>"101101011",
  15015=>"000011001",
  15016=>"111101110",
  15017=>"100110111",
  15018=>"011100011",
  15019=>"110011000",
  15020=>"000000001",
  15021=>"111100001",
  15022=>"001010010",
  15023=>"011010111",
  15024=>"001001111",
  15025=>"011001101",
  15026=>"110101000",
  15027=>"110000100",
  15028=>"000110110",
  15029=>"111111101",
  15030=>"111111010",
  15031=>"011100001",
  15032=>"011101110",
  15033=>"001101100",
  15034=>"110101101",
  15035=>"000001100",
  15036=>"011111011",
  15037=>"111100100",
  15038=>"111000001",
  15039=>"000011001",
  15040=>"101110000",
  15041=>"101100111",
  15042=>"111101110",
  15043=>"101100111",
  15044=>"101010110",
  15045=>"000110111",
  15046=>"010000100",
  15047=>"110110001",
  15048=>"010001100",
  15049=>"010001110",
  15050=>"101010100",
  15051=>"110100010",
  15052=>"101011010",
  15053=>"001011001",
  15054=>"010011101",
  15055=>"000101001",
  15056=>"110111101",
  15057=>"001111100",
  15058=>"111110110",
  15059=>"101000100",
  15060=>"010111110",
  15061=>"000111001",
  15062=>"101110100",
  15063=>"011010110",
  15064=>"000110010",
  15065=>"011101111",
  15066=>"111111101",
  15067=>"100011110",
  15068=>"010010111",
  15069=>"101001001",
  15070=>"001100011",
  15071=>"100111101",
  15072=>"110001000",
  15073=>"010111100",
  15074=>"101000101",
  15075=>"011001000",
  15076=>"110101100",
  15077=>"011010001",
  15078=>"001001100",
  15079=>"110001111",
  15080=>"010111011",
  15081=>"111000000",
  15082=>"101010111",
  15083=>"100001010",
  15084=>"001110000",
  15085=>"101101001",
  15086=>"101000010",
  15087=>"111111111",
  15088=>"011111000",
  15089=>"011001110",
  15090=>"100011100",
  15091=>"101100101",
  15092=>"000010011",
  15093=>"010101010",
  15094=>"100010111",
  15095=>"000011111",
  15096=>"010000010",
  15097=>"100111000",
  15098=>"110100100",
  15099=>"111001101",
  15100=>"111001001",
  15101=>"101001001",
  15102=>"110001110",
  15103=>"100011000",
  15104=>"001000110",
  15105=>"000010011",
  15106=>"010111100",
  15107=>"100011110",
  15108=>"111101000",
  15109=>"110000100",
  15110=>"110111010",
  15111=>"000011110",
  15112=>"100111000",
  15113=>"100110110",
  15114=>"101100010",
  15115=>"000100010",
  15116=>"001101111",
  15117=>"010000001",
  15118=>"000101101",
  15119=>"001001111",
  15120=>"101011010",
  15121=>"110001001",
  15122=>"011110000",
  15123=>"011000101",
  15124=>"110110101",
  15125=>"101101101",
  15126=>"101100111",
  15127=>"100100011",
  15128=>"001000010",
  15129=>"100111010",
  15130=>"111100110",
  15131=>"111100111",
  15132=>"010011001",
  15133=>"111010100",
  15134=>"010010001",
  15135=>"010010111",
  15136=>"000000101",
  15137=>"100001011",
  15138=>"110101111",
  15139=>"101100010",
  15140=>"000001001",
  15141=>"011110101",
  15142=>"100010010",
  15143=>"001010011",
  15144=>"110110010",
  15145=>"110000010",
  15146=>"111000111",
  15147=>"001000000",
  15148=>"110111000",
  15149=>"000100010",
  15150=>"111010001",
  15151=>"101000100",
  15152=>"010101110",
  15153=>"101010100",
  15154=>"010101010",
  15155=>"100110010",
  15156=>"010101000",
  15157=>"101101010",
  15158=>"001000100",
  15159=>"000001110",
  15160=>"000010011",
  15161=>"001000010",
  15162=>"000111100",
  15163=>"110010000",
  15164=>"110110100",
  15165=>"001010011",
  15166=>"010101011",
  15167=>"111011000",
  15168=>"001111101",
  15169=>"100111100",
  15170=>"011011010",
  15171=>"110001111",
  15172=>"000100011",
  15173=>"110001101",
  15174=>"111100100",
  15175=>"111100010",
  15176=>"000010000",
  15177=>"000011000",
  15178=>"000110111",
  15179=>"110000110",
  15180=>"101111010",
  15181=>"100011100",
  15182=>"001001110",
  15183=>"001111011",
  15184=>"000110010",
  15185=>"100100110",
  15186=>"111100011",
  15187=>"011110000",
  15188=>"101111110",
  15189=>"110001011",
  15190=>"011001000",
  15191=>"000000101",
  15192=>"111100110",
  15193=>"101101110",
  15194=>"000010101",
  15195=>"101010000",
  15196=>"110001001",
  15197=>"010000000",
  15198=>"100010110",
  15199=>"110001011",
  15200=>"001001101",
  15201=>"000010110",
  15202=>"010101100",
  15203=>"110000110",
  15204=>"100000100",
  15205=>"110001011",
  15206=>"110001000",
  15207=>"000000101",
  15208=>"011111100",
  15209=>"011001111",
  15210=>"010001110",
  15211=>"011011001",
  15212=>"010000011",
  15213=>"111000110",
  15214=>"000110100",
  15215=>"100110110",
  15216=>"011010001",
  15217=>"111010110",
  15218=>"100110000",
  15219=>"001001100",
  15220=>"010000011",
  15221=>"100110010",
  15222=>"001001101",
  15223=>"001100001",
  15224=>"111001101",
  15225=>"000001111",
  15226=>"100111010",
  15227=>"000011100",
  15228=>"111110000",
  15229=>"001010110",
  15230=>"001110111",
  15231=>"111101110",
  15232=>"010101111",
  15233=>"111001000",
  15234=>"000010110",
  15235=>"001111001",
  15236=>"111011010",
  15237=>"000100100",
  15238=>"100110001",
  15239=>"010000101",
  15240=>"111100010",
  15241=>"111100101",
  15242=>"000001110",
  15243=>"100000000",
  15244=>"101110111",
  15245=>"011110011",
  15246=>"100011101",
  15247=>"111001101",
  15248=>"001101001",
  15249=>"101101001",
  15250=>"011110001",
  15251=>"001000110",
  15252=>"100011111",
  15253=>"010101101",
  15254=>"001110100",
  15255=>"110100001",
  15256=>"101110101",
  15257=>"111010010",
  15258=>"000111110",
  15259=>"010011100",
  15260=>"111011011",
  15261=>"000100110",
  15262=>"110111111",
  15263=>"001011110",
  15264=>"000110001",
  15265=>"100000001",
  15266=>"010110100",
  15267=>"011000000",
  15268=>"001001100",
  15269=>"110011101",
  15270=>"001101010",
  15271=>"000111000",
  15272=>"011010101",
  15273=>"000010101",
  15274=>"111100010",
  15275=>"000010101",
  15276=>"011100010",
  15277=>"110100111",
  15278=>"101001100",
  15279=>"101100001",
  15280=>"100010111",
  15281=>"001101001",
  15282=>"110100011",
  15283=>"101111100",
  15284=>"010001111",
  15285=>"010011010",
  15286=>"111110001",
  15287=>"011101000",
  15288=>"001011000",
  15289=>"001001011",
  15290=>"010001000",
  15291=>"001010010",
  15292=>"110001000",
  15293=>"011111101",
  15294=>"000101000",
  15295=>"001101111",
  15296=>"110111011",
  15297=>"111101100",
  15298=>"011100111",
  15299=>"010000100",
  15300=>"000100101",
  15301=>"111100101",
  15302=>"011111111",
  15303=>"001010011",
  15304=>"111011110",
  15305=>"001111111",
  15306=>"111100111",
  15307=>"111101001",
  15308=>"001000101",
  15309=>"011110000",
  15310=>"011011100",
  15311=>"111011100",
  15312=>"011101000",
  15313=>"000110110",
  15314=>"011010000",
  15315=>"000100010",
  15316=>"100111011",
  15317=>"100111001",
  15318=>"011010100",
  15319=>"110100100",
  15320=>"011000101",
  15321=>"010010000",
  15322=>"010011111",
  15323=>"010001011",
  15324=>"001001000",
  15325=>"111101001",
  15326=>"000000100",
  15327=>"001010010",
  15328=>"101110111",
  15329=>"111001000",
  15330=>"011101110",
  15331=>"011010001",
  15332=>"110001100",
  15333=>"111110011",
  15334=>"000110101",
  15335=>"110111111",
  15336=>"110100010",
  15337=>"000011000",
  15338=>"001011001",
  15339=>"101101100",
  15340=>"000010010",
  15341=>"001110010",
  15342=>"011010110",
  15343=>"110000100",
  15344=>"100110000",
  15345=>"111001101",
  15346=>"110001001",
  15347=>"011010111",
  15348=>"100111110",
  15349=>"010110010",
  15350=>"101111110",
  15351=>"100100001",
  15352=>"111101001",
  15353=>"000100011",
  15354=>"100011010",
  15355=>"010010000",
  15356=>"100011001",
  15357=>"000001101",
  15358=>"111110011",
  15359=>"010111000",
  15360=>"001000111",
  15361=>"011100001",
  15362=>"101000111",
  15363=>"000010010",
  15364=>"000111101",
  15365=>"011010110",
  15366=>"100101110",
  15367=>"011100101",
  15368=>"111010011",
  15369=>"001101100",
  15370=>"000000100",
  15371=>"010010101",
  15372=>"101000100",
  15373=>"110001000",
  15374=>"010100101",
  15375=>"100101111",
  15376=>"011001100",
  15377=>"011001011",
  15378=>"111111111",
  15379=>"001110101",
  15380=>"110001010",
  15381=>"100011000",
  15382=>"010011110",
  15383=>"111111100",
  15384=>"101110100",
  15385=>"101110100",
  15386=>"110011111",
  15387=>"001011101",
  15388=>"000001101",
  15389=>"001011010",
  15390=>"111010010",
  15391=>"000111001",
  15392=>"110000000",
  15393=>"100111100",
  15394=>"001000001",
  15395=>"101101101",
  15396=>"000101101",
  15397=>"001000000",
  15398=>"101011111",
  15399=>"011011100",
  15400=>"100000010",
  15401=>"000110000",
  15402=>"011010100",
  15403=>"101110001",
  15404=>"100100100",
  15405=>"100001111",
  15406=>"001010011",
  15407=>"000111010",
  15408=>"100010000",
  15409=>"101101111",
  15410=>"111101101",
  15411=>"010010111",
  15412=>"110010001",
  15413=>"000000001",
  15414=>"100001000",
  15415=>"010011111",
  15416=>"101110000",
  15417=>"100010101",
  15418=>"010111101",
  15419=>"110100001",
  15420=>"000000110",
  15421=>"000110110",
  15422=>"010111101",
  15423=>"010001010",
  15424=>"001010000",
  15425=>"000011110",
  15426=>"001000000",
  15427=>"000011111",
  15428=>"111101111",
  15429=>"110011100",
  15430=>"010111101",
  15431=>"000001001",
  15432=>"111000001",
  15433=>"000010110",
  15434=>"110001111",
  15435=>"011011001",
  15436=>"010010010",
  15437=>"100101000",
  15438=>"001001000",
  15439=>"001100100",
  15440=>"000110111",
  15441=>"110110000",
  15442=>"101001110",
  15443=>"000011001",
  15444=>"100101110",
  15445=>"010010110",
  15446=>"110111001",
  15447=>"001000110",
  15448=>"111110111",
  15449=>"010010101",
  15450=>"001100100",
  15451=>"000011101",
  15452=>"001100001",
  15453=>"100111110",
  15454=>"111011000",
  15455=>"011001101",
  15456=>"000000110",
  15457=>"100011110",
  15458=>"100110010",
  15459=>"101010000",
  15460=>"100110000",
  15461=>"100010010",
  15462=>"111011000",
  15463=>"010110010",
  15464=>"100100110",
  15465=>"001000000",
  15466=>"011111010",
  15467=>"101110111",
  15468=>"000010100",
  15469=>"011010000",
  15470=>"100110100",
  15471=>"101110110",
  15472=>"100001000",
  15473=>"001111011",
  15474=>"100011000",
  15475=>"111110001",
  15476=>"011000101",
  15477=>"101101011",
  15478=>"111011111",
  15479=>"011010000",
  15480=>"000001110",
  15481=>"110010010",
  15482=>"111001001",
  15483=>"101110010",
  15484=>"111101111",
  15485=>"010100010",
  15486=>"010101101",
  15487=>"100000100",
  15488=>"000001110",
  15489=>"101111010",
  15490=>"001000101",
  15491=>"100000000",
  15492=>"000001010",
  15493=>"100011111",
  15494=>"000101111",
  15495=>"100000110",
  15496=>"111110001",
  15497=>"101001110",
  15498=>"000000001",
  15499=>"001011001",
  15500=>"001001111",
  15501=>"111011010",
  15502=>"100111000",
  15503=>"101110000",
  15504=>"100110000",
  15505=>"000010110",
  15506=>"000001111",
  15507=>"001000110",
  15508=>"010110101",
  15509=>"011011001",
  15510=>"100001001",
  15511=>"010100010",
  15512=>"000001101",
  15513=>"110000101",
  15514=>"111100001",
  15515=>"100001011",
  15516=>"000011000",
  15517=>"110110111",
  15518=>"011111010",
  15519=>"111000110",
  15520=>"110000101",
  15521=>"111011111",
  15522=>"001000011",
  15523=>"110100110",
  15524=>"100111011",
  15525=>"100111000",
  15526=>"111101011",
  15527=>"010010110",
  15528=>"011010000",
  15529=>"000000001",
  15530=>"101100110",
  15531=>"111101000",
  15532=>"010011100",
  15533=>"000101011",
  15534=>"100110101",
  15535=>"001010100",
  15536=>"100011001",
  15537=>"110011000",
  15538=>"001100110",
  15539=>"011010011",
  15540=>"100100000",
  15541=>"011100101",
  15542=>"111101110",
  15543=>"110111011",
  15544=>"010010010",
  15545=>"101101100",
  15546=>"011100010",
  15547=>"101100100",
  15548=>"110100000",
  15549=>"001010011",
  15550=>"011111000",
  15551=>"100000010",
  15552=>"100101011",
  15553=>"110100111",
  15554=>"010000000",
  15555=>"011010010",
  15556=>"110011100",
  15557=>"101111010",
  15558=>"111101010",
  15559=>"111110010",
  15560=>"011011000",
  15561=>"101110001",
  15562=>"111101111",
  15563=>"101110011",
  15564=>"110010100",
  15565=>"110010110",
  15566=>"011000101",
  15567=>"111101100",
  15568=>"001011100",
  15569=>"001101101",
  15570=>"100101010",
  15571=>"100101101",
  15572=>"111100100",
  15573=>"101001010",
  15574=>"111100001",
  15575=>"010100111",
  15576=>"111011111",
  15577=>"110110101",
  15578=>"111111011",
  15579=>"001101001",
  15580=>"100000011",
  15581=>"010111111",
  15582=>"001010000",
  15583=>"001110100",
  15584=>"100000110",
  15585=>"100100001",
  15586=>"110100110",
  15587=>"100100100",
  15588=>"111100010",
  15589=>"000111110",
  15590=>"010001101",
  15591=>"001011100",
  15592=>"111110000",
  15593=>"101001101",
  15594=>"100101011",
  15595=>"000100001",
  15596=>"100100110",
  15597=>"001000110",
  15598=>"000101011",
  15599=>"001010000",
  15600=>"001010010",
  15601=>"110110011",
  15602=>"010000000",
  15603=>"001101010",
  15604=>"100111101",
  15605=>"011101111",
  15606=>"111110100",
  15607=>"000011110",
  15608=>"100000010",
  15609=>"111100000",
  15610=>"100010111",
  15611=>"000010101",
  15612=>"101010111",
  15613=>"000000111",
  15614=>"000111010",
  15615=>"011011011",
  15616=>"101010001",
  15617=>"101111010",
  15618=>"011100011",
  15619=>"110011111",
  15620=>"001100000",
  15621=>"101010011",
  15622=>"000000111",
  15623=>"111110011",
  15624=>"011110011",
  15625=>"010101111",
  15626=>"101100001",
  15627=>"101111000",
  15628=>"110110101",
  15629=>"100001011",
  15630=>"100001110",
  15631=>"001110111",
  15632=>"010101011",
  15633=>"011100000",
  15634=>"111110101",
  15635=>"000011001",
  15636=>"110110110",
  15637=>"111011100",
  15638=>"011111010",
  15639=>"011001100",
  15640=>"111011111",
  15641=>"101101001",
  15642=>"011111100",
  15643=>"010010000",
  15644=>"100011010",
  15645=>"100000100",
  15646=>"010010010",
  15647=>"000010100",
  15648=>"001011110",
  15649=>"110101010",
  15650=>"010110110",
  15651=>"000001111",
  15652=>"111100100",
  15653=>"000111011",
  15654=>"100101110",
  15655=>"001110111",
  15656=>"101110110",
  15657=>"111110011",
  15658=>"010100100",
  15659=>"001000001",
  15660=>"011011100",
  15661=>"111001011",
  15662=>"100000011",
  15663=>"001001111",
  15664=>"011110110",
  15665=>"000000011",
  15666=>"100100010",
  15667=>"001111111",
  15668=>"101000101",
  15669=>"100100101",
  15670=>"010111101",
  15671=>"110010110",
  15672=>"101011110",
  15673=>"000111000",
  15674=>"101111110",
  15675=>"111110000",
  15676=>"111001001",
  15677=>"000100011",
  15678=>"111010111",
  15679=>"101001101",
  15680=>"111000011",
  15681=>"001000001",
  15682=>"100101101",
  15683=>"110101001",
  15684=>"111001100",
  15685=>"110111001",
  15686=>"000100000",
  15687=>"110101110",
  15688=>"010011101",
  15689=>"000000000",
  15690=>"010101110",
  15691=>"100100001",
  15692=>"100100111",
  15693=>"010001100",
  15694=>"110110011",
  15695=>"110110101",
  15696=>"010011000",
  15697=>"010001001",
  15698=>"100011010",
  15699=>"100101111",
  15700=>"011011010",
  15701=>"001011101",
  15702=>"010100011",
  15703=>"000111100",
  15704=>"110101001",
  15705=>"000100101",
  15706=>"000011010",
  15707=>"100000111",
  15708=>"000100011",
  15709=>"110000110",
  15710=>"111110000",
  15711=>"010100101",
  15712=>"000100101",
  15713=>"000000000",
  15714=>"001000101",
  15715=>"001100010",
  15716=>"100110001",
  15717=>"101011000",
  15718=>"111111001",
  15719=>"111001001",
  15720=>"111010010",
  15721=>"000101110",
  15722=>"101010100",
  15723=>"011011011",
  15724=>"001000110",
  15725=>"110000100",
  15726=>"100110100",
  15727=>"100111111",
  15728=>"000101110",
  15729=>"011011001",
  15730=>"000111010",
  15731=>"100111110",
  15732=>"111011110",
  15733=>"101001111",
  15734=>"110001000",
  15735=>"000001100",
  15736=>"000010111",
  15737=>"110010111",
  15738=>"000010111",
  15739=>"000000000",
  15740=>"110110101",
  15741=>"011111100",
  15742=>"011101000",
  15743=>"001110100",
  15744=>"101101011",
  15745=>"010010000",
  15746=>"011011000",
  15747=>"101011100",
  15748=>"110011101",
  15749=>"000001000",
  15750=>"111011001",
  15751=>"100111111",
  15752=>"010110000",
  15753=>"100000111",
  15754=>"100000011",
  15755=>"101000100",
  15756=>"000111100",
  15757=>"011011000",
  15758=>"001011110",
  15759=>"000000100",
  15760=>"111111101",
  15761=>"101000011",
  15762=>"000000111",
  15763=>"111001101",
  15764=>"111100001",
  15765=>"110110110",
  15766=>"100101000",
  15767=>"101100111",
  15768=>"001001010",
  15769=>"011110000",
  15770=>"111001101",
  15771=>"000000000",
  15772=>"100011100",
  15773=>"111010111",
  15774=>"011110000",
  15775=>"111010011",
  15776=>"010111111",
  15777=>"101000100",
  15778=>"101010000",
  15779=>"100111101",
  15780=>"111101111",
  15781=>"001000100",
  15782=>"000000001",
  15783=>"110011110",
  15784=>"111010011",
  15785=>"010001111",
  15786=>"100111111",
  15787=>"110101100",
  15788=>"110110000",
  15789=>"100100110",
  15790=>"100100110",
  15791=>"010001100",
  15792=>"100010101",
  15793=>"111000100",
  15794=>"110110000",
  15795=>"010110010",
  15796=>"001000000",
  15797=>"011100100",
  15798=>"111111110",
  15799=>"011000000",
  15800=>"101000101",
  15801=>"000111011",
  15802=>"001111111",
  15803=>"111010111",
  15804=>"000100100",
  15805=>"101010100",
  15806=>"110110011",
  15807=>"000111010",
  15808=>"101111000",
  15809=>"001011100",
  15810=>"001100011",
  15811=>"110001101",
  15812=>"101001000",
  15813=>"101000100",
  15814=>"000001000",
  15815=>"000000010",
  15816=>"000000001",
  15817=>"100001111",
  15818=>"100010011",
  15819=>"100011011",
  15820=>"111101110",
  15821=>"011011001",
  15822=>"001000101",
  15823=>"000101110",
  15824=>"111001001",
  15825=>"000110010",
  15826=>"101010000",
  15827=>"000111101",
  15828=>"110111110",
  15829=>"110111000",
  15830=>"111111000",
  15831=>"100111100",
  15832=>"011001000",
  15833=>"010000100",
  15834=>"101111010",
  15835=>"110000100",
  15836=>"001000000",
  15837=>"000010010",
  15838=>"010110000",
  15839=>"110000110",
  15840=>"100001111",
  15841=>"010100011",
  15842=>"001001000",
  15843=>"100011001",
  15844=>"111111101",
  15845=>"111111101",
  15846=>"110000010",
  15847=>"101100000",
  15848=>"000000111",
  15849=>"111100101",
  15850=>"010110001",
  15851=>"010010000",
  15852=>"100011000",
  15853=>"101010111",
  15854=>"101100000",
  15855=>"101110101",
  15856=>"000000001",
  15857=>"100000010",
  15858=>"001001001",
  15859=>"011000011",
  15860=>"100010100",
  15861=>"000110101",
  15862=>"000000100",
  15863=>"110100111",
  15864=>"000100111",
  15865=>"001010011",
  15866=>"110110001",
  15867=>"000000001",
  15868=>"000111011",
  15869=>"110011010",
  15870=>"110100101",
  15871=>"010010111",
  15872=>"110000111",
  15873=>"000011111",
  15874=>"111110110",
  15875=>"110110101",
  15876=>"011111010",
  15877=>"000100110",
  15878=>"110010111",
  15879=>"011000101",
  15880=>"111010010",
  15881=>"100000001",
  15882=>"000001010",
  15883=>"000000011",
  15884=>"000001011",
  15885=>"001111000",
  15886=>"101110000",
  15887=>"000001100",
  15888=>"001101100",
  15889=>"000101101",
  15890=>"110001110",
  15891=>"100111001",
  15892=>"110000101",
  15893=>"101000110",
  15894=>"110000111",
  15895=>"001111000",
  15896=>"100010001",
  15897=>"000010000",
  15898=>"000010000",
  15899=>"110000000",
  15900=>"100001101",
  15901=>"001000001",
  15902=>"010001011",
  15903=>"000000110",
  15904=>"110001000",
  15905=>"110001100",
  15906=>"010011101",
  15907=>"110010101",
  15908=>"101110100",
  15909=>"111010001",
  15910=>"000100001",
  15911=>"011100101",
  15912=>"100110011",
  15913=>"101100100",
  15914=>"101011001",
  15915=>"010000001",
  15916=>"011101110",
  15917=>"110001111",
  15918=>"101011110",
  15919=>"100100100",
  15920=>"000110001",
  15921=>"011101011",
  15922=>"000000001",
  15923=>"100010000",
  15924=>"010010101",
  15925=>"000010110",
  15926=>"010101111",
  15927=>"000001100",
  15928=>"100010010",
  15929=>"010101100",
  15930=>"000000001",
  15931=>"010010001",
  15932=>"001100001",
  15933=>"000010111",
  15934=>"000110001",
  15935=>"111111001",
  15936=>"100100111",
  15937=>"111010110",
  15938=>"110101111",
  15939=>"100100111",
  15940=>"010001011",
  15941=>"100000110",
  15942=>"111110111",
  15943=>"111110100",
  15944=>"100001111",
  15945=>"000000000",
  15946=>"111110000",
  15947=>"110100010",
  15948=>"101010100",
  15949=>"100000101",
  15950=>"111111111",
  15951=>"001110101",
  15952=>"111010011",
  15953=>"011100100",
  15954=>"010000010",
  15955=>"000111011",
  15956=>"101001001",
  15957=>"110101110",
  15958=>"001010001",
  15959=>"001011100",
  15960=>"100000110",
  15961=>"111100100",
  15962=>"101111101",
  15963=>"011001101",
  15964=>"110000000",
  15965=>"100000111",
  15966=>"100111101",
  15967=>"011110001",
  15968=>"000110010",
  15969=>"010110110",
  15970=>"101000000",
  15971=>"000000011",
  15972=>"111101010",
  15973=>"011100001",
  15974=>"111011100",
  15975=>"110100100",
  15976=>"000000001",
  15977=>"010111010",
  15978=>"111011010",
  15979=>"000100111",
  15980=>"100010111",
  15981=>"011110010",
  15982=>"001001011",
  15983=>"100001111",
  15984=>"101011010",
  15985=>"000000011",
  15986=>"001110000",
  15987=>"011011101",
  15988=>"100110011",
  15989=>"001000101",
  15990=>"100000111",
  15991=>"111110111",
  15992=>"111101001",
  15993=>"101100100",
  15994=>"111110011",
  15995=>"100100010",
  15996=>"011001011",
  15997=>"000000110",
  15998=>"110100111",
  15999=>"000111110",
  16000=>"001100110",
  16001=>"001110111",
  16002=>"110000100",
  16003=>"000000000",
  16004=>"000000101",
  16005=>"100010111",
  16006=>"000111000",
  16007=>"110001111",
  16008=>"001111101",
  16009=>"100000100",
  16010=>"111011011",
  16011=>"100000010",
  16012=>"111110100",
  16013=>"100101100",
  16014=>"111001110",
  16015=>"010110101",
  16016=>"010111101",
  16017=>"110010100",
  16018=>"101101111",
  16019=>"011100001",
  16020=>"000000000",
  16021=>"100000001",
  16022=>"101010110",
  16023=>"100000111",
  16024=>"010011101",
  16025=>"001101100",
  16026=>"000001110",
  16027=>"111111101",
  16028=>"011010110",
  16029=>"111011111",
  16030=>"011010100",
  16031=>"011000000",
  16032=>"000111010",
  16033=>"100001000",
  16034=>"000110110",
  16035=>"101000111",
  16036=>"001010101",
  16037=>"001110110",
  16038=>"111011000",
  16039=>"000010100",
  16040=>"000001011",
  16041=>"000100010",
  16042=>"010111011",
  16043=>"010100001",
  16044=>"000011000",
  16045=>"110011011",
  16046=>"011100010",
  16047=>"001001100",
  16048=>"010110010",
  16049=>"101100011",
  16050=>"011100000",
  16051=>"010101000",
  16052=>"111101011",
  16053=>"101000001",
  16054=>"000100101",
  16055=>"100101011",
  16056=>"111011100",
  16057=>"011001100",
  16058=>"101001110",
  16059=>"011011001",
  16060=>"011001011",
  16061=>"000110100",
  16062=>"100000111",
  16063=>"101001001",
  16064=>"111101010",
  16065=>"001101100",
  16066=>"100110000",
  16067=>"001000000",
  16068=>"001010001",
  16069=>"000000000",
  16070=>"110100011",
  16071=>"001000111",
  16072=>"111011101",
  16073=>"111100001",
  16074=>"011011101",
  16075=>"110010110",
  16076=>"000001100",
  16077=>"010001101",
  16078=>"101010101",
  16079=>"111001101",
  16080=>"010001111",
  16081=>"000110100",
  16082=>"010010010",
  16083=>"000000100",
  16084=>"111000100",
  16085=>"010000011",
  16086=>"111111100",
  16087=>"011111111",
  16088=>"100101110",
  16089=>"101101001",
  16090=>"110111001",
  16091=>"111000001",
  16092=>"101101011",
  16093=>"100100110",
  16094=>"111011101",
  16095=>"010111001",
  16096=>"011111011",
  16097=>"000000111",
  16098=>"011010110",
  16099=>"001011001",
  16100=>"100010011",
  16101=>"010001101",
  16102=>"010100101",
  16103=>"001010111",
  16104=>"001011110",
  16105=>"110011010",
  16106=>"010000110",
  16107=>"000100010",
  16108=>"001101111",
  16109=>"110100100",
  16110=>"001000001",
  16111=>"110100110",
  16112=>"111011001",
  16113=>"101100000",
  16114=>"111001011",
  16115=>"001110111",
  16116=>"001010001",
  16117=>"011000011",
  16118=>"110010101",
  16119=>"000110110",
  16120=>"111111101",
  16121=>"000100111",
  16122=>"001101001",
  16123=>"000000011",
  16124=>"011011001",
  16125=>"000000101",
  16126=>"110110000",
  16127=>"001010111",
  16128=>"000111000",
  16129=>"000001011",
  16130=>"110111000",
  16131=>"110111010",
  16132=>"011000001",
  16133=>"000100000",
  16134=>"010110001",
  16135=>"110011101",
  16136=>"100111011",
  16137=>"010110000",
  16138=>"011010110",
  16139=>"010001010",
  16140=>"001000000",
  16141=>"011101000",
  16142=>"111101001",
  16143=>"111011110",
  16144=>"001101111",
  16145=>"100100100",
  16146=>"011110101",
  16147=>"101100110",
  16148=>"110110101",
  16149=>"011110110",
  16150=>"101110000",
  16151=>"100101111",
  16152=>"000010110",
  16153=>"000001000",
  16154=>"110011111",
  16155=>"000010001",
  16156=>"101111000",
  16157=>"010110011",
  16158=>"100111001",
  16159=>"000001001",
  16160=>"110110111",
  16161=>"000001110",
  16162=>"001001011",
  16163=>"111100100",
  16164=>"100101101",
  16165=>"110111111",
  16166=>"000000111",
  16167=>"001101010",
  16168=>"100010010",
  16169=>"010000100",
  16170=>"010001100",
  16171=>"101000110",
  16172=>"111101111",
  16173=>"011111010",
  16174=>"010111011",
  16175=>"101010001",
  16176=>"100110101",
  16177=>"100110011",
  16178=>"100111000",
  16179=>"111110011",
  16180=>"111000100",
  16181=>"100100010",
  16182=>"000100000",
  16183=>"001100111",
  16184=>"100001111",
  16185=>"110101101",
  16186=>"001010111",
  16187=>"000000000",
  16188=>"100010000",
  16189=>"000000000",
  16190=>"001001100",
  16191=>"000111010",
  16192=>"000110011",
  16193=>"110001000",
  16194=>"000100010",
  16195=>"001110001",
  16196=>"111111101",
  16197=>"010010001",
  16198=>"100100111",
  16199=>"010000111",
  16200=>"001110010",
  16201=>"101110010",
  16202=>"100010111",
  16203=>"100011010",
  16204=>"010100001",
  16205=>"101111001",
  16206=>"000100011",
  16207=>"101010011",
  16208=>"100111011",
  16209=>"110111110",
  16210=>"100100000",
  16211=>"101010111",
  16212=>"001111001",
  16213=>"010011010",
  16214=>"011001111",
  16215=>"101111111",
  16216=>"111001111",
  16217=>"000010011",
  16218=>"010111010",
  16219=>"001000101",
  16220=>"111000111",
  16221=>"111000010",
  16222=>"001110011",
  16223=>"110011110",
  16224=>"101001001",
  16225=>"100100100",
  16226=>"000001010",
  16227=>"000100100",
  16228=>"101001100",
  16229=>"001100010",
  16230=>"011000001",
  16231=>"011100000",
  16232=>"000000001",
  16233=>"001001001",
  16234=>"100111111",
  16235=>"100010101",
  16236=>"000000111",
  16237=>"100000111",
  16238=>"101101101",
  16239=>"010100001",
  16240=>"101110110",
  16241=>"111100010",
  16242=>"101010110",
  16243=>"011100111",
  16244=>"100101111",
  16245=>"110011101",
  16246=>"010111110",
  16247=>"101010111",
  16248=>"001010100",
  16249=>"111000111",
  16250=>"010001010",
  16251=>"001010101",
  16252=>"000000000",
  16253=>"001000011",
  16254=>"001110111",
  16255=>"111011000",
  16256=>"001011010",
  16257=>"001001000",
  16258=>"000000011",
  16259=>"110101101",
  16260=>"110101110",
  16261=>"010111000",
  16262=>"000101111",
  16263=>"100010100",
  16264=>"010101101",
  16265=>"011011101",
  16266=>"111111100",
  16267=>"010100110",
  16268=>"000011111",
  16269=>"111111010",
  16270=>"100100001",
  16271=>"100111111",
  16272=>"100110111",
  16273=>"111110111",
  16274=>"100101001",
  16275=>"000011110",
  16276=>"001011011",
  16277=>"101010110",
  16278=>"111101100",
  16279=>"000010111",
  16280=>"101001111",
  16281=>"100100011",
  16282=>"011110111",
  16283=>"100100010",
  16284=>"101010010",
  16285=>"110010001",
  16286=>"010110001",
  16287=>"110101110",
  16288=>"000001001",
  16289=>"110000011",
  16290=>"000000101",
  16291=>"100001000",
  16292=>"011101001",
  16293=>"010111010",
  16294=>"011111011",
  16295=>"001001001",
  16296=>"100001100",
  16297=>"100000111",
  16298=>"011011001",
  16299=>"100100001",
  16300=>"001101100",
  16301=>"111001101",
  16302=>"111111101",
  16303=>"100001101",
  16304=>"010001010",
  16305=>"111000111",
  16306=>"100101011",
  16307=>"101000101",
  16308=>"111100111",
  16309=>"101000100",
  16310=>"000110010",
  16311=>"000001101",
  16312=>"110011000",
  16313=>"010101110",
  16314=>"000110101",
  16315=>"011110011",
  16316=>"000101011",
  16317=>"111110110",
  16318=>"000010111",
  16319=>"000000011",
  16320=>"111101101",
  16321=>"101010001",
  16322=>"000011010",
  16323=>"110011110",
  16324=>"000111010",
  16325=>"110001100",
  16326=>"110000011",
  16327=>"111000111",
  16328=>"000000010",
  16329=>"000100000",
  16330=>"010011111",
  16331=>"110111111",
  16332=>"111011010",
  16333=>"111011000",
  16334=>"111011110",
  16335=>"101001111",
  16336=>"100100001",
  16337=>"000101111",
  16338=>"010101101",
  16339=>"101010011",
  16340=>"110001010",
  16341=>"111010000",
  16342=>"001001010",
  16343=>"100001010",
  16344=>"101111100",
  16345=>"011000011",
  16346=>"100011001",
  16347=>"000011011",
  16348=>"110011000",
  16349=>"100011100",
  16350=>"010111110",
  16351=>"000101000",
  16352=>"111101011",
  16353=>"101001100",
  16354=>"110011011",
  16355=>"011000101",
  16356=>"010110000",
  16357=>"111011110",
  16358=>"001100011",
  16359=>"010110000",
  16360=>"000011001",
  16361=>"010011000",
  16362=>"111010110",
  16363=>"011111110",
  16364=>"010001000",
  16365=>"010100000",
  16366=>"000100011",
  16367=>"100110111",
  16368=>"110110111",
  16369=>"001111110",
  16370=>"111111001",
  16371=>"011100101",
  16372=>"111111000",
  16373=>"010110001",
  16374=>"011111110",
  16375=>"100001111",
  16376=>"011011100",
  16377=>"001100100",
  16378=>"101111000",
  16379=>"100101000",
  16380=>"100100101",
  16381=>"010100000",
  16382=>"001001111",
  16383=>"000110010",
  16384=>"111000001",
  16385=>"110111110",
  16386=>"001010101",
  16387=>"110001011",
  16388=>"111100110",
  16389=>"011001001",
  16390=>"011011110",
  16391=>"100111001",
  16392=>"101100010",
  16393=>"001000011",
  16394=>"111111101",
  16395=>"111100001",
  16396=>"010111000",
  16397=>"111100000",
  16398=>"101011001",
  16399=>"011100011",
  16400=>"100110111",
  16401=>"011011001",
  16402=>"000111110",
  16403=>"101111011",
  16404=>"010110111",
  16405=>"110001101",
  16406=>"110110000",
  16407=>"001111001",
  16408=>"001011001",
  16409=>"101011011",
  16410=>"110111110",
  16411=>"011010110",
  16412=>"100101110",
  16413=>"101100000",
  16414=>"011110100",
  16415=>"100111011",
  16416=>"111111111",
  16417=>"101111111",
  16418=>"101101001",
  16419=>"100100000",
  16420=>"110101000",
  16421=>"011101110",
  16422=>"000110100",
  16423=>"011110101",
  16424=>"000110010",
  16425=>"010000111",
  16426=>"111010000",
  16427=>"010101000",
  16428=>"110111000",
  16429=>"101110100",
  16430=>"000010100",
  16431=>"010110110",
  16432=>"100100100",
  16433=>"011000111",
  16434=>"100111111",
  16435=>"110111001",
  16436=>"101011100",
  16437=>"110011000",
  16438=>"000011010",
  16439=>"111100101",
  16440=>"001101111",
  16441=>"000110110",
  16442=>"111011011",
  16443=>"101010000",
  16444=>"111001010",
  16445=>"011111111",
  16446=>"100100111",
  16447=>"111101111",
  16448=>"001000000",
  16449=>"110000101",
  16450=>"000101110",
  16451=>"100001010",
  16452=>"110110100",
  16453=>"001101101",
  16454=>"110011000",
  16455=>"000100001",
  16456=>"000000000",
  16457=>"110110111",
  16458=>"000111101",
  16459=>"000010101",
  16460=>"101001110",
  16461=>"110110100",
  16462=>"110111111",
  16463=>"001010010",
  16464=>"100001111",
  16465=>"111001011",
  16466=>"011111111",
  16467=>"100011101",
  16468=>"011010011",
  16469=>"100000101",
  16470=>"011011011",
  16471=>"110001001",
  16472=>"111001110",
  16473=>"111100100",
  16474=>"011011001",
  16475=>"000000100",
  16476=>"100001101",
  16477=>"011001011",
  16478=>"101100110",
  16479=>"101001110",
  16480=>"011010101",
  16481=>"010100111",
  16482=>"100011000",
  16483=>"111001000",
  16484=>"100001100",
  16485=>"101001101",
  16486=>"000111111",
  16487=>"100000101",
  16488=>"110011011",
  16489=>"011010000",
  16490=>"000001001",
  16491=>"001111000",
  16492=>"110011001",
  16493=>"001000001",
  16494=>"100010010",
  16495=>"111000110",
  16496=>"110010011",
  16497=>"100011010",
  16498=>"110110101",
  16499=>"000111100",
  16500=>"111011110",
  16501=>"101001011",
  16502=>"100010110",
  16503=>"011111010",
  16504=>"000101111",
  16505=>"010101111",
  16506=>"010001110",
  16507=>"010001001",
  16508=>"001011110",
  16509=>"110010000",
  16510=>"000000101",
  16511=>"001100011",
  16512=>"011000100",
  16513=>"101011011",
  16514=>"111011100",
  16515=>"110000000",
  16516=>"100111100",
  16517=>"010101100",
  16518=>"001001011",
  16519=>"010111000",
  16520=>"000000000",
  16521=>"111000010",
  16522=>"011001001",
  16523=>"110010101",
  16524=>"101101111",
  16525=>"010101000",
  16526=>"010101111",
  16527=>"001101100",
  16528=>"011101111",
  16529=>"100111011",
  16530=>"110111011",
  16531=>"010111001",
  16532=>"101110110",
  16533=>"111110100",
  16534=>"010001010",
  16535=>"000100110",
  16536=>"010001111",
  16537=>"010101100",
  16538=>"000000100",
  16539=>"000001110",
  16540=>"010011011",
  16541=>"001110001",
  16542=>"010010001",
  16543=>"001010010",
  16544=>"001110101",
  16545=>"010111011",
  16546=>"110100000",
  16547=>"010111010",
  16548=>"010011000",
  16549=>"111101111",
  16550=>"011001011",
  16551=>"110101010",
  16552=>"110100110",
  16553=>"111111001",
  16554=>"001100110",
  16555=>"001011010",
  16556=>"011000000",
  16557=>"000000001",
  16558=>"000100100",
  16559=>"111110001",
  16560=>"001011111",
  16561=>"000101010",
  16562=>"010110000",
  16563=>"000101010",
  16564=>"110101101",
  16565=>"011110001",
  16566=>"100110010",
  16567=>"110011110",
  16568=>"110001100",
  16569=>"011010111",
  16570=>"000000001",
  16571=>"001000111",
  16572=>"011001111",
  16573=>"100101011",
  16574=>"000011110",
  16575=>"010000100",
  16576=>"101110011",
  16577=>"011011011",
  16578=>"010111101",
  16579=>"110100110",
  16580=>"101100000",
  16581=>"100010000",
  16582=>"100110101",
  16583=>"010001100",
  16584=>"110101011",
  16585=>"010010110",
  16586=>"000100000",
  16587=>"011010011",
  16588=>"010111100",
  16589=>"110100111",
  16590=>"100000000",
  16591=>"011011010",
  16592=>"011100010",
  16593=>"010010001",
  16594=>"010001101",
  16595=>"011111011",
  16596=>"101001111",
  16597=>"010101101",
  16598=>"100011111",
  16599=>"111001000",
  16600=>"110110111",
  16601=>"001010101",
  16602=>"101011010",
  16603=>"100000110",
  16604=>"001110001",
  16605=>"100100001",
  16606=>"001001111",
  16607=>"111011111",
  16608=>"101110100",
  16609=>"011011100",
  16610=>"101000100",
  16611=>"101000001",
  16612=>"100101101",
  16613=>"001011111",
  16614=>"001001011",
  16615=>"001111110",
  16616=>"110110100",
  16617=>"010111001",
  16618=>"101100010",
  16619=>"001001101",
  16620=>"101101001",
  16621=>"011100011",
  16622=>"110101100",
  16623=>"100110011",
  16624=>"001110100",
  16625=>"110000000",
  16626=>"110111111",
  16627=>"110001000",
  16628=>"110011001",
  16629=>"001111111",
  16630=>"111011100",
  16631=>"000000000",
  16632=>"011001110",
  16633=>"110001010",
  16634=>"011001100",
  16635=>"000000001",
  16636=>"000000001",
  16637=>"010110100",
  16638=>"100101011",
  16639=>"100010100",
  16640=>"111010000",
  16641=>"000110011",
  16642=>"100111100",
  16643=>"000110110",
  16644=>"000010110",
  16645=>"110110100",
  16646=>"101111101",
  16647=>"001110010",
  16648=>"000000110",
  16649=>"100000100",
  16650=>"000001000",
  16651=>"001010000",
  16652=>"101001111",
  16653=>"000011000",
  16654=>"101011011",
  16655=>"001101001",
  16656=>"010110100",
  16657=>"000001000",
  16658=>"011101111",
  16659=>"101101111",
  16660=>"101100000",
  16661=>"001111111",
  16662=>"001011111",
  16663=>"001101100",
  16664=>"111111100",
  16665=>"101001000",
  16666=>"101111011",
  16667=>"000001000",
  16668=>"101100110",
  16669=>"110111100",
  16670=>"000010010",
  16671=>"101000000",
  16672=>"011111010",
  16673=>"010101100",
  16674=>"100101110",
  16675=>"100010000",
  16676=>"111111001",
  16677=>"000011111",
  16678=>"000011101",
  16679=>"110010011",
  16680=>"111001111",
  16681=>"000011101",
  16682=>"000001000",
  16683=>"111011101",
  16684=>"100000110",
  16685=>"111101101",
  16686=>"000100101",
  16687=>"111111111",
  16688=>"010111101",
  16689=>"010001111",
  16690=>"000000101",
  16691=>"101010111",
  16692=>"000001011",
  16693=>"000010010",
  16694=>"011110001",
  16695=>"110100100",
  16696=>"100110111",
  16697=>"111101110",
  16698=>"000010001",
  16699=>"101010001",
  16700=>"011010000",
  16701=>"010000111",
  16702=>"000010001",
  16703=>"010101000",
  16704=>"011110101",
  16705=>"000101011",
  16706=>"011011111",
  16707=>"100110011",
  16708=>"110111011",
  16709=>"110000000",
  16710=>"111000010",
  16711=>"101100011",
  16712=>"001000110",
  16713=>"101101111",
  16714=>"101100110",
  16715=>"100110110",
  16716=>"110000000",
  16717=>"110011011",
  16718=>"001001000",
  16719=>"110000010",
  16720=>"111011010",
  16721=>"111110000",
  16722=>"011110011",
  16723=>"000110011",
  16724=>"101101101",
  16725=>"000110111",
  16726=>"111001110",
  16727=>"000011111",
  16728=>"000011111",
  16729=>"000110100",
  16730=>"000110011",
  16731=>"111100100",
  16732=>"100000000",
  16733=>"111001011",
  16734=>"000000110",
  16735=>"010100110",
  16736=>"001110000",
  16737=>"111011111",
  16738=>"111001100",
  16739=>"001000110",
  16740=>"000110000",
  16741=>"101111000",
  16742=>"000011011",
  16743=>"011001001",
  16744=>"101101111",
  16745=>"001101001",
  16746=>"100101010",
  16747=>"101010010",
  16748=>"000010010",
  16749=>"001010111",
  16750=>"101001010",
  16751=>"011001011",
  16752=>"000101111",
  16753=>"111000011",
  16754=>"101100001",
  16755=>"111001000",
  16756=>"110011000",
  16757=>"101011111",
  16758=>"010101110",
  16759=>"001100100",
  16760=>"100111011",
  16761=>"111010001",
  16762=>"110110000",
  16763=>"100111001",
  16764=>"111100011",
  16765=>"100010111",
  16766=>"101010110",
  16767=>"100000100",
  16768=>"010001111",
  16769=>"000110100",
  16770=>"111101000",
  16771=>"111011110",
  16772=>"011111111",
  16773=>"101100101",
  16774=>"110101101",
  16775=>"011010001",
  16776=>"010011011",
  16777=>"011000101",
  16778=>"001011111",
  16779=>"101001000",
  16780=>"111010001",
  16781=>"001111101",
  16782=>"110110001",
  16783=>"010100011",
  16784=>"000000000",
  16785=>"101010111",
  16786=>"010011111",
  16787=>"001110011",
  16788=>"100111100",
  16789=>"010001010",
  16790=>"100001000",
  16791=>"111011000",
  16792=>"001011011",
  16793=>"000011110",
  16794=>"001010111",
  16795=>"001100011",
  16796=>"111101011",
  16797=>"011001011",
  16798=>"111101100",
  16799=>"100100111",
  16800=>"100000110",
  16801=>"010000001",
  16802=>"011011010",
  16803=>"101110000",
  16804=>"000101110",
  16805=>"010110011",
  16806=>"000001011",
  16807=>"100110000",
  16808=>"101010001",
  16809=>"011000011",
  16810=>"000101111",
  16811=>"101001101",
  16812=>"011010011",
  16813=>"001111000",
  16814=>"001101100",
  16815=>"000000011",
  16816=>"111000001",
  16817=>"010010011",
  16818=>"000000101",
  16819=>"100111001",
  16820=>"100111010",
  16821=>"111111100",
  16822=>"011111101",
  16823=>"111110111",
  16824=>"011101000",
  16825=>"001001010",
  16826=>"011000100",
  16827=>"011100000",
  16828=>"010110000",
  16829=>"000001111",
  16830=>"011010110",
  16831=>"001000100",
  16832=>"011010100",
  16833=>"111011110",
  16834=>"111110101",
  16835=>"000101001",
  16836=>"001111101",
  16837=>"010100000",
  16838=>"110110101",
  16839=>"000000010",
  16840=>"100011100",
  16841=>"110100011",
  16842=>"100001001",
  16843=>"001100000",
  16844=>"001110111",
  16845=>"100110000",
  16846=>"101010010",
  16847=>"011011110",
  16848=>"110110000",
  16849=>"001001010",
  16850=>"011000100",
  16851=>"101001110",
  16852=>"010011101",
  16853=>"100010010",
  16854=>"111101010",
  16855=>"011010000",
  16856=>"010111010",
  16857=>"011000011",
  16858=>"001000100",
  16859=>"110011010",
  16860=>"010000100",
  16861=>"110000011",
  16862=>"010011111",
  16863=>"110110110",
  16864=>"000110101",
  16865=>"101110101",
  16866=>"011001001",
  16867=>"100111100",
  16868=>"111110111",
  16869=>"011100011",
  16870=>"101010001",
  16871=>"001001000",
  16872=>"011011110",
  16873=>"001011110",
  16874=>"100100000",
  16875=>"001110010",
  16876=>"100110000",
  16877=>"110010001",
  16878=>"110010100",
  16879=>"011000000",
  16880=>"110100111",
  16881=>"010010010",
  16882=>"111010011",
  16883=>"101110101",
  16884=>"000100000",
  16885=>"101010101",
  16886=>"100111000",
  16887=>"101001101",
  16888=>"001000111",
  16889=>"101101100",
  16890=>"111100010",
  16891=>"001101111",
  16892=>"111100111",
  16893=>"010101100",
  16894=>"001011010",
  16895=>"011000000",
  16896=>"000111100",
  16897=>"101100010",
  16898=>"011001011",
  16899=>"000100110",
  16900=>"111001010",
  16901=>"101000001",
  16902=>"101110100",
  16903=>"000001101",
  16904=>"111111011",
  16905=>"100011001",
  16906=>"000101101",
  16907=>"101001111",
  16908=>"101011000",
  16909=>"001101001",
  16910=>"011011111",
  16911=>"011101101",
  16912=>"011100101",
  16913=>"111101110",
  16914=>"110001100",
  16915=>"111001001",
  16916=>"010100100",
  16917=>"101011000",
  16918=>"000010010",
  16919=>"111100100",
  16920=>"010101111",
  16921=>"111101011",
  16922=>"010100000",
  16923=>"000100101",
  16924=>"000010100",
  16925=>"011010101",
  16926=>"101101000",
  16927=>"001100000",
  16928=>"111111111",
  16929=>"000110111",
  16930=>"110001101",
  16931=>"011001000",
  16932=>"100101100",
  16933=>"110100010",
  16934=>"001000110",
  16935=>"011001011",
  16936=>"001101110",
  16937=>"101000100",
  16938=>"101011111",
  16939=>"101111011",
  16940=>"011110011",
  16941=>"001100010",
  16942=>"010000010",
  16943=>"001000111",
  16944=>"100001000",
  16945=>"111110101",
  16946=>"000000011",
  16947=>"100000101",
  16948=>"110101001",
  16949=>"001101011",
  16950=>"101010110",
  16951=>"101101011",
  16952=>"110100110",
  16953=>"000010111",
  16954=>"110111111",
  16955=>"000000000",
  16956=>"010100101",
  16957=>"000000001",
  16958=>"110111010",
  16959=>"100100100",
  16960=>"001001001",
  16961=>"010011111",
  16962=>"011001001",
  16963=>"001000111",
  16964=>"001001000",
  16965=>"010111000",
  16966=>"100110101",
  16967=>"000001111",
  16968=>"101000010",
  16969=>"000011110",
  16970=>"101101110",
  16971=>"001011101",
  16972=>"100100000",
  16973=>"101110111",
  16974=>"001010100",
  16975=>"100001001",
  16976=>"101111001",
  16977=>"011110111",
  16978=>"110010010",
  16979=>"011001100",
  16980=>"011110110",
  16981=>"010110001",
  16982=>"011101000",
  16983=>"000111110",
  16984=>"101000000",
  16985=>"001010101",
  16986=>"111100111",
  16987=>"010101000",
  16988=>"111001111",
  16989=>"000100110",
  16990=>"100111101",
  16991=>"001000101",
  16992=>"110111111",
  16993=>"010110100",
  16994=>"010001111",
  16995=>"000101101",
  16996=>"111000111",
  16997=>"010001000",
  16998=>"001100000",
  16999=>"111000101",
  17000=>"010010000",
  17001=>"011110111",
  17002=>"111000111",
  17003=>"010100001",
  17004=>"101100110",
  17005=>"101010101",
  17006=>"001111001",
  17007=>"001110110",
  17008=>"000000000",
  17009=>"110101010",
  17010=>"010101101",
  17011=>"011000110",
  17012=>"001011111",
  17013=>"010000100",
  17014=>"010010111",
  17015=>"000111011",
  17016=>"110000100",
  17017=>"001111111",
  17018=>"100110010",
  17019=>"000001101",
  17020=>"100000001",
  17021=>"110101110",
  17022=>"000000000",
  17023=>"111010101",
  17024=>"011011111",
  17025=>"011111101",
  17026=>"011101111",
  17027=>"101000111",
  17028=>"111010101",
  17029=>"111001011",
  17030=>"010100101",
  17031=>"001110101",
  17032=>"001001010",
  17033=>"111001101",
  17034=>"111100001",
  17035=>"110001001",
  17036=>"000000010",
  17037=>"000010110",
  17038=>"010000010",
  17039=>"010101100",
  17040=>"011000010",
  17041=>"001111001",
  17042=>"010010111",
  17043=>"101110111",
  17044=>"001001001",
  17045=>"001110010",
  17046=>"111100100",
  17047=>"001101000",
  17048=>"010111010",
  17049=>"000010011",
  17050=>"100100101",
  17051=>"000110101",
  17052=>"011001011",
  17053=>"110011001",
  17054=>"111010001",
  17055=>"000000000",
  17056=>"111011111",
  17057=>"001110110",
  17058=>"000001110",
  17059=>"110010111",
  17060=>"001101001",
  17061=>"101111100",
  17062=>"010010110",
  17063=>"011111100",
  17064=>"111011111",
  17065=>"001000011",
  17066=>"000100010",
  17067=>"001010110",
  17068=>"101000110",
  17069=>"000001111",
  17070=>"000011110",
  17071=>"010110001",
  17072=>"101010110",
  17073=>"001110011",
  17074=>"101001011",
  17075=>"001011111",
  17076=>"101010011",
  17077=>"111010110",
  17078=>"110000111",
  17079=>"101000001",
  17080=>"001010010",
  17081=>"111001001",
  17082=>"000001001",
  17083=>"000001101",
  17084=>"000100000",
  17085=>"101101011",
  17086=>"110101001",
  17087=>"110101110",
  17088=>"000001010",
  17089=>"001011000",
  17090=>"011011000",
  17091=>"001101110",
  17092=>"000000001",
  17093=>"111001101",
  17094=>"111100000",
  17095=>"000001101",
  17096=>"100111000",
  17097=>"100010100",
  17098=>"111000110",
  17099=>"110000000",
  17100=>"111111111",
  17101=>"011101110",
  17102=>"010011011",
  17103=>"101011110",
  17104=>"101110111",
  17105=>"111010110",
  17106=>"100110010",
  17107=>"100011111",
  17108=>"010001100",
  17109=>"000000101",
  17110=>"111010010",
  17111=>"111011100",
  17112=>"011100011",
  17113=>"111100001",
  17114=>"001011011",
  17115=>"011001000",
  17116=>"001100001",
  17117=>"000000000",
  17118=>"101001010",
  17119=>"100101100",
  17120=>"110111000",
  17121=>"111001100",
  17122=>"101101010",
  17123=>"110010100",
  17124=>"000011011",
  17125=>"010000000",
  17126=>"100100000",
  17127=>"001111101",
  17128=>"111101110",
  17129=>"011101000",
  17130=>"111100101",
  17131=>"101111011",
  17132=>"010010110",
  17133=>"001111010",
  17134=>"100111001",
  17135=>"111011111",
  17136=>"110000001",
  17137=>"111111001",
  17138=>"001110100",
  17139=>"110001010",
  17140=>"110100000",
  17141=>"110010000",
  17142=>"110100001",
  17143=>"101110011",
  17144=>"111111010",
  17145=>"110111001",
  17146=>"011000010",
  17147=>"011100100",
  17148=>"100010010",
  17149=>"010111110",
  17150=>"110010011",
  17151=>"100011001",
  17152=>"000011011",
  17153=>"100001101",
  17154=>"000000000",
  17155=>"100001001",
  17156=>"001101000",
  17157=>"110101011",
  17158=>"101100000",
  17159=>"011011110",
  17160=>"110110011",
  17161=>"111111100",
  17162=>"011010010",
  17163=>"010001001",
  17164=>"100100001",
  17165=>"011110101",
  17166=>"001000001",
  17167=>"011001010",
  17168=>"100100110",
  17169=>"001001011",
  17170=>"111100001",
  17171=>"101001010",
  17172=>"101100100",
  17173=>"001001010",
  17174=>"111011011",
  17175=>"001000011",
  17176=>"111101111",
  17177=>"011011100",
  17178=>"101100010",
  17179=>"000101111",
  17180=>"010100001",
  17181=>"101100110",
  17182=>"000000001",
  17183=>"010100000",
  17184=>"011100100",
  17185=>"111010001",
  17186=>"101011000",
  17187=>"010000010",
  17188=>"000010011",
  17189=>"000011010",
  17190=>"101100000",
  17191=>"001111101",
  17192=>"100111110",
  17193=>"000110101",
  17194=>"110001100",
  17195=>"100000110",
  17196=>"111001110",
  17197=>"101101010",
  17198=>"101101110",
  17199=>"000001101",
  17200=>"001000111",
  17201=>"001011111",
  17202=>"000100100",
  17203=>"001000010",
  17204=>"101110011",
  17205=>"000000110",
  17206=>"000010001",
  17207=>"111110000",
  17208=>"010010101",
  17209=>"100001101",
  17210=>"100101101",
  17211=>"000111111",
  17212=>"001100010",
  17213=>"011110111",
  17214=>"100000001",
  17215=>"101100001",
  17216=>"100000101",
  17217=>"011011100",
  17218=>"011111101",
  17219=>"100000101",
  17220=>"100010111",
  17221=>"010110011",
  17222=>"011000010",
  17223=>"101101000",
  17224=>"001010011",
  17225=>"010100101",
  17226=>"111110010",
  17227=>"011101001",
  17228=>"101100001",
  17229=>"110100001",
  17230=>"000110100",
  17231=>"011111110",
  17232=>"110000000",
  17233=>"001000100",
  17234=>"011011111",
  17235=>"001101000",
  17236=>"100000010",
  17237=>"000110011",
  17238=>"111101101",
  17239=>"000011000",
  17240=>"000011111",
  17241=>"111100100",
  17242=>"010111111",
  17243=>"110010000",
  17244=>"111111101",
  17245=>"000101001",
  17246=>"011011011",
  17247=>"000100010",
  17248=>"110111010",
  17249=>"111100101",
  17250=>"101000111",
  17251=>"100101111",
  17252=>"000010000",
  17253=>"000101001",
  17254=>"100011010",
  17255=>"100000001",
  17256=>"011001100",
  17257=>"110101000",
  17258=>"001001000",
  17259=>"001000101",
  17260=>"100111100",
  17261=>"111010000",
  17262=>"000000100",
  17263=>"001011011",
  17264=>"000001001",
  17265=>"001100110",
  17266=>"101010010",
  17267=>"001001010",
  17268=>"010100111",
  17269=>"111001010",
  17270=>"011001100",
  17271=>"101100001",
  17272=>"111100100",
  17273=>"010010011",
  17274=>"101001000",
  17275=>"101110101",
  17276=>"000011011",
  17277=>"100000100",
  17278=>"011001001",
  17279=>"010110100",
  17280=>"110110110",
  17281=>"000111001",
  17282=>"100111111",
  17283=>"000000011",
  17284=>"011111100",
  17285=>"100100010",
  17286=>"001111011",
  17287=>"101111000",
  17288=>"110110000",
  17289=>"010010110",
  17290=>"011110111",
  17291=>"111011011",
  17292=>"100001000",
  17293=>"000110001",
  17294=>"111000100",
  17295=>"110100000",
  17296=>"011001011",
  17297=>"001010011",
  17298=>"000100000",
  17299=>"001101011",
  17300=>"111001111",
  17301=>"010011110",
  17302=>"010001111",
  17303=>"000001100",
  17304=>"101101010",
  17305=>"001011111",
  17306=>"110001011",
  17307=>"000011110",
  17308=>"100000100",
  17309=>"010010100",
  17310=>"101100000",
  17311=>"000110110",
  17312=>"000000101",
  17313=>"111011001",
  17314=>"010110010",
  17315=>"101100111",
  17316=>"100101000",
  17317=>"101110010",
  17318=>"010011001",
  17319=>"100110100",
  17320=>"000100001",
  17321=>"101110000",
  17322=>"100111100",
  17323=>"111000111",
  17324=>"100111100",
  17325=>"010000111",
  17326=>"111111101",
  17327=>"010110110",
  17328=>"111111001",
  17329=>"001111010",
  17330=>"111110000",
  17331=>"100011100",
  17332=>"010011111",
  17333=>"110111000",
  17334=>"111000011",
  17335=>"100010110",
  17336=>"011101001",
  17337=>"000011011",
  17338=>"010001000",
  17339=>"100011000",
  17340=>"110111100",
  17341=>"111000001",
  17342=>"100001011",
  17343=>"010010000",
  17344=>"010010000",
  17345=>"110101110",
  17346=>"011011110",
  17347=>"000000100",
  17348=>"010111101",
  17349=>"000111011",
  17350=>"110011011",
  17351=>"101011010",
  17352=>"001110110",
  17353=>"100010101",
  17354=>"001100100",
  17355=>"000100100",
  17356=>"101101011",
  17357=>"001010010",
  17358=>"000111011",
  17359=>"010101001",
  17360=>"000011010",
  17361=>"001101001",
  17362=>"001110110",
  17363=>"100101110",
  17364=>"011111111",
  17365=>"111110011",
  17366=>"011101011",
  17367=>"101010001",
  17368=>"011111110",
  17369=>"100111010",
  17370=>"101100000",
  17371=>"000010111",
  17372=>"001100111",
  17373=>"000100101",
  17374=>"001000101",
  17375=>"001001001",
  17376=>"010000111",
  17377=>"001001100",
  17378=>"001010101",
  17379=>"111001000",
  17380=>"010001001",
  17381=>"100001011",
  17382=>"000111110",
  17383=>"010000000",
  17384=>"001000111",
  17385=>"000100000",
  17386=>"010001000",
  17387=>"111000101",
  17388=>"011000001",
  17389=>"101001011",
  17390=>"000010001",
  17391=>"101101101",
  17392=>"001101110",
  17393=>"011111001",
  17394=>"001101101",
  17395=>"011111001",
  17396=>"000101111",
  17397=>"011000111",
  17398=>"011000101",
  17399=>"110010010",
  17400=>"000101000",
  17401=>"101010111",
  17402=>"101010100",
  17403=>"001001100",
  17404=>"011100111",
  17405=>"001110100",
  17406=>"110111110",
  17407=>"001000111",
  17408=>"110101100",
  17409=>"110001111",
  17410=>"010010100",
  17411=>"010110000",
  17412=>"010110110",
  17413=>"101101111",
  17414=>"001011111",
  17415=>"000001001",
  17416=>"000110110",
  17417=>"001000110",
  17418=>"001011000",
  17419=>"000010110",
  17420=>"101011001",
  17421=>"100111111",
  17422=>"100101011",
  17423=>"101011111",
  17424=>"010010011",
  17425=>"001110010",
  17426=>"000101100",
  17427=>"111001000",
  17428=>"111111010",
  17429=>"010101101",
  17430=>"111000111",
  17431=>"101001100",
  17432=>"000010100",
  17433=>"101001000",
  17434=>"101011011",
  17435=>"101010001",
  17436=>"011110100",
  17437=>"100110011",
  17438=>"001100000",
  17439=>"111000011",
  17440=>"011001111",
  17441=>"101111101",
  17442=>"000011110",
  17443=>"011100111",
  17444=>"101001101",
  17445=>"110000101",
  17446=>"101101001",
  17447=>"100011100",
  17448=>"100010100",
  17449=>"111101000",
  17450=>"000101001",
  17451=>"000010000",
  17452=>"000111011",
  17453=>"111101001",
  17454=>"100110110",
  17455=>"001011001",
  17456=>"010011111",
  17457=>"001000111",
  17458=>"111111010",
  17459=>"001100011",
  17460=>"101010000",
  17461=>"111100001",
  17462=>"100011111",
  17463=>"011011101",
  17464=>"000010100",
  17465=>"001000110",
  17466=>"011011111",
  17467=>"101000010",
  17468=>"111000101",
  17469=>"110101101",
  17470=>"100111001",
  17471=>"011101001",
  17472=>"111111111",
  17473=>"001100101",
  17474=>"000001110",
  17475=>"100010111",
  17476=>"000110110",
  17477=>"111110010",
  17478=>"100100000",
  17479=>"001100001",
  17480=>"001110011",
  17481=>"011110110",
  17482=>"011101000",
  17483=>"001000110",
  17484=>"011001110",
  17485=>"110011100",
  17486=>"110010001",
  17487=>"010000001",
  17488=>"010111100",
  17489=>"000001001",
  17490=>"101111011",
  17491=>"111001001",
  17492=>"000111111",
  17493=>"100001110",
  17494=>"011011010",
  17495=>"100001101",
  17496=>"111111111",
  17497=>"001011010",
  17498=>"001000110",
  17499=>"000110001",
  17500=>"110001111",
  17501=>"010111011",
  17502=>"000110111",
  17503=>"001101110",
  17504=>"000100001",
  17505=>"101010110",
  17506=>"001001010",
  17507=>"101100010",
  17508=>"100110001",
  17509=>"110010100",
  17510=>"111101100",
  17511=>"011101111",
  17512=>"101111110",
  17513=>"011011110",
  17514=>"100101111",
  17515=>"111001010",
  17516=>"101001110",
  17517=>"011010101",
  17518=>"111110011",
  17519=>"000111000",
  17520=>"110001010",
  17521=>"011000010",
  17522=>"101001011",
  17523=>"000100101",
  17524=>"000110011",
  17525=>"001010010",
  17526=>"011011001",
  17527=>"001100111",
  17528=>"011111100",
  17529=>"100001101",
  17530=>"011001111",
  17531=>"101100000",
  17532=>"100010101",
  17533=>"010000000",
  17534=>"101000111",
  17535=>"011001011",
  17536=>"001110010",
  17537=>"111111111",
  17538=>"110010111",
  17539=>"101011111",
  17540=>"011110111",
  17541=>"101100100",
  17542=>"000111000",
  17543=>"001100000",
  17544=>"111111101",
  17545=>"100100100",
  17546=>"000000001",
  17547=>"111111001",
  17548=>"010010010",
  17549=>"011001111",
  17550=>"111111111",
  17551=>"100000001",
  17552=>"110011001",
  17553=>"011110100",
  17554=>"000001111",
  17555=>"000111011",
  17556=>"100111001",
  17557=>"001000010",
  17558=>"101001001",
  17559=>"101100100",
  17560=>"101011000",
  17561=>"010101000",
  17562=>"001000111",
  17563=>"011010001",
  17564=>"100011101",
  17565=>"110100100",
  17566=>"000000011",
  17567=>"011011101",
  17568=>"111101001",
  17569=>"000100001",
  17570=>"000110111",
  17571=>"000011111",
  17572=>"101001110",
  17573=>"001100110",
  17574=>"101100100",
  17575=>"001000010",
  17576=>"000010011",
  17577=>"010010001",
  17578=>"000111101",
  17579=>"101101010",
  17580=>"101011100",
  17581=>"100110101",
  17582=>"010010100",
  17583=>"110000100",
  17584=>"100111000",
  17585=>"001010011",
  17586=>"110001100",
  17587=>"001011011",
  17588=>"011100001",
  17589=>"100100110",
  17590=>"100100000",
  17591=>"011101011",
  17592=>"100011110",
  17593=>"111000101",
  17594=>"010001010",
  17595=>"101101011",
  17596=>"000001000",
  17597=>"101000000",
  17598=>"000011001",
  17599=>"000001011",
  17600=>"000110001",
  17601=>"101011000",
  17602=>"001111010",
  17603=>"101011101",
  17604=>"001110000",
  17605=>"000000001",
  17606=>"000111001",
  17607=>"001000110",
  17608=>"000001100",
  17609=>"011101111",
  17610=>"011001001",
  17611=>"011101111",
  17612=>"110011001",
  17613=>"001110111",
  17614=>"000000101",
  17615=>"000001000",
  17616=>"011001110",
  17617=>"100011101",
  17618=>"100111110",
  17619=>"001100111",
  17620=>"000111111",
  17621=>"001001010",
  17622=>"000101000",
  17623=>"011110001",
  17624=>"110001001",
  17625=>"010111010",
  17626=>"100111110",
  17627=>"111010000",
  17628=>"011110000",
  17629=>"001010110",
  17630=>"111101110",
  17631=>"000111110",
  17632=>"101011101",
  17633=>"001001010",
  17634=>"111000010",
  17635=>"001101011",
  17636=>"001010110",
  17637=>"100100100",
  17638=>"110011101",
  17639=>"001110011",
  17640=>"111101001",
  17641=>"100011000",
  17642=>"011011101",
  17643=>"110101100",
  17644=>"000001111",
  17645=>"101000100",
  17646=>"101010010",
  17647=>"101111011",
  17648=>"110000001",
  17649=>"100110011",
  17650=>"100101000",
  17651=>"100010110",
  17652=>"101111110",
  17653=>"110101000",
  17654=>"101001110",
  17655=>"100100111",
  17656=>"001100011",
  17657=>"010010100",
  17658=>"010101101",
  17659=>"011000100",
  17660=>"011111001",
  17661=>"001110001",
  17662=>"101000111",
  17663=>"110111111",
  17664=>"110010011",
  17665=>"010110011",
  17666=>"110101101",
  17667=>"010011001",
  17668=>"101000001",
  17669=>"100010000",
  17670=>"110010010",
  17671=>"110100011",
  17672=>"101011101",
  17673=>"011001000",
  17674=>"010010111",
  17675=>"100000001",
  17676=>"100101110",
  17677=>"001111111",
  17678=>"100111101",
  17679=>"000001010",
  17680=>"111000000",
  17681=>"001101011",
  17682=>"100111101",
  17683=>"001100100",
  17684=>"011011000",
  17685=>"011101100",
  17686=>"001110001",
  17687=>"001011111",
  17688=>"110011010",
  17689=>"011101010",
  17690=>"001111110",
  17691=>"001001011",
  17692=>"001010100",
  17693=>"000110011",
  17694=>"010101001",
  17695=>"010100010",
  17696=>"000111111",
  17697=>"010101011",
  17698=>"101111001",
  17699=>"111000001",
  17700=>"101000000",
  17701=>"000100111",
  17702=>"011010011",
  17703=>"101111000",
  17704=>"110010010",
  17705=>"110001001",
  17706=>"011111101",
  17707=>"101111011",
  17708=>"101111001",
  17709=>"010111000",
  17710=>"010110010",
  17711=>"111001001",
  17712=>"101101101",
  17713=>"010110010",
  17714=>"101111000",
  17715=>"101101001",
  17716=>"101011111",
  17717=>"010101111",
  17718=>"111110000",
  17719=>"011111111",
  17720=>"011101101",
  17721=>"110011001",
  17722=>"001110011",
  17723=>"101111101",
  17724=>"000011110",
  17725=>"000111001",
  17726=>"110101000",
  17727=>"101111110",
  17728=>"100010101",
  17729=>"100000110",
  17730=>"000001100",
  17731=>"000001101",
  17732=>"010101010",
  17733=>"111101111",
  17734=>"010100010",
  17735=>"111011100",
  17736=>"111100100",
  17737=>"010100010",
  17738=>"110011000",
  17739=>"001011101",
  17740=>"100001000",
  17741=>"000110111",
  17742=>"110110001",
  17743=>"100110010",
  17744=>"000011001",
  17745=>"000010010",
  17746=>"010011010",
  17747=>"111111101",
  17748=>"001000011",
  17749=>"100110000",
  17750=>"011111011",
  17751=>"111000010",
  17752=>"010000100",
  17753=>"011000011",
  17754=>"010010100",
  17755=>"000011000",
  17756=>"101111111",
  17757=>"000010110",
  17758=>"000011011",
  17759=>"000110011",
  17760=>"101101100",
  17761=>"011000000",
  17762=>"000110101",
  17763=>"011111000",
  17764=>"000100101",
  17765=>"110001010",
  17766=>"011011101",
  17767=>"110110100",
  17768=>"111011011",
  17769=>"111000100",
  17770=>"000000000",
  17771=>"111000100",
  17772=>"100001000",
  17773=>"011011101",
  17774=>"010001101",
  17775=>"000111101",
  17776=>"100111101",
  17777=>"000001010",
  17778=>"110100110",
  17779=>"011010000",
  17780=>"110001100",
  17781=>"010111110",
  17782=>"000101010",
  17783=>"101111100",
  17784=>"000111000",
  17785=>"000001101",
  17786=>"111011100",
  17787=>"110111001",
  17788=>"000000111",
  17789=>"101010110",
  17790=>"011011111",
  17791=>"000011000",
  17792=>"101010111",
  17793=>"101000011",
  17794=>"100101111",
  17795=>"101111011",
  17796=>"001001100",
  17797=>"101101010",
  17798=>"110100111",
  17799=>"100001100",
  17800=>"011010010",
  17801=>"000100000",
  17802=>"010000110",
  17803=>"001110001",
  17804=>"110001011",
  17805=>"001101100",
  17806=>"101001011",
  17807=>"100011100",
  17808=>"000110000",
  17809=>"000000000",
  17810=>"100001011",
  17811=>"111110111",
  17812=>"000100100",
  17813=>"001110101",
  17814=>"010000100",
  17815=>"111111100",
  17816=>"000101010",
  17817=>"001000101",
  17818=>"111001111",
  17819=>"110000000",
  17820=>"011100001",
  17821=>"001100100",
  17822=>"110010110",
  17823=>"001101001",
  17824=>"110010010",
  17825=>"010000101",
  17826=>"011011101",
  17827=>"001001000",
  17828=>"100011100",
  17829=>"100100000",
  17830=>"110111101",
  17831=>"011000001",
  17832=>"000110100",
  17833=>"010000110",
  17834=>"011100111",
  17835=>"100010000",
  17836=>"001000000",
  17837=>"011100101",
  17838=>"011101100",
  17839=>"001001100",
  17840=>"101101111",
  17841=>"010111011",
  17842=>"000010011",
  17843=>"010010000",
  17844=>"000001111",
  17845=>"011000010",
  17846=>"110001111",
  17847=>"011100101",
  17848=>"010100110",
  17849=>"011011001",
  17850=>"011110111",
  17851=>"101001100",
  17852=>"000110000",
  17853=>"000101011",
  17854=>"110010111",
  17855=>"001101010",
  17856=>"110110000",
  17857=>"010101110",
  17858=>"010111001",
  17859=>"111000001",
  17860=>"000000001",
  17861=>"001000100",
  17862=>"000000101",
  17863=>"000001110",
  17864=>"101100010",
  17865=>"111111010",
  17866=>"111011010",
  17867=>"000000011",
  17868=>"001110011",
  17869=>"111000100",
  17870=>"011111100",
  17871=>"000010110",
  17872=>"010011011",
  17873=>"000011010",
  17874=>"111111111",
  17875=>"010101100",
  17876=>"101110110",
  17877=>"011111011",
  17878=>"011100000",
  17879=>"101111100",
  17880=>"010000110",
  17881=>"010000101",
  17882=>"101111011",
  17883=>"011111110",
  17884=>"000100101",
  17885=>"011111011",
  17886=>"011000110",
  17887=>"110000110",
  17888=>"111000000",
  17889=>"011111111",
  17890=>"010000000",
  17891=>"110000001",
  17892=>"101100000",
  17893=>"010010100",
  17894=>"011111110",
  17895=>"011001000",
  17896=>"010101001",
  17897=>"000110101",
  17898=>"011111000",
  17899=>"001010010",
  17900=>"111001110",
  17901=>"100110100",
  17902=>"010010100",
  17903=>"010101110",
  17904=>"011100101",
  17905=>"011010000",
  17906=>"101101101",
  17907=>"110000110",
  17908=>"011110010",
  17909=>"100010111",
  17910=>"011001001",
  17911=>"111010100",
  17912=>"010101011",
  17913=>"100110111",
  17914=>"001010111",
  17915=>"010101010",
  17916=>"110111101",
  17917=>"110110000",
  17918=>"011000001",
  17919=>"110010111",
  17920=>"010111011",
  17921=>"011001011",
  17922=>"110110111",
  17923=>"001011011",
  17924=>"111001000",
  17925=>"110100110",
  17926=>"110010110",
  17927=>"110011101",
  17928=>"100100011",
  17929=>"000101111",
  17930=>"011101100",
  17931=>"100001011",
  17932=>"000111111",
  17933=>"111100011",
  17934=>"110000001",
  17935=>"001101011",
  17936=>"010100110",
  17937=>"100010010",
  17938=>"111111001",
  17939=>"100011110",
  17940=>"001010101",
  17941=>"111110001",
  17942=>"101000111",
  17943=>"000101010",
  17944=>"011010000",
  17945=>"100011100",
  17946=>"001110001",
  17947=>"111000010",
  17948=>"100010010",
  17949=>"011111000",
  17950=>"111010001",
  17951=>"111001100",
  17952=>"010101001",
  17953=>"110110110",
  17954=>"100001000",
  17955=>"110000111",
  17956=>"111011110",
  17957=>"101100011",
  17958=>"011011101",
  17959=>"111100100",
  17960=>"001011011",
  17961=>"011011110",
  17962=>"111101000",
  17963=>"111101101",
  17964=>"110100101",
  17965=>"101111001",
  17966=>"111110110",
  17967=>"011001011",
  17968=>"111001010",
  17969=>"101111111",
  17970=>"100011110",
  17971=>"100011111",
  17972=>"000111101",
  17973=>"110011011",
  17974=>"011001001",
  17975=>"111001100",
  17976=>"100110011",
  17977=>"000110000",
  17978=>"111001110",
  17979=>"110100100",
  17980=>"001100011",
  17981=>"001100001",
  17982=>"001011111",
  17983=>"011010100",
  17984=>"101111111",
  17985=>"000000111",
  17986=>"100101101",
  17987=>"101000110",
  17988=>"001101100",
  17989=>"001110010",
  17990=>"101010010",
  17991=>"100111101",
  17992=>"010101001",
  17993=>"100000010",
  17994=>"011010111",
  17995=>"000110111",
  17996=>"110011110",
  17997=>"011001011",
  17998=>"000100101",
  17999=>"110000111",
  18000=>"110110010",
  18001=>"111101111",
  18002=>"110100101",
  18003=>"001110000",
  18004=>"110100111",
  18005=>"011000100",
  18006=>"101101100",
  18007=>"101011010",
  18008=>"001010000",
  18009=>"011110000",
  18010=>"101101101",
  18011=>"100101111",
  18012=>"001101011",
  18013=>"000100000",
  18014=>"101011101",
  18015=>"001111100",
  18016=>"111000011",
  18017=>"101101011",
  18018=>"101110111",
  18019=>"111101101",
  18020=>"110001101",
  18021=>"110111000",
  18022=>"100011100",
  18023=>"010111010",
  18024=>"110010111",
  18025=>"000110011",
  18026=>"110100010",
  18027=>"000001010",
  18028=>"010100011",
  18029=>"101000010",
  18030=>"000100001",
  18031=>"000000100",
  18032=>"100110110",
  18033=>"110001100",
  18034=>"000000111",
  18035=>"001100101",
  18036=>"011101111",
  18037=>"111100100",
  18038=>"101100011",
  18039=>"100110001",
  18040=>"101110110",
  18041=>"101101111",
  18042=>"011010101",
  18043=>"011100111",
  18044=>"100010100",
  18045=>"001001111",
  18046=>"111010110",
  18047=>"100111100",
  18048=>"011101100",
  18049=>"001111111",
  18050=>"011110000",
  18051=>"110100110",
  18052=>"101111111",
  18053=>"000000010",
  18054=>"011011111",
  18055=>"000111010",
  18056=>"001101111",
  18057=>"111101100",
  18058=>"000010000",
  18059=>"101100000",
  18060=>"101101010",
  18061=>"111111110",
  18062=>"001011010",
  18063=>"010111101",
  18064=>"010110011",
  18065=>"100101111",
  18066=>"000110011",
  18067=>"100111001",
  18068=>"000110011",
  18069=>"111100111",
  18070=>"111101100",
  18071=>"111010111",
  18072=>"000010011",
  18073=>"000000101",
  18074=>"110111000",
  18075=>"010010100",
  18076=>"001110010",
  18077=>"111000101",
  18078=>"001110000",
  18079=>"101000101",
  18080=>"110001100",
  18081=>"100101101",
  18082=>"110100011",
  18083=>"000101001",
  18084=>"001001001",
  18085=>"000110101",
  18086=>"110011101",
  18087=>"000100101",
  18088=>"110110110",
  18089=>"111000101",
  18090=>"010111011",
  18091=>"000100011",
  18092=>"011100100",
  18093=>"111100010",
  18094=>"101001001",
  18095=>"001011101",
  18096=>"111011001",
  18097=>"101100010",
  18098=>"111111000",
  18099=>"101000100",
  18100=>"111000110",
  18101=>"100001111",
  18102=>"000110110",
  18103=>"010001111",
  18104=>"111010010",
  18105=>"010000000",
  18106=>"010101101",
  18107=>"000001100",
  18108=>"011010100",
  18109=>"001001011",
  18110=>"011100000",
  18111=>"001100010",
  18112=>"110110010",
  18113=>"000000100",
  18114=>"101001110",
  18115=>"110111001",
  18116=>"001111011",
  18117=>"110010110",
  18118=>"100001000",
  18119=>"011110011",
  18120=>"101111110",
  18121=>"110001000",
  18122=>"111110001",
  18123=>"101010110",
  18124=>"011111111",
  18125=>"110110001",
  18126=>"010011110",
  18127=>"110001000",
  18128=>"001011101",
  18129=>"110110110",
  18130=>"000001110",
  18131=>"011001000",
  18132=>"011100101",
  18133=>"011101100",
  18134=>"111010101",
  18135=>"001011101",
  18136=>"100100100",
  18137=>"010111011",
  18138=>"100011011",
  18139=>"010010111",
  18140=>"000010100",
  18141=>"111100111",
  18142=>"011001011",
  18143=>"101011100",
  18144=>"010110000",
  18145=>"111110100",
  18146=>"101111001",
  18147=>"101011100",
  18148=>"111110110",
  18149=>"010111000",
  18150=>"111001100",
  18151=>"000110010",
  18152=>"001111000",
  18153=>"101000001",
  18154=>"100011100",
  18155=>"000111111",
  18156=>"000100011",
  18157=>"110111000",
  18158=>"101000011",
  18159=>"100111101",
  18160=>"000000100",
  18161=>"000110001",
  18162=>"100001111",
  18163=>"111100010",
  18164=>"100111100",
  18165=>"011101010",
  18166=>"000000111",
  18167=>"011001110",
  18168=>"011110100",
  18169=>"110111101",
  18170=>"011000011",
  18171=>"001110010",
  18172=>"001010000",
  18173=>"000001100",
  18174=>"010101110",
  18175=>"001110111",
  18176=>"101101010",
  18177=>"001100101",
  18178=>"101100110",
  18179=>"001000110",
  18180=>"000001010",
  18181=>"111100101",
  18182=>"000101101",
  18183=>"011000010",
  18184=>"110000111",
  18185=>"111101110",
  18186=>"101011011",
  18187=>"001111110",
  18188=>"011011001",
  18189=>"001110010",
  18190=>"111110101",
  18191=>"101001011",
  18192=>"101110100",
  18193=>"101100100",
  18194=>"000101010",
  18195=>"010100101",
  18196=>"110000110",
  18197=>"101110001",
  18198=>"010110101",
  18199=>"001010001",
  18200=>"110111111",
  18201=>"001111010",
  18202=>"010111011",
  18203=>"111000000",
  18204=>"111111110",
  18205=>"110101100",
  18206=>"011101101",
  18207=>"011001101",
  18208=>"100110011",
  18209=>"111010000",
  18210=>"110100101",
  18211=>"001111001",
  18212=>"011010101",
  18213=>"000110000",
  18214=>"010110110",
  18215=>"011000001",
  18216=>"001101001",
  18217=>"000100000",
  18218=>"111100011",
  18219=>"011011110",
  18220=>"110001110",
  18221=>"000001010",
  18222=>"101100101",
  18223=>"111111101",
  18224=>"001001110",
  18225=>"110100001",
  18226=>"101011000",
  18227=>"101011000",
  18228=>"000011110",
  18229=>"001011000",
  18230=>"100010000",
  18231=>"110010000",
  18232=>"001101001",
  18233=>"111010001",
  18234=>"100001000",
  18235=>"111101010",
  18236=>"011011000",
  18237=>"001101000",
  18238=>"101001110",
  18239=>"111110111",
  18240=>"011111011",
  18241=>"000011011",
  18242=>"111101000",
  18243=>"000000000",
  18244=>"101111101",
  18245=>"001000101",
  18246=>"000110001",
  18247=>"001000011",
  18248=>"011101111",
  18249=>"100111011",
  18250=>"011001101",
  18251=>"001110101",
  18252=>"000000011",
  18253=>"100010110",
  18254=>"111111011",
  18255=>"110010000",
  18256=>"110010111",
  18257=>"111100011",
  18258=>"001100001",
  18259=>"111000111",
  18260=>"110101000",
  18261=>"011010110",
  18262=>"101111100",
  18263=>"010111000",
  18264=>"100111110",
  18265=>"010111001",
  18266=>"001101111",
  18267=>"000100010",
  18268=>"110000111",
  18269=>"000100010",
  18270=>"111101101",
  18271=>"000100000",
  18272=>"000010001",
  18273=>"101000101",
  18274=>"001010110",
  18275=>"101110011",
  18276=>"110001110",
  18277=>"010001100",
  18278=>"100000001",
  18279=>"001010101",
  18280=>"000000100",
  18281=>"000111110",
  18282=>"111110100",
  18283=>"110000111",
  18284=>"100101111",
  18285=>"111010110",
  18286=>"100100011",
  18287=>"000000000",
  18288=>"100100001",
  18289=>"010011101",
  18290=>"000110111",
  18291=>"111011101",
  18292=>"101011110",
  18293=>"001101101",
  18294=>"000001100",
  18295=>"010000000",
  18296=>"001000111",
  18297=>"111011001",
  18298=>"010001011",
  18299=>"110110100",
  18300=>"000001011",
  18301=>"101001010",
  18302=>"011010110",
  18303=>"101011010",
  18304=>"010110101",
  18305=>"111111010",
  18306=>"100110001",
  18307=>"101011110",
  18308=>"000010101",
  18309=>"111001011",
  18310=>"100101010",
  18311=>"000001111",
  18312=>"001100111",
  18313=>"010000001",
  18314=>"010111101",
  18315=>"010011010",
  18316=>"100110001",
  18317=>"011000111",
  18318=>"111011101",
  18319=>"101110110",
  18320=>"111000011",
  18321=>"111110111",
  18322=>"111001011",
  18323=>"000011100",
  18324=>"001100111",
  18325=>"101110101",
  18326=>"001110100",
  18327=>"111010001",
  18328=>"001001001",
  18329=>"010101011",
  18330=>"011101001",
  18331=>"101010111",
  18332=>"011001001",
  18333=>"100100000",
  18334=>"101000001",
  18335=>"001011101",
  18336=>"110011100",
  18337=>"110000100",
  18338=>"011101101",
  18339=>"000011001",
  18340=>"101100100",
  18341=>"001100001",
  18342=>"000010010",
  18343=>"001111001",
  18344=>"100101111",
  18345=>"000011111",
  18346=>"100001100",
  18347=>"110101100",
  18348=>"110110100",
  18349=>"011001010",
  18350=>"011101111",
  18351=>"101100110",
  18352=>"010010111",
  18353=>"100011110",
  18354=>"011101101",
  18355=>"101000101",
  18356=>"101101100",
  18357=>"100000101",
  18358=>"111011000",
  18359=>"110111001",
  18360=>"100000000",
  18361=>"101011000",
  18362=>"010110110",
  18363=>"101000011",
  18364=>"001110110",
  18365=>"010001101",
  18366=>"000011011",
  18367=>"101101001",
  18368=>"110111010",
  18369=>"100111101",
  18370=>"101011100",
  18371=>"110011010",
  18372=>"010010100",
  18373=>"110000000",
  18374=>"101011110",
  18375=>"101100011",
  18376=>"111100010",
  18377=>"111011100",
  18378=>"010010011",
  18379=>"011010110",
  18380=>"010111110",
  18381=>"100000000",
  18382=>"101111010",
  18383=>"001100000",
  18384=>"101100011",
  18385=>"010110111",
  18386=>"010001010",
  18387=>"100000000",
  18388=>"000010011",
  18389=>"100110000",
  18390=>"100001101",
  18391=>"101011110",
  18392=>"000011110",
  18393=>"110111111",
  18394=>"000101001",
  18395=>"010001111",
  18396=>"000001100",
  18397=>"110100101",
  18398=>"101101011",
  18399=>"110011000",
  18400=>"000010000",
  18401=>"100011010",
  18402=>"011100010",
  18403=>"001001010",
  18404=>"000111000",
  18405=>"101111010",
  18406=>"000001110",
  18407=>"101111001",
  18408=>"001010000",
  18409=>"000010011",
  18410=>"110100000",
  18411=>"001101111",
  18412=>"000101010",
  18413=>"010010000",
  18414=>"010001110",
  18415=>"101111101",
  18416=>"000110111",
  18417=>"000110111",
  18418=>"001001000",
  18419=>"010111100",
  18420=>"110111001",
  18421=>"011001110",
  18422=>"100100001",
  18423=>"110011100",
  18424=>"011000110",
  18425=>"000010111",
  18426=>"101101010",
  18427=>"101100111",
  18428=>"001111101",
  18429=>"011111101",
  18430=>"010110101",
  18431=>"110110011",
  18432=>"101101111",
  18433=>"010000111",
  18434=>"010110101",
  18435=>"000000101",
  18436=>"101010100",
  18437=>"111100111",
  18438=>"111100000",
  18439=>"111010111",
  18440=>"110101011",
  18441=>"011101101",
  18442=>"100001100",
  18443=>"100100110",
  18444=>"110111100",
  18445=>"000011101",
  18446=>"011111010",
  18447=>"000101001",
  18448=>"010000110",
  18449=>"010000101",
  18450=>"111100110",
  18451=>"101000111",
  18452=>"111010011",
  18453=>"000000100",
  18454=>"110010101",
  18455=>"001100011",
  18456=>"011100010",
  18457=>"011110110",
  18458=>"010111010",
  18459=>"111111010",
  18460=>"011101010",
  18461=>"001000000",
  18462=>"011000100",
  18463=>"111111101",
  18464=>"110010001",
  18465=>"111010010",
  18466=>"011110011",
  18467=>"100001010",
  18468=>"010001111",
  18469=>"011101010",
  18470=>"100010111",
  18471=>"001000000",
  18472=>"000100111",
  18473=>"100010110",
  18474=>"000000100",
  18475=>"000100101",
  18476=>"010111110",
  18477=>"001111110",
  18478=>"111011000",
  18479=>"000000110",
  18480=>"010111000",
  18481=>"011010111",
  18482=>"101110110",
  18483=>"110111101",
  18484=>"011001110",
  18485=>"100110011",
  18486=>"111110100",
  18487=>"111000001",
  18488=>"110011001",
  18489=>"010001001",
  18490=>"001011111",
  18491=>"011001001",
  18492=>"010100001",
  18493=>"101011011",
  18494=>"010100100",
  18495=>"111111111",
  18496=>"110001100",
  18497=>"100011100",
  18498=>"000000100",
  18499=>"111001011",
  18500=>"100001000",
  18501=>"011000100",
  18502=>"100000110",
  18503=>"001010010",
  18504=>"000100000",
  18505=>"011011111",
  18506=>"000110010",
  18507=>"000000111",
  18508=>"111000110",
  18509=>"111111100",
  18510=>"001111110",
  18511=>"011101100",
  18512=>"001010100",
  18513=>"101110001",
  18514=>"111000111",
  18515=>"110111110",
  18516=>"110001110",
  18517=>"010010010",
  18518=>"100001100",
  18519=>"000000010",
  18520=>"011110101",
  18521=>"000011111",
  18522=>"001001110",
  18523=>"100010100",
  18524=>"100000100",
  18525=>"010001001",
  18526=>"101001000",
  18527=>"101001110",
  18528=>"011011101",
  18529=>"110101011",
  18530=>"100011001",
  18531=>"011011100",
  18532=>"010101011",
  18533=>"111111100",
  18534=>"011010110",
  18535=>"110110010",
  18536=>"111110011",
  18537=>"110001100",
  18538=>"100011001",
  18539=>"111001110",
  18540=>"101111111",
  18541=>"111101001",
  18542=>"110100011",
  18543=>"101001100",
  18544=>"000011000",
  18545=>"000100101",
  18546=>"111010111",
  18547=>"001101011",
  18548=>"011110001",
  18549=>"101110001",
  18550=>"100011101",
  18551=>"101010001",
  18552=>"100010000",
  18553=>"001111110",
  18554=>"010111100",
  18555=>"001100001",
  18556=>"011110011",
  18557=>"000010110",
  18558=>"110111011",
  18559=>"010111100",
  18560=>"111010000",
  18561=>"101101010",
  18562=>"111110101",
  18563=>"000011001",
  18564=>"010110101",
  18565=>"000011000",
  18566=>"011001001",
  18567=>"000000010",
  18568=>"110110101",
  18569=>"000110000",
  18570=>"001010111",
  18571=>"000010000",
  18572=>"011010111",
  18573=>"100011110",
  18574=>"001101001",
  18575=>"010001000",
  18576=>"010000001",
  18577=>"100111101",
  18578=>"100110000",
  18579=>"101000101",
  18580=>"100101000",
  18581=>"111111001",
  18582=>"001001101",
  18583=>"101010110",
  18584=>"010110000",
  18585=>"000011001",
  18586=>"010010000",
  18587=>"000111011",
  18588=>"100111001",
  18589=>"100101000",
  18590=>"000011011",
  18591=>"101001100",
  18592=>"111000100",
  18593=>"101110010",
  18594=>"011111000",
  18595=>"001110010",
  18596=>"111001101",
  18597=>"011010110",
  18598=>"100110000",
  18599=>"010000110",
  18600=>"111111010",
  18601=>"011011001",
  18602=>"011101110",
  18603=>"110001011",
  18604=>"101101011",
  18605=>"011110101",
  18606=>"000111100",
  18607=>"100110011",
  18608=>"101000110",
  18609=>"001101011",
  18610=>"111101011",
  18611=>"110010010",
  18612=>"110010110",
  18613=>"111111011",
  18614=>"011100110",
  18615=>"011000100",
  18616=>"001000000",
  18617=>"111111100",
  18618=>"001001110",
  18619=>"001011101",
  18620=>"111110111",
  18621=>"000001001",
  18622=>"100110011",
  18623=>"000001000",
  18624=>"010000110",
  18625=>"111100001",
  18626=>"011010010",
  18627=>"000110111",
  18628=>"000101111",
  18629=>"001001101",
  18630=>"110001110",
  18631=>"110010001",
  18632=>"001111110",
  18633=>"010110110",
  18634=>"111111000",
  18635=>"110101110",
  18636=>"001001100",
  18637=>"110101111",
  18638=>"011010100",
  18639=>"010000001",
  18640=>"100001010",
  18641=>"110101100",
  18642=>"111111101",
  18643=>"000001011",
  18644=>"000110111",
  18645=>"101111111",
  18646=>"011010100",
  18647=>"010010111",
  18648=>"101001001",
  18649=>"111000010",
  18650=>"000111110",
  18651=>"100101001",
  18652=>"010000000",
  18653=>"100110101",
  18654=>"001001010",
  18655=>"000001010",
  18656=>"110111101",
  18657=>"001010110",
  18658=>"101100101",
  18659=>"100110111",
  18660=>"000000010",
  18661=>"011001001",
  18662=>"111100111",
  18663=>"000110100",
  18664=>"001001010",
  18665=>"111110111",
  18666=>"001110010",
  18667=>"100110110",
  18668=>"011010110",
  18669=>"111010010",
  18670=>"110011100",
  18671=>"110000000",
  18672=>"011111101",
  18673=>"000010001",
  18674=>"010000110",
  18675=>"110100110",
  18676=>"110010000",
  18677=>"101101110",
  18678=>"001101000",
  18679=>"111001000",
  18680=>"011000001",
  18681=>"100100100",
  18682=>"101111111",
  18683=>"001100111",
  18684=>"111011100",
  18685=>"101111111",
  18686=>"101000110",
  18687=>"000111100",
  18688=>"111111001",
  18689=>"110000011",
  18690=>"010111010",
  18691=>"000100000",
  18692=>"000001010",
  18693=>"111000000",
  18694=>"000010000",
  18695=>"010111100",
  18696=>"101010101",
  18697=>"010001000",
  18698=>"001110000",
  18699=>"110111010",
  18700=>"111110101",
  18701=>"001111000",
  18702=>"000110011",
  18703=>"000000110",
  18704=>"011011110",
  18705=>"110100010",
  18706=>"011001100",
  18707=>"000011111",
  18708=>"110101000",
  18709=>"100001110",
  18710=>"001111111",
  18711=>"110100101",
  18712=>"101111100",
  18713=>"110000010",
  18714=>"101100111",
  18715=>"001100100",
  18716=>"000111100",
  18717=>"101000111",
  18718=>"100111110",
  18719=>"101111011",
  18720=>"100111101",
  18721=>"010111101",
  18722=>"010110001",
  18723=>"100010110",
  18724=>"000010001",
  18725=>"011101110",
  18726=>"111010011",
  18727=>"010011100",
  18728=>"000000111",
  18729=>"111000010",
  18730=>"110001101",
  18731=>"011101000",
  18732=>"100011111",
  18733=>"011000010",
  18734=>"011110001",
  18735=>"001100111",
  18736=>"101011101",
  18737=>"010011111",
  18738=>"011100111",
  18739=>"110110100",
  18740=>"100011010",
  18741=>"101001001",
  18742=>"100000101",
  18743=>"110110111",
  18744=>"001101100",
  18745=>"010011111",
  18746=>"100100101",
  18747=>"001011011",
  18748=>"100111001",
  18749=>"111101100",
  18750=>"110100001",
  18751=>"111001111",
  18752=>"001111100",
  18753=>"100110000",
  18754=>"010001111",
  18755=>"111000001",
  18756=>"110001001",
  18757=>"100101011",
  18758=>"000000100",
  18759=>"011111011",
  18760=>"001011110",
  18761=>"011010110",
  18762=>"111011010",
  18763=>"100101110",
  18764=>"111001100",
  18765=>"000011001",
  18766=>"111011110",
  18767=>"000111111",
  18768=>"010000110",
  18769=>"110011000",
  18770=>"011000011",
  18771=>"011100101",
  18772=>"010001111",
  18773=>"011011000",
  18774=>"110111111",
  18775=>"110111110",
  18776=>"111001111",
  18777=>"001110110",
  18778=>"011000001",
  18779=>"110110100",
  18780=>"011000011",
  18781=>"000100001",
  18782=>"111011100",
  18783=>"100011010",
  18784=>"001110111",
  18785=>"101111011",
  18786=>"110010011",
  18787=>"111111011",
  18788=>"010110100",
  18789=>"110101100",
  18790=>"110101011",
  18791=>"110101100",
  18792=>"001100111",
  18793=>"111101111",
  18794=>"100010001",
  18795=>"101111011",
  18796=>"010001111",
  18797=>"111110000",
  18798=>"101111001",
  18799=>"011100001",
  18800=>"100010001",
  18801=>"111101110",
  18802=>"001111001",
  18803=>"001111001",
  18804=>"010110111",
  18805=>"000111001",
  18806=>"111001011",
  18807=>"000110001",
  18808=>"110100010",
  18809=>"100011001",
  18810=>"001001001",
  18811=>"011001000",
  18812=>"100110100",
  18813=>"110101100",
  18814=>"111000000",
  18815=>"100011011",
  18816=>"111101100",
  18817=>"011101001",
  18818=>"001100100",
  18819=>"110001011",
  18820=>"101011101",
  18821=>"000111001",
  18822=>"100111011",
  18823=>"111111100",
  18824=>"011011010",
  18825=>"101100101",
  18826=>"000000000",
  18827=>"010000010",
  18828=>"111110001",
  18829=>"011011111",
  18830=>"001001110",
  18831=>"100010000",
  18832=>"011111000",
  18833=>"011111100",
  18834=>"100100100",
  18835=>"001110000",
  18836=>"110110110",
  18837=>"111001000",
  18838=>"101111100",
  18839=>"011001001",
  18840=>"001000110",
  18841=>"101110001",
  18842=>"100101001",
  18843=>"000101101",
  18844=>"110110011",
  18845=>"000100000",
  18846=>"010110111",
  18847=>"001011110",
  18848=>"100101100",
  18849=>"001100000",
  18850=>"010001110",
  18851=>"000110100",
  18852=>"100001100",
  18853=>"100110010",
  18854=>"110000100",
  18855=>"101110001",
  18856=>"011110100",
  18857=>"010111101",
  18858=>"100000100",
  18859=>"100011000",
  18860=>"101100010",
  18861=>"100101100",
  18862=>"101011011",
  18863=>"001110110",
  18864=>"110111011",
  18865=>"110010001",
  18866=>"001011000",
  18867=>"101111000",
  18868=>"000001001",
  18869=>"110011001",
  18870=>"110100000",
  18871=>"111101000",
  18872=>"110100101",
  18873=>"111011011",
  18874=>"101100100",
  18875=>"101100101",
  18876=>"000010010",
  18877=>"001011001",
  18878=>"000000011",
  18879=>"001111001",
  18880=>"111011010",
  18881=>"110101101",
  18882=>"001100011",
  18883=>"010111100",
  18884=>"001001100",
  18885=>"100101001",
  18886=>"010010001",
  18887=>"011000101",
  18888=>"111001011",
  18889=>"100111100",
  18890=>"010111110",
  18891=>"011110110",
  18892=>"000000011",
  18893=>"001100100",
  18894=>"100100000",
  18895=>"110000000",
  18896=>"100001010",
  18897=>"111111101",
  18898=>"111101111",
  18899=>"001100000",
  18900=>"110011110",
  18901=>"110010011",
  18902=>"110101001",
  18903=>"100010010",
  18904=>"111000101",
  18905=>"101000111",
  18906=>"100010010",
  18907=>"010111110",
  18908=>"101110100",
  18909=>"010000001",
  18910=>"001000110",
  18911=>"000100000",
  18912=>"110010101",
  18913=>"101110101",
  18914=>"010011000",
  18915=>"101110000",
  18916=>"110111010",
  18917=>"100000111",
  18918=>"110000100",
  18919=>"111001011",
  18920=>"101001111",
  18921=>"100100000",
  18922=>"001000111",
  18923=>"110110011",
  18924=>"000100111",
  18925=>"101010110",
  18926=>"011111010",
  18927=>"100011101",
  18928=>"100000000",
  18929=>"101111000",
  18930=>"101010011",
  18931=>"100010100",
  18932=>"011001010",
  18933=>"011010011",
  18934=>"101011101",
  18935=>"110001101",
  18936=>"100010000",
  18937=>"010000110",
  18938=>"101101001",
  18939=>"111000011",
  18940=>"011110111",
  18941=>"011111000",
  18942=>"110100111",
  18943=>"010000000",
  18944=>"110100011",
  18945=>"000011111",
  18946=>"111000101",
  18947=>"001001111",
  18948=>"111001000",
  18949=>"111100000",
  18950=>"001100010",
  18951=>"100110100",
  18952=>"001001001",
  18953=>"000101101",
  18954=>"110000110",
  18955=>"100001010",
  18956=>"111111000",
  18957=>"100001010",
  18958=>"111100000",
  18959=>"000001110",
  18960=>"010010100",
  18961=>"000110001",
  18962=>"111010000",
  18963=>"011101110",
  18964=>"011101011",
  18965=>"000000000",
  18966=>"000010000",
  18967=>"000001010",
  18968=>"000100010",
  18969=>"111000111",
  18970=>"001100010",
  18971=>"010000011",
  18972=>"101000101",
  18973=>"010000001",
  18974=>"000100110",
  18975=>"000110011",
  18976=>"001101101",
  18977=>"111100101",
  18978=>"110010000",
  18979=>"111010010",
  18980=>"100101110",
  18981=>"110100010",
  18982=>"001010000",
  18983=>"101000011",
  18984=>"011010101",
  18985=>"100111000",
  18986=>"101101101",
  18987=>"001100011",
  18988=>"000110001",
  18989=>"101000111",
  18990=>"111110111",
  18991=>"010000000",
  18992=>"110011010",
  18993=>"111011110",
  18994=>"000111110",
  18995=>"010000111",
  18996=>"011110110",
  18997=>"111100100",
  18998=>"110111110",
  18999=>"101011001",
  19000=>"101100100",
  19001=>"110100101",
  19002=>"111101111",
  19003=>"110000000",
  19004=>"010110101",
  19005=>"000100001",
  19006=>"011111111",
  19007=>"100011101",
  19008=>"101101101",
  19009=>"011111010",
  19010=>"001000001",
  19011=>"110010111",
  19012=>"001101101",
  19013=>"000010001",
  19014=>"111001101",
  19015=>"000101100",
  19016=>"000001011",
  19017=>"101010011",
  19018=>"010010000",
  19019=>"001101100",
  19020=>"110010011",
  19021=>"101000110",
  19022=>"101101011",
  19023=>"100001000",
  19024=>"110000010",
  19025=>"111101010",
  19026=>"111110100",
  19027=>"101011100",
  19028=>"001101111",
  19029=>"001011110",
  19030=>"000101110",
  19031=>"001000000",
  19032=>"100100010",
  19033=>"000111100",
  19034=>"111011000",
  19035=>"110001000",
  19036=>"111010101",
  19037=>"100111011",
  19038=>"110001110",
  19039=>"000101101",
  19040=>"111100010",
  19041=>"111110011",
  19042=>"111100110",
  19043=>"101001000",
  19044=>"001001111",
  19045=>"010010100",
  19046=>"010000011",
  19047=>"111000100",
  19048=>"100010111",
  19049=>"010011001",
  19050=>"111000001",
  19051=>"000101100",
  19052=>"100101111",
  19053=>"111110010",
  19054=>"101011101",
  19055=>"110000001",
  19056=>"100011000",
  19057=>"010100101",
  19058=>"111100111",
  19059=>"010110100",
  19060=>"101110111",
  19061=>"001111001",
  19062=>"101100101",
  19063=>"100101101",
  19064=>"010100010",
  19065=>"100111000",
  19066=>"001110100",
  19067=>"010110111",
  19068=>"000000110",
  19069=>"000111101",
  19070=>"110101011",
  19071=>"111111011",
  19072=>"011111010",
  19073=>"001111111",
  19074=>"101110001",
  19075=>"111100001",
  19076=>"011111101",
  19077=>"010110100",
  19078=>"101010110",
  19079=>"110111000",
  19080=>"101111000",
  19081=>"110101110",
  19082=>"010111101",
  19083=>"000101001",
  19084=>"010110100",
  19085=>"110011111",
  19086=>"001000000",
  19087=>"011000001",
  19088=>"010101001",
  19089=>"110110011",
  19090=>"001101101",
  19091=>"010010010",
  19092=>"000111001",
  19093=>"000000101",
  19094=>"111001100",
  19095=>"101001000",
  19096=>"000111111",
  19097=>"011101111",
  19098=>"011110100",
  19099=>"010001111",
  19100=>"111100100",
  19101=>"110000001",
  19102=>"010010000",
  19103=>"110010110",
  19104=>"110000101",
  19105=>"101010110",
  19106=>"011111000",
  19107=>"010111110",
  19108=>"111001111",
  19109=>"010110110",
  19110=>"110000001",
  19111=>"011000111",
  19112=>"110010110",
  19113=>"001011101",
  19114=>"110110111",
  19115=>"110001001",
  19116=>"100101110",
  19117=>"000001010",
  19118=>"001111010",
  19119=>"011101001",
  19120=>"111001001",
  19121=>"101001001",
  19122=>"111110010",
  19123=>"111101001",
  19124=>"111101010",
  19125=>"111100011",
  19126=>"000110000",
  19127=>"001101010",
  19128=>"011111000",
  19129=>"111111011",
  19130=>"011111100",
  19131=>"111010000",
  19132=>"110101101",
  19133=>"000001100",
  19134=>"101101000",
  19135=>"111101101",
  19136=>"101110101",
  19137=>"100001011",
  19138=>"101010100",
  19139=>"011001011",
  19140=>"000111101",
  19141=>"100001100",
  19142=>"100011000",
  19143=>"001111011",
  19144=>"000111001",
  19145=>"100011100",
  19146=>"000001000",
  19147=>"110111100",
  19148=>"011111001",
  19149=>"111100000",
  19150=>"011111100",
  19151=>"001100001",
  19152=>"010101101",
  19153=>"110110111",
  19154=>"000011111",
  19155=>"011101000",
  19156=>"000001000",
  19157=>"010000111",
  19158=>"000000101",
  19159=>"001100111",
  19160=>"111001001",
  19161=>"110101001",
  19162=>"110000110",
  19163=>"010101011",
  19164=>"000011000",
  19165=>"110100001",
  19166=>"010000011",
  19167=>"101101111",
  19168=>"110111010",
  19169=>"010100000",
  19170=>"100000100",
  19171=>"001101000",
  19172=>"001010100",
  19173=>"011001000",
  19174=>"100010100",
  19175=>"000011110",
  19176=>"010111000",
  19177=>"011001100",
  19178=>"010101000",
  19179=>"000101100",
  19180=>"000111000",
  19181=>"000100000",
  19182=>"100011001",
  19183=>"111111000",
  19184=>"110001000",
  19185=>"101110011",
  19186=>"101111110",
  19187=>"111110111",
  19188=>"000101011",
  19189=>"001101101",
  19190=>"010000100",
  19191=>"100001001",
  19192=>"001111000",
  19193=>"001111111",
  19194=>"001111100",
  19195=>"011111010",
  19196=>"001001000",
  19197=>"101001111",
  19198=>"101011001",
  19199=>"011110000",
  19200=>"001011000",
  19201=>"001010111",
  19202=>"011011101",
  19203=>"111010000",
  19204=>"100010110",
  19205=>"000001000",
  19206=>"011100010",
  19207=>"111011111",
  19208=>"001110110",
  19209=>"101101000",
  19210=>"111111000",
  19211=>"110001000",
  19212=>"000010101",
  19213=>"011000001",
  19214=>"100010000",
  19215=>"011001100",
  19216=>"011101111",
  19217=>"111111001",
  19218=>"000000111",
  19219=>"011111001",
  19220=>"110010011",
  19221=>"010011000",
  19222=>"100011000",
  19223=>"111101111",
  19224=>"101101100",
  19225=>"111100010",
  19226=>"000001110",
  19227=>"001101100",
  19228=>"001110001",
  19229=>"110111000",
  19230=>"100101100",
  19231=>"010111110",
  19232=>"110001001",
  19233=>"000100001",
  19234=>"110010001",
  19235=>"111010011",
  19236=>"011110011",
  19237=>"010111011",
  19238=>"001001001",
  19239=>"111010010",
  19240=>"111011001",
  19241=>"000111100",
  19242=>"111101011",
  19243=>"000011001",
  19244=>"010110011",
  19245=>"000000100",
  19246=>"101011101",
  19247=>"100000001",
  19248=>"101100011",
  19249=>"100111000",
  19250=>"110111000",
  19251=>"010001010",
  19252=>"000111101",
  19253=>"011010000",
  19254=>"011000010",
  19255=>"110100001",
  19256=>"110011000",
  19257=>"111100001",
  19258=>"010110110",
  19259=>"001010100",
  19260=>"100011000",
  19261=>"010000010",
  19262=>"101010111",
  19263=>"101110001",
  19264=>"100110101",
  19265=>"110001100",
  19266=>"100010010",
  19267=>"110111001",
  19268=>"101101100",
  19269=>"011101100",
  19270=>"010101101",
  19271=>"101011011",
  19272=>"011001100",
  19273=>"101001010",
  19274=>"000111100",
  19275=>"000101110",
  19276=>"010100101",
  19277=>"110110000",
  19278=>"101010000",
  19279=>"001001110",
  19280=>"100000100",
  19281=>"001100110",
  19282=>"001111111",
  19283=>"101100010",
  19284=>"111110111",
  19285=>"110101111",
  19286=>"011111010",
  19287=>"100001100",
  19288=>"010111001",
  19289=>"110110111",
  19290=>"101110100",
  19291=>"010101100",
  19292=>"101101001",
  19293=>"111000000",
  19294=>"000000000",
  19295=>"001011100",
  19296=>"011001010",
  19297=>"010011000",
  19298=>"000110001",
  19299=>"011000000",
  19300=>"111011101",
  19301=>"001010011",
  19302=>"011011101",
  19303=>"000001001",
  19304=>"011000000",
  19305=>"011000010",
  19306=>"100101011",
  19307=>"101100111",
  19308=>"101111101",
  19309=>"101101000",
  19310=>"100110111",
  19311=>"101110000",
  19312=>"010011001",
  19313=>"111110000",
  19314=>"111101111",
  19315=>"101101000",
  19316=>"101101000",
  19317=>"111110001",
  19318=>"001100011",
  19319=>"101111000",
  19320=>"010000000",
  19321=>"110000010",
  19322=>"000110010",
  19323=>"000000010",
  19324=>"000111000",
  19325=>"000100110",
  19326=>"100110111",
  19327=>"110111010",
  19328=>"111001101",
  19329=>"000000001",
  19330=>"111011100",
  19331=>"010101010",
  19332=>"111000010",
  19333=>"100110001",
  19334=>"001110101",
  19335=>"101000101",
  19336=>"100001110",
  19337=>"111011010",
  19338=>"100101010",
  19339=>"100111010",
  19340=>"010100010",
  19341=>"111000001",
  19342=>"111111110",
  19343=>"101110011",
  19344=>"101111110",
  19345=>"110111001",
  19346=>"100101110",
  19347=>"110000000",
  19348=>"010011101",
  19349=>"110000110",
  19350=>"000000111",
  19351=>"100000011",
  19352=>"100011011",
  19353=>"100001111",
  19354=>"100001100",
  19355=>"011100110",
  19356=>"000011110",
  19357=>"101011100",
  19358=>"000000001",
  19359=>"101111111",
  19360=>"111111011",
  19361=>"000000101",
  19362=>"101111000",
  19363=>"000111000",
  19364=>"001000000",
  19365=>"111010110",
  19366=>"001100100",
  19367=>"111001000",
  19368=>"011100000",
  19369=>"110000110",
  19370=>"011010010",
  19371=>"110000110",
  19372=>"100010010",
  19373=>"011110001",
  19374=>"101101101",
  19375=>"010011111",
  19376=>"110000110",
  19377=>"101101011",
  19378=>"110011100",
  19379=>"110111000",
  19380=>"110110110",
  19381=>"010000010",
  19382=>"010100100",
  19383=>"110100110",
  19384=>"101111111",
  19385=>"111101011",
  19386=>"010001101",
  19387=>"100101000",
  19388=>"101110010",
  19389=>"010101101",
  19390=>"010110000",
  19391=>"001001111",
  19392=>"101101101",
  19393=>"000010000",
  19394=>"011011000",
  19395=>"111000010",
  19396=>"101110111",
  19397=>"010000110",
  19398=>"110111101",
  19399=>"000101011",
  19400=>"110010010",
  19401=>"010101011",
  19402=>"001100000",
  19403=>"011110101",
  19404=>"011101101",
  19405=>"110111100",
  19406=>"110011100",
  19407=>"101101100",
  19408=>"001111101",
  19409=>"000011100",
  19410=>"101001101",
  19411=>"110100000",
  19412=>"111001011",
  19413=>"110001111",
  19414=>"000101001",
  19415=>"011111110",
  19416=>"100111100",
  19417=>"011000111",
  19418=>"001010001",
  19419=>"001011111",
  19420=>"011001000",
  19421=>"011100111",
  19422=>"110110001",
  19423=>"011100100",
  19424=>"110100010",
  19425=>"111010101",
  19426=>"111011101",
  19427=>"001100100",
  19428=>"000101011",
  19429=>"000010000",
  19430=>"101000000",
  19431=>"000001110",
  19432=>"011101101",
  19433=>"001000010",
  19434=>"011010000",
  19435=>"100110110",
  19436=>"001000010",
  19437=>"100001101",
  19438=>"100001000",
  19439=>"000111100",
  19440=>"011000000",
  19441=>"001010001",
  19442=>"010100001",
  19443=>"111011111",
  19444=>"100000000",
  19445=>"010001011",
  19446=>"110011011",
  19447=>"000100001",
  19448=>"110100011",
  19449=>"110100101",
  19450=>"101111001",
  19451=>"000000011",
  19452=>"110011111",
  19453=>"110000111",
  19454=>"010001111",
  19455=>"001101001",
  19456=>"110001110",
  19457=>"010010011",
  19458=>"111101100",
  19459=>"100101100",
  19460=>"100100101",
  19461=>"101001001",
  19462=>"111110000",
  19463=>"111110100",
  19464=>"101001010",
  19465=>"100010100",
  19466=>"000001100",
  19467=>"001110000",
  19468=>"001010100",
  19469=>"000000010",
  19470=>"000101111",
  19471=>"111000110",
  19472=>"000001111",
  19473=>"111001001",
  19474=>"110010010",
  19475=>"101110111",
  19476=>"100100000",
  19477=>"111010001",
  19478=>"101010111",
  19479=>"001100111",
  19480=>"111001111",
  19481=>"111111011",
  19482=>"010010100",
  19483=>"010101110",
  19484=>"110000100",
  19485=>"100011111",
  19486=>"111010011",
  19487=>"110111000",
  19488=>"111011011",
  19489=>"100100000",
  19490=>"001000000",
  19491=>"010000101",
  19492=>"110011011",
  19493=>"110100110",
  19494=>"110110001",
  19495=>"000111010",
  19496=>"101111110",
  19497=>"001000110",
  19498=>"011001110",
  19499=>"110111100",
  19500=>"000100100",
  19501=>"000100000",
  19502=>"011101100",
  19503=>"001111001",
  19504=>"010111100",
  19505=>"010010001",
  19506=>"101001100",
  19507=>"111001010",
  19508=>"010011100",
  19509=>"101001001",
  19510=>"000111011",
  19511=>"101010100",
  19512=>"000101011",
  19513=>"000100111",
  19514=>"101101011",
  19515=>"101101010",
  19516=>"110000110",
  19517=>"010100110",
  19518=>"101101100",
  19519=>"001101111",
  19520=>"100001100",
  19521=>"011111111",
  19522=>"111100110",
  19523=>"011100000",
  19524=>"010000100",
  19525=>"100001110",
  19526=>"000011010",
  19527=>"001001000",
  19528=>"101100000",
  19529=>"000001010",
  19530=>"000100010",
  19531=>"011100100",
  19532=>"100100011",
  19533=>"110000011",
  19534=>"001100001",
  19535=>"010010101",
  19536=>"001101001",
  19537=>"101011000",
  19538=>"100110101",
  19539=>"101000000",
  19540=>"000101010",
  19541=>"011101111",
  19542=>"010100100",
  19543=>"111111010",
  19544=>"101011101",
  19545=>"101100101",
  19546=>"110001111",
  19547=>"111010101",
  19548=>"010000000",
  19549=>"000011101",
  19550=>"001011110",
  19551=>"100100101",
  19552=>"110001011",
  19553=>"101001010",
  19554=>"011110010",
  19555=>"101101110",
  19556=>"011001101",
  19557=>"100010111",
  19558=>"000110000",
  19559=>"000011100",
  19560=>"110010110",
  19561=>"111111101",
  19562=>"100010010",
  19563=>"010000111",
  19564=>"101000111",
  19565=>"100001011",
  19566=>"101100011",
  19567=>"000001101",
  19568=>"100000111",
  19569=>"010000001",
  19570=>"000111011",
  19571=>"010100011",
  19572=>"111100101",
  19573=>"000000001",
  19574=>"111111100",
  19575=>"110111001",
  19576=>"101111110",
  19577=>"101110001",
  19578=>"000010011",
  19579=>"000100010",
  19580=>"100100000",
  19581=>"011011000",
  19582=>"100011001",
  19583=>"001000000",
  19584=>"010001011",
  19585=>"011101111",
  19586=>"101100011",
  19587=>"011100011",
  19588=>"101000001",
  19589=>"001101011",
  19590=>"100100010",
  19591=>"110010000",
  19592=>"100111001",
  19593=>"011001010",
  19594=>"100001111",
  19595=>"110010010",
  19596=>"001000100",
  19597=>"110111101",
  19598=>"111101111",
  19599=>"010110000",
  19600=>"011101001",
  19601=>"101100111",
  19602=>"010111001",
  19603=>"111011111",
  19604=>"101000100",
  19605=>"010101110",
  19606=>"101110111",
  19607=>"111110111",
  19608=>"110001010",
  19609=>"101000111",
  19610=>"111110111",
  19611=>"101101001",
  19612=>"011011010",
  19613=>"011010100",
  19614=>"101100100",
  19615=>"111010111",
  19616=>"111101101",
  19617=>"110011111",
  19618=>"101000110",
  19619=>"011001010",
  19620=>"100000000",
  19621=>"001111100",
  19622=>"011000001",
  19623=>"100110001",
  19624=>"111111001",
  19625=>"000000110",
  19626=>"000000000",
  19627=>"111010010",
  19628=>"111000101",
  19629=>"100100101",
  19630=>"010110000",
  19631=>"111101111",
  19632=>"001011000",
  19633=>"000010100",
  19634=>"001010110",
  19635=>"010100101",
  19636=>"011001011",
  19637=>"011010000",
  19638=>"010101001",
  19639=>"010001010",
  19640=>"110001011",
  19641=>"101101101",
  19642=>"100111111",
  19643=>"101110010",
  19644=>"010101100",
  19645=>"110110000",
  19646=>"010000100",
  19647=>"011011111",
  19648=>"011001110",
  19649=>"110000001",
  19650=>"100001100",
  19651=>"101001001",
  19652=>"010010100",
  19653=>"100001000",
  19654=>"011101110",
  19655=>"011110100",
  19656=>"011010001",
  19657=>"100100110",
  19658=>"000100000",
  19659=>"000100010",
  19660=>"011001110",
  19661=>"101110011",
  19662=>"100100010",
  19663=>"111100110",
  19664=>"111101001",
  19665=>"100100100",
  19666=>"111011000",
  19667=>"000011001",
  19668=>"110001001",
  19669=>"110111110",
  19670=>"110101110",
  19671=>"010011100",
  19672=>"010000001",
  19673=>"000010110",
  19674=>"010100111",
  19675=>"001101011",
  19676=>"010110100",
  19677=>"110011110",
  19678=>"111100111",
  19679=>"011010011",
  19680=>"000100111",
  19681=>"000101110",
  19682=>"111111111",
  19683=>"010001100",
  19684=>"110001101",
  19685=>"100101110",
  19686=>"100001100",
  19687=>"100001010",
  19688=>"111101101",
  19689=>"100000001",
  19690=>"110000000",
  19691=>"000101010",
  19692=>"000001001",
  19693=>"000101110",
  19694=>"100010010",
  19695=>"101100000",
  19696=>"011100011",
  19697=>"000001101",
  19698=>"100001001",
  19699=>"110010110",
  19700=>"001100110",
  19701=>"111110011",
  19702=>"001010100",
  19703=>"101000000",
  19704=>"000011001",
  19705=>"111001100",
  19706=>"001000001",
  19707=>"000110000",
  19708=>"011100110",
  19709=>"100011100",
  19710=>"010111011",
  19711=>"111111011",
  19712=>"110111111",
  19713=>"111110011",
  19714=>"000111100",
  19715=>"001111100",
  19716=>"000110110",
  19717=>"101100110",
  19718=>"001010100",
  19719=>"110100110",
  19720=>"001001011",
  19721=>"011110110",
  19722=>"011110110",
  19723=>"110110110",
  19724=>"000000000",
  19725=>"101001111",
  19726=>"100000001",
  19727=>"010011101",
  19728=>"111001100",
  19729=>"100011001",
  19730=>"000010111",
  19731=>"001100001",
  19732=>"011000001",
  19733=>"010000110",
  19734=>"101000000",
  19735=>"001101110",
  19736=>"111110111",
  19737=>"010000011",
  19738=>"110000101",
  19739=>"111110001",
  19740=>"001110111",
  19741=>"000000011",
  19742=>"111101011",
  19743=>"000001100",
  19744=>"000100010",
  19745=>"111011010",
  19746=>"011101101",
  19747=>"000101101",
  19748=>"010000000",
  19749=>"110111100",
  19750=>"100000100",
  19751=>"011010111",
  19752=>"111010011",
  19753=>"000000100",
  19754=>"011001100",
  19755=>"110000010",
  19756=>"011010000",
  19757=>"101000100",
  19758=>"001101010",
  19759=>"010100011",
  19760=>"010111111",
  19761=>"001110100",
  19762=>"010010110",
  19763=>"101111000",
  19764=>"101000001",
  19765=>"100111001",
  19766=>"000001001",
  19767=>"001010001",
  19768=>"000001100",
  19769=>"101001111",
  19770=>"011001001",
  19771=>"010011001",
  19772=>"111001100",
  19773=>"110000010",
  19774=>"011000000",
  19775=>"100000000",
  19776=>"011001000",
  19777=>"011111111",
  19778=>"111010100",
  19779=>"101100100",
  19780=>"011010100",
  19781=>"010010101",
  19782=>"011111110",
  19783=>"100010110",
  19784=>"010000100",
  19785=>"000000000",
  19786=>"001001110",
  19787=>"101100000",
  19788=>"111000111",
  19789=>"010011101",
  19790=>"110011100",
  19791=>"010111011",
  19792=>"101000110",
  19793=>"010001010",
  19794=>"011000111",
  19795=>"000010100",
  19796=>"101011010",
  19797=>"000110110",
  19798=>"101000101",
  19799=>"000001000",
  19800=>"100111111",
  19801=>"101001111",
  19802=>"010000001",
  19803=>"001000001",
  19804=>"101101001",
  19805=>"000000000",
  19806=>"110011100",
  19807=>"000000101",
  19808=>"110110111",
  19809=>"101011101",
  19810=>"000101110",
  19811=>"001010101",
  19812=>"111011011",
  19813=>"001100100",
  19814=>"101010111",
  19815=>"000011100",
  19816=>"010011100",
  19817=>"100000011",
  19818=>"000010010",
  19819=>"001111110",
  19820=>"010011001",
  19821=>"110011110",
  19822=>"000101011",
  19823=>"101010100",
  19824=>"000011101",
  19825=>"011001111",
  19826=>"100001001",
  19827=>"100110000",
  19828=>"000100010",
  19829=>"011110100",
  19830=>"001011111",
  19831=>"110010010",
  19832=>"000101100",
  19833=>"110000110",
  19834=>"101101100",
  19835=>"110100010",
  19836=>"110011010",
  19837=>"111100111",
  19838=>"001011111",
  19839=>"111111110",
  19840=>"010111010",
  19841=>"101001010",
  19842=>"100100111",
  19843=>"000000111",
  19844=>"111111010",
  19845=>"001000111",
  19846=>"111011111",
  19847=>"100010001",
  19848=>"111010000",
  19849=>"101111001",
  19850=>"010100110",
  19851=>"111111111",
  19852=>"010000001",
  19853=>"010111110",
  19854=>"001101110",
  19855=>"000000000",
  19856=>"011010010",
  19857=>"000001010",
  19858=>"101010110",
  19859=>"010101100",
  19860=>"011010100",
  19861=>"001111000",
  19862=>"101001001",
  19863=>"010110011",
  19864=>"101100111",
  19865=>"000110010",
  19866=>"000010101",
  19867=>"111110100",
  19868=>"111000011",
  19869=>"101010101",
  19870=>"111101100",
  19871=>"110010001",
  19872=>"010001011",
  19873=>"001000010",
  19874=>"111101010",
  19875=>"100001010",
  19876=>"010100110",
  19877=>"000001000",
  19878=>"000000100",
  19879=>"100000001",
  19880=>"101101011",
  19881=>"010010000",
  19882=>"110110011",
  19883=>"100010010",
  19884=>"010110101",
  19885=>"011111000",
  19886=>"000010000",
  19887=>"001001101",
  19888=>"011111010",
  19889=>"001111111",
  19890=>"011010101",
  19891=>"100001110",
  19892=>"110011100",
  19893=>"101011010",
  19894=>"101011111",
  19895=>"011010011",
  19896=>"110000101",
  19897=>"000111111",
  19898=>"000000001",
  19899=>"110111111",
  19900=>"110001000",
  19901=>"011101101",
  19902=>"011111010",
  19903=>"101001011",
  19904=>"001000011",
  19905=>"110010011",
  19906=>"011001011",
  19907=>"111011000",
  19908=>"001111001",
  19909=>"110111110",
  19910=>"101111001",
  19911=>"000000100",
  19912=>"100001110",
  19913=>"000101110",
  19914=>"001100000",
  19915=>"101010000",
  19916=>"110000101",
  19917=>"011111010",
  19918=>"100011111",
  19919=>"111011000",
  19920=>"110011000",
  19921=>"111100000",
  19922=>"100010001",
  19923=>"111101010",
  19924=>"111011011",
  19925=>"000100110",
  19926=>"000100101",
  19927=>"000111100",
  19928=>"101100111",
  19929=>"010000011",
  19930=>"111001111",
  19931=>"001011001",
  19932=>"011101011",
  19933=>"111111001",
  19934=>"011111001",
  19935=>"010011001",
  19936=>"010110101",
  19937=>"011011111",
  19938=>"001100010",
  19939=>"111110011",
  19940=>"000011111",
  19941=>"000111111",
  19942=>"011000100",
  19943=>"000001001",
  19944=>"000111001",
  19945=>"110110001",
  19946=>"010000101",
  19947=>"010011111",
  19948=>"010011001",
  19949=>"001101011",
  19950=>"100101000",
  19951=>"111101101",
  19952=>"110000010",
  19953=>"000001011",
  19954=>"111001100",
  19955=>"111000110",
  19956=>"001101111",
  19957=>"111011010",
  19958=>"110001000",
  19959=>"110000111",
  19960=>"000000000",
  19961=>"110111000",
  19962=>"100100100",
  19963=>"100111001",
  19964=>"100011000",
  19965=>"101010000",
  19966=>"110011010",
  19967=>"110110110",
  19968=>"101101100",
  19969=>"110110000",
  19970=>"001100010",
  19971=>"110000110",
  19972=>"001101000",
  19973=>"001111000",
  19974=>"100011110",
  19975=>"010101101",
  19976=>"001000111",
  19977=>"111111111",
  19978=>"100110111",
  19979=>"010000110",
  19980=>"011101100",
  19981=>"100011100",
  19982=>"001101000",
  19983=>"011010011",
  19984=>"111001011",
  19985=>"010010101",
  19986=>"011000011",
  19987=>"101010001",
  19988=>"010111101",
  19989=>"010101011",
  19990=>"011011000",
  19991=>"101010111",
  19992=>"100011111",
  19993=>"010000111",
  19994=>"111000001",
  19995=>"100111100",
  19996=>"000100011",
  19997=>"010001100",
  19998=>"001111001",
  19999=>"111100100",
  20000=>"001110010",
  20001=>"011010011",
  20002=>"110000010",
  20003=>"100101101",
  20004=>"111110000",
  20005=>"000011011",
  20006=>"110110001",
  20007=>"011110001",
  20008=>"101101101",
  20009=>"100110011",
  20010=>"101000100",
  20011=>"010101100",
  20012=>"101101101",
  20013=>"110110011",
  20014=>"101100000",
  20015=>"111011101",
  20016=>"110011111",
  20017=>"110011110",
  20018=>"011011010",
  20019=>"110000111",
  20020=>"000000001",
  20021=>"100000010",
  20022=>"011001110",
  20023=>"110010111",
  20024=>"101001100",
  20025=>"111101110",
  20026=>"000111100",
  20027=>"011101101",
  20028=>"111111111",
  20029=>"100010010",
  20030=>"110100001",
  20031=>"101111110",
  20032=>"011110010",
  20033=>"111111100",
  20034=>"010010100",
  20035=>"010111001",
  20036=>"110100110",
  20037=>"011010110",
  20038=>"000101110",
  20039=>"101010000",
  20040=>"100111000",
  20041=>"010001010",
  20042=>"110000010",
  20043=>"001110110",
  20044=>"111111011",
  20045=>"011011010",
  20046=>"101000000",
  20047=>"000111110",
  20048=>"011000000",
  20049=>"110010001",
  20050=>"000110111",
  20051=>"001111011",
  20052=>"100110011",
  20053=>"000001010",
  20054=>"000010001",
  20055=>"111001100",
  20056=>"000011101",
  20057=>"001100000",
  20058=>"001010001",
  20059=>"000001011",
  20060=>"101111110",
  20061=>"010100110",
  20062=>"001101011",
  20063=>"000101101",
  20064=>"111101010",
  20065=>"001100000",
  20066=>"110010110",
  20067=>"100100000",
  20068=>"110101110",
  20069=>"011010011",
  20070=>"100111001",
  20071=>"000000000",
  20072=>"001000101",
  20073=>"110101000",
  20074=>"111100001",
  20075=>"111110000",
  20076=>"001111110",
  20077=>"000001101",
  20078=>"100011001",
  20079=>"011100000",
  20080=>"000010010",
  20081=>"000011010",
  20082=>"101011000",
  20083=>"100110101",
  20084=>"011001100",
  20085=>"000000010",
  20086=>"110101100",
  20087=>"011010100",
  20088=>"110011000",
  20089=>"101101010",
  20090=>"011100010",
  20091=>"110111011",
  20092=>"100011011",
  20093=>"101010100",
  20094=>"111011000",
  20095=>"011011011",
  20096=>"111011100",
  20097=>"110001001",
  20098=>"010001000",
  20099=>"011111011",
  20100=>"111001000",
  20101=>"001101111",
  20102=>"011110110",
  20103=>"000110001",
  20104=>"000001000",
  20105=>"001101000",
  20106=>"110101110",
  20107=>"110011000",
  20108=>"111011110",
  20109=>"000110000",
  20110=>"101011101",
  20111=>"110110010",
  20112=>"111101011",
  20113=>"001111001",
  20114=>"101010111",
  20115=>"110111111",
  20116=>"000010011",
  20117=>"100110011",
  20118=>"010101000",
  20119=>"011010010",
  20120=>"011111100",
  20121=>"010111010",
  20122=>"010110111",
  20123=>"111000000",
  20124=>"110001101",
  20125=>"000111001",
  20126=>"111111001",
  20127=>"101101001",
  20128=>"000110000",
  20129=>"010100010",
  20130=>"000011010",
  20131=>"111100111",
  20132=>"001100001",
  20133=>"011001101",
  20134=>"100100000",
  20135=>"000000000",
  20136=>"101010110",
  20137=>"011101010",
  20138=>"010000001",
  20139=>"101101000",
  20140=>"110000100",
  20141=>"100100010",
  20142=>"011000100",
  20143=>"010111111",
  20144=>"011101100",
  20145=>"000010001",
  20146=>"010000111",
  20147=>"011110001",
  20148=>"010011010",
  20149=>"110010100",
  20150=>"010011100",
  20151=>"001011010",
  20152=>"101011100",
  20153=>"110100001",
  20154=>"100111010",
  20155=>"110110111",
  20156=>"101111010",
  20157=>"010011100",
  20158=>"001001000",
  20159=>"000010000",
  20160=>"001011001",
  20161=>"111100110",
  20162=>"111101010",
  20163=>"011000000",
  20164=>"000000100",
  20165=>"001001000",
  20166=>"110010100",
  20167=>"000011001",
  20168=>"010110001",
  20169=>"110101111",
  20170=>"010010000",
  20171=>"100110110",
  20172=>"001100011",
  20173=>"000100101",
  20174=>"011100001",
  20175=>"111111110",
  20176=>"110011010",
  20177=>"011000011",
  20178=>"101110110",
  20179=>"000001111",
  20180=>"110101000",
  20181=>"001010111",
  20182=>"001000010",
  20183=>"001000010",
  20184=>"000010000",
  20185=>"011000111",
  20186=>"100010100",
  20187=>"010011101",
  20188=>"001101011",
  20189=>"010000000",
  20190=>"100111011",
  20191=>"011110101",
  20192=>"111110011",
  20193=>"010010011",
  20194=>"011110111",
  20195=>"100110011",
  20196=>"010001010",
  20197=>"100100000",
  20198=>"000001011",
  20199=>"110000010",
  20200=>"000110000",
  20201=>"011010101",
  20202=>"110010010",
  20203=>"100000001",
  20204=>"100001110",
  20205=>"000010010",
  20206=>"100110010",
  20207=>"001011010",
  20208=>"011110001",
  20209=>"010100101",
  20210=>"001111111",
  20211=>"101101111",
  20212=>"111011100",
  20213=>"010001111",
  20214=>"100111011",
  20215=>"111100010",
  20216=>"011011111",
  20217=>"110010101",
  20218=>"011011010",
  20219=>"101100011",
  20220=>"110001110",
  20221=>"001010111",
  20222=>"001111011",
  20223=>"010001110",
  20224=>"111010110",
  20225=>"101011011",
  20226=>"010000110",
  20227=>"110101000",
  20228=>"110101111",
  20229=>"100100111",
  20230=>"011101110",
  20231=>"110011111",
  20232=>"001101110",
  20233=>"101010100",
  20234=>"100011000",
  20235=>"111101111",
  20236=>"110111001",
  20237=>"001011001",
  20238=>"010001100",
  20239=>"110001101",
  20240=>"100000011",
  20241=>"100111110",
  20242=>"010001000",
  20243=>"111001110",
  20244=>"111011100",
  20245=>"100111101",
  20246=>"110001110",
  20247=>"101101000",
  20248=>"001111110",
  20249=>"110000100",
  20250=>"100110101",
  20251=>"011011001",
  20252=>"110011000",
  20253=>"001111000",
  20254=>"011100100",
  20255=>"110001101",
  20256=>"010100001",
  20257=>"010111011",
  20258=>"000011100",
  20259=>"101111100",
  20260=>"110111001",
  20261=>"000010000",
  20262=>"001110001",
  20263=>"010101001",
  20264=>"001110011",
  20265=>"100101100",
  20266=>"110100111",
  20267=>"100001100",
  20268=>"101110010",
  20269=>"100100000",
  20270=>"010110010",
  20271=>"110010010",
  20272=>"011010110",
  20273=>"011000100",
  20274=>"101111010",
  20275=>"111111100",
  20276=>"001001011",
  20277=>"100101110",
  20278=>"010000100",
  20279=>"110100011",
  20280=>"100111100",
  20281=>"001101000",
  20282=>"100110100",
  20283=>"010000010",
  20284=>"011001011",
  20285=>"010000111",
  20286=>"110001000",
  20287=>"010000101",
  20288=>"110000001",
  20289=>"101100111",
  20290=>"010001101",
  20291=>"011001001",
  20292=>"010000001",
  20293=>"110001011",
  20294=>"000011111",
  20295=>"101011010",
  20296=>"000100011",
  20297=>"101010001",
  20298=>"001111111",
  20299=>"010101000",
  20300=>"001010101",
  20301=>"010010111",
  20302=>"100010000",
  20303=>"111101101",
  20304=>"101111110",
  20305=>"110110000",
  20306=>"000100001",
  20307=>"000111110",
  20308=>"000101110",
  20309=>"011000101",
  20310=>"100010110",
  20311=>"001010000",
  20312=>"011001000",
  20313=>"110111100",
  20314=>"010010101",
  20315=>"100001010",
  20316=>"100101011",
  20317=>"101000000",
  20318=>"111111111",
  20319=>"000011111",
  20320=>"110011000",
  20321=>"111000001",
  20322=>"000110101",
  20323=>"100111010",
  20324=>"101011010",
  20325=>"001000100",
  20326=>"110001100",
  20327=>"000100000",
  20328=>"010010011",
  20329=>"111101010",
  20330=>"000000100",
  20331=>"011100111",
  20332=>"101010000",
  20333=>"000000010",
  20334=>"110000010",
  20335=>"001100111",
  20336=>"011111100",
  20337=>"010011110",
  20338=>"011011011",
  20339=>"000010100",
  20340=>"100000010",
  20341=>"010011101",
  20342=>"110011101",
  20343=>"001011101",
  20344=>"101010000",
  20345=>"010111101",
  20346=>"100000010",
  20347=>"001101001",
  20348=>"011011100",
  20349=>"100110001",
  20350=>"110101011",
  20351=>"111001110",
  20352=>"010111010",
  20353=>"111011110",
  20354=>"000101110",
  20355=>"000101001",
  20356=>"100011101",
  20357=>"110001001",
  20358=>"101010010",
  20359=>"011101101",
  20360=>"001101000",
  20361=>"100101000",
  20362=>"101011101",
  20363=>"010001001",
  20364=>"001010100",
  20365=>"011100000",
  20366=>"101111010",
  20367=>"100101001",
  20368=>"000001110",
  20369=>"101101111",
  20370=>"011111110",
  20371=>"101011011",
  20372=>"010010100",
  20373=>"110000000",
  20374=>"000010111",
  20375=>"011110001",
  20376=>"110011001",
  20377=>"000100010",
  20378=>"000001101",
  20379=>"101111011",
  20380=>"000000001",
  20381=>"000111111",
  20382=>"001000001",
  20383=>"011011010",
  20384=>"100001110",
  20385=>"101110111",
  20386=>"100111011",
  20387=>"110000011",
  20388=>"100100110",
  20389=>"010001110",
  20390=>"001100001",
  20391=>"000001001",
  20392=>"011000011",
  20393=>"111001111",
  20394=>"011111110",
  20395=>"110110001",
  20396=>"101001101",
  20397=>"001111100",
  20398=>"101111100",
  20399=>"000000000",
  20400=>"100110110",
  20401=>"100111101",
  20402=>"011110000",
  20403=>"011010001",
  20404=>"000010010",
  20405=>"100110100",
  20406=>"111000001",
  20407=>"011011011",
  20408=>"101101010",
  20409=>"011010110",
  20410=>"011100000",
  20411=>"011010000",
  20412=>"000101010",
  20413=>"010110000",
  20414=>"001010001",
  20415=>"011100011",
  20416=>"001110001",
  20417=>"100010101",
  20418=>"110100100",
  20419=>"100100010",
  20420=>"110011111",
  20421=>"101101001",
  20422=>"000111100",
  20423=>"010001000",
  20424=>"010111110",
  20425=>"001011000",
  20426=>"101001011",
  20427=>"001011101",
  20428=>"110111010",
  20429=>"110000001",
  20430=>"101111110",
  20431=>"011100111",
  20432=>"011111001",
  20433=>"111110001",
  20434=>"010111011",
  20435=>"110110010",
  20436=>"011000001",
  20437=>"011100010",
  20438=>"100111001",
  20439=>"111111000",
  20440=>"100010010",
  20441=>"100010110",
  20442=>"110001010",
  20443=>"100111001",
  20444=>"111111001",
  20445=>"110111101",
  20446=>"101111000",
  20447=>"000000000",
  20448=>"101111100",
  20449=>"000010111",
  20450=>"000001010",
  20451=>"100000000",
  20452=>"000011100",
  20453=>"111101000",
  20454=>"001010001",
  20455=>"100110000",
  20456=>"100100101",
  20457=>"100110110",
  20458=>"111111111",
  20459=>"010010110",
  20460=>"110000010",
  20461=>"111111000",
  20462=>"000011011",
  20463=>"001110100",
  20464=>"000011011",
  20465=>"001010011",
  20466=>"011111111",
  20467=>"011010100",
  20468=>"001110110",
  20469=>"101101011",
  20470=>"101110110",
  20471=>"100111111",
  20472=>"001011101",
  20473=>"101101010",
  20474=>"100101001",
  20475=>"011111011",
  20476=>"011001110",
  20477=>"101110011",
  20478=>"101000000",
  20479=>"011011111",
  20480=>"111101101",
  20481=>"011101110",
  20482=>"100010110",
  20483=>"110101001",
  20484=>"000111010",
  20485=>"001100101",
  20486=>"001010001",
  20487=>"000001000",
  20488=>"111110100",
  20489=>"010000101",
  20490=>"010110111",
  20491=>"101110011",
  20492=>"001111110",
  20493=>"100100100",
  20494=>"001001101",
  20495=>"011011111",
  20496=>"110111011",
  20497=>"110110101",
  20498=>"100001100",
  20499=>"100010111",
  20500=>"100111111",
  20501=>"101111100",
  20502=>"110011011",
  20503=>"110011101",
  20504=>"010010011",
  20505=>"001001100",
  20506=>"000111110",
  20507=>"110010010",
  20508=>"011010000",
  20509=>"110011101",
  20510=>"101111011",
  20511=>"010000000",
  20512=>"010010111",
  20513=>"111010101",
  20514=>"100010100",
  20515=>"001100001",
  20516=>"001011110",
  20517=>"001110001",
  20518=>"101001000",
  20519=>"001011010",
  20520=>"010010010",
  20521=>"010001110",
  20522=>"110001110",
  20523=>"110001010",
  20524=>"111000100",
  20525=>"011110110",
  20526=>"110101110",
  20527=>"001111111",
  20528=>"011011100",
  20529=>"000110101",
  20530=>"101111111",
  20531=>"000100101",
  20532=>"000000001",
  20533=>"100000010",
  20534=>"101001011",
  20535=>"000110010",
  20536=>"000110001",
  20537=>"000101010",
  20538=>"111111110",
  20539=>"110010010",
  20540=>"110001110",
  20541=>"011010101",
  20542=>"101000000",
  20543=>"110011100",
  20544=>"110110111",
  20545=>"011010011",
  20546=>"000100101",
  20547=>"101000010",
  20548=>"000011100",
  20549=>"100011111",
  20550=>"100101101",
  20551=>"000001000",
  20552=>"001110001",
  20553=>"110000110",
  20554=>"001001110",
  20555=>"111111111",
  20556=>"111111100",
  20557=>"000111010",
  20558=>"010011000",
  20559=>"100101110",
  20560=>"001001100",
  20561=>"011010011",
  20562=>"010011010",
  20563=>"000111000",
  20564=>"110111100",
  20565=>"000010100",
  20566=>"111010001",
  20567=>"100100011",
  20568=>"100101000",
  20569=>"000011110",
  20570=>"010011111",
  20571=>"010001101",
  20572=>"000000010",
  20573=>"001001111",
  20574=>"100011101",
  20575=>"000000111",
  20576=>"001100011",
  20577=>"011100101",
  20578=>"111011010",
  20579=>"111100011",
  20580=>"001010100",
  20581=>"000110111",
  20582=>"001001011",
  20583=>"001010011",
  20584=>"110100010",
  20585=>"110000001",
  20586=>"010101111",
  20587=>"101101001",
  20588=>"101110000",
  20589=>"110111010",
  20590=>"100100111",
  20591=>"011111111",
  20592=>"110111111",
  20593=>"001100101",
  20594=>"110110011",
  20595=>"000101011",
  20596=>"100011011",
  20597=>"110100000",
  20598=>"111011011",
  20599=>"011011010",
  20600=>"110101100",
  20601=>"010001011",
  20602=>"011101000",
  20603=>"011001010",
  20604=>"001100011",
  20605=>"010010011",
  20606=>"000011011",
  20607=>"101001000",
  20608=>"101101011",
  20609=>"000001000",
  20610=>"010111010",
  20611=>"010011101",
  20612=>"000100011",
  20613=>"101010101",
  20614=>"010000101",
  20615=>"011100001",
  20616=>"001000111",
  20617=>"000010101",
  20618=>"101101001",
  20619=>"101010110",
  20620=>"000110010",
  20621=>"110000111",
  20622=>"001010001",
  20623=>"001101101",
  20624=>"000001110",
  20625=>"110100000",
  20626=>"101111111",
  20627=>"101000111",
  20628=>"101000010",
  20629=>"110101111",
  20630=>"001110101",
  20631=>"000001101",
  20632=>"000010111",
  20633=>"101001001",
  20634=>"000100000",
  20635=>"000101011",
  20636=>"100101010",
  20637=>"011001001",
  20638=>"110010100",
  20639=>"011000001",
  20640=>"101110111",
  20641=>"001100001",
  20642=>"110100100",
  20643=>"000001100",
  20644=>"110111011",
  20645=>"111001110",
  20646=>"011001100",
  20647=>"111110010",
  20648=>"101000010",
  20649=>"000000000",
  20650=>"010000101",
  20651=>"001001110",
  20652=>"011100111",
  20653=>"011011101",
  20654=>"100010111",
  20655=>"000110100",
  20656=>"001101111",
  20657=>"000100111",
  20658=>"010101011",
  20659=>"010110001",
  20660=>"010010011",
  20661=>"111000100",
  20662=>"001000011",
  20663=>"001011010",
  20664=>"110001100",
  20665=>"110100101",
  20666=>"001110111",
  20667=>"000110000",
  20668=>"011011010",
  20669=>"111110001",
  20670=>"101010010",
  20671=>"100100100",
  20672=>"111111110",
  20673=>"111000001",
  20674=>"011011101",
  20675=>"100110111",
  20676=>"000110000",
  20677=>"001011000",
  20678=>"111110001",
  20679=>"001001011",
  20680=>"101101111",
  20681=>"111011110",
  20682=>"110100111",
  20683=>"101011110",
  20684=>"110100001",
  20685=>"101101001",
  20686=>"010000110",
  20687=>"011110111",
  20688=>"111001000",
  20689=>"100011111",
  20690=>"010001011",
  20691=>"101010101",
  20692=>"100110000",
  20693=>"000101111",
  20694=>"000011110",
  20695=>"111101101",
  20696=>"000011000",
  20697=>"011100001",
  20698=>"011010000",
  20699=>"001010001",
  20700=>"110111110",
  20701=>"000100110",
  20702=>"101000100",
  20703=>"010111110",
  20704=>"110111011",
  20705=>"001111011",
  20706=>"110110001",
  20707=>"000001100",
  20708=>"010100011",
  20709=>"100100000",
  20710=>"000010101",
  20711=>"000001001",
  20712=>"011100010",
  20713=>"000001000",
  20714=>"110000001",
  20715=>"001010111",
  20716=>"001011011",
  20717=>"111011110",
  20718=>"111111010",
  20719=>"010001000",
  20720=>"010110111",
  20721=>"101110101",
  20722=>"011001101",
  20723=>"000101100",
  20724=>"001110111",
  20725=>"100111100",
  20726=>"001011101",
  20727=>"000000010",
  20728=>"011000010",
  20729=>"000101000",
  20730=>"110110101",
  20731=>"011000111",
  20732=>"010001111",
  20733=>"010010110",
  20734=>"010010111",
  20735=>"011001100",
  20736=>"101111001",
  20737=>"000001100",
  20738=>"000101111",
  20739=>"111101101",
  20740=>"001001010",
  20741=>"111011000",
  20742=>"111100111",
  20743=>"011101100",
  20744=>"000001100",
  20745=>"111110111",
  20746=>"100101000",
  20747=>"010011101",
  20748=>"101110010",
  20749=>"111001000",
  20750=>"000001111",
  20751=>"000110110",
  20752=>"100011111",
  20753=>"101110001",
  20754=>"010101110",
  20755=>"000100100",
  20756=>"100110110",
  20757=>"000101011",
  20758=>"011110000",
  20759=>"011111101",
  20760=>"001011101",
  20761=>"001001111",
  20762=>"110001111",
  20763=>"110111000",
  20764=>"011000001",
  20765=>"100100101",
  20766=>"101000110",
  20767=>"000000010",
  20768=>"111111001",
  20769=>"100111001",
  20770=>"001110111",
  20771=>"000011101",
  20772=>"110110100",
  20773=>"100100010",
  20774=>"010100101",
  20775=>"100010001",
  20776=>"101110000",
  20777=>"111100001",
  20778=>"000000011",
  20779=>"001010010",
  20780=>"011001000",
  20781=>"100010010",
  20782=>"101111111",
  20783=>"010011000",
  20784=>"110101000",
  20785=>"101111110",
  20786=>"000001011",
  20787=>"010011111",
  20788=>"011011101",
  20789=>"011100111",
  20790=>"001000010",
  20791=>"000111110",
  20792=>"100100111",
  20793=>"001111011",
  20794=>"110010011",
  20795=>"001011111",
  20796=>"111011110",
  20797=>"001101000",
  20798=>"001000111",
  20799=>"011000001",
  20800=>"001101000",
  20801=>"100011001",
  20802=>"011100000",
  20803=>"011011010",
  20804=>"010011100",
  20805=>"001000101",
  20806=>"011101110",
  20807=>"110101001",
  20808=>"111011110",
  20809=>"010111011",
  20810=>"100000110",
  20811=>"010010100",
  20812=>"101101001",
  20813=>"100001111",
  20814=>"100000000",
  20815=>"100110111",
  20816=>"011110001",
  20817=>"110010001",
  20818=>"010100110",
  20819=>"000111110",
  20820=>"111111100",
  20821=>"001110100",
  20822=>"000011000",
  20823=>"000101010",
  20824=>"110111010",
  20825=>"010111100",
  20826=>"011000000",
  20827=>"101000110",
  20828=>"011111001",
  20829=>"001111110",
  20830=>"010111101",
  20831=>"011000000",
  20832=>"011111000",
  20833=>"000001110",
  20834=>"000010101",
  20835=>"010011000",
  20836=>"000101111",
  20837=>"101010110",
  20838=>"011110100",
  20839=>"111111001",
  20840=>"111100101",
  20841=>"010011110",
  20842=>"110001100",
  20843=>"000000101",
  20844=>"101101111",
  20845=>"001001101",
  20846=>"010010111",
  20847=>"010110110",
  20848=>"001010000",
  20849=>"111100110",
  20850=>"010011010",
  20851=>"001111001",
  20852=>"011001110",
  20853=>"010001100",
  20854=>"100100010",
  20855=>"001100110",
  20856=>"000110100",
  20857=>"110001000",
  20858=>"110010111",
  20859=>"110011001",
  20860=>"001101101",
  20861=>"110101101",
  20862=>"011110010",
  20863=>"001110100",
  20864=>"100111100",
  20865=>"100010101",
  20866=>"011010111",
  20867=>"111111001",
  20868=>"111000001",
  20869=>"111100011",
  20870=>"001111110",
  20871=>"110000010",
  20872=>"111110111",
  20873=>"100110101",
  20874=>"100110001",
  20875=>"110100111",
  20876=>"000001000",
  20877=>"101001111",
  20878=>"001110101",
  20879=>"010101110",
  20880=>"111000110",
  20881=>"110010000",
  20882=>"111010111",
  20883=>"010000001",
  20884=>"101111101",
  20885=>"000001111",
  20886=>"001100111",
  20887=>"010100010",
  20888=>"100011110",
  20889=>"111011000",
  20890=>"101001101",
  20891=>"111101010",
  20892=>"010001111",
  20893=>"010110001",
  20894=>"010100100",
  20895=>"111110011",
  20896=>"010100111",
  20897=>"011000000",
  20898=>"111110111",
  20899=>"111100110",
  20900=>"111111001",
  20901=>"101010010",
  20902=>"100000110",
  20903=>"100001111",
  20904=>"101010011",
  20905=>"101011010",
  20906=>"011110010",
  20907=>"110000011",
  20908=>"001011100",
  20909=>"111100100",
  20910=>"101001001",
  20911=>"111001001",
  20912=>"000101000",
  20913=>"111011001",
  20914=>"111100110",
  20915=>"011000110",
  20916=>"000100000",
  20917=>"000000110",
  20918=>"101011001",
  20919=>"101110000",
  20920=>"001000100",
  20921=>"110011001",
  20922=>"011101110",
  20923=>"110001111",
  20924=>"110100101",
  20925=>"010111111",
  20926=>"001100001",
  20927=>"110111101",
  20928=>"100110001",
  20929=>"010001111",
  20930=>"011001110",
  20931=>"011001000",
  20932=>"111110110",
  20933=>"101000001",
  20934=>"011010011",
  20935=>"100000100",
  20936=>"100011101",
  20937=>"111010000",
  20938=>"001000011",
  20939=>"101010000",
  20940=>"101110100",
  20941=>"001010011",
  20942=>"010100110",
  20943=>"110010100",
  20944=>"010100101",
  20945=>"000111110",
  20946=>"001100111",
  20947=>"000010010",
  20948=>"101101111",
  20949=>"010001111",
  20950=>"011010001",
  20951=>"100110001",
  20952=>"000010110",
  20953=>"111010110",
  20954=>"001101011",
  20955=>"101000101",
  20956=>"101001100",
  20957=>"011111011",
  20958=>"001110100",
  20959=>"111110110",
  20960=>"110000110",
  20961=>"000000100",
  20962=>"010110010",
  20963=>"110100100",
  20964=>"010010001",
  20965=>"000110101",
  20966=>"011000100",
  20967=>"100001011",
  20968=>"110000010",
  20969=>"111000011",
  20970=>"000000101",
  20971=>"100101110",
  20972=>"101011011",
  20973=>"110111111",
  20974=>"000101011",
  20975=>"111001011",
  20976=>"100011101",
  20977=>"100010010",
  20978=>"010011100",
  20979=>"100010100",
  20980=>"001100000",
  20981=>"000001001",
  20982=>"000110100",
  20983=>"010011111",
  20984=>"010000001",
  20985=>"010001001",
  20986=>"101001101",
  20987=>"100100011",
  20988=>"010001110",
  20989=>"010100100",
  20990=>"101000110",
  20991=>"110100000",
  20992=>"001101001",
  20993=>"000111101",
  20994=>"111011000",
  20995=>"111101101",
  20996=>"000100000",
  20997=>"100111101",
  20998=>"111101000",
  20999=>"110110111",
  21000=>"011011001",
  21001=>"000111100",
  21002=>"000111101",
  21003=>"101001000",
  21004=>"011011011",
  21005=>"001011001",
  21006=>"011000010",
  21007=>"100100111",
  21008=>"110011110",
  21009=>"101010001",
  21010=>"000010111",
  21011=>"100101100",
  21012=>"000111110",
  21013=>"011111100",
  21014=>"011110100",
  21015=>"001101001",
  21016=>"000100110",
  21017=>"000100011",
  21018=>"100010111",
  21019=>"001011001",
  21020=>"111101011",
  21021=>"101010010",
  21022=>"110100101",
  21023=>"010000100",
  21024=>"001010001",
  21025=>"111111111",
  21026=>"011100011",
  21027=>"001011011",
  21028=>"101111011",
  21029=>"110110010",
  21030=>"110000100",
  21031=>"110100100",
  21032=>"011000000",
  21033=>"010100000",
  21034=>"101100110",
  21035=>"001011110",
  21036=>"010100001",
  21037=>"100111011",
  21038=>"100001111",
  21039=>"000010110",
  21040=>"011101001",
  21041=>"110000111",
  21042=>"110011001",
  21043=>"011101101",
  21044=>"100011110",
  21045=>"101100000",
  21046=>"001101011",
  21047=>"111110010",
  21048=>"101001111",
  21049=>"001100100",
  21050=>"111010001",
  21051=>"000001101",
  21052=>"101111110",
  21053=>"100111111",
  21054=>"001110000",
  21055=>"101110001",
  21056=>"010010111",
  21057=>"101000011",
  21058=>"101011001",
  21059=>"110000101",
  21060=>"010010000",
  21061=>"000000110",
  21062=>"111111101",
  21063=>"110100101",
  21064=>"100001000",
  21065=>"111001010",
  21066=>"110000110",
  21067=>"110001000",
  21068=>"011010111",
  21069=>"111000101",
  21070=>"111010111",
  21071=>"010011010",
  21072=>"010001000",
  21073=>"100110000",
  21074=>"111010000",
  21075=>"000110001",
  21076=>"000100110",
  21077=>"000001111",
  21078=>"111000111",
  21079=>"100110101",
  21080=>"001000000",
  21081=>"100110001",
  21082=>"010010101",
  21083=>"000010100",
  21084=>"001001111",
  21085=>"000100101",
  21086=>"011101100",
  21087=>"001000000",
  21088=>"010111011",
  21089=>"010110010",
  21090=>"101011100",
  21091=>"100000100",
  21092=>"101001100",
  21093=>"010111011",
  21094=>"011011111",
  21095=>"011000010",
  21096=>"100011000",
  21097=>"001110110",
  21098=>"110011001",
  21099=>"000110001",
  21100=>"101001010",
  21101=>"111101010",
  21102=>"101101011",
  21103=>"110010001",
  21104=>"101111111",
  21105=>"111011000",
  21106=>"011111011",
  21107=>"001011011",
  21108=>"111101010",
  21109=>"010010010",
  21110=>"110110010",
  21111=>"001010111",
  21112=>"101000000",
  21113=>"010100111",
  21114=>"101001011",
  21115=>"101010111",
  21116=>"011000111",
  21117=>"111101000",
  21118=>"010001000",
  21119=>"000100110",
  21120=>"101000111",
  21121=>"101110111",
  21122=>"001111000",
  21123=>"011001111",
  21124=>"011000000",
  21125=>"101011011",
  21126=>"010011110",
  21127=>"111101001",
  21128=>"101111101",
  21129=>"000001001",
  21130=>"000110000",
  21131=>"111010000",
  21132=>"000101101",
  21133=>"011100011",
  21134=>"000011010",
  21135=>"000100111",
  21136=>"010101110",
  21137=>"101100111",
  21138=>"011101110",
  21139=>"000011011",
  21140=>"001001001",
  21141=>"001100111",
  21142=>"110101101",
  21143=>"101110010",
  21144=>"001001100",
  21145=>"010110000",
  21146=>"101010011",
  21147=>"100100101",
  21148=>"100100001",
  21149=>"000000000",
  21150=>"011100000",
  21151=>"111100111",
  21152=>"101100110",
  21153=>"011101101",
  21154=>"001100111",
  21155=>"111111101",
  21156=>"101001011",
  21157=>"001000001",
  21158=>"110010101",
  21159=>"010010101",
  21160=>"001010000",
  21161=>"000111001",
  21162=>"011001000",
  21163=>"100000110",
  21164=>"110001000",
  21165=>"001110010",
  21166=>"001111000",
  21167=>"100101000",
  21168=>"100001100",
  21169=>"000111001",
  21170=>"101010010",
  21171=>"011100111",
  21172=>"100011100",
  21173=>"010010010",
  21174=>"000101010",
  21175=>"011100010",
  21176=>"110111011",
  21177=>"010100111",
  21178=>"110110111",
  21179=>"000000101",
  21180=>"001101000",
  21181=>"001011110",
  21182=>"100000111",
  21183=>"101111100",
  21184=>"111100110",
  21185=>"001110000",
  21186=>"101000011",
  21187=>"010110001",
  21188=>"110100110",
  21189=>"010000010",
  21190=>"110000011",
  21191=>"000010010",
  21192=>"111110101",
  21193=>"001110000",
  21194=>"000010010",
  21195=>"100111100",
  21196=>"001111001",
  21197=>"110001011",
  21198=>"111100001",
  21199=>"110000110",
  21200=>"101111001",
  21201=>"100100000",
  21202=>"101011001",
  21203=>"110010110",
  21204=>"010101001",
  21205=>"001111001",
  21206=>"111001111",
  21207=>"100100011",
  21208=>"101000000",
  21209=>"110111010",
  21210=>"011101101",
  21211=>"011000100",
  21212=>"001100101",
  21213=>"101000101",
  21214=>"110111110",
  21215=>"111000111",
  21216=>"011111111",
  21217=>"111101001",
  21218=>"010000111",
  21219=>"100000101",
  21220=>"100000010",
  21221=>"001100001",
  21222=>"100010001",
  21223=>"100000110",
  21224=>"110100110",
  21225=>"101011011",
  21226=>"001010010",
  21227=>"111100100",
  21228=>"110101111",
  21229=>"100011011",
  21230=>"001110010",
  21231=>"000101111",
  21232=>"011101111",
  21233=>"001001111",
  21234=>"110101110",
  21235=>"001100111",
  21236=>"111001100",
  21237=>"110110100",
  21238=>"100111101",
  21239=>"001110000",
  21240=>"001001110",
  21241=>"111001000",
  21242=>"011011111",
  21243=>"000000110",
  21244=>"111101000",
  21245=>"000110010",
  21246=>"011000001",
  21247=>"001110111",
  21248=>"001001101",
  21249=>"010000001",
  21250=>"010000110",
  21251=>"001110001",
  21252=>"011111101",
  21253=>"001100000",
  21254=>"010011001",
  21255=>"111101101",
  21256=>"011000001",
  21257=>"111010100",
  21258=>"111001001",
  21259=>"001101110",
  21260=>"001100110",
  21261=>"101101110",
  21262=>"000100101",
  21263=>"000001001",
  21264=>"010111100",
  21265=>"111101110",
  21266=>"000110010",
  21267=>"111100001",
  21268=>"110000010",
  21269=>"011000001",
  21270=>"101000110",
  21271=>"010110010",
  21272=>"001000010",
  21273=>"111011000",
  21274=>"110101001",
  21275=>"001001011",
  21276=>"100010101",
  21277=>"101101011",
  21278=>"111110000",
  21279=>"000000000",
  21280=>"101110110",
  21281=>"000011011",
  21282=>"001000111",
  21283=>"111101011",
  21284=>"111101101",
  21285=>"100100011",
  21286=>"110001110",
  21287=>"001001111",
  21288=>"110010101",
  21289=>"010110110",
  21290=>"110101001",
  21291=>"101110101",
  21292=>"011111010",
  21293=>"100111111",
  21294=>"110111011",
  21295=>"111010000",
  21296=>"011000100",
  21297=>"001010000",
  21298=>"101000001",
  21299=>"010100100",
  21300=>"101101100",
  21301=>"111011100",
  21302=>"100111000",
  21303=>"001111010",
  21304=>"101101000",
  21305=>"000000111",
  21306=>"010000110",
  21307=>"110101000",
  21308=>"001011000",
  21309=>"100111001",
  21310=>"111010010",
  21311=>"000001011",
  21312=>"101001010",
  21313=>"001010100",
  21314=>"111110001",
  21315=>"000000000",
  21316=>"000001100",
  21317=>"001110011",
  21318=>"100000010",
  21319=>"110011100",
  21320=>"101011100",
  21321=>"100100100",
  21322=>"111011001",
  21323=>"001011110",
  21324=>"001100000",
  21325=>"010110000",
  21326=>"010100111",
  21327=>"110011111",
  21328=>"111001111",
  21329=>"001000001",
  21330=>"000011001",
  21331=>"011110000",
  21332=>"011110010",
  21333=>"101011101",
  21334=>"111011100",
  21335=>"011011010",
  21336=>"000111101",
  21337=>"000110001",
  21338=>"000101011",
  21339=>"011101010",
  21340=>"101011110",
  21341=>"110010101",
  21342=>"010000010",
  21343=>"000011010",
  21344=>"101100111",
  21345=>"100101011",
  21346=>"001101011",
  21347=>"110011111",
  21348=>"001101110",
  21349=>"110110101",
  21350=>"001001110",
  21351=>"111111010",
  21352=>"101001010",
  21353=>"000001110",
  21354=>"101110101",
  21355=>"101100000",
  21356=>"001011100",
  21357=>"111100101",
  21358=>"110100001",
  21359=>"011101001",
  21360=>"001011010",
  21361=>"110101101",
  21362=>"001000010",
  21363=>"001100101",
  21364=>"000001110",
  21365=>"000101111",
  21366=>"111001110",
  21367=>"100101011",
  21368=>"011110111",
  21369=>"000001101",
  21370=>"000001100",
  21371=>"110101011",
  21372=>"001010110",
  21373=>"001110001",
  21374=>"010001011",
  21375=>"010001100",
  21376=>"111000010",
  21377=>"001001011",
  21378=>"000110010",
  21379=>"100101100",
  21380=>"011100001",
  21381=>"110111110",
  21382=>"110001001",
  21383=>"010011001",
  21384=>"100001010",
  21385=>"101000001",
  21386=>"111000110",
  21387=>"110101101",
  21388=>"111110111",
  21389=>"001111111",
  21390=>"111110010",
  21391=>"011101110",
  21392=>"110011110",
  21393=>"111110000",
  21394=>"001100000",
  21395=>"010111011",
  21396=>"111100100",
  21397=>"100101110",
  21398=>"101011010",
  21399=>"011000100",
  21400=>"011011111",
  21401=>"001100010",
  21402=>"111100111",
  21403=>"101011111",
  21404=>"100010000",
  21405=>"110111010",
  21406=>"101011001",
  21407=>"001111011",
  21408=>"111100101",
  21409=>"110100010",
  21410=>"000001111",
  21411=>"000010001",
  21412=>"101000001",
  21413=>"111001101",
  21414=>"111101111",
  21415=>"101010000",
  21416=>"111000100",
  21417=>"001011101",
  21418=>"100011000",
  21419=>"010101010",
  21420=>"110100000",
  21421=>"010010110",
  21422=>"011111101",
  21423=>"100100010",
  21424=>"100110011",
  21425=>"101100111",
  21426=>"011000100",
  21427=>"000010110",
  21428=>"001111010",
  21429=>"100011010",
  21430=>"000111101",
  21431=>"000000000",
  21432=>"001000001",
  21433=>"110001011",
  21434=>"100110011",
  21435=>"101100001",
  21436=>"010010110",
  21437=>"101000011",
  21438=>"111101011",
  21439=>"000000000",
  21440=>"000110100",
  21441=>"110000100",
  21442=>"010110011",
  21443=>"100011110",
  21444=>"100111111",
  21445=>"010110110",
  21446=>"000111000",
  21447=>"111010111",
  21448=>"001011101",
  21449=>"000000000",
  21450=>"110000010",
  21451=>"000010101",
  21452=>"010110001",
  21453=>"111000011",
  21454=>"000101101",
  21455=>"001101101",
  21456=>"011101100",
  21457=>"011101100",
  21458=>"001101100",
  21459=>"100001011",
  21460=>"101010001",
  21461=>"101101000",
  21462=>"100110000",
  21463=>"000111010",
  21464=>"001011100",
  21465=>"110100100",
  21466=>"010111100",
  21467=>"001111011",
  21468=>"010101100",
  21469=>"000101111",
  21470=>"001110001",
  21471=>"111000010",
  21472=>"110001111",
  21473=>"111000111",
  21474=>"100110010",
  21475=>"000001100",
  21476=>"010001001",
  21477=>"001011011",
  21478=>"001111101",
  21479=>"101111101",
  21480=>"100000010",
  21481=>"110100011",
  21482=>"111001001",
  21483=>"111000011",
  21484=>"111111111",
  21485=>"011011000",
  21486=>"001000010",
  21487=>"110010111",
  21488=>"000011010",
  21489=>"100111000",
  21490=>"100111101",
  21491=>"101110011",
  21492=>"010111010",
  21493=>"100011010",
  21494=>"011111000",
  21495=>"010110001",
  21496=>"110011110",
  21497=>"011100010",
  21498=>"010000110",
  21499=>"001010101",
  21500=>"110100110",
  21501=>"000001101",
  21502=>"111011111",
  21503=>"011101001",
  21504=>"101101111",
  21505=>"100101000",
  21506=>"001000001",
  21507=>"111101000",
  21508=>"101000110",
  21509=>"101111010",
  21510=>"010011000",
  21511=>"000101011",
  21512=>"001111011",
  21513=>"001010000",
  21514=>"001010110",
  21515=>"000001100",
  21516=>"100001111",
  21517=>"101001111",
  21518=>"000110101",
  21519=>"100011000",
  21520=>"101111100",
  21521=>"110001111",
  21522=>"111101011",
  21523=>"100111110",
  21524=>"111100100",
  21525=>"010111010",
  21526=>"011100110",
  21527=>"111100010",
  21528=>"111000010",
  21529=>"000001001",
  21530=>"001010010",
  21531=>"110010110",
  21532=>"010110101",
  21533=>"101001001",
  21534=>"100110101",
  21535=>"010101101",
  21536=>"011011010",
  21537=>"011111111",
  21538=>"111011100",
  21539=>"000010111",
  21540=>"110011110",
  21541=>"111101010",
  21542=>"101110001",
  21543=>"001111001",
  21544=>"100011101",
  21545=>"100101100",
  21546=>"011111100",
  21547=>"111010011",
  21548=>"110101010",
  21549=>"111010010",
  21550=>"101110011",
  21551=>"000001111",
  21552=>"101000011",
  21553=>"010111001",
  21554=>"010101111",
  21555=>"011001101",
  21556=>"110100010",
  21557=>"010100010",
  21558=>"010101100",
  21559=>"010010010",
  21560=>"101111001",
  21561=>"011110110",
  21562=>"000110010",
  21563=>"011011010",
  21564=>"110101010",
  21565=>"011000111",
  21566=>"111110100",
  21567=>"000101111",
  21568=>"111000011",
  21569=>"000100100",
  21570=>"110000000",
  21571=>"000111111",
  21572=>"010101101",
  21573=>"001000000",
  21574=>"011110111",
  21575=>"101111001",
  21576=>"101000011",
  21577=>"101001010",
  21578=>"000010011",
  21579=>"101100110",
  21580=>"011110110",
  21581=>"011000100",
  21582=>"111100100",
  21583=>"111001010",
  21584=>"001011000",
  21585=>"010110010",
  21586=>"011111011",
  21587=>"110001000",
  21588=>"001011100",
  21589=>"111111101",
  21590=>"011111011",
  21591=>"001100000",
  21592=>"011100100",
  21593=>"111110011",
  21594=>"011111010",
  21595=>"100001110",
  21596=>"110110000",
  21597=>"011011011",
  21598=>"100010010",
  21599=>"111101000",
  21600=>"000000010",
  21601=>"100110101",
  21602=>"001110111",
  21603=>"011100011",
  21604=>"110011000",
  21605=>"011011011",
  21606=>"111010011",
  21607=>"111010100",
  21608=>"101110110",
  21609=>"001110010",
  21610=>"101010100",
  21611=>"111001001",
  21612=>"111111110",
  21613=>"110100000",
  21614=>"100000101",
  21615=>"001001011",
  21616=>"111001100",
  21617=>"011011111",
  21618=>"000110110",
  21619=>"111010000",
  21620=>"001000010",
  21621=>"111010010",
  21622=>"000101111",
  21623=>"001110111",
  21624=>"111100111",
  21625=>"000010000",
  21626=>"010101100",
  21627=>"111111011",
  21628=>"011010110",
  21629=>"100100001",
  21630=>"110110101",
  21631=>"001000011",
  21632=>"101101010",
  21633=>"100000100",
  21634=>"010001010",
  21635=>"001000110",
  21636=>"110001011",
  21637=>"000000100",
  21638=>"111110100",
  21639=>"011000111",
  21640=>"000111111",
  21641=>"001011011",
  21642=>"001101110",
  21643=>"001101100",
  21644=>"110010110",
  21645=>"111100101",
  21646=>"011010001",
  21647=>"000111000",
  21648=>"100111100",
  21649=>"010001111",
  21650=>"001110000",
  21651=>"111001000",
  21652=>"001100111",
  21653=>"111011110",
  21654=>"010011100",
  21655=>"001110001",
  21656=>"110101011",
  21657=>"110010010",
  21658=>"011001010",
  21659=>"010110101",
  21660=>"100001100",
  21661=>"111110000",
  21662=>"100001101",
  21663=>"101011101",
  21664=>"000111100",
  21665=>"001001100",
  21666=>"010010110",
  21667=>"100101110",
  21668=>"111110000",
  21669=>"011001000",
  21670=>"100111110",
  21671=>"011011111",
  21672=>"110010110",
  21673=>"101001000",
  21674=>"011010010",
  21675=>"110111110",
  21676=>"111010110",
  21677=>"000001101",
  21678=>"000011010",
  21679=>"000001110",
  21680=>"001001101",
  21681=>"001000010",
  21682=>"001000100",
  21683=>"100101110",
  21684=>"100011000",
  21685=>"001111000",
  21686=>"010100001",
  21687=>"010001101",
  21688=>"011110001",
  21689=>"001000111",
  21690=>"100110010",
  21691=>"100101111",
  21692=>"000100001",
  21693=>"010011100",
  21694=>"110101100",
  21695=>"011001000",
  21696=>"111100100",
  21697=>"110010011",
  21698=>"001010011",
  21699=>"000000110",
  21700=>"010000100",
  21701=>"110110001",
  21702=>"001110010",
  21703=>"001010000",
  21704=>"110111101",
  21705=>"001111110",
  21706=>"011100010",
  21707=>"110001001",
  21708=>"011111001",
  21709=>"100010110",
  21710=>"000011110",
  21711=>"111100111",
  21712=>"111010000",
  21713=>"111101111",
  21714=>"110100100",
  21715=>"110000010",
  21716=>"000011110",
  21717=>"100110011",
  21718=>"001110011",
  21719=>"011001000",
  21720=>"000011110",
  21721=>"111111101",
  21722=>"111011100",
  21723=>"011111001",
  21724=>"010010101",
  21725=>"101010011",
  21726=>"000011011",
  21727=>"000100000",
  21728=>"101011000",
  21729=>"110011011",
  21730=>"010010000",
  21731=>"111000110",
  21732=>"100010010",
  21733=>"001110011",
  21734=>"100110101",
  21735=>"100111000",
  21736=>"000011100",
  21737=>"011010111",
  21738=>"111000101",
  21739=>"110111010",
  21740=>"111101101",
  21741=>"111001010",
  21742=>"000011010",
  21743=>"100100100",
  21744=>"010000001",
  21745=>"100111010",
  21746=>"101010011",
  21747=>"001100001",
  21748=>"010100010",
  21749=>"011010010",
  21750=>"100000101",
  21751=>"111101000",
  21752=>"111101100",
  21753=>"010000011",
  21754=>"110000011",
  21755=>"100011011",
  21756=>"100110111",
  21757=>"000010011",
  21758=>"100100100",
  21759=>"001010000",
  21760=>"101000111",
  21761=>"011101011",
  21762=>"001111111",
  21763=>"000011001",
  21764=>"000001100",
  21765=>"111010011",
  21766=>"101101001",
  21767=>"101001110",
  21768=>"101111101",
  21769=>"100100011",
  21770=>"100111010",
  21771=>"101100010",
  21772=>"010111101",
  21773=>"011111010",
  21774=>"110111110",
  21775=>"000011110",
  21776=>"001000101",
  21777=>"101011100",
  21778=>"010000101",
  21779=>"000100001",
  21780=>"001101001",
  21781=>"000011101",
  21782=>"110101001",
  21783=>"100111010",
  21784=>"001101100",
  21785=>"101010111",
  21786=>"011110001",
  21787=>"010011110",
  21788=>"000110000",
  21789=>"011001001",
  21790=>"100001100",
  21791=>"100111110",
  21792=>"010000000",
  21793=>"111001000",
  21794=>"001110101",
  21795=>"000011100",
  21796=>"001100010",
  21797=>"111001111",
  21798=>"110110100",
  21799=>"101101010",
  21800=>"101001100",
  21801=>"101110000",
  21802=>"100001111",
  21803=>"111101101",
  21804=>"100100111",
  21805=>"000001001",
  21806=>"101010111",
  21807=>"010000001",
  21808=>"110100010",
  21809=>"111110111",
  21810=>"111000011",
  21811=>"111001101",
  21812=>"101001110",
  21813=>"101111101",
  21814=>"010100111",
  21815=>"101110000",
  21816=>"110110011",
  21817=>"110010111",
  21818=>"110000010",
  21819=>"100110010",
  21820=>"000001011",
  21821=>"101010101",
  21822=>"111001111",
  21823=>"101100100",
  21824=>"101111101",
  21825=>"011110010",
  21826=>"000010010",
  21827=>"011101011",
  21828=>"000101000",
  21829=>"111101111",
  21830=>"111010100",
  21831=>"111010011",
  21832=>"000011110",
  21833=>"101010110",
  21834=>"111100111",
  21835=>"011101101",
  21836=>"110001110",
  21837=>"110011010",
  21838=>"111011001",
  21839=>"101101000",
  21840=>"010010101",
  21841=>"101100011",
  21842=>"110100101",
  21843=>"001101011",
  21844=>"011100101",
  21845=>"111010001",
  21846=>"111000010",
  21847=>"100101000",
  21848=>"111100101",
  21849=>"010011111",
  21850=>"011111110",
  21851=>"100010111",
  21852=>"010011000",
  21853=>"111100101",
  21854=>"101110111",
  21855=>"111000000",
  21856=>"000000010",
  21857=>"011010010",
  21858=>"100011101",
  21859=>"011110000",
  21860=>"000111110",
  21861=>"111110110",
  21862=>"110110111",
  21863=>"011101010",
  21864=>"110111011",
  21865=>"011100000",
  21866=>"011111100",
  21867=>"000001010",
  21868=>"111101011",
  21869=>"011110011",
  21870=>"110100101",
  21871=>"101000010",
  21872=>"100000010",
  21873=>"001011001",
  21874=>"011101001",
  21875=>"101011100",
  21876=>"101010001",
  21877=>"010100101",
  21878=>"010101111",
  21879=>"000001001",
  21880=>"000010010",
  21881=>"110111111",
  21882=>"001111101",
  21883=>"101110111",
  21884=>"100100010",
  21885=>"110111000",
  21886=>"000011000",
  21887=>"000110010",
  21888=>"010011100",
  21889=>"011101111",
  21890=>"110001001",
  21891=>"100011101",
  21892=>"011100011",
  21893=>"010000000",
  21894=>"111111111",
  21895=>"001101101",
  21896=>"011111011",
  21897=>"100000111",
  21898=>"000100001",
  21899=>"000101100",
  21900=>"000001101",
  21901=>"111101110",
  21902=>"000001001",
  21903=>"100001011",
  21904=>"100101011",
  21905=>"111110101",
  21906=>"001011101",
  21907=>"101100111",
  21908=>"111110111",
  21909=>"100000000",
  21910=>"010001001",
  21911=>"100000010",
  21912=>"100100101",
  21913=>"000001110",
  21914=>"111001101",
  21915=>"011110100",
  21916=>"111010101",
  21917=>"001010110",
  21918=>"010000110",
  21919=>"110000100",
  21920=>"110000000",
  21921=>"100110010",
  21922=>"000101000",
  21923=>"001000110",
  21924=>"101110001",
  21925=>"011000101",
  21926=>"101101111",
  21927=>"010111010",
  21928=>"011010101",
  21929=>"001001100",
  21930=>"110001101",
  21931=>"000001001",
  21932=>"100000101",
  21933=>"110101111",
  21934=>"001110000",
  21935=>"000110111",
  21936=>"011101010",
  21937=>"111100001",
  21938=>"100100000",
  21939=>"001100000",
  21940=>"000100100",
  21941=>"100111111",
  21942=>"000010000",
  21943=>"110000011",
  21944=>"000101001",
  21945=>"111101110",
  21946=>"111010000",
  21947=>"101010100",
  21948=>"110000000",
  21949=>"100100001",
  21950=>"010011010",
  21951=>"010100100",
  21952=>"001110010",
  21953=>"101111101",
  21954=>"000100001",
  21955=>"111100110",
  21956=>"000010001",
  21957=>"101000101",
  21958=>"111101101",
  21959=>"110011011",
  21960=>"011010011",
  21961=>"011001001",
  21962=>"100100001",
  21963=>"101101010",
  21964=>"110001011",
  21965=>"101101011",
  21966=>"000000010",
  21967=>"110111111",
  21968=>"100111111",
  21969=>"111111101",
  21970=>"110000100",
  21971=>"001111111",
  21972=>"110001011",
  21973=>"010001111",
  21974=>"000000001",
  21975=>"100011101",
  21976=>"001010010",
  21977=>"100111111",
  21978=>"110011100",
  21979=>"001000111",
  21980=>"111010100",
  21981=>"100011111",
  21982=>"000110001",
  21983=>"101100011",
  21984=>"100110110",
  21985=>"111011101",
  21986=>"011101111",
  21987=>"110101010",
  21988=>"100111101",
  21989=>"010011010",
  21990=>"001001001",
  21991=>"001110001",
  21992=>"101011100",
  21993=>"000100101",
  21994=>"011001010",
  21995=>"010110101",
  21996=>"001010000",
  21997=>"101001010",
  21998=>"110111111",
  21999=>"111101100",
  22000=>"101001010",
  22001=>"001010000",
  22002=>"001010110",
  22003=>"001100001",
  22004=>"010011010",
  22005=>"001101111",
  22006=>"100001111",
  22007=>"000111011",
  22008=>"110001000",
  22009=>"010101011",
  22010=>"001011010",
  22011=>"100010101",
  22012=>"101100001",
  22013=>"100101101",
  22014=>"000101010",
  22015=>"011000010",
  22016=>"001100110",
  22017=>"100001110",
  22018=>"110011100",
  22019=>"100110000",
  22020=>"000111100",
  22021=>"100100101",
  22022=>"100101111",
  22023=>"001110110",
  22024=>"100111111",
  22025=>"110100000",
  22026=>"010100010",
  22027=>"001101001",
  22028=>"110111010",
  22029=>"000000110",
  22030=>"001010100",
  22031=>"111111110",
  22032=>"110100110",
  22033=>"110111111",
  22034=>"100001110",
  22035=>"001100111",
  22036=>"101000001",
  22037=>"110011110",
  22038=>"011000110",
  22039=>"010110001",
  22040=>"001000010",
  22041=>"000001010",
  22042=>"010001001",
  22043=>"111000001",
  22044=>"111111110",
  22045=>"111100001",
  22046=>"000101110",
  22047=>"000101110",
  22048=>"110101101",
  22049=>"000001001",
  22050=>"011010110",
  22051=>"000011010",
  22052=>"011001100",
  22053=>"000000110",
  22054=>"001000010",
  22055=>"101111001",
  22056=>"101110001",
  22057=>"011001000",
  22058=>"010101010",
  22059=>"011110101",
  22060=>"010101010",
  22061=>"000010100",
  22062=>"000100001",
  22063=>"010011011",
  22064=>"000001111",
  22065=>"110000001",
  22066=>"111001101",
  22067=>"111001101",
  22068=>"101110001",
  22069=>"101010100",
  22070=>"011011101",
  22071=>"001011011",
  22072=>"110110001",
  22073=>"110001111",
  22074=>"000111100",
  22075=>"110001010",
  22076=>"111110110",
  22077=>"011100011",
  22078=>"111000111",
  22079=>"000110011",
  22080=>"111100100",
  22081=>"100010110",
  22082=>"000010100",
  22083=>"011111110",
  22084=>"100001111",
  22085=>"000111101",
  22086=>"001001001",
  22087=>"111111011",
  22088=>"001111011",
  22089=>"101110100",
  22090=>"000110110",
  22091=>"110111100",
  22092=>"101010110",
  22093=>"001001101",
  22094=>"010000001",
  22095=>"100100000",
  22096=>"110011100",
  22097=>"110100011",
  22098=>"011011001",
  22099=>"110010001",
  22100=>"011000001",
  22101=>"000000110",
  22102=>"100111110",
  22103=>"101100011",
  22104=>"111101000",
  22105=>"101101010",
  22106=>"111111111",
  22107=>"111101001",
  22108=>"000001111",
  22109=>"111010111",
  22110=>"111101110",
  22111=>"010110011",
  22112=>"111100101",
  22113=>"110000010",
  22114=>"001001100",
  22115=>"000100000",
  22116=>"101110011",
  22117=>"010101001",
  22118=>"000101001",
  22119=>"011100000",
  22120=>"000011111",
  22121=>"100011001",
  22122=>"111100011",
  22123=>"100010001",
  22124=>"011000011",
  22125=>"100101100",
  22126=>"101100101",
  22127=>"111111000",
  22128=>"011011100",
  22129=>"100101011",
  22130=>"001000110",
  22131=>"001101010",
  22132=>"010001111",
  22133=>"010101101",
  22134=>"101111001",
  22135=>"101011000",
  22136=>"011111011",
  22137=>"100010001",
  22138=>"000001001",
  22139=>"111111111",
  22140=>"010011000",
  22141=>"001101000",
  22142=>"111010010",
  22143=>"101001000",
  22144=>"000011011",
  22145=>"000011110",
  22146=>"101011100",
  22147=>"000101001",
  22148=>"100000010",
  22149=>"001000001",
  22150=>"001100101",
  22151=>"111100111",
  22152=>"010010001",
  22153=>"010001111",
  22154=>"011110100",
  22155=>"110000010",
  22156=>"111101000",
  22157=>"101101100",
  22158=>"110001110",
  22159=>"001100110",
  22160=>"101111011",
  22161=>"101111100",
  22162=>"101101001",
  22163=>"111101111",
  22164=>"000001011",
  22165=>"111110101",
  22166=>"110100101",
  22167=>"011001101",
  22168=>"001101100",
  22169=>"001111001",
  22170=>"010100100",
  22171=>"001000001",
  22172=>"100000101",
  22173=>"010011110",
  22174=>"100000111",
  22175=>"010100101",
  22176=>"100111010",
  22177=>"110000010",
  22178=>"100011100",
  22179=>"100011110",
  22180=>"010011010",
  22181=>"101000011",
  22182=>"101000111",
  22183=>"101101000",
  22184=>"010111111",
  22185=>"110111001",
  22186=>"010000010",
  22187=>"111001110",
  22188=>"111000110",
  22189=>"001111001",
  22190=>"001111000",
  22191=>"100011000",
  22192=>"100100000",
  22193=>"101011111",
  22194=>"001110101",
  22195=>"100000011",
  22196=>"101010001",
  22197=>"100000001",
  22198=>"011001001",
  22199=>"101111110",
  22200=>"101101100",
  22201=>"000110111",
  22202=>"101111011",
  22203=>"101001111",
  22204=>"100110010",
  22205=>"110100111",
  22206=>"001101011",
  22207=>"100001001",
  22208=>"101100110",
  22209=>"011010000",
  22210=>"011000010",
  22211=>"011011111",
  22212=>"101010110",
  22213=>"110011010",
  22214=>"001001100",
  22215=>"100100000",
  22216=>"100001000",
  22217=>"010110000",
  22218=>"101111111",
  22219=>"010110100",
  22220=>"011100110",
  22221=>"110010000",
  22222=>"011011001",
  22223=>"011101111",
  22224=>"011001010",
  22225=>"111011101",
  22226=>"101011001",
  22227=>"001100111",
  22228=>"000000000",
  22229=>"100011100",
  22230=>"101000000",
  22231=>"110011100",
  22232=>"011101110",
  22233=>"000101000",
  22234=>"111000010",
  22235=>"101100010",
  22236=>"111000011",
  22237=>"000001101",
  22238=>"100011110",
  22239=>"101011010",
  22240=>"101000000",
  22241=>"001101001",
  22242=>"001000001",
  22243=>"110000010",
  22244=>"010110010",
  22245=>"001001111",
  22246=>"010111110",
  22247=>"010001001",
  22248=>"111000101",
  22249=>"000010101",
  22250=>"011111100",
  22251=>"110110000",
  22252=>"111011000",
  22253=>"110100000",
  22254=>"101110000",
  22255=>"001111000",
  22256=>"000010100",
  22257=>"100101001",
  22258=>"110000010",
  22259=>"110111100",
  22260=>"011110011",
  22261=>"111011011",
  22262=>"110001011",
  22263=>"111011000",
  22264=>"001111101",
  22265=>"011101001",
  22266=>"111111111",
  22267=>"011010010",
  22268=>"100101000",
  22269=>"101100111",
  22270=>"010110110",
  22271=>"101011000",
  22272=>"010001101",
  22273=>"011100111",
  22274=>"011011111",
  22275=>"010101011",
  22276=>"111111001",
  22277=>"100001101",
  22278=>"100010110",
  22279=>"101010110",
  22280=>"010100010",
  22281=>"001101101",
  22282=>"100001000",
  22283=>"100111110",
  22284=>"011000011",
  22285=>"010111011",
  22286=>"110000010",
  22287=>"011111000",
  22288=>"100001101",
  22289=>"011100001",
  22290=>"110011000",
  22291=>"100011000",
  22292=>"110111111",
  22293=>"010100000",
  22294=>"010110010",
  22295=>"111110101",
  22296=>"000100010",
  22297=>"000001010",
  22298=>"110001000",
  22299=>"111111011",
  22300=>"011101010",
  22301=>"111010011",
  22302=>"010101100",
  22303=>"110111010",
  22304=>"010010111",
  22305=>"001100001",
  22306=>"101010001",
  22307=>"000111110",
  22308=>"010010110",
  22309=>"011110011",
  22310=>"010001110",
  22311=>"010110110",
  22312=>"011011010",
  22313=>"000100010",
  22314=>"100001001",
  22315=>"001000000",
  22316=>"010110001",
  22317=>"000101000",
  22318=>"000110110",
  22319=>"011100010",
  22320=>"001000100",
  22321=>"111110100",
  22322=>"101111111",
  22323=>"101111010",
  22324=>"111000010",
  22325=>"110000111",
  22326=>"000001100",
  22327=>"100101100",
  22328=>"111011101",
  22329=>"000101011",
  22330=>"001100101",
  22331=>"111101010",
  22332=>"001100000",
  22333=>"101110001",
  22334=>"101011101",
  22335=>"111111110",
  22336=>"001001011",
  22337=>"000010000",
  22338=>"100100010",
  22339=>"001100000",
  22340=>"011000100",
  22341=>"100001110",
  22342=>"101101100",
  22343=>"101101110",
  22344=>"100111001",
  22345=>"110001111",
  22346=>"100110011",
  22347=>"000000101",
  22348=>"010110010",
  22349=>"010011001",
  22350=>"110001101",
  22351=>"000011100",
  22352=>"111011010",
  22353=>"111000001",
  22354=>"000000111",
  22355=>"000001001",
  22356=>"101000101",
  22357=>"000110110",
  22358=>"101101100",
  22359=>"010011111",
  22360=>"010010101",
  22361=>"100010100",
  22362=>"101111010",
  22363=>"100001000",
  22364=>"011011011",
  22365=>"010111110",
  22366=>"010100110",
  22367=>"101011010",
  22368=>"100010100",
  22369=>"011101010",
  22370=>"000110100",
  22371=>"111100111",
  22372=>"001011010",
  22373=>"011000000",
  22374=>"000010000",
  22375=>"011100111",
  22376=>"011000001",
  22377=>"000000110",
  22378=>"011100110",
  22379=>"111001111",
  22380=>"000000110",
  22381=>"010011111",
  22382=>"101110001",
  22383=>"100101101",
  22384=>"010101101",
  22385=>"111101011",
  22386=>"101000110",
  22387=>"011101111",
  22388=>"111011101",
  22389=>"001100101",
  22390=>"111011011",
  22391=>"100111111",
  22392=>"001010010",
  22393=>"111000110",
  22394=>"100000000",
  22395=>"011100111",
  22396=>"110001100",
  22397=>"011010101",
  22398=>"001000001",
  22399=>"010100000",
  22400=>"001001010",
  22401=>"101010011",
  22402=>"111000101",
  22403=>"010010001",
  22404=>"110000110",
  22405=>"111011001",
  22406=>"100100110",
  22407=>"001110011",
  22408=>"110100010",
  22409=>"101001000",
  22410=>"000010111",
  22411=>"011110111",
  22412=>"001111011",
  22413=>"101000000",
  22414=>"001001100",
  22415=>"110101111",
  22416=>"000101001",
  22417=>"010100111",
  22418=>"100111011",
  22419=>"100000001",
  22420=>"010000001",
  22421=>"110101011",
  22422=>"111111010",
  22423=>"001010101",
  22424=>"001000100",
  22425=>"000000111",
  22426=>"101110000",
  22427=>"000001111",
  22428=>"010000110",
  22429=>"000000111",
  22430=>"001101100",
  22431=>"000011010",
  22432=>"101110011",
  22433=>"011101111",
  22434=>"100001010",
  22435=>"011011011",
  22436=>"110010010",
  22437=>"011001100",
  22438=>"011011010",
  22439=>"111000100",
  22440=>"101000100",
  22441=>"111111101",
  22442=>"100000011",
  22443=>"111100001",
  22444=>"101010110",
  22445=>"111101000",
  22446=>"001010101",
  22447=>"010001111",
  22448=>"010111011",
  22449=>"110100010",
  22450=>"111101100",
  22451=>"000000100",
  22452=>"111001000",
  22453=>"100111110",
  22454=>"010100001",
  22455=>"010000001",
  22456=>"010000110",
  22457=>"101100110",
  22458=>"000110110",
  22459=>"111010001",
  22460=>"110111011",
  22461=>"111111011",
  22462=>"010000011",
  22463=>"110111110",
  22464=>"010111101",
  22465=>"000100110",
  22466=>"110100110",
  22467=>"100100101",
  22468=>"101011101",
  22469=>"111100001",
  22470=>"100010010",
  22471=>"010101011",
  22472=>"110101111",
  22473=>"100100100",
  22474=>"000110011",
  22475=>"101100100",
  22476=>"011010100",
  22477=>"110011100",
  22478=>"011111100",
  22479=>"110011100",
  22480=>"010010010",
  22481=>"011110011",
  22482=>"000001001",
  22483=>"000001110",
  22484=>"010001111",
  22485=>"001000001",
  22486=>"011010001",
  22487=>"110111010",
  22488=>"100101101",
  22489=>"110011110",
  22490=>"011100111",
  22491=>"111111011",
  22492=>"001010001",
  22493=>"011010100",
  22494=>"000010000",
  22495=>"101000110",
  22496=>"100000100",
  22497=>"011111110",
  22498=>"111010101",
  22499=>"011000011",
  22500=>"000111000",
  22501=>"101001101",
  22502=>"101101001",
  22503=>"111010001",
  22504=>"100000010",
  22505=>"100000011",
  22506=>"110000101",
  22507=>"011111010",
  22508=>"001000101",
  22509=>"110110100",
  22510=>"001000100",
  22511=>"100110110",
  22512=>"000100100",
  22513=>"110001100",
  22514=>"001011110",
  22515=>"110011110",
  22516=>"110110110",
  22517=>"001101011",
  22518=>"000101001",
  22519=>"010001100",
  22520=>"011111001",
  22521=>"111111111",
  22522=>"101111101",
  22523=>"010100101",
  22524=>"001000001",
  22525=>"010100011",
  22526=>"111101111",
  22527=>"000011010",
  22528=>"010010001",
  22529=>"001010011",
  22530=>"111100011",
  22531=>"111011110",
  22532=>"101101001",
  22533=>"111011101",
  22534=>"100100101",
  22535=>"011111101",
  22536=>"001010010",
  22537=>"110001111",
  22538=>"110111111",
  22539=>"011100100",
  22540=>"011000101",
  22541=>"001010001",
  22542=>"001110110",
  22543=>"111100100",
  22544=>"010001100",
  22545=>"111100010",
  22546=>"111111011",
  22547=>"100011000",
  22548=>"110010100",
  22549=>"010001111",
  22550=>"000011111",
  22551=>"001001100",
  22552=>"011010001",
  22553=>"010111111",
  22554=>"001011001",
  22555=>"000100110",
  22556=>"110011100",
  22557=>"101011011",
  22558=>"011110001",
  22559=>"011011010",
  22560=>"011000010",
  22561=>"000110110",
  22562=>"011110111",
  22563=>"011100111",
  22564=>"110101001",
  22565=>"000100011",
  22566=>"100011001",
  22567=>"110010000",
  22568=>"001001011",
  22569=>"101010100",
  22570=>"001001000",
  22571=>"010101001",
  22572=>"101111110",
  22573=>"111000100",
  22574=>"001011100",
  22575=>"001001010",
  22576=>"110011110",
  22577=>"000001110",
  22578=>"101101010",
  22579=>"000011000",
  22580=>"001001100",
  22581=>"001111010",
  22582=>"000000010",
  22583=>"100100111",
  22584=>"001000001",
  22585=>"101011111",
  22586=>"100000001",
  22587=>"111001111",
  22588=>"100101000",
  22589=>"101111110",
  22590=>"000110011",
  22591=>"001101111",
  22592=>"000100010",
  22593=>"100100100",
  22594=>"111110011",
  22595=>"111101010",
  22596=>"001001100",
  22597=>"111011000",
  22598=>"100001000",
  22599=>"000000100",
  22600=>"111010001",
  22601=>"101111001",
  22602=>"111101000",
  22603=>"111001011",
  22604=>"110000000",
  22605=>"111001101",
  22606=>"110100101",
  22607=>"010100010",
  22608=>"111000011",
  22609=>"100010011",
  22610=>"100011111",
  22611=>"101010101",
  22612=>"100111010",
  22613=>"001111011",
  22614=>"101100000",
  22615=>"100111100",
  22616=>"110101010",
  22617=>"110111100",
  22618=>"111111101",
  22619=>"000001001",
  22620=>"111101110",
  22621=>"101111011",
  22622=>"000110111",
  22623=>"100101101",
  22624=>"010001001",
  22625=>"100101100",
  22626=>"101101101",
  22627=>"011001000",
  22628=>"011001001",
  22629=>"001110111",
  22630=>"011001110",
  22631=>"101000101",
  22632=>"010000011",
  22633=>"011111011",
  22634=>"010001100",
  22635=>"001010011",
  22636=>"010001010",
  22637=>"110111010",
  22638=>"110100001",
  22639=>"101000101",
  22640=>"001100001",
  22641=>"001101111",
  22642=>"100111011",
  22643=>"111111011",
  22644=>"011010101",
  22645=>"110100100",
  22646=>"000101010",
  22647=>"010111111",
  22648=>"110001100",
  22649=>"010001001",
  22650=>"010110110",
  22651=>"100101110",
  22652=>"100110011",
  22653=>"001001101",
  22654=>"011010011",
  22655=>"110011100",
  22656=>"000110101",
  22657=>"000100111",
  22658=>"100000111",
  22659=>"001010011",
  22660=>"100101101",
  22661=>"010101110",
  22662=>"101011000",
  22663=>"011010001",
  22664=>"001000001",
  22665=>"000011001",
  22666=>"101010000",
  22667=>"011010110",
  22668=>"001101001",
  22669=>"010101101",
  22670=>"101010111",
  22671=>"111011001",
  22672=>"010111011",
  22673=>"110111011",
  22674=>"000000111",
  22675=>"110011100",
  22676=>"011010000",
  22677=>"101000110",
  22678=>"111000100",
  22679=>"101100101",
  22680=>"011010011",
  22681=>"000001010",
  22682=>"100011111",
  22683=>"000100111",
  22684=>"010101010",
  22685=>"100100001",
  22686=>"001000001",
  22687=>"110010110",
  22688=>"110111011",
  22689=>"000000100",
  22690=>"110000100",
  22691=>"111001110",
  22692=>"101110111",
  22693=>"101000011",
  22694=>"000100011",
  22695=>"001001011",
  22696=>"110011100",
  22697=>"011000111",
  22698=>"001100110",
  22699=>"000010010",
  22700=>"011001011",
  22701=>"111010011",
  22702=>"011001101",
  22703=>"111000001",
  22704=>"010000110",
  22705=>"011101011",
  22706=>"000000111",
  22707=>"000101000",
  22708=>"000010000",
  22709=>"111000111",
  22710=>"000100101",
  22711=>"101100101",
  22712=>"100000110",
  22713=>"000100101",
  22714=>"101001110",
  22715=>"111111111",
  22716=>"110011010",
  22717=>"010010100",
  22718=>"111010101",
  22719=>"110111111",
  22720=>"011101101",
  22721=>"001001100",
  22722=>"101000000",
  22723=>"010000010",
  22724=>"111111000",
  22725=>"010001010",
  22726=>"101101111",
  22727=>"111010100",
  22728=>"100100111",
  22729=>"000110011",
  22730=>"010010111",
  22731=>"011110111",
  22732=>"011110000",
  22733=>"010011101",
  22734=>"000001010",
  22735=>"000000001",
  22736=>"000011101",
  22737=>"010100000",
  22738=>"000001100",
  22739=>"011010001",
  22740=>"000010011",
  22741=>"000101011",
  22742=>"111011011",
  22743=>"001000010",
  22744=>"110100001",
  22745=>"100101111",
  22746=>"010100111",
  22747=>"110010011",
  22748=>"111001101",
  22749=>"100010000",
  22750=>"101101000",
  22751=>"010111100",
  22752=>"010001010",
  22753=>"001111000",
  22754=>"011110111",
  22755=>"001011111",
  22756=>"101111101",
  22757=>"110111011",
  22758=>"001000011",
  22759=>"100111010",
  22760=>"100010100",
  22761=>"001010000",
  22762=>"001101010",
  22763=>"100001111",
  22764=>"101010000",
  22765=>"000001101",
  22766=>"101100111",
  22767=>"000000100",
  22768=>"110011100",
  22769=>"111111101",
  22770=>"000110000",
  22771=>"011100010",
  22772=>"111100100",
  22773=>"110000001",
  22774=>"100011101",
  22775=>"000001010",
  22776=>"011110000",
  22777=>"000001000",
  22778=>"101000010",
  22779=>"000001100",
  22780=>"000001110",
  22781=>"000111010",
  22782=>"000110101",
  22783=>"101101100",
  22784=>"101100001",
  22785=>"000010101",
  22786=>"100010110",
  22787=>"101111001",
  22788=>"001000010",
  22789=>"101101101",
  22790=>"100000000",
  22791=>"011100000",
  22792=>"000000010",
  22793=>"101000111",
  22794=>"010111110",
  22795=>"110001001",
  22796=>"011110101",
  22797=>"110000000",
  22798=>"011010101",
  22799=>"000110001",
  22800=>"011000111",
  22801=>"111000100",
  22802=>"010101110",
  22803=>"000110010",
  22804=>"100001000",
  22805=>"000100111",
  22806=>"110111000",
  22807=>"110101111",
  22808=>"110110000",
  22809=>"101110010",
  22810=>"101000101",
  22811=>"000100010",
  22812=>"001011101",
  22813=>"111001110",
  22814=>"011111001",
  22815=>"101000100",
  22816=>"000110011",
  22817=>"001110001",
  22818=>"011001001",
  22819=>"001100010",
  22820=>"101000010",
  22821=>"001111111",
  22822=>"110000010",
  22823=>"101110001",
  22824=>"110011001",
  22825=>"011010001",
  22826=>"001100110",
  22827=>"100011010",
  22828=>"010001111",
  22829=>"000011100",
  22830=>"100100000",
  22831=>"101010011",
  22832=>"000111010",
  22833=>"010010011",
  22834=>"110000101",
  22835=>"100101001",
  22836=>"100000011",
  22837=>"101100001",
  22838=>"101010101",
  22839=>"100001110",
  22840=>"010100000",
  22841=>"011110101",
  22842=>"100111101",
  22843=>"110100001",
  22844=>"100000001",
  22845=>"010010010",
  22846=>"100011101",
  22847=>"111111100",
  22848=>"100111101",
  22849=>"100000010",
  22850=>"010000110",
  22851=>"110111000",
  22852=>"010111010",
  22853=>"110111111",
  22854=>"001000000",
  22855=>"111110110",
  22856=>"110101110",
  22857=>"001010001",
  22858=>"100101011",
  22859=>"100111110",
  22860=>"111101101",
  22861=>"110101101",
  22862=>"111011001",
  22863=>"001010010",
  22864=>"101000010",
  22865=>"111001100",
  22866=>"110111001",
  22867=>"101001101",
  22868=>"010101000",
  22869=>"100110011",
  22870=>"010110011",
  22871=>"110111101",
  22872=>"100100001",
  22873=>"000011110",
  22874=>"000101110",
  22875=>"111100101",
  22876=>"111100000",
  22877=>"111010010",
  22878=>"101000011",
  22879=>"000110010",
  22880=>"101010010",
  22881=>"001010100",
  22882=>"000000100",
  22883=>"000100011",
  22884=>"111111111",
  22885=>"011100101",
  22886=>"101001010",
  22887=>"011000100",
  22888=>"000001010",
  22889=>"000001000",
  22890=>"001101100",
  22891=>"101011011",
  22892=>"011001101",
  22893=>"000110011",
  22894=>"100110001",
  22895=>"001000100",
  22896=>"000011101",
  22897=>"100100100",
  22898=>"010010111",
  22899=>"111001111",
  22900=>"001000111",
  22901=>"111011100",
  22902=>"011100100",
  22903=>"001100110",
  22904=>"110111111",
  22905=>"101110111",
  22906=>"000010001",
  22907=>"010110111",
  22908=>"011010011",
  22909=>"101101110",
  22910=>"010000011",
  22911=>"010100111",
  22912=>"110101001",
  22913=>"111101001",
  22914=>"011011011",
  22915=>"000010100",
  22916=>"011000001",
  22917=>"101100100",
  22918=>"011101011",
  22919=>"000001011",
  22920=>"011110100",
  22921=>"011010111",
  22922=>"110000110",
  22923=>"101001111",
  22924=>"000010011",
  22925=>"111000111",
  22926=>"011001010",
  22927=>"000100001",
  22928=>"001010101",
  22929=>"001101101",
  22930=>"110011011",
  22931=>"001010111",
  22932=>"010100101",
  22933=>"111001101",
  22934=>"001010000",
  22935=>"000001001",
  22936=>"110000011",
  22937=>"110000000",
  22938=>"011111110",
  22939=>"000011000",
  22940=>"100001001",
  22941=>"100111010",
  22942=>"100100000",
  22943=>"110001011",
  22944=>"000001001",
  22945=>"010000000",
  22946=>"111011111",
  22947=>"000000111",
  22948=>"100101110",
  22949=>"000000001",
  22950=>"101111110",
  22951=>"110100101",
  22952=>"000110011",
  22953=>"111001000",
  22954=>"010010111",
  22955=>"011000101",
  22956=>"000000011",
  22957=>"011011111",
  22958=>"100001010",
  22959=>"010011101",
  22960=>"101100010",
  22961=>"001100110",
  22962=>"110000011",
  22963=>"001100111",
  22964=>"100001011",
  22965=>"111110001",
  22966=>"010010110",
  22967=>"100100100",
  22968=>"111000101",
  22969=>"000111111",
  22970=>"000110101",
  22971=>"111001111",
  22972=>"011000110",
  22973=>"111011000",
  22974=>"100011010",
  22975=>"110001011",
  22976=>"001010010",
  22977=>"101000001",
  22978=>"011111101",
  22979=>"000101111",
  22980=>"111011001",
  22981=>"000000011",
  22982=>"111100011",
  22983=>"011001001",
  22984=>"111100000",
  22985=>"000101111",
  22986=>"011110100",
  22987=>"001000001",
  22988=>"001100100",
  22989=>"111101000",
  22990=>"101010111",
  22991=>"011111000",
  22992=>"100100100",
  22993=>"110100101",
  22994=>"011100010",
  22995=>"001100100",
  22996=>"011001001",
  22997=>"100000100",
  22998=>"110111001",
  22999=>"101001100",
  23000=>"111101110",
  23001=>"110001110",
  23002=>"001111101",
  23003=>"010101010",
  23004=>"010011001",
  23005=>"101010011",
  23006=>"100111110",
  23007=>"100000001",
  23008=>"111100110",
  23009=>"011011100",
  23010=>"000100000",
  23011=>"100001000",
  23012=>"101110101",
  23013=>"011000100",
  23014=>"111111011",
  23015=>"111100000",
  23016=>"111111101",
  23017=>"100111110",
  23018=>"111010110",
  23019=>"100011101",
  23020=>"010110101",
  23021=>"100110110",
  23022=>"001010100",
  23023=>"111111110",
  23024=>"110100010",
  23025=>"101111111",
  23026=>"111111001",
  23027=>"101110001",
  23028=>"110000101",
  23029=>"011000000",
  23030=>"111101001",
  23031=>"010100000",
  23032=>"000010010",
  23033=>"100101110",
  23034=>"111100101",
  23035=>"101110011",
  23036=>"011101000",
  23037=>"001011101",
  23038=>"010100101",
  23039=>"111100001",
  23040=>"000001010",
  23041=>"111111110",
  23042=>"000100011",
  23043=>"101111110",
  23044=>"001110010",
  23045=>"011010111",
  23046=>"111000001",
  23047=>"101011101",
  23048=>"010010011",
  23049=>"100100010",
  23050=>"101011110",
  23051=>"010100010",
  23052=>"001000111",
  23053=>"001111111",
  23054=>"001000101",
  23055=>"100111111",
  23056=>"001011010",
  23057=>"110101110",
  23058=>"001000000",
  23059=>"001100011",
  23060=>"011011101",
  23061=>"101110100",
  23062=>"011111010",
  23063=>"111101010",
  23064=>"001110101",
  23065=>"101101001",
  23066=>"011000010",
  23067=>"100100100",
  23068=>"000000011",
  23069=>"100100001",
  23070=>"111000000",
  23071=>"010000000",
  23072=>"010010000",
  23073=>"111100101",
  23074=>"001100011",
  23075=>"110111110",
  23076=>"011010001",
  23077=>"111000101",
  23078=>"011001110",
  23079=>"011100001",
  23080=>"110100111",
  23081=>"001010001",
  23082=>"001000000",
  23083=>"110011110",
  23084=>"110111101",
  23085=>"001110111",
  23086=>"010111110",
  23087=>"100101011",
  23088=>"011110011",
  23089=>"111110100",
  23090=>"000110111",
  23091=>"010001011",
  23092=>"011000111",
  23093=>"000010000",
  23094=>"100010100",
  23095=>"100101011",
  23096=>"001110101",
  23097=>"010110100",
  23098=>"100101010",
  23099=>"110011010",
  23100=>"001100010",
  23101=>"100000001",
  23102=>"000100110",
  23103=>"011110111",
  23104=>"000011111",
  23105=>"000110001",
  23106=>"001011011",
  23107=>"100000110",
  23108=>"011010011",
  23109=>"110000010",
  23110=>"111010101",
  23111=>"010001001",
  23112=>"010100100",
  23113=>"001011101",
  23114=>"101000111",
  23115=>"110011011",
  23116=>"110011010",
  23117=>"100101011",
  23118=>"111101111",
  23119=>"011011110",
  23120=>"111111011",
  23121=>"101110000",
  23122=>"111000111",
  23123=>"000101100",
  23124=>"100100010",
  23125=>"000110010",
  23126=>"010000000",
  23127=>"000111000",
  23128=>"010000100",
  23129=>"100000010",
  23130=>"101110011",
  23131=>"000001000",
  23132=>"000100110",
  23133=>"101010100",
  23134=>"100111100",
  23135=>"101010001",
  23136=>"101000111",
  23137=>"000000101",
  23138=>"101110101",
  23139=>"000001110",
  23140=>"111110111",
  23141=>"000110110",
  23142=>"111111011",
  23143=>"010001011",
  23144=>"010010100",
  23145=>"000011110",
  23146=>"010110011",
  23147=>"101010000",
  23148=>"001000100",
  23149=>"001000000",
  23150=>"010100011",
  23151=>"100100110",
  23152=>"101111000",
  23153=>"100010011",
  23154=>"000011011",
  23155=>"001100101",
  23156=>"011011011",
  23157=>"010100001",
  23158=>"111100010",
  23159=>"101101110",
  23160=>"101111111",
  23161=>"110101101",
  23162=>"111101001",
  23163=>"110111100",
  23164=>"011011010",
  23165=>"000111111",
  23166=>"010011011",
  23167=>"101011111",
  23168=>"000001100",
  23169=>"001011110",
  23170=>"001010011",
  23171=>"011101011",
  23172=>"100011101",
  23173=>"011101001",
  23174=>"011011101",
  23175=>"101100100",
  23176=>"000101110",
  23177=>"001100111",
  23178=>"010101010",
  23179=>"100111101",
  23180=>"110001110",
  23181=>"100100000",
  23182=>"100100001",
  23183=>"101001101",
  23184=>"111110011",
  23185=>"110010010",
  23186=>"010100110",
  23187=>"000000111",
  23188=>"011100011",
  23189=>"110101110",
  23190=>"011000000",
  23191=>"000000101",
  23192=>"000110100",
  23193=>"100111000",
  23194=>"001000010",
  23195=>"111010010",
  23196=>"000000110",
  23197=>"101100110",
  23198=>"100000111",
  23199=>"001010100",
  23200=>"100010001",
  23201=>"000111011",
  23202=>"010011000",
  23203=>"001011100",
  23204=>"111001100",
  23205=>"001110100",
  23206=>"100110100",
  23207=>"001000000",
  23208=>"101001111",
  23209=>"111100001",
  23210=>"011010100",
  23211=>"000100010",
  23212=>"000100100",
  23213=>"001000000",
  23214=>"100011000",
  23215=>"011100101",
  23216=>"001001010",
  23217=>"011100011",
  23218=>"110000101",
  23219=>"011001100",
  23220=>"111011110",
  23221=>"011001100",
  23222=>"100010010",
  23223=>"111000110",
  23224=>"111010011",
  23225=>"100101010",
  23226=>"010011000",
  23227=>"011000101",
  23228=>"010101101",
  23229=>"011110101",
  23230=>"001100010",
  23231=>"011110011",
  23232=>"000011100",
  23233=>"011001110",
  23234=>"110011001",
  23235=>"110111110",
  23236=>"011110010",
  23237=>"100011000",
  23238=>"001010111",
  23239=>"101000010",
  23240=>"100001000",
  23241=>"110000100",
  23242=>"111110011",
  23243=>"001001000",
  23244=>"100000001",
  23245=>"101111110",
  23246=>"000001011",
  23247=>"110111111",
  23248=>"000010010",
  23249=>"111001001",
  23250=>"011011000",
  23251=>"111000010",
  23252=>"011101111",
  23253=>"100100101",
  23254=>"011101110",
  23255=>"111101100",
  23256=>"010001001",
  23257=>"110001011",
  23258=>"100100110",
  23259=>"010100000",
  23260=>"101100101",
  23261=>"000001011",
  23262=>"111110010",
  23263=>"110111000",
  23264=>"100101011",
  23265=>"101010100",
  23266=>"110000111",
  23267=>"110100001",
  23268=>"101101100",
  23269=>"001101111",
  23270=>"000011000",
  23271=>"001001010",
  23272=>"001001110",
  23273=>"001011010",
  23274=>"001100000",
  23275=>"110111100",
  23276=>"110100111",
  23277=>"001011010",
  23278=>"001110100",
  23279=>"000110010",
  23280=>"100110000",
  23281=>"000000001",
  23282=>"110010100",
  23283=>"110000000",
  23284=>"010001010",
  23285=>"100100101",
  23286=>"000001000",
  23287=>"111110000",
  23288=>"011111011",
  23289=>"000011011",
  23290=>"001011111",
  23291=>"000001011",
  23292=>"110011000",
  23293=>"101001011",
  23294=>"100101111",
  23295=>"111111010",
  23296=>"101111100",
  23297=>"101000110",
  23298=>"111101010",
  23299=>"000101011",
  23300=>"111001000",
  23301=>"111100101",
  23302=>"100001101",
  23303=>"011110100",
  23304=>"111100101",
  23305=>"000010111",
  23306=>"001100010",
  23307=>"111100101",
  23308=>"100100001",
  23309=>"101111101",
  23310=>"011100001",
  23311=>"111100110",
  23312=>"101110111",
  23313=>"001110100",
  23314=>"100111100",
  23315=>"110010100",
  23316=>"101100001",
  23317=>"001010000",
  23318=>"100010010",
  23319=>"111111101",
  23320=>"001101101",
  23321=>"111101010",
  23322=>"100100011",
  23323=>"100000000",
  23324=>"011010000",
  23325=>"101011110",
  23326=>"011111100",
  23327=>"000010101",
  23328=>"000011011",
  23329=>"110110011",
  23330=>"011000001",
  23331=>"100010001",
  23332=>"101000100",
  23333=>"100000010",
  23334=>"000111101",
  23335=>"101101010",
  23336=>"101111101",
  23337=>"111110000",
  23338=>"001000100",
  23339=>"111100010",
  23340=>"110101001",
  23341=>"111100101",
  23342=>"101110110",
  23343=>"100100001",
  23344=>"000101110",
  23345=>"101011111",
  23346=>"101001000",
  23347=>"100111101",
  23348=>"111101111",
  23349=>"001000111",
  23350=>"011011110",
  23351=>"000100010",
  23352=>"100111011",
  23353=>"001100100",
  23354=>"011100000",
  23355=>"000101100",
  23356=>"011111011",
  23357=>"110000010",
  23358=>"110000000",
  23359=>"011110011",
  23360=>"100110000",
  23361=>"001011000",
  23362=>"011010011",
  23363=>"010010110",
  23364=>"110111111",
  23365=>"010110000",
  23366=>"111111000",
  23367=>"011101001",
  23368=>"100111101",
  23369=>"010011001",
  23370=>"101110111",
  23371=>"010110001",
  23372=>"100100011",
  23373=>"110101001",
  23374=>"110100101",
  23375=>"100101111",
  23376=>"111110101",
  23377=>"010100101",
  23378=>"011101001",
  23379=>"011011100",
  23380=>"001010111",
  23381=>"000101110",
  23382=>"110100110",
  23383=>"001100011",
  23384=>"110100101",
  23385=>"110011100",
  23386=>"011010001",
  23387=>"000000110",
  23388=>"100010101",
  23389=>"100100101",
  23390=>"100011011",
  23391=>"100001111",
  23392=>"001101010",
  23393=>"010011111",
  23394=>"001100011",
  23395=>"000101101",
  23396=>"011010011",
  23397=>"000001000",
  23398=>"011010011",
  23399=>"101101000",
  23400=>"010100000",
  23401=>"010000001",
  23402=>"110001001",
  23403=>"001100100",
  23404=>"010001010",
  23405=>"010010010",
  23406=>"110101001",
  23407=>"110010000",
  23408=>"001011110",
  23409=>"111011100",
  23410=>"000010001",
  23411=>"011010000",
  23412=>"111101111",
  23413=>"000110000",
  23414=>"111010001",
  23415=>"001101001",
  23416=>"101001011",
  23417=>"101010110",
  23418=>"111110111",
  23419=>"011000110",
  23420=>"110010011",
  23421=>"001101011",
  23422=>"111111100",
  23423=>"011011110",
  23424=>"110010001",
  23425=>"011100100",
  23426=>"010000101",
  23427=>"010111101",
  23428=>"100011100",
  23429=>"110010000",
  23430=>"100010010",
  23431=>"110001000",
  23432=>"101100100",
  23433=>"010001001",
  23434=>"001100011",
  23435=>"100000100",
  23436=>"111001100",
  23437=>"101110010",
  23438=>"110010011",
  23439=>"111000011",
  23440=>"111110111",
  23441=>"111011010",
  23442=>"010101000",
  23443=>"010111001",
  23444=>"110011010",
  23445=>"110100101",
  23446=>"010011010",
  23447=>"001101110",
  23448=>"110000111",
  23449=>"101011100",
  23450=>"100011011",
  23451=>"011110001",
  23452=>"010010100",
  23453=>"100000110",
  23454=>"111110010",
  23455=>"111000100",
  23456=>"001010000",
  23457=>"101111111",
  23458=>"100011100",
  23459=>"000101111",
  23460=>"101010000",
  23461=>"111011111",
  23462=>"000110011",
  23463=>"100101100",
  23464=>"100001000",
  23465=>"101011001",
  23466=>"110111001",
  23467=>"111100000",
  23468=>"001111101",
  23469=>"001000010",
  23470=>"110000000",
  23471=>"000001001",
  23472=>"011100000",
  23473=>"010011111",
  23474=>"011110010",
  23475=>"010110011",
  23476=>"100101100",
  23477=>"111101011",
  23478=>"001001111",
  23479=>"110010010",
  23480=>"111110100",
  23481=>"000110111",
  23482=>"100011001",
  23483=>"001110010",
  23484=>"000101111",
  23485=>"111110011",
  23486=>"010000001",
  23487=>"001110010",
  23488=>"011101011",
  23489=>"001000001",
  23490=>"100111001",
  23491=>"100000110",
  23492=>"000100011",
  23493=>"101000110",
  23494=>"101011111",
  23495=>"111011010",
  23496=>"000110110",
  23497=>"100010110",
  23498=>"110111010",
  23499=>"010110111",
  23500=>"001111101",
  23501=>"010100110",
  23502=>"000111111",
  23503=>"110110000",
  23504=>"111110101",
  23505=>"111010001",
  23506=>"011110010",
  23507=>"100101001",
  23508=>"111010010",
  23509=>"000000001",
  23510=>"101111011",
  23511=>"000110101",
  23512=>"100101010",
  23513=>"011000100",
  23514=>"010000110",
  23515=>"100001010",
  23516=>"101000100",
  23517=>"001011001",
  23518=>"110111101",
  23519=>"101101100",
  23520=>"101000001",
  23521=>"110001011",
  23522=>"111100100",
  23523=>"010101010",
  23524=>"011010000",
  23525=>"010001100",
  23526=>"000111001",
  23527=>"111100010",
  23528=>"101000000",
  23529=>"001001011",
  23530=>"110111010",
  23531=>"100010100",
  23532=>"001110111",
  23533=>"100000011",
  23534=>"001101110",
  23535=>"111010101",
  23536=>"111011111",
  23537=>"101100000",
  23538=>"010101110",
  23539=>"101001010",
  23540=>"101000001",
  23541=>"010000111",
  23542=>"000101010",
  23543=>"011000011",
  23544=>"011101111",
  23545=>"111110000",
  23546=>"010001000",
  23547=>"001111011",
  23548=>"100011001",
  23549=>"010111100",
  23550=>"000011001",
  23551=>"011111010",
  23552=>"011111100",
  23553=>"100111010",
  23554=>"001101001",
  23555=>"110011011",
  23556=>"100110111",
  23557=>"111111010",
  23558=>"000110110",
  23559=>"101011101",
  23560=>"001011101",
  23561=>"110100000",
  23562=>"100000110",
  23563=>"111010011",
  23564=>"111000001",
  23565=>"110110011",
  23566=>"001010001",
  23567=>"101001000",
  23568=>"111110110",
  23569=>"111111001",
  23570=>"111100000",
  23571=>"111000111",
  23572=>"001000100",
  23573=>"110000000",
  23574=>"110001110",
  23575=>"000001010",
  23576=>"000100001",
  23577=>"011000111",
  23578=>"101101100",
  23579=>"111010111",
  23580=>"010110111",
  23581=>"010101010",
  23582=>"011000000",
  23583=>"100000101",
  23584=>"111110111",
  23585=>"101101111",
  23586=>"010111000",
  23587=>"010011000",
  23588=>"101001101",
  23589=>"011110000",
  23590=>"110110000",
  23591=>"010101111",
  23592=>"111100000",
  23593=>"000000110",
  23594=>"000011001",
  23595=>"011110110",
  23596=>"111110101",
  23597=>"110101100",
  23598=>"111010010",
  23599=>"011100000",
  23600=>"010100100",
  23601=>"001110100",
  23602=>"100100001",
  23603=>"101000010",
  23604=>"011100011",
  23605=>"101010000",
  23606=>"100110110",
  23607=>"001101111",
  23608=>"100101001",
  23609=>"111111110",
  23610=>"101100111",
  23611=>"101011101",
  23612=>"110001010",
  23613=>"010100000",
  23614=>"110010110",
  23615=>"000100110",
  23616=>"001000010",
  23617=>"000010000",
  23618=>"111001111",
  23619=>"010001000",
  23620=>"100001111",
  23621=>"001001000",
  23622=>"110101011",
  23623=>"001011010",
  23624=>"111010110",
  23625=>"010100101",
  23626=>"000000110",
  23627=>"100011110",
  23628=>"010000111",
  23629=>"001110111",
  23630=>"010101111",
  23631=>"101101011",
  23632=>"011111000",
  23633=>"000111000",
  23634=>"000111110",
  23635=>"010001110",
  23636=>"000111010",
  23637=>"101101001",
  23638=>"000000010",
  23639=>"000000100",
  23640=>"100000100",
  23641=>"111111011",
  23642=>"000101110",
  23643=>"111100100",
  23644=>"110001100",
  23645=>"000000100",
  23646=>"101111001",
  23647=>"000101000",
  23648=>"101000001",
  23649=>"011101100",
  23650=>"011011011",
  23651=>"011010111",
  23652=>"101011100",
  23653=>"100101101",
  23654=>"010110110",
  23655=>"000000101",
  23656=>"100010110",
  23657=>"101000111",
  23658=>"000011101",
  23659=>"100110000",
  23660=>"010100011",
  23661=>"001100010",
  23662=>"000110001",
  23663=>"011101111",
  23664=>"000001110",
  23665=>"000000101",
  23666=>"001001101",
  23667=>"111101000",
  23668=>"101000110",
  23669=>"101111010",
  23670=>"110100110",
  23671=>"010000011",
  23672=>"000100111",
  23673=>"010111111",
  23674=>"000010110",
  23675=>"100010100",
  23676=>"110101011",
  23677=>"000000011",
  23678=>"101001000",
  23679=>"001101111",
  23680=>"100001100",
  23681=>"101010010",
  23682=>"011001001",
  23683=>"011010100",
  23684=>"000110100",
  23685=>"101001110",
  23686=>"110010010",
  23687=>"010101110",
  23688=>"111101110",
  23689=>"001011100",
  23690=>"001010011",
  23691=>"100010100",
  23692=>"001010100",
  23693=>"111010100",
  23694=>"111000111",
  23695=>"111010001",
  23696=>"001101101",
  23697=>"100010101",
  23698=>"010011000",
  23699=>"010101101",
  23700=>"010010110",
  23701=>"001110000",
  23702=>"111010010",
  23703=>"000000101",
  23704=>"010010010",
  23705=>"011110110",
  23706=>"100011001",
  23707=>"111011001",
  23708=>"000111111",
  23709=>"100111101",
  23710=>"111000000",
  23711=>"110000010",
  23712=>"010100000",
  23713=>"000111100",
  23714=>"001001100",
  23715=>"110010011",
  23716=>"111101011",
  23717=>"000010010",
  23718=>"011110101",
  23719=>"000100110",
  23720=>"100001100",
  23721=>"010000111",
  23722=>"000001101",
  23723=>"011101011",
  23724=>"010110110",
  23725=>"001110100",
  23726=>"000110000",
  23727=>"011011000",
  23728=>"011011001",
  23729=>"011111100",
  23730=>"011110110",
  23731=>"000000101",
  23732=>"101110000",
  23733=>"101000110",
  23734=>"000010111",
  23735=>"111110101",
  23736=>"100000101",
  23737=>"000001110",
  23738=>"011101100",
  23739=>"000010011",
  23740=>"111010111",
  23741=>"000111110",
  23742=>"000001010",
  23743=>"101000011",
  23744=>"101010101",
  23745=>"110011000",
  23746=>"110110101",
  23747=>"110101010",
  23748=>"110010111",
  23749=>"100010111",
  23750=>"100100001",
  23751=>"000000111",
  23752=>"111101111",
  23753=>"100101000",
  23754=>"010010101",
  23755=>"010000000",
  23756=>"100011111",
  23757=>"010011000",
  23758=>"111110011",
  23759=>"011111011",
  23760=>"101001111",
  23761=>"011000101",
  23762=>"001111100",
  23763=>"100000011",
  23764=>"110001001",
  23765=>"111100010",
  23766=>"011101111",
  23767=>"000100110",
  23768=>"110010000",
  23769=>"110110100",
  23770=>"000001101",
  23771=>"101110000",
  23772=>"110000110",
  23773=>"111011111",
  23774=>"101101011",
  23775=>"111100000",
  23776=>"010011101",
  23777=>"011111100",
  23778=>"100011011",
  23779=>"010100010",
  23780=>"100100001",
  23781=>"101010010",
  23782=>"011100001",
  23783=>"100100011",
  23784=>"010010111",
  23785=>"101001101",
  23786=>"001011011",
  23787=>"001001110",
  23788=>"100100001",
  23789=>"101000110",
  23790=>"011000010",
  23791=>"100110001",
  23792=>"111001110",
  23793=>"101111100",
  23794=>"001011111",
  23795=>"110101010",
  23796=>"011110110",
  23797=>"000111001",
  23798=>"001001010",
  23799=>"001000001",
  23800=>"011001110",
  23801=>"101110111",
  23802=>"111111101",
  23803=>"101110000",
  23804=>"010000011",
  23805=>"111001101",
  23806=>"110010100",
  23807=>"001111000",
  23808=>"011101100",
  23809=>"000011000",
  23810=>"111000100",
  23811=>"000000000",
  23812=>"011001110",
  23813=>"011111111",
  23814=>"010010000",
  23815=>"111111111",
  23816=>"000010011",
  23817=>"101100110",
  23818=>"000111100",
  23819=>"010111100",
  23820=>"111110001",
  23821=>"100100010",
  23822=>"001011100",
  23823=>"101010100",
  23824=>"111101110",
  23825=>"100101010",
  23826=>"101001001",
  23827=>"101011101",
  23828=>"100110001",
  23829=>"110011011",
  23830=>"110100100",
  23831=>"010111110",
  23832=>"011110011",
  23833=>"111110100",
  23834=>"010000110",
  23835=>"111100010",
  23836=>"100111000",
  23837=>"100010010",
  23838=>"011001101",
  23839=>"111011110",
  23840=>"100101100",
  23841=>"010011010",
  23842=>"001001111",
  23843=>"010100100",
  23844=>"011110101",
  23845=>"111110011",
  23846=>"111010010",
  23847=>"101010111",
  23848=>"100110000",
  23849=>"100101001",
  23850=>"010100001",
  23851=>"011011010",
  23852=>"111111000",
  23853=>"010100100",
  23854=>"011010011",
  23855=>"000110010",
  23856=>"001000100",
  23857=>"110001111",
  23858=>"110101010",
  23859=>"100100010",
  23860=>"110000010",
  23861=>"101001001",
  23862=>"001111010",
  23863=>"011010111",
  23864=>"000000001",
  23865=>"010100000",
  23866=>"001001100",
  23867=>"110100010",
  23868=>"101111101",
  23869=>"010010011",
  23870=>"111011000",
  23871=>"000101110",
  23872=>"011011001",
  23873=>"000000101",
  23874=>"110111111",
  23875=>"001110111",
  23876=>"110001111",
  23877=>"101101011",
  23878=>"110101010",
  23879=>"110000000",
  23880=>"101000110",
  23881=>"100111000",
  23882=>"010111110",
  23883=>"100000100",
  23884=>"100010010",
  23885=>"011011000",
  23886=>"001010110",
  23887=>"010100010",
  23888=>"111111100",
  23889=>"001111101",
  23890=>"110100011",
  23891=>"110001101",
  23892=>"101110101",
  23893=>"010010110",
  23894=>"010101100",
  23895=>"000110010",
  23896=>"000010000",
  23897=>"010110110",
  23898=>"101111011",
  23899=>"001001111",
  23900=>"010011111",
  23901=>"100000100",
  23902=>"111111010",
  23903=>"010011011",
  23904=>"101110110",
  23905=>"010100011",
  23906=>"111100001",
  23907=>"101111011",
  23908=>"000010101",
  23909=>"110110011",
  23910=>"111001000",
  23911=>"110100010",
  23912=>"000100110",
  23913=>"011100011",
  23914=>"111011000",
  23915=>"101100000",
  23916=>"000010101",
  23917=>"011101010",
  23918=>"001010001",
  23919=>"110010100",
  23920=>"100000000",
  23921=>"100010001",
  23922=>"010000011",
  23923=>"100100010",
  23924=>"000111100",
  23925=>"101101000",
  23926=>"011011110",
  23927=>"101111001",
  23928=>"001101000",
  23929=>"001011100",
  23930=>"100111111",
  23931=>"110110010",
  23932=>"101101100",
  23933=>"011101111",
  23934=>"100100110",
  23935=>"100010011",
  23936=>"000111001",
  23937=>"010100010",
  23938=>"100000000",
  23939=>"111000110",
  23940=>"010011010",
  23941=>"101100110",
  23942=>"111110110",
  23943=>"100110010",
  23944=>"101110100",
  23945=>"011101000",
  23946=>"110011000",
  23947=>"010000010",
  23948=>"000101010",
  23949=>"110111110",
  23950=>"011100100",
  23951=>"011110101",
  23952=>"100110001",
  23953=>"101000100",
  23954=>"101010000",
  23955=>"100010110",
  23956=>"011010111",
  23957=>"000000110",
  23958=>"000010000",
  23959=>"111011010",
  23960=>"001100011",
  23961=>"001101011",
  23962=>"101101100",
  23963=>"000101001",
  23964=>"000110111",
  23965=>"010100110",
  23966=>"001110101",
  23967=>"011011111",
  23968=>"101100001",
  23969=>"100001000",
  23970=>"000011111",
  23971=>"110110001",
  23972=>"010011100",
  23973=>"000000000",
  23974=>"000101011",
  23975=>"100110001",
  23976=>"111110010",
  23977=>"111100010",
  23978=>"000100000",
  23979=>"100001001",
  23980=>"101000100",
  23981=>"100000001",
  23982=>"111101111",
  23983=>"111100001",
  23984=>"001110110",
  23985=>"001010110",
  23986=>"001100110",
  23987=>"111001010",
  23988=>"010101000",
  23989=>"101111111",
  23990=>"100010110",
  23991=>"010101010",
  23992=>"100101001",
  23993=>"111000110",
  23994=>"111010010",
  23995=>"101011011",
  23996=>"001011000",
  23997=>"100101001",
  23998=>"011001001",
  23999=>"010100100",
  24000=>"101010001",
  24001=>"000111100",
  24002=>"001011111",
  24003=>"011111110",
  24004=>"001000101",
  24005=>"111100100",
  24006=>"010011111",
  24007=>"100101011",
  24008=>"010001000",
  24009=>"100110100",
  24010=>"101000000",
  24011=>"100110111",
  24012=>"111111011",
  24013=>"001001010",
  24014=>"011111100",
  24015=>"110000011",
  24016=>"010101111",
  24017=>"010010000",
  24018=>"000100111",
  24019=>"100100101",
  24020=>"000001111",
  24021=>"000101101",
  24022=>"001111100",
  24023=>"010001000",
  24024=>"001011101",
  24025=>"001000110",
  24026=>"011101001",
  24027=>"010011101",
  24028=>"111110010",
  24029=>"111001111",
  24030=>"000001101",
  24031=>"001000010",
  24032=>"000010001",
  24033=>"110110111",
  24034=>"001111011",
  24035=>"111011001",
  24036=>"111010101",
  24037=>"000101111",
  24038=>"100100000",
  24039=>"001000001",
  24040=>"000010001",
  24041=>"001011101",
  24042=>"111000100",
  24043=>"101100001",
  24044=>"010101011",
  24045=>"100011011",
  24046=>"010111001",
  24047=>"111100001",
  24048=>"111001011",
  24049=>"011000111",
  24050=>"000111100",
  24051=>"000011101",
  24052=>"010110000",
  24053=>"010110110",
  24054=>"110111000",
  24055=>"011000100",
  24056=>"101000100",
  24057=>"010001100",
  24058=>"101011110",
  24059=>"000111100",
  24060=>"001001110",
  24061=>"110001000",
  24062=>"101101001",
  24063=>"111101000",
  24064=>"010011001",
  24065=>"101000101",
  24066=>"101011001",
  24067=>"010111111",
  24068=>"000000000",
  24069=>"001011000",
  24070=>"001010101",
  24071=>"111101100",
  24072=>"000000010",
  24073=>"100001110",
  24074=>"000100110",
  24075=>"010010101",
  24076=>"001101000",
  24077=>"100001101",
  24078=>"101000111",
  24079=>"110100001",
  24080=>"001110001",
  24081=>"100100100",
  24082=>"101101011",
  24083=>"101010011",
  24084=>"010011010",
  24085=>"101001100",
  24086=>"001010011",
  24087=>"010001001",
  24088=>"100011001",
  24089=>"011000101",
  24090=>"101001110",
  24091=>"110011011",
  24092=>"101001001",
  24093=>"111010101",
  24094=>"111110010",
  24095=>"010110110",
  24096=>"100000001",
  24097=>"000101011",
  24098=>"011010110",
  24099=>"010000100",
  24100=>"111110111",
  24101=>"100010100",
  24102=>"011001011",
  24103=>"111010000",
  24104=>"001010001",
  24105=>"100101110",
  24106=>"000011100",
  24107=>"100110110",
  24108=>"000111010",
  24109=>"101100110",
  24110=>"110001001",
  24111=>"101101001",
  24112=>"100101100",
  24113=>"101000011",
  24114=>"010100001",
  24115=>"000001111",
  24116=>"000000010",
  24117=>"001000010",
  24118=>"100011111",
  24119=>"101100101",
  24120=>"110010100",
  24121=>"000110101",
  24122=>"000001100",
  24123=>"100100100",
  24124=>"100101011",
  24125=>"111000001",
  24126=>"100100000",
  24127=>"101111110",
  24128=>"110001111",
  24129=>"111110100",
  24130=>"011000011",
  24131=>"011011110",
  24132=>"001111110",
  24133=>"101000111",
  24134=>"101100000",
  24135=>"000001000",
  24136=>"110010111",
  24137=>"010011111",
  24138=>"001001101",
  24139=>"001001001",
  24140=>"000000110",
  24141=>"001001101",
  24142=>"100001011",
  24143=>"010100000",
  24144=>"111101000",
  24145=>"100110001",
  24146=>"111100100",
  24147=>"111001111",
  24148=>"100101001",
  24149=>"100001010",
  24150=>"110001101",
  24151=>"101010111",
  24152=>"011000000",
  24153=>"010001100",
  24154=>"001111100",
  24155=>"111100101",
  24156=>"111110001",
  24157=>"100000001",
  24158=>"101111001",
  24159=>"010100101",
  24160=>"010101000",
  24161=>"001010010",
  24162=>"010010010",
  24163=>"001100101",
  24164=>"010110000",
  24165=>"011011011",
  24166=>"110011000",
  24167=>"001100010",
  24168=>"000101100",
  24169=>"101011100",
  24170=>"000110110",
  24171=>"110101000",
  24172=>"101011001",
  24173=>"011000001",
  24174=>"011101101",
  24175=>"100100000",
  24176=>"010110101",
  24177=>"101110111",
  24178=>"100111011",
  24179=>"110011011",
  24180=>"100001000",
  24181=>"111010000",
  24182=>"011011011",
  24183=>"000011001",
  24184=>"000111010",
  24185=>"100010011",
  24186=>"010100100",
  24187=>"110111110",
  24188=>"101011010",
  24189=>"011001000",
  24190=>"100010000",
  24191=>"001111111",
  24192=>"011101000",
  24193=>"000001101",
  24194=>"111011110",
  24195=>"101011001",
  24196=>"110101001",
  24197=>"110001101",
  24198=>"100011011",
  24199=>"010111101",
  24200=>"101110100",
  24201=>"101010101",
  24202=>"100011010",
  24203=>"000011001",
  24204=>"011101011",
  24205=>"111000111",
  24206=>"000111001",
  24207=>"001001000",
  24208=>"101110000",
  24209=>"111110101",
  24210=>"101000000",
  24211=>"001001011",
  24212=>"001111010",
  24213=>"010001111",
  24214=>"100001001",
  24215=>"111111110",
  24216=>"010100011",
  24217=>"011111111",
  24218=>"010011111",
  24219=>"010100111",
  24220=>"001100001",
  24221=>"101001111",
  24222=>"101001011",
  24223=>"101000000",
  24224=>"111001010",
  24225=>"001111001",
  24226=>"001100100",
  24227=>"100011100",
  24228=>"110111011",
  24229=>"011010110",
  24230=>"111100001",
  24231=>"000011100",
  24232=>"011110111",
  24233=>"111101110",
  24234=>"101001111",
  24235=>"000101010",
  24236=>"100110010",
  24237=>"000011100",
  24238=>"100011110",
  24239=>"010010111",
  24240=>"100111101",
  24241=>"000010000",
  24242=>"000010010",
  24243=>"110111000",
  24244=>"010100010",
  24245=>"111111001",
  24246=>"111100111",
  24247=>"011111010",
  24248=>"111110110",
  24249=>"100001100",
  24250=>"011111100",
  24251=>"100111111",
  24252=>"010000011",
  24253=>"000010011",
  24254=>"101000000",
  24255=>"010111001",
  24256=>"111000111",
  24257=>"111010111",
  24258=>"111111100",
  24259=>"011000010",
  24260=>"010000110",
  24261=>"001110110",
  24262=>"101010100",
  24263=>"100110111",
  24264=>"010001000",
  24265=>"010111000",
  24266=>"001110111",
  24267=>"001111001",
  24268=>"101111110",
  24269=>"011101011",
  24270=>"111011011",
  24271=>"111011000",
  24272=>"100010110",
  24273=>"100010101",
  24274=>"101011001",
  24275=>"101000100",
  24276=>"110100110",
  24277=>"101100010",
  24278=>"010100111",
  24279=>"101011010",
  24280=>"000000001",
  24281=>"010001011",
  24282=>"111101101",
  24283=>"111100111",
  24284=>"011101101",
  24285=>"111001010",
  24286=>"010111100",
  24287=>"001101110",
  24288=>"110000010",
  24289=>"000010111",
  24290=>"000100101",
  24291=>"000010111",
  24292=>"011100110",
  24293=>"100010111",
  24294=>"000100000",
  24295=>"111101110",
  24296=>"000100110",
  24297=>"111110111",
  24298=>"011001111",
  24299=>"001100111",
  24300=>"010000110",
  24301=>"000000111",
  24302=>"001000100",
  24303=>"110010101",
  24304=>"110100101",
  24305=>"000011110",
  24306=>"001010000",
  24307=>"111110001",
  24308=>"101011110",
  24309=>"111110010",
  24310=>"000010010",
  24311=>"111101010",
  24312=>"011100110",
  24313=>"101100010",
  24314=>"001111110",
  24315=>"100110110",
  24316=>"000100001",
  24317=>"100100110",
  24318=>"001000000",
  24319=>"011101110",
  24320=>"010100011",
  24321=>"000101101",
  24322=>"101111100",
  24323=>"000100101",
  24324=>"011001101",
  24325=>"111000000",
  24326=>"110001000",
  24327=>"111111101",
  24328=>"100101110",
  24329=>"011011110",
  24330=>"100000011",
  24331=>"110100101",
  24332=>"001100010",
  24333=>"111001011",
  24334=>"011000010",
  24335=>"101111000",
  24336=>"110111010",
  24337=>"011000100",
  24338=>"100010000",
  24339=>"001011100",
  24340=>"010000101",
  24341=>"000110101",
  24342=>"010111001",
  24343=>"010111101",
  24344=>"010000000",
  24345=>"110100111",
  24346=>"100010011",
  24347=>"011111011",
  24348=>"001111010",
  24349=>"010001101",
  24350=>"110111110",
  24351=>"011101111",
  24352=>"000001100",
  24353=>"110001001",
  24354=>"100010110",
  24355=>"100110010",
  24356=>"000011000",
  24357=>"101011101",
  24358=>"001100010",
  24359=>"100000001",
  24360=>"000010110",
  24361=>"100111111",
  24362=>"100110011",
  24363=>"100101100",
  24364=>"100110001",
  24365=>"000001101",
  24366=>"011001011",
  24367=>"000100101",
  24368=>"000000000",
  24369=>"100000000",
  24370=>"110100011",
  24371=>"111110000",
  24372=>"111001110",
  24373=>"110010010",
  24374=>"101011100",
  24375=>"111000100",
  24376=>"101111001",
  24377=>"100000110",
  24378=>"111001111",
  24379=>"111001001",
  24380=>"010101000",
  24381=>"101100101",
  24382=>"001101111",
  24383=>"110111110",
  24384=>"111111001",
  24385=>"110010011",
  24386=>"100101101",
  24387=>"110100101",
  24388=>"100011110",
  24389=>"000111011",
  24390=>"010101010",
  24391=>"110001111",
  24392=>"110010110",
  24393=>"011010010",
  24394=>"111000111",
  24395=>"001000100",
  24396=>"101001101",
  24397=>"001100011",
  24398=>"100101010",
  24399=>"111111010",
  24400=>"000001101",
  24401=>"000101011",
  24402=>"101000101",
  24403=>"111100111",
  24404=>"101001101",
  24405=>"001001001",
  24406=>"100111011",
  24407=>"001001010",
  24408=>"100000011",
  24409=>"011101111",
  24410=>"101010110",
  24411=>"100011001",
  24412=>"110011011",
  24413=>"001101000",
  24414=>"100110100",
  24415=>"001000001",
  24416=>"111111110",
  24417=>"100011011",
  24418=>"001100000",
  24419=>"011010110",
  24420=>"101111011",
  24421=>"010101010",
  24422=>"100100101",
  24423=>"011001100",
  24424=>"110010000",
  24425=>"010110001",
  24426=>"001101110",
  24427=>"111000011",
  24428=>"000100001",
  24429=>"000001110",
  24430=>"111000101",
  24431=>"110100011",
  24432=>"011001100",
  24433=>"000011001",
  24434=>"010011001",
  24435=>"100000010",
  24436=>"001001011",
  24437=>"111100001",
  24438=>"010000111",
  24439=>"011111001",
  24440=>"000101100",
  24441=>"000000001",
  24442=>"000000011",
  24443=>"111010010",
  24444=>"011011010",
  24445=>"010100011",
  24446=>"000000000",
  24447=>"000111010",
  24448=>"001011110",
  24449=>"010001001",
  24450=>"000110110",
  24451=>"011000000",
  24452=>"000110010",
  24453=>"101010111",
  24454=>"010110101",
  24455=>"110000010",
  24456=>"010010110",
  24457=>"010111000",
  24458=>"100001111",
  24459=>"011101111",
  24460=>"011110001",
  24461=>"111111100",
  24462=>"010000100",
  24463=>"001000100",
  24464=>"100101011",
  24465=>"111010100",
  24466=>"111101101",
  24467=>"110100100",
  24468=>"111110111",
  24469=>"101111010",
  24470=>"011001010",
  24471=>"000011000",
  24472=>"011011101",
  24473=>"000101000",
  24474=>"010010000",
  24475=>"001001000",
  24476=>"000101001",
  24477=>"010111111",
  24478=>"101000010",
  24479=>"011111010",
  24480=>"000100110",
  24481=>"100100111",
  24482=>"000000110",
  24483=>"110100100",
  24484=>"011011001",
  24485=>"100010110",
  24486=>"010000100",
  24487=>"111001110",
  24488=>"010011101",
  24489=>"010100010",
  24490=>"010000010",
  24491=>"101000100",
  24492=>"000110000",
  24493=>"110011110",
  24494=>"111011011",
  24495=>"111111110",
  24496=>"000111111",
  24497=>"110100111",
  24498=>"101000100",
  24499=>"010010000",
  24500=>"001111111",
  24501=>"100100100",
  24502=>"000110100",
  24503=>"011110010",
  24504=>"100101001",
  24505=>"011111011",
  24506=>"101011110",
  24507=>"001000011",
  24508=>"111101000",
  24509=>"011100101",
  24510=>"111111111",
  24511=>"000000001",
  24512=>"010101100",
  24513=>"100000101",
  24514=>"101001110",
  24515=>"000100001",
  24516=>"111111111",
  24517=>"101001001",
  24518=>"111100101",
  24519=>"001010111",
  24520=>"111000110",
  24521=>"111110110",
  24522=>"100000100",
  24523=>"011000100",
  24524=>"101000100",
  24525=>"001001110",
  24526=>"001010110",
  24527=>"101101100",
  24528=>"010111000",
  24529=>"101011011",
  24530=>"000100001",
  24531=>"011001011",
  24532=>"101000111",
  24533=>"101010000",
  24534=>"100000111",
  24535=>"101001011",
  24536=>"000010010",
  24537=>"000011110",
  24538=>"011100000",
  24539=>"111000110",
  24540=>"010010101",
  24541=>"101100111",
  24542=>"100011011",
  24543=>"000001111",
  24544=>"100100010",
  24545=>"110000110",
  24546=>"000011000",
  24547=>"000010011",
  24548=>"010011010",
  24549=>"010000001",
  24550=>"100010010",
  24551=>"111100101",
  24552=>"011001001",
  24553=>"001100001",
  24554=>"101101001",
  24555=>"000010101",
  24556=>"001101101",
  24557=>"100100110",
  24558=>"011011011",
  24559=>"101111000",
  24560=>"110110010",
  24561=>"001010111",
  24562=>"110000010",
  24563=>"010010010",
  24564=>"111110011",
  24565=>"000100011",
  24566=>"100100110",
  24567=>"110110100",
  24568=>"111010011",
  24569=>"101001100",
  24570=>"101001111",
  24571=>"111001010",
  24572=>"100000100",
  24573=>"110111001",
  24574=>"101000011",
  24575=>"110000001",
  24576=>"101101111",
  24577=>"001101111",
  24578=>"010011011",
  24579=>"110111111",
  24580=>"011000100",
  24581=>"011001000",
  24582=>"110100101",
  24583=>"000000000",
  24584=>"001010011",
  24585=>"111010011",
  24586=>"101101011",
  24587=>"010111010",
  24588=>"100010111",
  24589=>"001101010",
  24590=>"011000000",
  24591=>"110000010",
  24592=>"011011101",
  24593=>"110110110",
  24594=>"000001010",
  24595=>"011000101",
  24596=>"001111011",
  24597=>"000101010",
  24598=>"011111001",
  24599=>"001101111",
  24600=>"101011000",
  24601=>"110101010",
  24602=>"110000100",
  24603=>"100010111",
  24604=>"100010000",
  24605=>"011001101",
  24606=>"000000001",
  24607=>"100000110",
  24608=>"100000010",
  24609=>"110110100",
  24610=>"010111000",
  24611=>"011010111",
  24612=>"010110100",
  24613=>"000110001",
  24614=>"111111100",
  24615=>"100001100",
  24616=>"110100000",
  24617=>"001101111",
  24618=>"111101111",
  24619=>"100010110",
  24620=>"110001111",
  24621=>"011000010",
  24622=>"110100111",
  24623=>"100001101",
  24624=>"001010010",
  24625=>"010111100",
  24626=>"011000010",
  24627=>"000010001",
  24628=>"101111000",
  24629=>"011010001",
  24630=>"010101110",
  24631=>"010000111",
  24632=>"001101111",
  24633=>"011101010",
  24634=>"101010100",
  24635=>"110100110",
  24636=>"010111111",
  24637=>"111110100",
  24638=>"100001100",
  24639=>"111001010",
  24640=>"011000100",
  24641=>"010010011",
  24642=>"000000010",
  24643=>"100101110",
  24644=>"101000110",
  24645=>"010111111",
  24646=>"001111110",
  24647=>"001100000",
  24648=>"100101011",
  24649=>"111110110",
  24650=>"111100100",
  24651=>"000001001",
  24652=>"101001111",
  24653=>"011011110",
  24654=>"000001101",
  24655=>"110011111",
  24656=>"110010001",
  24657=>"101000010",
  24658=>"001000001",
  24659=>"101111001",
  24660=>"001111100",
  24661=>"101000110",
  24662=>"011011101",
  24663=>"111001101",
  24664=>"101110111",
  24665=>"110110001",
  24666=>"010111110",
  24667=>"011111110",
  24668=>"100110010",
  24669=>"100100101",
  24670=>"111110011",
  24671=>"110010111",
  24672=>"110000011",
  24673=>"011001011",
  24674=>"111010001",
  24675=>"010001101",
  24676=>"010100101",
  24677=>"011101001",
  24678=>"111010101",
  24679=>"111110000",
  24680=>"001001100",
  24681=>"011100100",
  24682=>"010101000",
  24683=>"111000101",
  24684=>"110101101",
  24685=>"110010111",
  24686=>"101010001",
  24687=>"011011000",
  24688=>"101111111",
  24689=>"110100000",
  24690=>"110100000",
  24691=>"100111001",
  24692=>"101000100",
  24693=>"010010100",
  24694=>"110111110",
  24695=>"111011101",
  24696=>"010010001",
  24697=>"100110001",
  24698=>"101111111",
  24699=>"011000010",
  24700=>"111100101",
  24701=>"001110011",
  24702=>"111110110",
  24703=>"001111111",
  24704=>"101100110",
  24705=>"001010111",
  24706=>"111011101",
  24707=>"110000010",
  24708=>"001110000",
  24709=>"111000001",
  24710=>"010101010",
  24711=>"100111001",
  24712=>"111100111",
  24713=>"100100100",
  24714=>"101001010",
  24715=>"001111011",
  24716=>"001001010",
  24717=>"010111101",
  24718=>"000101101",
  24719=>"000101111",
  24720=>"111101001",
  24721=>"001100100",
  24722=>"001010100",
  24723=>"001110100",
  24724=>"111011110",
  24725=>"001111010",
  24726=>"010000110",
  24727=>"011100110",
  24728=>"110010101",
  24729=>"110010100",
  24730=>"000010101",
  24731=>"000110101",
  24732=>"010111011",
  24733=>"100100111",
  24734=>"010010110",
  24735=>"100110110",
  24736=>"001000011",
  24737=>"110111100",
  24738=>"000001010",
  24739=>"010001010",
  24740=>"000110100",
  24741=>"001101000",
  24742=>"101110111",
  24743=>"010000110",
  24744=>"101101000",
  24745=>"000000111",
  24746=>"011111111",
  24747=>"000010101",
  24748=>"111110011",
  24749=>"110111101",
  24750=>"100010011",
  24751=>"110101000",
  24752=>"000011001",
  24753=>"110000001",
  24754=>"111100110",
  24755=>"101011000",
  24756=>"001101110",
  24757=>"011000111",
  24758=>"000101101",
  24759=>"001010110",
  24760=>"000010100",
  24761=>"010101001",
  24762=>"010001100",
  24763=>"011110000",
  24764=>"000110100",
  24765=>"010001001",
  24766=>"100101101",
  24767=>"000010101",
  24768=>"100011011",
  24769=>"010010001",
  24770=>"011100101",
  24771=>"011001010",
  24772=>"100110111",
  24773=>"000001001",
  24774=>"000000001",
  24775=>"100001000",
  24776=>"101010011",
  24777=>"110101000",
  24778=>"011000111",
  24779=>"001110001",
  24780=>"000100010",
  24781=>"001100010",
  24782=>"101001011",
  24783=>"001011110",
  24784=>"100010000",
  24785=>"101111100",
  24786=>"101010100",
  24787=>"110001000",
  24788=>"010111000",
  24789=>"111011110",
  24790=>"010111110",
  24791=>"111110001",
  24792=>"100000101",
  24793=>"000110101",
  24794=>"101100000",
  24795=>"111100100",
  24796=>"111100111",
  24797=>"010011110",
  24798=>"000011011",
  24799=>"000000100",
  24800=>"100110111",
  24801=>"000110100",
  24802=>"101101101",
  24803=>"010010100",
  24804=>"100010101",
  24805=>"011010101",
  24806=>"101100011",
  24807=>"000010100",
  24808=>"110000001",
  24809=>"001010110",
  24810=>"111111110",
  24811=>"111101111",
  24812=>"101110110",
  24813=>"101100010",
  24814=>"010101011",
  24815=>"001001010",
  24816=>"011000100",
  24817=>"010010101",
  24818=>"001000000",
  24819=>"100001110",
  24820=>"000000111",
  24821=>"110111101",
  24822=>"101011110",
  24823=>"011110101",
  24824=>"100111000",
  24825=>"100000000",
  24826=>"100010011",
  24827=>"000110000",
  24828=>"011000000",
  24829=>"101101111",
  24830=>"010010110",
  24831=>"000000111",
  24832=>"111001001",
  24833=>"010111001",
  24834=>"001101011",
  24835=>"010110101",
  24836=>"101100100",
  24837=>"100111011",
  24838=>"110111011",
  24839=>"011101010",
  24840=>"110011000",
  24841=>"101101110",
  24842=>"110001110",
  24843=>"001000100",
  24844=>"000001111",
  24845=>"001110110",
  24846=>"000110001",
  24847=>"111010000",
  24848=>"010101110",
  24849=>"000000110",
  24850=>"001101100",
  24851=>"011111101",
  24852=>"111101011",
  24853=>"101011111",
  24854=>"000101000",
  24855=>"101001101",
  24856=>"110101111",
  24857=>"111011110",
  24858=>"010010000",
  24859=>"101010111",
  24860=>"100111101",
  24861=>"011101011",
  24862=>"111101011",
  24863=>"001000000",
  24864=>"010111111",
  24865=>"000101000",
  24866=>"011001100",
  24867=>"110111101",
  24868=>"100001100",
  24869=>"011101001",
  24870=>"000010110",
  24871=>"001011100",
  24872=>"010001011",
  24873=>"110100110",
  24874=>"101111001",
  24875=>"011000011",
  24876=>"010010000",
  24877=>"011010111",
  24878=>"101110111",
  24879=>"000110011",
  24880=>"011000001",
  24881=>"000101111",
  24882=>"011011000",
  24883=>"101011101",
  24884=>"001010100",
  24885=>"110011100",
  24886=>"101010000",
  24887=>"100000111",
  24888=>"101011011",
  24889=>"011111111",
  24890=>"101101010",
  24891=>"001011000",
  24892=>"111110000",
  24893=>"111000100",
  24894=>"111111111",
  24895=>"010111010",
  24896=>"010010011",
  24897=>"010001100",
  24898=>"110110100",
  24899=>"111100000",
  24900=>"001100111",
  24901=>"001101000",
  24902=>"101110000",
  24903=>"111110010",
  24904=>"011110111",
  24905=>"101011101",
  24906=>"010011011",
  24907=>"000001011",
  24908=>"010100001",
  24909=>"000011000",
  24910=>"101001011",
  24911=>"011110011",
  24912=>"000101111",
  24913=>"001100100",
  24914=>"000001011",
  24915=>"111101010",
  24916=>"101011011",
  24917=>"101011101",
  24918=>"010000100",
  24919=>"000011000",
  24920=>"011000111",
  24921=>"001101010",
  24922=>"100011101",
  24923=>"001011000",
  24924=>"011001110",
  24925=>"100100000",
  24926=>"101000011",
  24927=>"000001001",
  24928=>"101000010",
  24929=>"111010111",
  24930=>"100101110",
  24931=>"111000010",
  24932=>"000111111",
  24933=>"111001100",
  24934=>"101110010",
  24935=>"011111101",
  24936=>"101010101",
  24937=>"101110001",
  24938=>"110111100",
  24939=>"000010000",
  24940=>"010000001",
  24941=>"000000111",
  24942=>"010000011",
  24943=>"111001000",
  24944=>"110111101",
  24945=>"011001001",
  24946=>"010010010",
  24947=>"111000000",
  24948=>"011000000",
  24949=>"101011110",
  24950=>"101011010",
  24951=>"101100000",
  24952=>"101001011",
  24953=>"100100110",
  24954=>"000100011",
  24955=>"110111011",
  24956=>"000111001",
  24957=>"101011011",
  24958=>"110000101",
  24959=>"011111011",
  24960=>"101100101",
  24961=>"010001000",
  24962=>"010001110",
  24963=>"101000001",
  24964=>"010101100",
  24965=>"110101101",
  24966=>"011111001",
  24967=>"000001110",
  24968=>"011000001",
  24969=>"111000110",
  24970=>"110110100",
  24971=>"111101111",
  24972=>"111011111",
  24973=>"010000000",
  24974=>"111011111",
  24975=>"101110111",
  24976=>"011011100",
  24977=>"000110111",
  24978=>"000001001",
  24979=>"111100000",
  24980=>"110101010",
  24981=>"000000111",
  24982=>"111001011",
  24983=>"010110010",
  24984=>"000100010",
  24985=>"110011011",
  24986=>"101010000",
  24987=>"000100111",
  24988=>"001110101",
  24989=>"000010100",
  24990=>"111111000",
  24991=>"100110100",
  24992=>"001111010",
  24993=>"010100111",
  24994=>"111101111",
  24995=>"011111100",
  24996=>"010010111",
  24997=>"100010000",
  24998=>"000100100",
  24999=>"111100000",
  25000=>"010011001",
  25001=>"010101100",
  25002=>"110110010",
  25003=>"110100000",
  25004=>"011111011",
  25005=>"001110110",
  25006=>"101100010",
  25007=>"111110010",
  25008=>"111010100",
  25009=>"001001011",
  25010=>"101010100",
  25011=>"011001010",
  25012=>"011011001",
  25013=>"111111010",
  25014=>"111101101",
  25015=>"000111011",
  25016=>"110111100",
  25017=>"010010000",
  25018=>"101101101",
  25019=>"100100110",
  25020=>"101000111",
  25021=>"010110001",
  25022=>"001110100",
  25023=>"000000000",
  25024=>"101101001",
  25025=>"001011001",
  25026=>"000001001",
  25027=>"110111110",
  25028=>"110000000",
  25029=>"000011101",
  25030=>"010100011",
  25031=>"010000001",
  25032=>"011000111",
  25033=>"001010110",
  25034=>"110100000",
  25035=>"110110011",
  25036=>"001110001",
  25037=>"010000100",
  25038=>"000000111",
  25039=>"010001110",
  25040=>"110110001",
  25041=>"001100101",
  25042=>"001001101",
  25043=>"111110111",
  25044=>"010100110",
  25045=>"010111001",
  25046=>"110011101",
  25047=>"011111011",
  25048=>"001000010",
  25049=>"000111101",
  25050=>"110111110",
  25051=>"011101010",
  25052=>"100000100",
  25053=>"110110011",
  25054=>"101001101",
  25055=>"101001000",
  25056=>"100010011",
  25057=>"011001000",
  25058=>"110110110",
  25059=>"100100100",
  25060=>"101110100",
  25061=>"001101100",
  25062=>"011010100",
  25063=>"110011110",
  25064=>"001110001",
  25065=>"001011000",
  25066=>"011011000",
  25067=>"001110101",
  25068=>"111010011",
  25069=>"001101110",
  25070=>"011110111",
  25071=>"100010001",
  25072=>"111010011",
  25073=>"100111011",
  25074=>"000000110",
  25075=>"101111011",
  25076=>"010100011",
  25077=>"000101010",
  25078=>"001011100",
  25079=>"100010010",
  25080=>"000000111",
  25081=>"011101110",
  25082=>"111011001",
  25083=>"000101111",
  25084=>"001011100",
  25085=>"011001101",
  25086=>"110010111",
  25087=>"000011001",
  25088=>"101110000",
  25089=>"011000010",
  25090=>"111100001",
  25091=>"001001001",
  25092=>"111001010",
  25093=>"011011111",
  25094=>"110100101",
  25095=>"010101111",
  25096=>"010010000",
  25097=>"101101111",
  25098=>"010001000",
  25099=>"111000100",
  25100=>"011001111",
  25101=>"001111010",
  25102=>"010000000",
  25103=>"101000011",
  25104=>"111100001",
  25105=>"001000101",
  25106=>"011111000",
  25107=>"100111011",
  25108=>"101110110",
  25109=>"101011010",
  25110=>"000000000",
  25111=>"100110011",
  25112=>"110111110",
  25113=>"000100111",
  25114=>"010100110",
  25115=>"011100001",
  25116=>"101111101",
  25117=>"001100100",
  25118=>"000000011",
  25119=>"111000101",
  25120=>"011010101",
  25121=>"001101010",
  25122=>"011001010",
  25123=>"010101101",
  25124=>"100001011",
  25125=>"000010101",
  25126=>"100100100",
  25127=>"110010110",
  25128=>"100101100",
  25129=>"001111101",
  25130=>"001011000",
  25131=>"110011101",
  25132=>"001101011",
  25133=>"110110100",
  25134=>"010110010",
  25135=>"110011001",
  25136=>"001110100",
  25137=>"011000101",
  25138=>"001010011",
  25139=>"011110110",
  25140=>"010110001",
  25141=>"000001101",
  25142=>"010110110",
  25143=>"100111001",
  25144=>"110110000",
  25145=>"001101010",
  25146=>"110111011",
  25147=>"101010100",
  25148=>"110010001",
  25149=>"110000000",
  25150=>"101011001",
  25151=>"110111011",
  25152=>"100011000",
  25153=>"110100110",
  25154=>"111001100",
  25155=>"100000110",
  25156=>"110100101",
  25157=>"000111000",
  25158=>"010110001",
  25159=>"010100001",
  25160=>"100100001",
  25161=>"001011000",
  25162=>"000000111",
  25163=>"000110101",
  25164=>"001000111",
  25165=>"100001101",
  25166=>"011000011",
  25167=>"011101101",
  25168=>"001110010",
  25169=>"010110110",
  25170=>"110000000",
  25171=>"101101101",
  25172=>"100001101",
  25173=>"011011101",
  25174=>"000100010",
  25175=>"100011101",
  25176=>"000010101",
  25177=>"000000001",
  25178=>"111101011",
  25179=>"101110100",
  25180=>"100111100",
  25181=>"011100001",
  25182=>"001110100",
  25183=>"000001110",
  25184=>"010100100",
  25185=>"011111111",
  25186=>"110110000",
  25187=>"100010110",
  25188=>"111000110",
  25189=>"101001011",
  25190=>"101011000",
  25191=>"110010110",
  25192=>"010001011",
  25193=>"011111010",
  25194=>"001111100",
  25195=>"000001010",
  25196=>"111101011",
  25197=>"100011001",
  25198=>"101100000",
  25199=>"010111101",
  25200=>"111000110",
  25201=>"010000000",
  25202=>"100000011",
  25203=>"100111111",
  25204=>"001000001",
  25205=>"101100101",
  25206=>"101100100",
  25207=>"001000100",
  25208=>"001110110",
  25209=>"010101110",
  25210=>"111101111",
  25211=>"100001001",
  25212=>"010011111",
  25213=>"101101001",
  25214=>"010011100",
  25215=>"000100010",
  25216=>"011000000",
  25217=>"100010110",
  25218=>"010001100",
  25219=>"100110110",
  25220=>"010100011",
  25221=>"101111011",
  25222=>"101100110",
  25223=>"100111101",
  25224=>"010001000",
  25225=>"100010110",
  25226=>"110001011",
  25227=>"010001110",
  25228=>"011101111",
  25229=>"100001010",
  25230=>"010011000",
  25231=>"011101011",
  25232=>"101101111",
  25233=>"100100101",
  25234=>"110010110",
  25235=>"010111001",
  25236=>"100010101",
  25237=>"010111011",
  25238=>"011011000",
  25239=>"111101001",
  25240=>"111000101",
  25241=>"100001111",
  25242=>"010111000",
  25243=>"010000110",
  25244=>"100110101",
  25245=>"100000000",
  25246=>"001001111",
  25247=>"101100011",
  25248=>"111010000",
  25249=>"111011101",
  25250=>"011010010",
  25251=>"010111100",
  25252=>"111010100",
  25253=>"111011000",
  25254=>"001001000",
  25255=>"011110001",
  25256=>"001101001",
  25257=>"101101110",
  25258=>"000101011",
  25259=>"010000000",
  25260=>"101111011",
  25261=>"000010010",
  25262=>"000110101",
  25263=>"001001111",
  25264=>"101001001",
  25265=>"010111010",
  25266=>"010111001",
  25267=>"101001101",
  25268=>"110101010",
  25269=>"111111010",
  25270=>"111101110",
  25271=>"011010001",
  25272=>"000011011",
  25273=>"111010001",
  25274=>"110001000",
  25275=>"100000110",
  25276=>"110101111",
  25277=>"110011010",
  25278=>"101101011",
  25279=>"110101010",
  25280=>"111001110",
  25281=>"110000100",
  25282=>"101010010",
  25283=>"010010000",
  25284=>"100011000",
  25285=>"000110010",
  25286=>"000111101",
  25287=>"101100100",
  25288=>"001001101",
  25289=>"011100111",
  25290=>"110110010",
  25291=>"001111000",
  25292=>"010100000",
  25293=>"100110100",
  25294=>"010111010",
  25295=>"010010110",
  25296=>"000000110",
  25297=>"011110110",
  25298=>"001101101",
  25299=>"101011100",
  25300=>"001111100",
  25301=>"000110000",
  25302=>"101100011",
  25303=>"010010011",
  25304=>"100110110",
  25305=>"101000111",
  25306=>"010101101",
  25307=>"110110101",
  25308=>"101111111",
  25309=>"100000000",
  25310=>"001001000",
  25311=>"000100001",
  25312=>"110001111",
  25313=>"100001011",
  25314=>"110100111",
  25315=>"001010001",
  25316=>"010110011",
  25317=>"111000101",
  25318=>"110000100",
  25319=>"011100101",
  25320=>"100110000",
  25321=>"101000001",
  25322=>"101001111",
  25323=>"111011101",
  25324=>"101000101",
  25325=>"000110101",
  25326=>"111000111",
  25327=>"010001110",
  25328=>"011011111",
  25329=>"111110001",
  25330=>"001000001",
  25331=>"010100001",
  25332=>"111101010",
  25333=>"100011111",
  25334=>"011101010",
  25335=>"010011000",
  25336=>"110000101",
  25337=>"001000001",
  25338=>"000010100",
  25339=>"001100100",
  25340=>"000101111",
  25341=>"011100001",
  25342=>"010001111",
  25343=>"110000101",
  25344=>"000110110",
  25345=>"111100011",
  25346=>"111101101",
  25347=>"010111011",
  25348=>"011110001",
  25349=>"110101100",
  25350=>"000000110",
  25351=>"100011000",
  25352=>"110001101",
  25353=>"000110010",
  25354=>"011111100",
  25355=>"101010001",
  25356=>"110110101",
  25357=>"011100010",
  25358=>"100000101",
  25359=>"000001000",
  25360=>"001000100",
  25361=>"100101100",
  25362=>"000111111",
  25363=>"110001000",
  25364=>"100010101",
  25365=>"000000101",
  25366=>"100100100",
  25367=>"110111100",
  25368=>"011000010",
  25369=>"011001100",
  25370=>"100110010",
  25371=>"110000001",
  25372=>"001111110",
  25373=>"000010011",
  25374=>"011000110",
  25375=>"010101100",
  25376=>"111001011",
  25377=>"010000111",
  25378=>"001011101",
  25379=>"011011111",
  25380=>"101111111",
  25381=>"010011101",
  25382=>"010000000",
  25383=>"100110101",
  25384=>"101011010",
  25385=>"001011001",
  25386=>"110100000",
  25387=>"010001010",
  25388=>"000011101",
  25389=>"011010111",
  25390=>"101111100",
  25391=>"000010110",
  25392=>"111101000",
  25393=>"110000000",
  25394=>"001000000",
  25395=>"100101001",
  25396=>"011011111",
  25397=>"000101100",
  25398=>"111101000",
  25399=>"111111111",
  25400=>"110000100",
  25401=>"000001010",
  25402=>"010111110",
  25403=>"111111001",
  25404=>"110001011",
  25405=>"101001000",
  25406=>"000101101",
  25407=>"001111000",
  25408=>"101001000",
  25409=>"110101100",
  25410=>"100101001",
  25411=>"111001011",
  25412=>"000101111",
  25413=>"110110111",
  25414=>"010101111",
  25415=>"101111111",
  25416=>"110000100",
  25417=>"010110110",
  25418=>"000100101",
  25419=>"001010101",
  25420=>"001000100",
  25421=>"001100000",
  25422=>"000000010",
  25423=>"111110000",
  25424=>"011100001",
  25425=>"100100011",
  25426=>"100000001",
  25427=>"001111101",
  25428=>"011001101",
  25429=>"101110110",
  25430=>"000101111",
  25431=>"010001001",
  25432=>"110011000",
  25433=>"001101000",
  25434=>"010101110",
  25435=>"001101101",
  25436=>"001000100",
  25437=>"111110011",
  25438=>"110000011",
  25439=>"101010011",
  25440=>"010101001",
  25441=>"111101110",
  25442=>"111101010",
  25443=>"011001001",
  25444=>"000001101",
  25445=>"000100011",
  25446=>"010100000",
  25447=>"110100100",
  25448=>"100011001",
  25449=>"011110101",
  25450=>"101001001",
  25451=>"000010101",
  25452=>"000001101",
  25453=>"001010011",
  25454=>"101101110",
  25455=>"001000011",
  25456=>"000110001",
  25457=>"101000010",
  25458=>"110000001",
  25459=>"001010001",
  25460=>"011000111",
  25461=>"010100011",
  25462=>"111000001",
  25463=>"111011100",
  25464=>"001000101",
  25465=>"000110001",
  25466=>"110001111",
  25467=>"001011100",
  25468=>"010111010",
  25469=>"111000111",
  25470=>"111111101",
  25471=>"001101101",
  25472=>"110100011",
  25473=>"011000100",
  25474=>"100101111",
  25475=>"010001010",
  25476=>"000001110",
  25477=>"111000010",
  25478=>"101110010",
  25479=>"101010111",
  25480=>"111110010",
  25481=>"010011011",
  25482=>"111011000",
  25483=>"000011111",
  25484=>"110000110",
  25485=>"111111000",
  25486=>"100001011",
  25487=>"110100100",
  25488=>"010000111",
  25489=>"001110101",
  25490=>"101011010",
  25491=>"100010011",
  25492=>"011001011",
  25493=>"011001101",
  25494=>"010001100",
  25495=>"100110000",
  25496=>"010111001",
  25497=>"000011001",
  25498=>"111110001",
  25499=>"000000110",
  25500=>"000110011",
  25501=>"101101101",
  25502=>"100100001",
  25503=>"000011110",
  25504=>"011100111",
  25505=>"111000101",
  25506=>"001110111",
  25507=>"001000001",
  25508=>"001110101",
  25509=>"111100001",
  25510=>"100111010",
  25511=>"100001000",
  25512=>"101011011",
  25513=>"011100011",
  25514=>"001011100",
  25515=>"011101010",
  25516=>"110101010",
  25517=>"101110001",
  25518=>"000100011",
  25519=>"101001011",
  25520=>"011000010",
  25521=>"001001110",
  25522=>"101000000",
  25523=>"101100000",
  25524=>"000110111",
  25525=>"000001010",
  25526=>"011011000",
  25527=>"010001010",
  25528=>"100111101",
  25529=>"101010100",
  25530=>"111001001",
  25531=>"111010101",
  25532=>"000010100",
  25533=>"101110111",
  25534=>"000001101",
  25535=>"000000010",
  25536=>"110110110",
  25537=>"100111111",
  25538=>"110010010",
  25539=>"101010100",
  25540=>"000111000",
  25541=>"100000110",
  25542=>"000010001",
  25543=>"000000000",
  25544=>"000100000",
  25545=>"000110111",
  25546=>"010001111",
  25547=>"011010000",
  25548=>"101010011",
  25549=>"000010010",
  25550=>"111111001",
  25551=>"001100000",
  25552=>"100101011",
  25553=>"100100101",
  25554=>"111000001",
  25555=>"110010001",
  25556=>"011101001",
  25557=>"010010111",
  25558=>"011111001",
  25559=>"110011101",
  25560=>"111101000",
  25561=>"001001010",
  25562=>"001110011",
  25563=>"010000000",
  25564=>"110100101",
  25565=>"001001100",
  25566=>"100100001",
  25567=>"000111011",
  25568=>"101000001",
  25569=>"101010111",
  25570=>"011001010",
  25571=>"111101111",
  25572=>"100010000",
  25573=>"011101001",
  25574=>"000110101",
  25575=>"101011101",
  25576=>"110011110",
  25577=>"100111111",
  25578=>"111101011",
  25579=>"000001101",
  25580=>"101111011",
  25581=>"011001000",
  25582=>"101111100",
  25583=>"110000100",
  25584=>"101101110",
  25585=>"000011100",
  25586=>"100110000",
  25587=>"111111101",
  25588=>"010001101",
  25589=>"001001000",
  25590=>"000111011",
  25591=>"101101100",
  25592=>"000101000",
  25593=>"010110001",
  25594=>"110010011",
  25595=>"111001111",
  25596=>"100111111",
  25597=>"010001011",
  25598=>"011010010",
  25599=>"110100011",
  25600=>"111011111",
  25601=>"100011111",
  25602=>"000111110",
  25603=>"011010000",
  25604=>"010100110",
  25605=>"000010110",
  25606=>"011011010",
  25607=>"100010010",
  25608=>"111110100",
  25609=>"111100110",
  25610=>"000110001",
  25611=>"001110110",
  25612=>"100000001",
  25613=>"100111101",
  25614=>"011101111",
  25615=>"100101101",
  25616=>"110010101",
  25617=>"000000101",
  25618=>"110110111",
  25619=>"101111100",
  25620=>"001011111",
  25621=>"101101111",
  25622=>"010100110",
  25623=>"001011110",
  25624=>"100011110",
  25625=>"101010011",
  25626=>"100001110",
  25627=>"100000000",
  25628=>"001010100",
  25629=>"011011110",
  25630=>"001110110",
  25631=>"000000000",
  25632=>"001110011",
  25633=>"101011011",
  25634=>"001001010",
  25635=>"010000110",
  25636=>"010100011",
  25637=>"010101110",
  25638=>"111101001",
  25639=>"101000001",
  25640=>"111010111",
  25641=>"010000001",
  25642=>"000010111",
  25643=>"100111011",
  25644=>"110110000",
  25645=>"011110111",
  25646=>"001101110",
  25647=>"000001111",
  25648=>"110001011",
  25649=>"010011111",
  25650=>"001000000",
  25651=>"000100100",
  25652=>"110001001",
  25653=>"100100000",
  25654=>"111011010",
  25655=>"001110110",
  25656=>"101101010",
  25657=>"100101101",
  25658=>"100111001",
  25659=>"000010101",
  25660=>"111101001",
  25661=>"111100101",
  25662=>"110010011",
  25663=>"011100000",
  25664=>"000100111",
  25665=>"101000101",
  25666=>"111101010",
  25667=>"000100001",
  25668=>"100001110",
  25669=>"100100101",
  25670=>"000001111",
  25671=>"100000010",
  25672=>"000001110",
  25673=>"101101110",
  25674=>"010000000",
  25675=>"000100111",
  25676=>"000000111",
  25677=>"100101100",
  25678=>"011111110",
  25679=>"001011100",
  25680=>"101101110",
  25681=>"111100010",
  25682=>"011010100",
  25683=>"111111111",
  25684=>"001101011",
  25685=>"000111011",
  25686=>"101101111",
  25687=>"000110101",
  25688=>"001111010",
  25689=>"101111011",
  25690=>"001001010",
  25691=>"101001110",
  25692=>"011111100",
  25693=>"011110010",
  25694=>"001111110",
  25695=>"111001000",
  25696=>"110000100",
  25697=>"000110110",
  25698=>"100111110",
  25699=>"010000100",
  25700=>"100111001",
  25701=>"010101101",
  25702=>"001010110",
  25703=>"111001000",
  25704=>"011110001",
  25705=>"011100011",
  25706=>"001100000",
  25707=>"011100000",
  25708=>"111100101",
  25709=>"110101101",
  25710=>"100010100",
  25711=>"011011000",
  25712=>"111001111",
  25713=>"001010001",
  25714=>"100001000",
  25715=>"110010101",
  25716=>"000110100",
  25717=>"110100011",
  25718=>"000101001",
  25719=>"110011110",
  25720=>"100000101",
  25721=>"010110101",
  25722=>"111101011",
  25723=>"100111010",
  25724=>"011010011",
  25725=>"010111101",
  25726=>"100001101",
  25727=>"010011111",
  25728=>"110111111",
  25729=>"011110010",
  25730=>"010111011",
  25731=>"111010111",
  25732=>"001010011",
  25733=>"011100001",
  25734=>"101101010",
  25735=>"000111101",
  25736=>"010100101",
  25737=>"000001011",
  25738=>"101100101",
  25739=>"000000100",
  25740=>"001001000",
  25741=>"101110111",
  25742=>"110000111",
  25743=>"101011110",
  25744=>"100101101",
  25745=>"100000100",
  25746=>"101110011",
  25747=>"011001100",
  25748=>"010111001",
  25749=>"010111100",
  25750=>"100101100",
  25751=>"000000110",
  25752=>"001100011",
  25753=>"100101011",
  25754=>"000010101",
  25755=>"010111011",
  25756=>"010011110",
  25757=>"111010110",
  25758=>"010101011",
  25759=>"110100011",
  25760=>"000011010",
  25761=>"111110010",
  25762=>"010110100",
  25763=>"110110101",
  25764=>"011010100",
  25765=>"110011000",
  25766=>"101001011",
  25767=>"011101100",
  25768=>"011000000",
  25769=>"011111110",
  25770=>"010101101",
  25771=>"110111000",
  25772=>"111101000",
  25773=>"011101001",
  25774=>"101111110",
  25775=>"101110010",
  25776=>"100100101",
  25777=>"000000010",
  25778=>"111111011",
  25779=>"000110011",
  25780=>"100110100",
  25781=>"100010101",
  25782=>"010001100",
  25783=>"100100100",
  25784=>"010110011",
  25785=>"010101001",
  25786=>"111010011",
  25787=>"111101011",
  25788=>"011000010",
  25789=>"001001011",
  25790=>"010000010",
  25791=>"110101100",
  25792=>"011001100",
  25793=>"101010111",
  25794=>"110010000",
  25795=>"001001011",
  25796=>"011010101",
  25797=>"110110111",
  25798=>"110000100",
  25799=>"011110110",
  25800=>"111000101",
  25801=>"110110110",
  25802=>"101000000",
  25803=>"110100101",
  25804=>"110010101",
  25805=>"110011000",
  25806=>"010101100",
  25807=>"000000000",
  25808=>"010010101",
  25809=>"000011010",
  25810=>"111111000",
  25811=>"110100110",
  25812=>"000000000",
  25813=>"010011111",
  25814=>"111111001",
  25815=>"000001001",
  25816=>"111000100",
  25817=>"000011000",
  25818=>"110111000",
  25819=>"111011001",
  25820=>"110110111",
  25821=>"110011111",
  25822=>"111101000",
  25823=>"010100111",
  25824=>"011001111",
  25825=>"100011011",
  25826=>"111010100",
  25827=>"000101110",
  25828=>"100010000",
  25829=>"000000100",
  25830=>"111100101",
  25831=>"100011001",
  25832=>"010011001",
  25833=>"110011101",
  25834=>"100101110",
  25835=>"111100000",
  25836=>"100110111",
  25837=>"010000010",
  25838=>"011101000",
  25839=>"101001101",
  25840=>"101100101",
  25841=>"101100011",
  25842=>"101000010",
  25843=>"000100010",
  25844=>"101100000",
  25845=>"110010011",
  25846=>"000001111",
  25847=>"000101011",
  25848=>"110110011",
  25849=>"111101101",
  25850=>"011010000",
  25851=>"111011000",
  25852=>"100100011",
  25853=>"101111111",
  25854=>"101111100",
  25855=>"111100111",
  25856=>"001100100",
  25857=>"010110000",
  25858=>"010100001",
  25859=>"100100101",
  25860=>"010110101",
  25861=>"100100000",
  25862=>"001110111",
  25863=>"111000010",
  25864=>"101001000",
  25865=>"101111011",
  25866=>"011101011",
  25867=>"101010001",
  25868=>"001011110",
  25869=>"110100001",
  25870=>"010001110",
  25871=>"011111001",
  25872=>"111011001",
  25873=>"011110011",
  25874=>"111110001",
  25875=>"111111011",
  25876=>"111100100",
  25877=>"001100001",
  25878=>"000000001",
  25879=>"000100100",
  25880=>"010011011",
  25881=>"100011001",
  25882=>"100110001",
  25883=>"101001111",
  25884=>"110101100",
  25885=>"010011111",
  25886=>"100110100",
  25887=>"000111001",
  25888=>"100011111",
  25889=>"000000010",
  25890=>"101001000",
  25891=>"101101100",
  25892=>"110000000",
  25893=>"111100000",
  25894=>"000101010",
  25895=>"010101000",
  25896=>"101000001",
  25897=>"011110000",
  25898=>"011010000",
  25899=>"000001000",
  25900=>"010010101",
  25901=>"010111000",
  25902=>"010100010",
  25903=>"011001100",
  25904=>"101100111",
  25905=>"110100010",
  25906=>"001101100",
  25907=>"110100101",
  25908=>"111001101",
  25909=>"111001000",
  25910=>"100110011",
  25911=>"000000111",
  25912=>"000011010",
  25913=>"010001100",
  25914=>"111111000",
  25915=>"011100101",
  25916=>"010111000",
  25917=>"110000100",
  25918=>"100100100",
  25919=>"101011110",
  25920=>"000000101",
  25921=>"001000111",
  25922=>"101101010",
  25923=>"000110000",
  25924=>"001101101",
  25925=>"111110011",
  25926=>"001101001",
  25927=>"101000000",
  25928=>"010011100",
  25929=>"001011110",
  25930=>"100110001",
  25931=>"101111100",
  25932=>"100111011",
  25933=>"100101001",
  25934=>"011000110",
  25935=>"111100001",
  25936=>"000101001",
  25937=>"100000010",
  25938=>"011101111",
  25939=>"100101110",
  25940=>"110111010",
  25941=>"011000010",
  25942=>"101010000",
  25943=>"001001010",
  25944=>"110000100",
  25945=>"110101100",
  25946=>"111101101",
  25947=>"010110011",
  25948=>"001100101",
  25949=>"010110110",
  25950=>"010100000",
  25951=>"101010100",
  25952=>"001001010",
  25953=>"000010010",
  25954=>"010100101",
  25955=>"100110111",
  25956=>"110101000",
  25957=>"001010101",
  25958=>"010010000",
  25959=>"001011110",
  25960=>"010000110",
  25961=>"001111111",
  25962=>"001001001",
  25963=>"100100010",
  25964=>"011010111",
  25965=>"110101011",
  25966=>"111001100",
  25967=>"101110100",
  25968=>"000001000",
  25969=>"001000111",
  25970=>"100001111",
  25971=>"011000001",
  25972=>"011100100",
  25973=>"000111011",
  25974=>"110010000",
  25975=>"001110110",
  25976=>"110000100",
  25977=>"100111101",
  25978=>"000110001",
  25979=>"101110000",
  25980=>"110111001",
  25981=>"001000001",
  25982=>"100110010",
  25983=>"100010111",
  25984=>"101001001",
  25985=>"010101110",
  25986=>"000011101",
  25987=>"100011111",
  25988=>"011101111",
  25989=>"111101111",
  25990=>"101001110",
  25991=>"000010100",
  25992=>"000000100",
  25993=>"101000100",
  25994=>"100001100",
  25995=>"101010110",
  25996=>"110001111",
  25997=>"010100110",
  25998=>"101100111",
  25999=>"101111010",
  26000=>"110111111",
  26001=>"100000001",
  26002=>"011101111",
  26003=>"001100110",
  26004=>"111010010",
  26005=>"100000101",
  26006=>"110000101",
  26007=>"000011011",
  26008=>"010111001",
  26009=>"011111110",
  26010=>"100000010",
  26011=>"011111011",
  26012=>"110000000",
  26013=>"000010100",
  26014=>"110011111",
  26015=>"110000000",
  26016=>"000111101",
  26017=>"010111110",
  26018=>"101000100",
  26019=>"000011000",
  26020=>"001000111",
  26021=>"010010100",
  26022=>"000100110",
  26023=>"001101001",
  26024=>"001001100",
  26025=>"000010001",
  26026=>"111111111",
  26027=>"010110100",
  26028=>"010110001",
  26029=>"011111001",
  26030=>"100111111",
  26031=>"101111100",
  26032=>"001110100",
  26033=>"010111100",
  26034=>"010010101",
  26035=>"101000101",
  26036=>"011010101",
  26037=>"100110111",
  26038=>"100110010",
  26039=>"111010101",
  26040=>"010000011",
  26041=>"110110100",
  26042=>"111100100",
  26043=>"000000111",
  26044=>"110100111",
  26045=>"000111011",
  26046=>"000010100",
  26047=>"011110011",
  26048=>"001011001",
  26049=>"111110000",
  26050=>"110100011",
  26051=>"010001000",
  26052=>"101110111",
  26053=>"110101000",
  26054=>"001011101",
  26055=>"100111100",
  26056=>"111011110",
  26057=>"010101100",
  26058=>"000010011",
  26059=>"111111100",
  26060=>"111101110",
  26061=>"001110001",
  26062=>"101101010",
  26063=>"110011001",
  26064=>"001001000",
  26065=>"000001111",
  26066=>"111100100",
  26067=>"111011100",
  26068=>"100101111",
  26069=>"001001010",
  26070=>"100100000",
  26071=>"110000011",
  26072=>"011011101",
  26073=>"111100000",
  26074=>"111110111",
  26075=>"011110001",
  26076=>"010010111",
  26077=>"100011001",
  26078=>"101000101",
  26079=>"011011101",
  26080=>"101011111",
  26081=>"111000111",
  26082=>"010111111",
  26083=>"101101001",
  26084=>"101010001",
  26085=>"000001001",
  26086=>"101100110",
  26087=>"111011001",
  26088=>"110001101",
  26089=>"110010100",
  26090=>"010000110",
  26091=>"110111101",
  26092=>"010001010",
  26093=>"111010110",
  26094=>"111011000",
  26095=>"000010001",
  26096=>"001110101",
  26097=>"111010010",
  26098=>"100111001",
  26099=>"111000110",
  26100=>"110100011",
  26101=>"011000000",
  26102=>"001111101",
  26103=>"100100010",
  26104=>"000011001",
  26105=>"101000100",
  26106=>"011001101",
  26107=>"101010001",
  26108=>"111100100",
  26109=>"000000101",
  26110=>"101110010",
  26111=>"000110111",
  26112=>"101011110",
  26113=>"101111011",
  26114=>"000100000",
  26115=>"000100000",
  26116=>"001110001",
  26117=>"111001111",
  26118=>"110001011",
  26119=>"101111111",
  26120=>"110011101",
  26121=>"011011011",
  26122=>"101001000",
  26123=>"010110010",
  26124=>"110001011",
  26125=>"100101001",
  26126=>"010111111",
  26127=>"011011001",
  26128=>"000100010",
  26129=>"110110110",
  26130=>"100011001",
  26131=>"111010000",
  26132=>"011001001",
  26133=>"100111101",
  26134=>"101110000",
  26135=>"101110101",
  26136=>"100000110",
  26137=>"110011111",
  26138=>"001010111",
  26139=>"010001010",
  26140=>"110100011",
  26141=>"000011011",
  26142=>"000010011",
  26143=>"101010111",
  26144=>"010001001",
  26145=>"000011010",
  26146=>"111010101",
  26147=>"000110010",
  26148=>"000111010",
  26149=>"001111100",
  26150=>"001001001",
  26151=>"100101001",
  26152=>"100100100",
  26153=>"000001001",
  26154=>"010110011",
  26155=>"111010010",
  26156=>"000111101",
  26157=>"000000001",
  26158=>"100010010",
  26159=>"001100010",
  26160=>"010000111",
  26161=>"111101011",
  26162=>"110110101",
  26163=>"101101010",
  26164=>"000000101",
  26165=>"111001100",
  26166=>"011010010",
  26167=>"111000010",
  26168=>"000100110",
  26169=>"111101100",
  26170=>"100000100",
  26171=>"010111010",
  26172=>"011101001",
  26173=>"011110101",
  26174=>"000101111",
  26175=>"111110011",
  26176=>"000100111",
  26177=>"011011010",
  26178=>"101111011",
  26179=>"000010111",
  26180=>"101111101",
  26181=>"110111000",
  26182=>"111101111",
  26183=>"001011001",
  26184=>"110010001",
  26185=>"110011101",
  26186=>"110000100",
  26187=>"000100101",
  26188=>"110111110",
  26189=>"010000010",
  26190=>"111000110",
  26191=>"100100101",
  26192=>"000100011",
  26193=>"010111011",
  26194=>"101101011",
  26195=>"011001110",
  26196=>"101000000",
  26197=>"000010000",
  26198=>"000110010",
  26199=>"010000111",
  26200=>"010100100",
  26201=>"000110011",
  26202=>"001100010",
  26203=>"101110100",
  26204=>"011010100",
  26205=>"111100001",
  26206=>"000111010",
  26207=>"100011111",
  26208=>"000101111",
  26209=>"011000010",
  26210=>"101111100",
  26211=>"100000010",
  26212=>"000010110",
  26213=>"011000101",
  26214=>"001111100",
  26215=>"011101100",
  26216=>"101001000",
  26217=>"001111100",
  26218=>"101110010",
  26219=>"011001011",
  26220=>"010101001",
  26221=>"110011110",
  26222=>"001100011",
  26223=>"110100010",
  26224=>"111010101",
  26225=>"000101100",
  26226=>"111111001",
  26227=>"000000110",
  26228=>"100111000",
  26229=>"001000101",
  26230=>"001100101",
  26231=>"010010110",
  26232=>"011110011",
  26233=>"000111111",
  26234=>"010111101",
  26235=>"010001011",
  26236=>"011110000",
  26237=>"001011000",
  26238=>"011110100",
  26239=>"110011111",
  26240=>"110011100",
  26241=>"000001111",
  26242=>"110001000",
  26243=>"010110000",
  26244=>"100110101",
  26245=>"101010101",
  26246=>"000001000",
  26247=>"001000101",
  26248=>"100000100",
  26249=>"010101000",
  26250=>"110001111",
  26251=>"101100011",
  26252=>"011110101",
  26253=>"100100100",
  26254=>"010010111",
  26255=>"111110001",
  26256=>"111100010",
  26257=>"011100100",
  26258=>"011011101",
  26259=>"011111110",
  26260=>"010011011",
  26261=>"010110100",
  26262=>"001100100",
  26263=>"111010000",
  26264=>"001010000",
  26265=>"101111010",
  26266=>"010101001",
  26267=>"010111110",
  26268=>"000110001",
  26269=>"010011000",
  26270=>"010100011",
  26271=>"111010011",
  26272=>"010001100",
  26273=>"001010111",
  26274=>"111110100",
  26275=>"111001001",
  26276=>"011101110",
  26277=>"101000001",
  26278=>"010001011",
  26279=>"100000010",
  26280=>"100001011",
  26281=>"100001010",
  26282=>"011110001",
  26283=>"010011010",
  26284=>"110100010",
  26285=>"110011011",
  26286=>"010001111",
  26287=>"011010010",
  26288=>"111110110",
  26289=>"111101100",
  26290=>"111100001",
  26291=>"010101000",
  26292=>"100101010",
  26293=>"010001111",
  26294=>"000100011",
  26295=>"001110100",
  26296=>"111111111",
  26297=>"101101000",
  26298=>"011000011",
  26299=>"001010101",
  26300=>"001111111",
  26301=>"011000011",
  26302=>"010101111",
  26303=>"000000100",
  26304=>"110011100",
  26305=>"001111001",
  26306=>"000111110",
  26307=>"000100100",
  26308=>"100100101",
  26309=>"000111000",
  26310=>"111010110",
  26311=>"101101100",
  26312=>"011000110",
  26313=>"101101101",
  26314=>"011100000",
  26315=>"101110110",
  26316=>"110111111",
  26317=>"001110101",
  26318=>"111010111",
  26319=>"100010010",
  26320=>"101101111",
  26321=>"110111111",
  26322=>"110010110",
  26323=>"111110110",
  26324=>"100001001",
  26325=>"010111110",
  26326=>"001000010",
  26327=>"010000111",
  26328=>"100011100",
  26329=>"100111110",
  26330=>"111011000",
  26331=>"111100101",
  26332=>"010000001",
  26333=>"010011011",
  26334=>"101010001",
  26335=>"000010011",
  26336=>"101101001",
  26337=>"001101000",
  26338=>"000110001",
  26339=>"000101101",
  26340=>"000001100",
  26341=>"111010111",
  26342=>"111000111",
  26343=>"001111010",
  26344=>"110110000",
  26345=>"010001011",
  26346=>"111011111",
  26347=>"111000100",
  26348=>"000000001",
  26349=>"101110100",
  26350=>"000001100",
  26351=>"111110101",
  26352=>"011100000",
  26353=>"111111111",
  26354=>"101010101",
  26355=>"100101100",
  26356=>"101101000",
  26357=>"111010011",
  26358=>"101001000",
  26359=>"110001000",
  26360=>"000000011",
  26361=>"011000001",
  26362=>"001001111",
  26363=>"011010000",
  26364=>"101101010",
  26365=>"110110011",
  26366=>"101011011",
  26367=>"111100111",
  26368=>"100101010",
  26369=>"100100100",
  26370=>"100001001",
  26371=>"001110110",
  26372=>"100100010",
  26373=>"110100111",
  26374=>"010010100",
  26375=>"000111100",
  26376=>"001100111",
  26377=>"100111111",
  26378=>"110110001",
  26379=>"010101011",
  26380=>"110011101",
  26381=>"000001001",
  26382=>"011001011",
  26383=>"101001100",
  26384=>"110001100",
  26385=>"100011010",
  26386=>"101110100",
  26387=>"011011110",
  26388=>"010001101",
  26389=>"111001000",
  26390=>"011100001",
  26391=>"001010101",
  26392=>"000000101",
  26393=>"001101001",
  26394=>"100110111",
  26395=>"001010000",
  26396=>"010100101",
  26397=>"110001011",
  26398=>"100001001",
  26399=>"110111110",
  26400=>"011000010",
  26401=>"100010111",
  26402=>"100111111",
  26403=>"011010011",
  26404=>"100001011",
  26405=>"100100110",
  26406=>"101101101",
  26407=>"010110111",
  26408=>"010111111",
  26409=>"000110100",
  26410=>"000100001",
  26411=>"111010010",
  26412=>"111011011",
  26413=>"011010101",
  26414=>"101110010",
  26415=>"101110000",
  26416=>"001010101",
  26417=>"011111111",
  26418=>"111100100",
  26419=>"010001000",
  26420=>"011100110",
  26421=>"000110100",
  26422=>"000010100",
  26423=>"000010010",
  26424=>"100000101",
  26425=>"101000110",
  26426=>"100011111",
  26427=>"100001000",
  26428=>"000010011",
  26429=>"000101100",
  26430=>"010011111",
  26431=>"001010100",
  26432=>"001010101",
  26433=>"100010001",
  26434=>"111100001",
  26435=>"101110111",
  26436=>"010100000",
  26437=>"010101101",
  26438=>"110111100",
  26439=>"100101000",
  26440=>"100101100",
  26441=>"101101010",
  26442=>"011111100",
  26443=>"100100011",
  26444=>"010110100",
  26445=>"000111100",
  26446=>"010011111",
  26447=>"001011001",
  26448=>"110011000",
  26449=>"010010000",
  26450=>"000000111",
  26451=>"011011110",
  26452=>"101000110",
  26453=>"111001001",
  26454=>"000000010",
  26455=>"101010101",
  26456=>"010111010",
  26457=>"110101000",
  26458=>"001001001",
  26459=>"111111010",
  26460=>"001011111",
  26461=>"011111011",
  26462=>"010101111",
  26463=>"000111101",
  26464=>"111101110",
  26465=>"011010111",
  26466=>"000100100",
  26467=>"010101101",
  26468=>"110010100",
  26469=>"011000101",
  26470=>"111111011",
  26471=>"111110000",
  26472=>"001000011",
  26473=>"011110111",
  26474=>"110100100",
  26475=>"000111000",
  26476=>"101001001",
  26477=>"000011110",
  26478=>"100001110",
  26479=>"001111100",
  26480=>"101001101",
  26481=>"000101001",
  26482=>"011101010",
  26483=>"110011001",
  26484=>"100101011",
  26485=>"101001100",
  26486=>"111101010",
  26487=>"111110110",
  26488=>"110100100",
  26489=>"011010000",
  26490=>"011011101",
  26491=>"110010001",
  26492=>"010100010",
  26493=>"101101100",
  26494=>"101001111",
  26495=>"001011100",
  26496=>"101110010",
  26497=>"010001001",
  26498=>"011110010",
  26499=>"101111111",
  26500=>"101100011",
  26501=>"110001110",
  26502=>"001010000",
  26503=>"000010010",
  26504=>"011011001",
  26505=>"010111110",
  26506=>"111001011",
  26507=>"010100100",
  26508=>"010110000",
  26509=>"110010110",
  26510=>"100000100",
  26511=>"011010111",
  26512=>"100001101",
  26513=>"000110000",
  26514=>"000100010",
  26515=>"001000111",
  26516=>"001100000",
  26517=>"000100111",
  26518=>"111001000",
  26519=>"001111100",
  26520=>"100111000",
  26521=>"101101000",
  26522=>"101011100",
  26523=>"100010110",
  26524=>"010000011",
  26525=>"011011010",
  26526=>"011011111",
  26527=>"000011100",
  26528=>"100010110",
  26529=>"100001101",
  26530=>"100001000",
  26531=>"111010011",
  26532=>"010000010",
  26533=>"010100000",
  26534=>"100000101",
  26535=>"111110001",
  26536=>"111100100",
  26537=>"100001101",
  26538=>"001110000",
  26539=>"111100101",
  26540=>"111011101",
  26541=>"010110110",
  26542=>"001000001",
  26543=>"101101010",
  26544=>"011010110",
  26545=>"110001111",
  26546=>"111110001",
  26547=>"101000000",
  26548=>"100110000",
  26549=>"111010100",
  26550=>"010011001",
  26551=>"100010010",
  26552=>"010000111",
  26553=>"010100101",
  26554=>"010000100",
  26555=>"110100001",
  26556=>"001111001",
  26557=>"011101111",
  26558=>"000010010",
  26559=>"110010111",
  26560=>"110001010",
  26561=>"111101000",
  26562=>"000111011",
  26563=>"000100011",
  26564=>"110010100",
  26565=>"100000111",
  26566=>"101001101",
  26567=>"100001101",
  26568=>"100111111",
  26569=>"111111010",
  26570=>"110110110",
  26571=>"111111100",
  26572=>"010010000",
  26573=>"100101010",
  26574=>"110111000",
  26575=>"110000011",
  26576=>"110101100",
  26577=>"100111100",
  26578=>"110110010",
  26579=>"011110011",
  26580=>"101110111",
  26581=>"000100001",
  26582=>"011111010",
  26583=>"111111000",
  26584=>"010001111",
  26585=>"110101011",
  26586=>"111000001",
  26587=>"000101001",
  26588=>"101111111",
  26589=>"111010111",
  26590=>"110011111",
  26591=>"011000101",
  26592=>"111100110",
  26593=>"011000000",
  26594=>"000011010",
  26595=>"010010100",
  26596=>"111001001",
  26597=>"001111000",
  26598=>"100001100",
  26599=>"011010011",
  26600=>"101100001",
  26601=>"001010010",
  26602=>"001110010",
  26603=>"100001010",
  26604=>"001010111",
  26605=>"000010101",
  26606=>"000101001",
  26607=>"110111110",
  26608=>"110110001",
  26609=>"001110000",
  26610=>"011000100",
  26611=>"001111100",
  26612=>"100110011",
  26613=>"110000101",
  26614=>"010110001",
  26615=>"000011100",
  26616=>"001111011",
  26617=>"010101011",
  26618=>"010010010",
  26619=>"011100000",
  26620=>"110000010",
  26621=>"010001000",
  26622=>"010001010",
  26623=>"110111001",
  26624=>"011011111",
  26625=>"000011001",
  26626=>"101110110",
  26627=>"101100011",
  26628=>"001110101",
  26629=>"110100100",
  26630=>"011010100",
  26631=>"111010011",
  26632=>"110111101",
  26633=>"111001000",
  26634=>"010011001",
  26635=>"010010010",
  26636=>"001001001",
  26637=>"100101100",
  26638=>"011001010",
  26639=>"001000100",
  26640=>"101101100",
  26641=>"011001101",
  26642=>"111001010",
  26643=>"011100011",
  26644=>"111111101",
  26645=>"000010111",
  26646=>"110001111",
  26647=>"111110000",
  26648=>"110100101",
  26649=>"001111111",
  26650=>"110100001",
  26651=>"001001101",
  26652=>"100000001",
  26653=>"101000101",
  26654=>"111111001",
  26655=>"000010011",
  26656=>"001001010",
  26657=>"111110100",
  26658=>"011011001",
  26659=>"110000010",
  26660=>"000110111",
  26661=>"101000100",
  26662=>"101110001",
  26663=>"111011100",
  26664=>"111011011",
  26665=>"100011101",
  26666=>"001010000",
  26667=>"010010011",
  26668=>"010010000",
  26669=>"101011011",
  26670=>"000101011",
  26671=>"110000100",
  26672=>"100100111",
  26673=>"110110110",
  26674=>"111101111",
  26675=>"011110101",
  26676=>"110010110",
  26677=>"100001110",
  26678=>"111000010",
  26679=>"000010001",
  26680=>"100011000",
  26681=>"110110110",
  26682=>"000010010",
  26683=>"100110010",
  26684=>"110010111",
  26685=>"101011001",
  26686=>"111101110",
  26687=>"010111101",
  26688=>"110100000",
  26689=>"010001110",
  26690=>"001011101",
  26691=>"101110010",
  26692=>"100111110",
  26693=>"101101110",
  26694=>"001011111",
  26695=>"110000010",
  26696=>"011000000",
  26697=>"110001001",
  26698=>"100110001",
  26699=>"000100111",
  26700=>"100000111",
  26701=>"111010101",
  26702=>"001110011",
  26703=>"101100110",
  26704=>"101101100",
  26705=>"000001000",
  26706=>"110101000",
  26707=>"001011001",
  26708=>"110101010",
  26709=>"101110101",
  26710=>"111101011",
  26711=>"000010101",
  26712=>"100101110",
  26713=>"111110001",
  26714=>"001001001",
  26715=>"010011111",
  26716=>"001100111",
  26717=>"000000111",
  26718=>"111111011",
  26719=>"010100110",
  26720=>"001011110",
  26721=>"100110101",
  26722=>"111010011",
  26723=>"100001110",
  26724=>"100010111",
  26725=>"010101111",
  26726=>"001110011",
  26727=>"011111111",
  26728=>"100101100",
  26729=>"101101001",
  26730=>"100100001",
  26731=>"110010101",
  26732=>"111111100",
  26733=>"000000111",
  26734=>"000111111",
  26735=>"111101110",
  26736=>"111100010",
  26737=>"000000000",
  26738=>"000001111",
  26739=>"101110010",
  26740=>"001111100",
  26741=>"000011110",
  26742=>"011101011",
  26743=>"001100100",
  26744=>"010001110",
  26745=>"000011100",
  26746=>"001001010",
  26747=>"010010000",
  26748=>"100011111",
  26749=>"010110000",
  26750=>"000011100",
  26751=>"000000101",
  26752=>"001011100",
  26753=>"110110100",
  26754=>"100000011",
  26755=>"001011001",
  26756=>"111111011",
  26757=>"100100101",
  26758=>"110101101",
  26759=>"010111110",
  26760=>"011100010",
  26761=>"000100011",
  26762=>"000111011",
  26763=>"100011010",
  26764=>"111010110",
  26765=>"000101101",
  26766=>"000101010",
  26767=>"100110000",
  26768=>"000100110",
  26769=>"101011000",
  26770=>"001001101",
  26771=>"101001010",
  26772=>"001000001",
  26773=>"100001110",
  26774=>"001011010",
  26775=>"001000011",
  26776=>"010010110",
  26777=>"001101001",
  26778=>"001111011",
  26779=>"101010010",
  26780=>"011100111",
  26781=>"011110111",
  26782=>"111100011",
  26783=>"001000000",
  26784=>"010111010",
  26785=>"111111110",
  26786=>"111111000",
  26787=>"001111110",
  26788=>"000100110",
  26789=>"000100111",
  26790=>"110011111",
  26791=>"000110010",
  26792=>"000011100",
  26793=>"110101001",
  26794=>"000010011",
  26795=>"110101110",
  26796=>"100001100",
  26797=>"001011001",
  26798=>"100100000",
  26799=>"011111100",
  26800=>"101011111",
  26801=>"000001101",
  26802=>"100100111",
  26803=>"010101000",
  26804=>"101010001",
  26805=>"011010100",
  26806=>"111100010",
  26807=>"000100000",
  26808=>"001000011",
  26809=>"000111110",
  26810=>"010000101",
  26811=>"110011100",
  26812=>"011000011",
  26813=>"001010101",
  26814=>"111111001",
  26815=>"100100110",
  26816=>"100111001",
  26817=>"100001011",
  26818=>"111001101",
  26819=>"101011100",
  26820=>"111100110",
  26821=>"110110000",
  26822=>"000111001",
  26823=>"101001001",
  26824=>"000000011",
  26825=>"101111001",
  26826=>"110010100",
  26827=>"000011101",
  26828=>"100010001",
  26829=>"000111000",
  26830=>"100111011",
  26831=>"000010010",
  26832=>"100101110",
  26833=>"100010000",
  26834=>"011000001",
  26835=>"101101001",
  26836=>"111010111",
  26837=>"000001011",
  26838=>"001010101",
  26839=>"111111110",
  26840=>"110000001",
  26841=>"011111110",
  26842=>"111111000",
  26843=>"110001011",
  26844=>"100001001",
  26845=>"011010101",
  26846=>"001001110",
  26847=>"111100110",
  26848=>"001000101",
  26849=>"010000100",
  26850=>"001100101",
  26851=>"101011100",
  26852=>"001001001",
  26853=>"100000110",
  26854=>"000100101",
  26855=>"101110111",
  26856=>"001000010",
  26857=>"111111101",
  26858=>"010100111",
  26859=>"110111000",
  26860=>"101000001",
  26861=>"000101000",
  26862=>"000001001",
  26863=>"111010110",
  26864=>"000000000",
  26865=>"111111111",
  26866=>"000000100",
  26867=>"001000010",
  26868=>"101000110",
  26869=>"010000010",
  26870=>"111011011",
  26871=>"000101110",
  26872=>"000001000",
  26873=>"011100001",
  26874=>"101000100",
  26875=>"000011011",
  26876=>"010000101",
  26877=>"011101100",
  26878=>"101001010",
  26879=>"011000001",
  26880=>"000011100",
  26881=>"100011101",
  26882=>"111101101",
  26883=>"001011000",
  26884=>"010011101",
  26885=>"001111001",
  26886=>"001000110",
  26887=>"100100010",
  26888=>"100100000",
  26889=>"011010111",
  26890=>"011000010",
  26891=>"000000111",
  26892=>"000010110",
  26893=>"111111001",
  26894=>"011111100",
  26895=>"000000110",
  26896=>"111100010",
  26897=>"101110001",
  26898=>"000010011",
  26899=>"110101000",
  26900=>"001100001",
  26901=>"101001111",
  26902=>"000110111",
  26903=>"110111100",
  26904=>"010111100",
  26905=>"011111011",
  26906=>"000111010",
  26907=>"011011100",
  26908=>"010100001",
  26909=>"011001011",
  26910=>"111011101",
  26911=>"000010000",
  26912=>"001001001",
  26913=>"110100101",
  26914=>"000100001",
  26915=>"001110101",
  26916=>"001101111",
  26917=>"100111011",
  26918=>"111110110",
  26919=>"110110001",
  26920=>"001100001",
  26921=>"000111101",
  26922=>"110101011",
  26923=>"000000100",
  26924=>"110011000",
  26925=>"000000011",
  26926=>"001001010",
  26927=>"101011110",
  26928=>"001100000",
  26929=>"010010111",
  26930=>"100010110",
  26931=>"110111111",
  26932=>"011101110",
  26933=>"000100000",
  26934=>"000011000",
  26935=>"110000111",
  26936=>"110111110",
  26937=>"011011000",
  26938=>"110000000",
  26939=>"000011111",
  26940=>"010001101",
  26941=>"110111010",
  26942=>"101110110",
  26943=>"010101101",
  26944=>"100001010",
  26945=>"011001011",
  26946=>"000110110",
  26947=>"101110100",
  26948=>"111111111",
  26949=>"100011000",
  26950=>"001011011",
  26951=>"001010010",
  26952=>"100010111",
  26953=>"100101010",
  26954=>"011110100",
  26955=>"001000011",
  26956=>"011001110",
  26957=>"011111110",
  26958=>"101000010",
  26959=>"010101001",
  26960=>"001000000",
  26961=>"111010011",
  26962=>"001110111",
  26963=>"001010110",
  26964=>"100000001",
  26965=>"111111111",
  26966=>"001010010",
  26967=>"010110010",
  26968=>"001010100",
  26969=>"101001001",
  26970=>"110100111",
  26971=>"000111010",
  26972=>"010110000",
  26973=>"011101001",
  26974=>"011101011",
  26975=>"110101001",
  26976=>"001110001",
  26977=>"011101011",
  26978=>"101111011",
  26979=>"110101001",
  26980=>"001011011",
  26981=>"101001101",
  26982=>"000110000",
  26983=>"111000111",
  26984=>"111001111",
  26985=>"001000000",
  26986=>"110101000",
  26987=>"000000111",
  26988=>"010101101",
  26989=>"110001001",
  26990=>"010001100",
  26991=>"000001000",
  26992=>"110110111",
  26993=>"111001101",
  26994=>"000010111",
  26995=>"011000101",
  26996=>"110110000",
  26997=>"110101100",
  26998=>"111000111",
  26999=>"101111000",
  27000=>"001101010",
  27001=>"111111110",
  27002=>"111101101",
  27003=>"001110111",
  27004=>"001000001",
  27005=>"011010101",
  27006=>"010001001",
  27007=>"111111001",
  27008=>"111010101",
  27009=>"111101011",
  27010=>"111111010",
  27011=>"101010010",
  27012=>"000000011",
  27013=>"001010000",
  27014=>"001000011",
  27015=>"111100111",
  27016=>"111010101",
  27017=>"000010001",
  27018=>"000011000",
  27019=>"111001110",
  27020=>"100111110",
  27021=>"010100101",
  27022=>"101011100",
  27023=>"001010101",
  27024=>"001000011",
  27025=>"110101111",
  27026=>"011101011",
  27027=>"110110000",
  27028=>"110001010",
  27029=>"101010001",
  27030=>"011010111",
  27031=>"111001111",
  27032=>"010111000",
  27033=>"110110000",
  27034=>"001101110",
  27035=>"001101000",
  27036=>"011111000",
  27037=>"011110111",
  27038=>"010110010",
  27039=>"001101100",
  27040=>"101100011",
  27041=>"000101101",
  27042=>"010011011",
  27043=>"110010111",
  27044=>"111101010",
  27045=>"011110000",
  27046=>"101110100",
  27047=>"111111001",
  27048=>"110010110",
  27049=>"010010100",
  27050=>"000100001",
  27051=>"100100010",
  27052=>"001111111",
  27053=>"011100100",
  27054=>"011010101",
  27055=>"110100110",
  27056=>"101101011",
  27057=>"010011101",
  27058=>"010111001",
  27059=>"000100111",
  27060=>"010100100",
  27061=>"100111100",
  27062=>"011101010",
  27063=>"001001001",
  27064=>"100101110",
  27065=>"111110110",
  27066=>"010001001",
  27067=>"110000000",
  27068=>"000010100",
  27069=>"001011111",
  27070=>"001110111",
  27071=>"001111111",
  27072=>"010110000",
  27073=>"111001011",
  27074=>"110001010",
  27075=>"010111001",
  27076=>"010000000",
  27077=>"110001000",
  27078=>"010111110",
  27079=>"011000000",
  27080=>"000001100",
  27081=>"111001011",
  27082=>"100010001",
  27083=>"111010101",
  27084=>"100100100",
  27085=>"001111111",
  27086=>"000100000",
  27087=>"101110110",
  27088=>"000000101",
  27089=>"101100110",
  27090=>"100000010",
  27091=>"111110101",
  27092=>"011011100",
  27093=>"111111000",
  27094=>"101011101",
  27095=>"001111101",
  27096=>"101101101",
  27097=>"111110101",
  27098=>"001011010",
  27099=>"111100100",
  27100=>"011000111",
  27101=>"100111010",
  27102=>"011110110",
  27103=>"110010010",
  27104=>"100000110",
  27105=>"001001011",
  27106=>"000111011",
  27107=>"001111100",
  27108=>"111100110",
  27109=>"110000010",
  27110=>"010010001",
  27111=>"011011001",
  27112=>"000110110",
  27113=>"010001011",
  27114=>"011010000",
  27115=>"100111010",
  27116=>"000110010",
  27117=>"101110100",
  27118=>"000001101",
  27119=>"110111110",
  27120=>"100111111",
  27121=>"101001100",
  27122=>"010000010",
  27123=>"000010110",
  27124=>"001010000",
  27125=>"011011111",
  27126=>"100001001",
  27127=>"000100010",
  27128=>"010010101",
  27129=>"011001000",
  27130=>"001001011",
  27131=>"101000110",
  27132=>"010001100",
  27133=>"110100001",
  27134=>"000011101",
  27135=>"011000111",
  27136=>"100000010",
  27137=>"101011100",
  27138=>"100000011",
  27139=>"000001000",
  27140=>"011100110",
  27141=>"010101011",
  27142=>"111011010",
  27143=>"001110010",
  27144=>"001001101",
  27145=>"000000101",
  27146=>"101101001",
  27147=>"001110101",
  27148=>"001011100",
  27149=>"001011110",
  27150=>"100010000",
  27151=>"000100010",
  27152=>"111011101",
  27153=>"101011111",
  27154=>"100100011",
  27155=>"101100100",
  27156=>"000100000",
  27157=>"010100000",
  27158=>"000000110",
  27159=>"101111101",
  27160=>"001000000",
  27161=>"111111001",
  27162=>"011101011",
  27163=>"101010001",
  27164=>"110001111",
  27165=>"011000010",
  27166=>"110111100",
  27167=>"111100100",
  27168=>"111001100",
  27169=>"001011101",
  27170=>"101010110",
  27171=>"111011001",
  27172=>"110101110",
  27173=>"111011001",
  27174=>"101011101",
  27175=>"101011111",
  27176=>"010010011",
  27177=>"000110110",
  27178=>"010000010",
  27179=>"101001110",
  27180=>"110111110",
  27181=>"100111010",
  27182=>"010010000",
  27183=>"110011100",
  27184=>"000111110",
  27185=>"011011100",
  27186=>"000100111",
  27187=>"100000010",
  27188=>"110101011",
  27189=>"000011110",
  27190=>"100101001",
  27191=>"110100011",
  27192=>"011010011",
  27193=>"110110110",
  27194=>"011000100",
  27195=>"001011111",
  27196=>"110010111",
  27197=>"000011101",
  27198=>"010000101",
  27199=>"110000110",
  27200=>"000111110",
  27201=>"011011001",
  27202=>"101111001",
  27203=>"000100011",
  27204=>"111010110",
  27205=>"000011001",
  27206=>"101011101",
  27207=>"111111010",
  27208=>"010100011",
  27209=>"110000110",
  27210=>"111110000",
  27211=>"100111111",
  27212=>"111110010",
  27213=>"111111100",
  27214=>"111110000",
  27215=>"111001000",
  27216=>"110000111",
  27217=>"100101101",
  27218=>"100000011",
  27219=>"111010011",
  27220=>"011000000",
  27221=>"001101000",
  27222=>"011001101",
  27223=>"101111011",
  27224=>"000110101",
  27225=>"111100000",
  27226=>"111011110",
  27227=>"110001100",
  27228=>"111111000",
  27229=>"010100000",
  27230=>"101011100",
  27231=>"000000110",
  27232=>"101111000",
  27233=>"100001001",
  27234=>"011000001",
  27235=>"101010111",
  27236=>"110111000",
  27237=>"011110010",
  27238=>"001001111",
  27239=>"111100110",
  27240=>"010011000",
  27241=>"111101100",
  27242=>"101000100",
  27243=>"010010111",
  27244=>"110000000",
  27245=>"001010001",
  27246=>"001111100",
  27247=>"101111001",
  27248=>"000110111",
  27249=>"010100001",
  27250=>"001001001",
  27251=>"100111010",
  27252=>"000010011",
  27253=>"101101010",
  27254=>"000000010",
  27255=>"011001000",
  27256=>"010111101",
  27257=>"011011001",
  27258=>"001101011",
  27259=>"010101101",
  27260=>"011010100",
  27261=>"100011010",
  27262=>"001011000",
  27263=>"000101010",
  27264=>"110101111",
  27265=>"010101110",
  27266=>"000110101",
  27267=>"011100001",
  27268=>"010100111",
  27269=>"110011101",
  27270=>"110100011",
  27271=>"111011111",
  27272=>"111010001",
  27273=>"000101001",
  27274=>"011101000",
  27275=>"110000001",
  27276=>"111010111",
  27277=>"010000100",
  27278=>"011111100",
  27279=>"000100111",
  27280=>"000010001",
  27281=>"100011000",
  27282=>"100001100",
  27283=>"101111111",
  27284=>"001000001",
  27285=>"010001110",
  27286=>"100110001",
  27287=>"001000010",
  27288=>"011010101",
  27289=>"010000000",
  27290=>"110010011",
  27291=>"000100000",
  27292=>"010101100",
  27293=>"000011101",
  27294=>"101011101",
  27295=>"000100000",
  27296=>"101100010",
  27297=>"000111000",
  27298=>"111110000",
  27299=>"111101111",
  27300=>"000001100",
  27301=>"001100101",
  27302=>"100010010",
  27303=>"100111011",
  27304=>"111000011",
  27305=>"011000010",
  27306=>"101000111",
  27307=>"001000100",
  27308=>"011110000",
  27309=>"100101101",
  27310=>"101110010",
  27311=>"110011010",
  27312=>"101000100",
  27313=>"111010001",
  27314=>"010001111",
  27315=>"010011111",
  27316=>"010000011",
  27317=>"011110001",
  27318=>"010100011",
  27319=>"011010001",
  27320=>"000100100",
  27321=>"010010111",
  27322=>"111010011",
  27323=>"101100110",
  27324=>"101000011",
  27325=>"101110010",
  27326=>"010110111",
  27327=>"000100101",
  27328=>"011011111",
  27329=>"111101110",
  27330=>"101111110",
  27331=>"000110111",
  27332=>"001110010",
  27333=>"101000110",
  27334=>"110110010",
  27335=>"000110100",
  27336=>"010100001",
  27337=>"010000100",
  27338=>"001101101",
  27339=>"010000100",
  27340=>"111101010",
  27341=>"100111100",
  27342=>"110010101",
  27343=>"011101001",
  27344=>"000001100",
  27345=>"110110101",
  27346=>"011111011",
  27347=>"111000111",
  27348=>"011101010",
  27349=>"010110111",
  27350=>"010110101",
  27351=>"100011011",
  27352=>"111010110",
  27353=>"111101010",
  27354=>"001101101",
  27355=>"000001011",
  27356=>"110000001",
  27357=>"111010110",
  27358=>"000000111",
  27359=>"010110010",
  27360=>"010100110",
  27361=>"101110010",
  27362=>"001101000",
  27363=>"101100010",
  27364=>"001100011",
  27365=>"000101101",
  27366=>"111010100",
  27367=>"001010000",
  27368=>"010010111",
  27369=>"010011110",
  27370=>"010001010",
  27371=>"001111101",
  27372=>"110101101",
  27373=>"011101101",
  27374=>"011110000",
  27375=>"010111001",
  27376=>"010100110",
  27377=>"001000100",
  27378=>"001010110",
  27379=>"010010010",
  27380=>"001101000",
  27381=>"001110011",
  27382=>"000000101",
  27383=>"011001011",
  27384=>"110001100",
  27385=>"100111001",
  27386=>"000000100",
  27387=>"000000111",
  27388=>"001101001",
  27389=>"111101010",
  27390=>"101111000",
  27391=>"001100010",
  27392=>"001011101",
  27393=>"100110010",
  27394=>"010111110",
  27395=>"000010011",
  27396=>"011110101",
  27397=>"010111111",
  27398=>"010000001",
  27399=>"110011000",
  27400=>"000101001",
  27401=>"000010001",
  27402=>"111101000",
  27403=>"011011110",
  27404=>"001011010",
  27405=>"101100010",
  27406=>"100001111",
  27407=>"100101100",
  27408=>"101010100",
  27409=>"000101000",
  27410=>"011101001",
  27411=>"010000011",
  27412=>"101100101",
  27413=>"110101000",
  27414=>"110011000",
  27415=>"011000011",
  27416=>"111100110",
  27417=>"110111001",
  27418=>"001010001",
  27419=>"000010000",
  27420=>"101111010",
  27421=>"000101111",
  27422=>"011101111",
  27423=>"011010010",
  27424=>"010110010",
  27425=>"000111010",
  27426=>"001001010",
  27427=>"000001011",
  27428=>"001100110",
  27429=>"100010111",
  27430=>"001101100",
  27431=>"110100000",
  27432=>"000111001",
  27433=>"001011101",
  27434=>"100100010",
  27435=>"100011111",
  27436=>"011101100",
  27437=>"001011110",
  27438=>"101010000",
  27439=>"000100000",
  27440=>"111101111",
  27441=>"000101100",
  27442=>"111011000",
  27443=>"010100010",
  27444=>"101010100",
  27445=>"110010010",
  27446=>"101011100",
  27447=>"100000000",
  27448=>"000010110",
  27449=>"010110001",
  27450=>"011011111",
  27451=>"001000111",
  27452=>"011101010",
  27453=>"101000000",
  27454=>"100000111",
  27455=>"111100011",
  27456=>"000101110",
  27457=>"011011000",
  27458=>"011000111",
  27459=>"100101111",
  27460=>"100000110",
  27461=>"100110111",
  27462=>"100001111",
  27463=>"011000101",
  27464=>"001101010",
  27465=>"111001101",
  27466=>"001010100",
  27467=>"101100000",
  27468=>"000101010",
  27469=>"001011110",
  27470=>"111111000",
  27471=>"100011001",
  27472=>"010101001",
  27473=>"111000110",
  27474=>"110001011",
  27475=>"100010110",
  27476=>"111010000",
  27477=>"101111011",
  27478=>"100011101",
  27479=>"101110100",
  27480=>"100010001",
  27481=>"011100110",
  27482=>"000100110",
  27483=>"000000110",
  27484=>"111110101",
  27485=>"000111001",
  27486=>"011110001",
  27487=>"000101000",
  27488=>"011101000",
  27489=>"000000100",
  27490=>"000111101",
  27491=>"110000011",
  27492=>"000011111",
  27493=>"011011001",
  27494=>"100001111",
  27495=>"111110101",
  27496=>"010100101",
  27497=>"111010000",
  27498=>"010110100",
  27499=>"110000100",
  27500=>"110101111",
  27501=>"001001000",
  27502=>"011001101",
  27503=>"101001010",
  27504=>"001110010",
  27505=>"000111111",
  27506=>"000101101",
  27507=>"011001101",
  27508=>"111001110",
  27509=>"111111110",
  27510=>"000110011",
  27511=>"011011110",
  27512=>"110000110",
  27513=>"001010101",
  27514=>"110000001",
  27515=>"111000110",
  27516=>"101111101",
  27517=>"110011101",
  27518=>"100101010",
  27519=>"100100010",
  27520=>"000101111",
  27521=>"111100110",
  27522=>"110010010",
  27523=>"110101101",
  27524=>"100010101",
  27525=>"001100100",
  27526=>"011100101",
  27527=>"011001111",
  27528=>"110111111",
  27529=>"101100001",
  27530=>"101111000",
  27531=>"011111000",
  27532=>"101000001",
  27533=>"110110101",
  27534=>"101100111",
  27535=>"110101111",
  27536=>"110011010",
  27537=>"001110100",
  27538=>"110110010",
  27539=>"101111100",
  27540=>"110000110",
  27541=>"000000110",
  27542=>"011000001",
  27543=>"010110110",
  27544=>"010000110",
  27545=>"010011100",
  27546=>"100110010",
  27547=>"001111011",
  27548=>"010010101",
  27549=>"101000000",
  27550=>"101110111",
  27551=>"111100000",
  27552=>"011011010",
  27553=>"000101001",
  27554=>"010110101",
  27555=>"010010000",
  27556=>"101110000",
  27557=>"000011110",
  27558=>"100000101",
  27559=>"010110101",
  27560=>"101100001",
  27561=>"111001111",
  27562=>"000101110",
  27563=>"100011011",
  27564=>"100001100",
  27565=>"011000011",
  27566=>"100001000",
  27567=>"010000011",
  27568=>"111010101",
  27569=>"001100100",
  27570=>"111101000",
  27571=>"001000000",
  27572=>"111111100",
  27573=>"101011011",
  27574=>"100110001",
  27575=>"000011110",
  27576=>"100100011",
  27577=>"110011011",
  27578=>"110110100",
  27579=>"001111100",
  27580=>"010101010",
  27581=>"011111001",
  27582=>"000010000",
  27583=>"001100000",
  27584=>"000010001",
  27585=>"000100010",
  27586=>"100111001",
  27587=>"111010001",
  27588=>"000001001",
  27589=>"111100010",
  27590=>"000011110",
  27591=>"000111011",
  27592=>"100101110",
  27593=>"000010010",
  27594=>"110000000",
  27595=>"001100110",
  27596=>"110001000",
  27597=>"110100100",
  27598=>"010001011",
  27599=>"111001010",
  27600=>"001010101",
  27601=>"100000110",
  27602=>"011100010",
  27603=>"001000101",
  27604=>"000100011",
  27605=>"000100111",
  27606=>"001001000",
  27607=>"111001000",
  27608=>"001001010",
  27609=>"100110010",
  27610=>"100110111",
  27611=>"111100000",
  27612=>"111101111",
  27613=>"000111010",
  27614=>"000010010",
  27615=>"001100000",
  27616=>"100000100",
  27617=>"000111101",
  27618=>"000001000",
  27619=>"000100001",
  27620=>"010011010",
  27621=>"010101011",
  27622=>"011110110",
  27623=>"011111111",
  27624=>"001101101",
  27625=>"000011001",
  27626=>"001001100",
  27627=>"001000110",
  27628=>"011011010",
  27629=>"001011100",
  27630=>"100100100",
  27631=>"100011111",
  27632=>"000101011",
  27633=>"011011000",
  27634=>"001111101",
  27635=>"010000100",
  27636=>"100001110",
  27637=>"110100000",
  27638=>"000110001",
  27639=>"011010111",
  27640=>"010000101",
  27641=>"101110010",
  27642=>"100001011",
  27643=>"110011000",
  27644=>"100001011",
  27645=>"001111100",
  27646=>"111001101",
  27647=>"001000100",
  27648=>"000001101",
  27649=>"101111111",
  27650=>"101000010",
  27651=>"101010000",
  27652=>"001111111",
  27653=>"111001011",
  27654=>"000111001",
  27655=>"110010001",
  27656=>"111110110",
  27657=>"010000000",
  27658=>"011010011",
  27659=>"010011110",
  27660=>"110010010",
  27661=>"001110010",
  27662=>"010010000",
  27663=>"010000001",
  27664=>"111000111",
  27665=>"000000010",
  27666=>"000101010",
  27667=>"001010110",
  27668=>"101000111",
  27669=>"000010000",
  27670=>"000110010",
  27671=>"010001000",
  27672=>"001100101",
  27673=>"110001110",
  27674=>"111000001",
  27675=>"101100110",
  27676=>"001101011",
  27677=>"101001101",
  27678=>"011000000",
  27679=>"001000000",
  27680=>"100110110",
  27681=>"011000011",
  27682=>"100100111",
  27683=>"100111111",
  27684=>"000110011",
  27685=>"101101111",
  27686=>"101011111",
  27687=>"010111000",
  27688=>"000000111",
  27689=>"000000100",
  27690=>"101000111",
  27691=>"011010110",
  27692=>"101010110",
  27693=>"011000110",
  27694=>"000100011",
  27695=>"010101010",
  27696=>"010101100",
  27697=>"111011101",
  27698=>"111100111",
  27699=>"110100001",
  27700=>"100101000",
  27701=>"101100110",
  27702=>"111001100",
  27703=>"000010010",
  27704=>"010110011",
  27705=>"000100110",
  27706=>"100111110",
  27707=>"001101001",
  27708=>"011100000",
  27709=>"011000110",
  27710=>"011101100",
  27711=>"011010111",
  27712=>"101001110",
  27713=>"011001100",
  27714=>"110100100",
  27715=>"001101100",
  27716=>"110100000",
  27717=>"001001001",
  27718=>"110010010",
  27719=>"100001111",
  27720=>"111101100",
  27721=>"010011011",
  27722=>"110110000",
  27723=>"111001100",
  27724=>"100100000",
  27725=>"111100100",
  27726=>"100101101",
  27727=>"101110011",
  27728=>"110011100",
  27729=>"010011001",
  27730=>"001101101",
  27731=>"101000100",
  27732=>"000010111",
  27733=>"010100111",
  27734=>"001010100",
  27735=>"110101000",
  27736=>"101001011",
  27737=>"110101011",
  27738=>"001011001",
  27739=>"110000010",
  27740=>"100011001",
  27741=>"100001010",
  27742=>"011011001",
  27743=>"101001110",
  27744=>"010001111",
  27745=>"011111111",
  27746=>"000011011",
  27747=>"001011100",
  27748=>"110001100",
  27749=>"010100011",
  27750=>"101100001",
  27751=>"001001000",
  27752=>"000100101",
  27753=>"000000110",
  27754=>"111101001",
  27755=>"000110101",
  27756=>"000010010",
  27757=>"110100101",
  27758=>"110100111",
  27759=>"111001010",
  27760=>"000001000",
  27761=>"110001111",
  27762=>"011011100",
  27763=>"000101101",
  27764=>"111110001",
  27765=>"010111001",
  27766=>"000111010",
  27767=>"111101001",
  27768=>"100001101",
  27769=>"111111100",
  27770=>"101100010",
  27771=>"101110101",
  27772=>"110101100",
  27773=>"011111001",
  27774=>"110011100",
  27775=>"101010111",
  27776=>"000100011",
  27777=>"010001100",
  27778=>"101001111",
  27779=>"000001000",
  27780=>"001001001",
  27781=>"110000010",
  27782=>"011010011",
  27783=>"010001000",
  27784=>"100100011",
  27785=>"010101100",
  27786=>"010110101",
  27787=>"101000111",
  27788=>"100110010",
  27789=>"110011111",
  27790=>"111010100",
  27791=>"011111010",
  27792=>"011000011",
  27793=>"001001000",
  27794=>"000100000",
  27795=>"001110011",
  27796=>"001001100",
  27797=>"000110001",
  27798=>"101110101",
  27799=>"100100000",
  27800=>"111001110",
  27801=>"100111100",
  27802=>"110000100",
  27803=>"110010000",
  27804=>"010011010",
  27805=>"100001000",
  27806=>"000101101",
  27807=>"011111000",
  27808=>"100100100",
  27809=>"111110001",
  27810=>"100100011",
  27811=>"011000111",
  27812=>"110000001",
  27813=>"101011001",
  27814=>"111110001",
  27815=>"010010011",
  27816=>"001111000",
  27817=>"010001111",
  27818=>"110111111",
  27819=>"011101101",
  27820=>"011100000",
  27821=>"110111100",
  27822=>"100011100",
  27823=>"111000110",
  27824=>"011111100",
  27825=>"010001000",
  27826=>"000010110",
  27827=>"110010111",
  27828=>"000100001",
  27829=>"010011000",
  27830=>"010110101",
  27831=>"101110101",
  27832=>"010111010",
  27833=>"100010110",
  27834=>"000101000",
  27835=>"110001000",
  27836=>"101000100",
  27837=>"001110001",
  27838=>"111100001",
  27839=>"101101100",
  27840=>"010011100",
  27841=>"101000110",
  27842=>"011110010",
  27843=>"011011010",
  27844=>"111111100",
  27845=>"111101111",
  27846=>"100010101",
  27847=>"001110010",
  27848=>"000010000",
  27849=>"010111000",
  27850=>"000100100",
  27851=>"001100001",
  27852=>"011111001",
  27853=>"111011110",
  27854=>"000110111",
  27855=>"000010010",
  27856=>"110010001",
  27857=>"111101011",
  27858=>"010000010",
  27859=>"101001111",
  27860=>"011101001",
  27861=>"001010001",
  27862=>"110001010",
  27863=>"101000001",
  27864=>"000001111",
  27865=>"001010001",
  27866=>"100101110",
  27867=>"001010101",
  27868=>"001011111",
  27869=>"010111111",
  27870=>"101011100",
  27871=>"101110011",
  27872=>"111111110",
  27873=>"011010001",
  27874=>"111010001",
  27875=>"000110110",
  27876=>"100001010",
  27877=>"101110011",
  27878=>"001000101",
  27879=>"011001111",
  27880=>"011101111",
  27881=>"110100101",
  27882=>"111010100",
  27883=>"011000111",
  27884=>"100000100",
  27885=>"010110100",
  27886=>"000000110",
  27887=>"000000101",
  27888=>"101001011",
  27889=>"101111000",
  27890=>"001110101",
  27891=>"000100100",
  27892=>"110001000",
  27893=>"101000100",
  27894=>"010011011",
  27895=>"101000000",
  27896=>"001100001",
  27897=>"101110010",
  27898=>"101010000",
  27899=>"000011000",
  27900=>"010101000",
  27901=>"011001011",
  27902=>"011000110",
  27903=>"111110011",
  27904=>"000101011",
  27905=>"011100011",
  27906=>"111100000",
  27907=>"000110101",
  27908=>"011010110",
  27909=>"000011110",
  27910=>"011010001",
  27911=>"110000000",
  27912=>"001111011",
  27913=>"110011100",
  27914=>"111101111",
  27915=>"010000000",
  27916=>"000101111",
  27917=>"101010101",
  27918=>"000000001",
  27919=>"100011010",
  27920=>"001101001",
  27921=>"110001100",
  27922=>"000011111",
  27923=>"000101011",
  27924=>"000100010",
  27925=>"000110001",
  27926=>"111111000",
  27927=>"100110111",
  27928=>"110001101",
  27929=>"001100100",
  27930=>"010111100",
  27931=>"000100001",
  27932=>"111010110",
  27933=>"011001111",
  27934=>"010011111",
  27935=>"101011001",
  27936=>"000100100",
  27937=>"010001001",
  27938=>"101111100",
  27939=>"011011011",
  27940=>"100010011",
  27941=>"000100010",
  27942=>"111011110",
  27943=>"100100001",
  27944=>"011000001",
  27945=>"010000011",
  27946=>"011010000",
  27947=>"001011000",
  27948=>"001010001",
  27949=>"111011000",
  27950=>"111111100",
  27951=>"000111011",
  27952=>"000001011",
  27953=>"010101101",
  27954=>"011000111",
  27955=>"111100111",
  27956=>"100100101",
  27957=>"101001111",
  27958=>"111100001",
  27959=>"001000111",
  27960=>"101010010",
  27961=>"110101111",
  27962=>"101100110",
  27963=>"101000001",
  27964=>"011110101",
  27965=>"111010110",
  27966=>"101101101",
  27967=>"111100101",
  27968=>"010001001",
  27969=>"000101100",
  27970=>"110110010",
  27971=>"010010001",
  27972=>"000111011",
  27973=>"001001011",
  27974=>"010101001",
  27975=>"010110010",
  27976=>"110001011",
  27977=>"110000101",
  27978=>"101101111",
  27979=>"010101100",
  27980=>"001101010",
  27981=>"100100111",
  27982=>"111110010",
  27983=>"001011010",
  27984=>"011010110",
  27985=>"101110011",
  27986=>"010001000",
  27987=>"010011100",
  27988=>"101100111",
  27989=>"111101111",
  27990=>"100000000",
  27991=>"000101001",
  27992=>"010010100",
  27993=>"000010100",
  27994=>"101000010",
  27995=>"011101100",
  27996=>"101001101",
  27997=>"001111100",
  27998=>"101001001",
  27999=>"000101010",
  28000=>"001111111",
  28001=>"101111000",
  28002=>"101101011",
  28003=>"000001110",
  28004=>"001111001",
  28005=>"100000101",
  28006=>"100001100",
  28007=>"010100111",
  28008=>"010010001",
  28009=>"100110001",
  28010=>"000110110",
  28011=>"101111101",
  28012=>"011011000",
  28013=>"101110101",
  28014=>"111100000",
  28015=>"000110101",
  28016=>"111100100",
  28017=>"101110110",
  28018=>"111101011",
  28019=>"001000001",
  28020=>"010111001",
  28021=>"110000100",
  28022=>"111010100",
  28023=>"000101000",
  28024=>"011110110",
  28025=>"100101001",
  28026=>"000001110",
  28027=>"111001111",
  28028=>"100100000",
  28029=>"100000111",
  28030=>"110100000",
  28031=>"001110010",
  28032=>"000010100",
  28033=>"001011011",
  28034=>"101111101",
  28035=>"110010000",
  28036=>"000011011",
  28037=>"100101011",
  28038=>"110111001",
  28039=>"101100101",
  28040=>"001100010",
  28041=>"010011001",
  28042=>"101111111",
  28043=>"100011010",
  28044=>"001101101",
  28045=>"111100010",
  28046=>"011100010",
  28047=>"011000011",
  28048=>"111010001",
  28049=>"101101110",
  28050=>"010011001",
  28051=>"001100010",
  28052=>"100111001",
  28053=>"110010001",
  28054=>"000110111",
  28055=>"011011001",
  28056=>"110110010",
  28057=>"010011010",
  28058=>"111111011",
  28059=>"001111010",
  28060=>"010000100",
  28061=>"000000110",
  28062=>"110000111",
  28063=>"101001001",
  28064=>"100111110",
  28065=>"110001000",
  28066=>"001001101",
  28067=>"010011100",
  28068=>"100111110",
  28069=>"100101101",
  28070=>"100110001",
  28071=>"100010010",
  28072=>"010000101",
  28073=>"001000111",
  28074=>"110010111",
  28075=>"010001000",
  28076=>"001101001",
  28077=>"001111100",
  28078=>"000000110",
  28079=>"100001111",
  28080=>"100110010",
  28081=>"011011111",
  28082=>"110100001",
  28083=>"100111011",
  28084=>"000001011",
  28085=>"100110110",
  28086=>"111011100",
  28087=>"111001110",
  28088=>"101100110",
  28089=>"001011100",
  28090=>"010111101",
  28091=>"100101100",
  28092=>"101100110",
  28093=>"010100000",
  28094=>"000100000",
  28095=>"011010011",
  28096=>"111111010",
  28097=>"110111011",
  28098=>"000110111",
  28099=>"000011101",
  28100=>"110111001",
  28101=>"100111110",
  28102=>"111110011",
  28103=>"010000000",
  28104=>"001001111",
  28105=>"010011101",
  28106=>"100001100",
  28107=>"010011101",
  28108=>"111101110",
  28109=>"111000011",
  28110=>"000111011",
  28111=>"101001011",
  28112=>"111101110",
  28113=>"001110101",
  28114=>"000001011",
  28115=>"110011100",
  28116=>"101100111",
  28117=>"110000110",
  28118=>"110100010",
  28119=>"011000000",
  28120=>"000011000",
  28121=>"101011010",
  28122=>"011111100",
  28123=>"101011011",
  28124=>"001011011",
  28125=>"000000000",
  28126=>"100001110",
  28127=>"111001011",
  28128=>"111101100",
  28129=>"001001010",
  28130=>"001011001",
  28131=>"000100010",
  28132=>"111110001",
  28133=>"010110010",
  28134=>"101100000",
  28135=>"110100000",
  28136=>"110101110",
  28137=>"100000110",
  28138=>"101010111",
  28139=>"110100011",
  28140=>"100001001",
  28141=>"000101110",
  28142=>"101101100",
  28143=>"101000100",
  28144=>"001111010",
  28145=>"101100010",
  28146=>"010000010",
  28147=>"000011101",
  28148=>"000110111",
  28149=>"100101010",
  28150=>"010111001",
  28151=>"001100101",
  28152=>"011100001",
  28153=>"001111101",
  28154=>"010110000",
  28155=>"101110011",
  28156=>"001100111",
  28157=>"000100001",
  28158=>"110001100",
  28159=>"000111111",
  28160=>"100100000",
  28161=>"001010011",
  28162=>"010111100",
  28163=>"011000100",
  28164=>"011111000",
  28165=>"111110110",
  28166=>"010111100",
  28167=>"010111011",
  28168=>"111010000",
  28169=>"000111100",
  28170=>"000000100",
  28171=>"101000000",
  28172=>"111011010",
  28173=>"101010000",
  28174=>"011111001",
  28175=>"101101001",
  28176=>"000001010",
  28177=>"001100110",
  28178=>"000010001",
  28179=>"001010101",
  28180=>"001101010",
  28181=>"100110111",
  28182=>"000110100",
  28183=>"011010110",
  28184=>"111011111",
  28185=>"001001001",
  28186=>"111000100",
  28187=>"101011101",
  28188=>"000110001",
  28189=>"010010010",
  28190=>"000100110",
  28191=>"000011011",
  28192=>"001001010",
  28193=>"010101110",
  28194=>"001110101",
  28195=>"001011000",
  28196=>"110001010",
  28197=>"011000010",
  28198=>"010001101",
  28199=>"100101000",
  28200=>"010010000",
  28201=>"100101111",
  28202=>"100000101",
  28203=>"101101111",
  28204=>"100001001",
  28205=>"011100110",
  28206=>"111101111",
  28207=>"000111000",
  28208=>"100111000",
  28209=>"101110011",
  28210=>"110110011",
  28211=>"000001110",
  28212=>"001110110",
  28213=>"100001000",
  28214=>"000001011",
  28215=>"000001011",
  28216=>"000111111",
  28217=>"100010001",
  28218=>"111111111",
  28219=>"011001101",
  28220=>"101000001",
  28221=>"111111000",
  28222=>"010000001",
  28223=>"001111100",
  28224=>"111011001",
  28225=>"101010001",
  28226=>"000100110",
  28227=>"000111100",
  28228=>"100001110",
  28229=>"010100001",
  28230=>"011100100",
  28231=>"101010101",
  28232=>"010110010",
  28233=>"110100001",
  28234=>"100110010",
  28235=>"010100110",
  28236=>"110011100",
  28237=>"100111100",
  28238=>"000101000",
  28239=>"011111110",
  28240=>"101000011",
  28241=>"000010100",
  28242=>"000110001",
  28243=>"000111011",
  28244=>"001001000",
  28245=>"011010011",
  28246=>"000000101",
  28247=>"111011001",
  28248=>"000101010",
  28249=>"110000111",
  28250=>"101010110",
  28251=>"000101000",
  28252=>"101001010",
  28253=>"010101010",
  28254=>"110110101",
  28255=>"001101101",
  28256=>"110100111",
  28257=>"001100110",
  28258=>"000100011",
  28259=>"011100100",
  28260=>"110101001",
  28261=>"000100100",
  28262=>"000011100",
  28263=>"101100011",
  28264=>"110100001",
  28265=>"001000011",
  28266=>"010010111",
  28267=>"011111010",
  28268=>"100000010",
  28269=>"101110110",
  28270=>"110010111",
  28271=>"011001110",
  28272=>"010101010",
  28273=>"101001000",
  28274=>"110100000",
  28275=>"000001000",
  28276=>"101100110",
  28277=>"000111000",
  28278=>"010111100",
  28279=>"000101010",
  28280=>"001010000",
  28281=>"011100010",
  28282=>"000011000",
  28283=>"111100111",
  28284=>"101100100",
  28285=>"010000000",
  28286=>"001000101",
  28287=>"010010111",
  28288=>"000010000",
  28289=>"101001100",
  28290=>"000100110",
  28291=>"000100011",
  28292=>"101110010",
  28293=>"011010111",
  28294=>"010111110",
  28295=>"010001011",
  28296=>"000000001",
  28297=>"001110001",
  28298=>"000111001",
  28299=>"011111000",
  28300=>"100111001",
  28301=>"010000111",
  28302=>"011000000",
  28303=>"011001111",
  28304=>"011111111",
  28305=>"010000101",
  28306=>"011011111",
  28307=>"100011011",
  28308=>"111110000",
  28309=>"111100010",
  28310=>"101000111",
  28311=>"011110011",
  28312=>"110111100",
  28313=>"001001110",
  28314=>"001011010",
  28315=>"101111110",
  28316=>"111110011",
  28317=>"010011011",
  28318=>"101000000",
  28319=>"010011000",
  28320=>"010011100",
  28321=>"100101000",
  28322=>"110111101",
  28323=>"001101111",
  28324=>"111010000",
  28325=>"011000001",
  28326=>"011100110",
  28327=>"000101100",
  28328=>"101010110",
  28329=>"000101101",
  28330=>"100010010",
  28331=>"000101000",
  28332=>"100101001",
  28333=>"100100010",
  28334=>"011101111",
  28335=>"000100001",
  28336=>"100110101",
  28337=>"010010100",
  28338=>"100110100",
  28339=>"011001010",
  28340=>"011000010",
  28341=>"000101110",
  28342=>"011110011",
  28343=>"101010011",
  28344=>"010101001",
  28345=>"101100000",
  28346=>"110100011",
  28347=>"111100111",
  28348=>"011010100",
  28349=>"011010101",
  28350=>"100000110",
  28351=>"010010100",
  28352=>"111001000",
  28353=>"111011001",
  28354=>"101110110",
  28355=>"100000010",
  28356=>"001001000",
  28357=>"110101000",
  28358=>"111110001",
  28359=>"011011000",
  28360=>"111011111",
  28361=>"001111111",
  28362=>"011010000",
  28363=>"101011110",
  28364=>"010000010",
  28365=>"001110010",
  28366=>"111010100",
  28367=>"010000000",
  28368=>"110111111",
  28369=>"010110000",
  28370=>"010000010",
  28371=>"100011111",
  28372=>"111011111",
  28373=>"011101110",
  28374=>"111011001",
  28375=>"001010101",
  28376=>"110010001",
  28377=>"111000110",
  28378=>"110111110",
  28379=>"101111010",
  28380=>"001010111",
  28381=>"010010110",
  28382=>"001111010",
  28383=>"100010000",
  28384=>"100000111",
  28385=>"000011001",
  28386=>"110001111",
  28387=>"011011000",
  28388=>"000001110",
  28389=>"110011110",
  28390=>"000111010",
  28391=>"011111100",
  28392=>"001011100",
  28393=>"110011010",
  28394=>"000100010",
  28395=>"000001101",
  28396=>"011011010",
  28397=>"011101110",
  28398=>"000000010",
  28399=>"111111111",
  28400=>"011101111",
  28401=>"101101111",
  28402=>"000001010",
  28403=>"110010100",
  28404=>"111010001",
  28405=>"000111011",
  28406=>"101010111",
  28407=>"001101000",
  28408=>"111011110",
  28409=>"010001100",
  28410=>"100001110",
  28411=>"000000001",
  28412=>"001100001",
  28413=>"100011101",
  28414=>"001100100",
  28415=>"101101001",
  28416=>"100100100",
  28417=>"100011010",
  28418=>"000101101",
  28419=>"111000111",
  28420=>"010000011",
  28421=>"100110001",
  28422=>"111000010",
  28423=>"101000001",
  28424=>"010011111",
  28425=>"111101111",
  28426=>"111101000",
  28427=>"110010101",
  28428=>"111010100",
  28429=>"001000101",
  28430=>"110111001",
  28431=>"111101011",
  28432=>"000001010",
  28433=>"010101101",
  28434=>"101010100",
  28435=>"101010011",
  28436=>"011001000",
  28437=>"000110111",
  28438=>"110000011",
  28439=>"001000101",
  28440=>"001101100",
  28441=>"010101110",
  28442=>"100010110",
  28443=>"110000101",
  28444=>"101101010",
  28445=>"110000000",
  28446=>"001111011",
  28447=>"111101000",
  28448=>"101001010",
  28449=>"111100110",
  28450=>"000001010",
  28451=>"111011000",
  28452=>"111011111",
  28453=>"101110010",
  28454=>"111011011",
  28455=>"011010111",
  28456=>"010001100",
  28457=>"100001111",
  28458=>"110010010",
  28459=>"110010111",
  28460=>"010111110",
  28461=>"000000110",
  28462=>"001011000",
  28463=>"110101100",
  28464=>"110111010",
  28465=>"011011001",
  28466=>"111011100",
  28467=>"000110110",
  28468=>"110101111",
  28469=>"111000011",
  28470=>"100010011",
  28471=>"000110110",
  28472=>"100000000",
  28473=>"111111110",
  28474=>"111110011",
  28475=>"011010010",
  28476=>"010111010",
  28477=>"011110010",
  28478=>"010001000",
  28479=>"001011111",
  28480=>"110010100",
  28481=>"011001101",
  28482=>"100101111",
  28483=>"000101000",
  28484=>"000100111",
  28485=>"111111110",
  28486=>"100111111",
  28487=>"110010100",
  28488=>"110001011",
  28489=>"000010010",
  28490=>"011010011",
  28491=>"111101010",
  28492=>"011110000",
  28493=>"110111001",
  28494=>"000010010",
  28495=>"011011111",
  28496=>"111111101",
  28497=>"111001110",
  28498=>"100010111",
  28499=>"101101010",
  28500=>"110011110",
  28501=>"110011000",
  28502=>"001110000",
  28503=>"101100010",
  28504=>"001001000",
  28505=>"011111011",
  28506=>"001111101",
  28507=>"000011100",
  28508=>"010100011",
  28509=>"001111111",
  28510=>"001011101",
  28511=>"011010100",
  28512=>"010010110",
  28513=>"101010011",
  28514=>"100000010",
  28515=>"011111001",
  28516=>"000010101",
  28517=>"110110101",
  28518=>"001110110",
  28519=>"000100100",
  28520=>"001100000",
  28521=>"110100001",
  28522=>"110100010",
  28523=>"110111000",
  28524=>"110110100",
  28525=>"011001101",
  28526=>"111100001",
  28527=>"011010011",
  28528=>"110110100",
  28529=>"111001110",
  28530=>"101101001",
  28531=>"010001101",
  28532=>"011010001",
  28533=>"100100111",
  28534=>"011001101",
  28535=>"100010001",
  28536=>"100000101",
  28537=>"011110101",
  28538=>"010000110",
  28539=>"100101111",
  28540=>"000100001",
  28541=>"101111110",
  28542=>"000011001",
  28543=>"100001100",
  28544=>"000001000",
  28545=>"100001000",
  28546=>"110000111",
  28547=>"001000010",
  28548=>"010010110",
  28549=>"011110111",
  28550=>"010110000",
  28551=>"111011000",
  28552=>"111001110",
  28553=>"010010110",
  28554=>"111010010",
  28555=>"101011011",
  28556=>"010000100",
  28557=>"001011111",
  28558=>"000001101",
  28559=>"010110000",
  28560=>"101101000",
  28561=>"000001001",
  28562=>"100110101",
  28563=>"000011100",
  28564=>"011110100",
  28565=>"001001110",
  28566=>"110111001",
  28567=>"111000100",
  28568=>"111010011",
  28569=>"011101110",
  28570=>"010100110",
  28571=>"000000011",
  28572=>"111010000",
  28573=>"011001111",
  28574=>"011110001",
  28575=>"100100100",
  28576=>"010000010",
  28577=>"100100011",
  28578=>"110011100",
  28579=>"010000110",
  28580=>"101011111",
  28581=>"101111011",
  28582=>"011011010",
  28583=>"111100011",
  28584=>"011011010",
  28585=>"110011010",
  28586=>"000011010",
  28587=>"000010101",
  28588=>"101101010",
  28589=>"100000110",
  28590=>"010111110",
  28591=>"110101101",
  28592=>"011011011",
  28593=>"100011001",
  28594=>"111010011",
  28595=>"000101110",
  28596=>"000100000",
  28597=>"000100001",
  28598=>"111110011",
  28599=>"101001101",
  28600=>"010011101",
  28601=>"110110101",
  28602=>"101000011",
  28603=>"000111010",
  28604=>"111000101",
  28605=>"000000000",
  28606=>"100100000",
  28607=>"000000000",
  28608=>"100011000",
  28609=>"111111110",
  28610=>"000101111",
  28611=>"100110000",
  28612=>"110011000",
  28613=>"010011100",
  28614=>"101000111",
  28615=>"011011110",
  28616=>"000000001",
  28617=>"000110101",
  28618=>"100000000",
  28619=>"101111010",
  28620=>"101111100",
  28621=>"010100011",
  28622=>"000000000",
  28623=>"001110011",
  28624=>"101111010",
  28625=>"110000101",
  28626=>"111110101",
  28627=>"100001001",
  28628=>"110000011",
  28629=>"111100111",
  28630=>"100111101",
  28631=>"101010010",
  28632=>"101010110",
  28633=>"111110000",
  28634=>"100010010",
  28635=>"000110010",
  28636=>"000010000",
  28637=>"010101110",
  28638=>"111110111",
  28639=>"011010101",
  28640=>"010101010",
  28641=>"001100000",
  28642=>"010011101",
  28643=>"100101100",
  28644=>"101010100",
  28645=>"111100110",
  28646=>"101101110",
  28647=>"110111010",
  28648=>"101110001",
  28649=>"000110001",
  28650=>"110111000",
  28651=>"110000111",
  28652=>"100010100",
  28653=>"000110101",
  28654=>"110011011",
  28655=>"111111100",
  28656=>"010000110",
  28657=>"011011010",
  28658=>"101010110",
  28659=>"010110101",
  28660=>"000100101",
  28661=>"001010010",
  28662=>"111100000",
  28663=>"011001010",
  28664=>"000011001",
  28665=>"000010010",
  28666=>"011100100",
  28667=>"110101011",
  28668=>"101000110",
  28669=>"011001001",
  28670=>"110000101",
  28671=>"101101110",
  28672=>"101011001",
  28673=>"110100101",
  28674=>"011110000",
  28675=>"011010011",
  28676=>"100111000",
  28677=>"000100101",
  28678=>"010011000",
  28679=>"110001100",
  28680=>"101110111",
  28681=>"101100110",
  28682=>"100011101",
  28683=>"011101110",
  28684=>"111001110",
  28685=>"111101000",
  28686=>"101100101",
  28687=>"111110010",
  28688=>"000101001",
  28689=>"000010111",
  28690=>"110001001",
  28691=>"010111101",
  28692=>"101110111",
  28693=>"011101011",
  28694=>"101101011",
  28695=>"110000001",
  28696=>"000000101",
  28697=>"011101100",
  28698=>"000111100",
  28699=>"001110111",
  28700=>"110111010",
  28701=>"010010010",
  28702=>"111011000",
  28703=>"010110101",
  28704=>"011010110",
  28705=>"000011000",
  28706=>"111011111",
  28707=>"110110001",
  28708=>"101001011",
  28709=>"010011001",
  28710=>"011110100",
  28711=>"110111111",
  28712=>"101000111",
  28713=>"111011011",
  28714=>"000000111",
  28715=>"001000000",
  28716=>"000011001",
  28717=>"000001101",
  28718=>"001000100",
  28719=>"011011011",
  28720=>"101000001",
  28721=>"100101101",
  28722=>"100001110",
  28723=>"001001101",
  28724=>"010100000",
  28725=>"011011010",
  28726=>"001011011",
  28727=>"011010110",
  28728=>"111000010",
  28729=>"111000010",
  28730=>"110000100",
  28731=>"000001010",
  28732=>"001011010",
  28733=>"010110010",
  28734=>"111110100",
  28735=>"010011100",
  28736=>"100110011",
  28737=>"001010111",
  28738=>"011110110",
  28739=>"100000110",
  28740=>"101011001",
  28741=>"100000111",
  28742=>"010100111",
  28743=>"001001011",
  28744=>"010010110",
  28745=>"111001000",
  28746=>"111010000",
  28747=>"010000001",
  28748=>"011000001",
  28749=>"110101111",
  28750=>"010111101",
  28751=>"110111110",
  28752=>"110110010",
  28753=>"110101001",
  28754=>"110111000",
  28755=>"010010101",
  28756=>"110011110",
  28757=>"000110010",
  28758=>"000000110",
  28759=>"001011111",
  28760=>"000100000",
  28761=>"010101011",
  28762=>"100111101",
  28763=>"100011110",
  28764=>"011001101",
  28765=>"010011000",
  28766=>"111111110",
  28767=>"110111110",
  28768=>"010011010",
  28769=>"101110101",
  28770=>"001111111",
  28771=>"100011010",
  28772=>"010111110",
  28773=>"010000010",
  28774=>"001111111",
  28775=>"000110001",
  28776=>"110000010",
  28777=>"111001101",
  28778=>"111101100",
  28779=>"001101100",
  28780=>"011011111",
  28781=>"101101011",
  28782=>"110110010",
  28783=>"011010000",
  28784=>"111110110",
  28785=>"010010010",
  28786=>"101100000",
  28787=>"000100101",
  28788=>"110011000",
  28789=>"101110110",
  28790=>"100111010",
  28791=>"000001011",
  28792=>"000010000",
  28793=>"011110110",
  28794=>"000100011",
  28795=>"000000000",
  28796=>"111111110",
  28797=>"111101110",
  28798=>"000100000",
  28799=>"111010100",
  28800=>"111101100",
  28801=>"010110101",
  28802=>"110110111",
  28803=>"111100000",
  28804=>"000110100",
  28805=>"111111100",
  28806=>"011101000",
  28807=>"011111100",
  28808=>"111010100",
  28809=>"000000010",
  28810=>"000100001",
  28811=>"011011010",
  28812=>"110101000",
  28813=>"010010000",
  28814=>"011111000",
  28815=>"111000101",
  28816=>"111011010",
  28817=>"001000110",
  28818=>"100001100",
  28819=>"101000010",
  28820=>"010010010",
  28821=>"101000000",
  28822=>"011011100",
  28823=>"000010010",
  28824=>"001010011",
  28825=>"001001100",
  28826=>"000101101",
  28827=>"000010100",
  28828=>"000110000",
  28829=>"101011110",
  28830=>"000000011",
  28831=>"111010011",
  28832=>"010010100",
  28833=>"111100101",
  28834=>"010011001",
  28835=>"000100111",
  28836=>"111111110",
  28837=>"101010101",
  28838=>"011001010",
  28839=>"010000001",
  28840=>"100011100",
  28841=>"011001101",
  28842=>"111110110",
  28843=>"011111011",
  28844=>"111011011",
  28845=>"101110000",
  28846=>"011011100",
  28847=>"110000111",
  28848=>"000011011",
  28849=>"000110101",
  28850=>"000110010",
  28851=>"010000000",
  28852=>"010011110",
  28853=>"111111010",
  28854=>"000111011",
  28855=>"000110110",
  28856=>"101001111",
  28857=>"111111111",
  28858=>"110001100",
  28859=>"101011011",
  28860=>"111110010",
  28861=>"011101111",
  28862=>"000100001",
  28863=>"000000110",
  28864=>"101001101",
  28865=>"110100100",
  28866=>"000010010",
  28867=>"011010011",
  28868=>"111101000",
  28869=>"100100000",
  28870=>"001000011",
  28871=>"000011001",
  28872=>"110110010",
  28873=>"010010001",
  28874=>"101101001",
  28875=>"110101100",
  28876=>"000001011",
  28877=>"101100010",
  28878=>"010000000",
  28879=>"011100101",
  28880=>"110010000",
  28881=>"010100001",
  28882=>"011111010",
  28883=>"000100011",
  28884=>"001110011",
  28885=>"011110100",
  28886=>"001111001",
  28887=>"010011011",
  28888=>"110011010",
  28889=>"100101110",
  28890=>"011011011",
  28891=>"010111001",
  28892=>"100010110",
  28893=>"011001001",
  28894=>"100000101",
  28895=>"101100000",
  28896=>"010110000",
  28897=>"011110001",
  28898=>"000011010",
  28899=>"011111110",
  28900=>"100010100",
  28901=>"010101001",
  28902=>"101011100",
  28903=>"101000111",
  28904=>"000000000",
  28905=>"100001000",
  28906=>"111011110",
  28907=>"000100011",
  28908=>"001100000",
  28909=>"100000101",
  28910=>"101000101",
  28911=>"011111110",
  28912=>"010001101",
  28913=>"000100111",
  28914=>"011010011",
  28915=>"010011000",
  28916=>"001101000",
  28917=>"111001011",
  28918=>"011110010",
  28919=>"000000101",
  28920=>"001100100",
  28921=>"000101000",
  28922=>"110110011",
  28923=>"000111011",
  28924=>"100000000",
  28925=>"111110101",
  28926=>"111111011",
  28927=>"000101011",
  28928=>"100100011",
  28929=>"010111001",
  28930=>"011000001",
  28931=>"100010010",
  28932=>"000001001",
  28933=>"011111001",
  28934=>"111101101",
  28935=>"000011001",
  28936=>"010011011",
  28937=>"001110011",
  28938=>"101100010",
  28939=>"101100100",
  28940=>"011010111",
  28941=>"010111110",
  28942=>"001111000",
  28943=>"011001011",
  28944=>"000111010",
  28945=>"001001001",
  28946=>"111111010",
  28947=>"011100000",
  28948=>"101100101",
  28949=>"110010000",
  28950=>"110010010",
  28951=>"010011010",
  28952=>"100001011",
  28953=>"110001111",
  28954=>"100010000",
  28955=>"001001010",
  28956=>"101011011",
  28957=>"000011111",
  28958=>"011011010",
  28959=>"010000100",
  28960=>"111001110",
  28961=>"000101000",
  28962=>"010011101",
  28963=>"100111100",
  28964=>"011000110",
  28965=>"001001011",
  28966=>"001110101",
  28967=>"101110000",
  28968=>"110001000",
  28969=>"100101110",
  28970=>"011000101",
  28971=>"011011001",
  28972=>"010000010",
  28973=>"000110110",
  28974=>"110100101",
  28975=>"010100011",
  28976=>"000001100",
  28977=>"110010110",
  28978=>"001001101",
  28979=>"110011100",
  28980=>"011011011",
  28981=>"010010010",
  28982=>"100111000",
  28983=>"111111010",
  28984=>"010101111",
  28985=>"001010100",
  28986=>"111010101",
  28987=>"000001101",
  28988=>"101000011",
  28989=>"111110011",
  28990=>"011000011",
  28991=>"111111110",
  28992=>"100110011",
  28993=>"001001011",
  28994=>"101011110",
  28995=>"110000100",
  28996=>"110110100",
  28997=>"001001011",
  28998=>"101100011",
  28999=>"010111001",
  29000=>"001001011",
  29001=>"010111011",
  29002=>"111100100",
  29003=>"101101010",
  29004=>"000100011",
  29005=>"110111000",
  29006=>"000110001",
  29007=>"010010110",
  29008=>"101011110",
  29009=>"100100001",
  29010=>"000100000",
  29011=>"110010110",
  29012=>"111100101",
  29013=>"100111010",
  29014=>"010011111",
  29015=>"111100100",
  29016=>"111001100",
  29017=>"001011110",
  29018=>"101001110",
  29019=>"000100000",
  29020=>"011001110",
  29021=>"100011011",
  29022=>"100110011",
  29023=>"000101010",
  29024=>"011010101",
  29025=>"011101101",
  29026=>"000010011",
  29027=>"010010100",
  29028=>"110011111",
  29029=>"000001000",
  29030=>"100110010",
  29031=>"000000101",
  29032=>"001011001",
  29033=>"010110011",
  29034=>"001010100",
  29035=>"101111011",
  29036=>"111111000",
  29037=>"000001111",
  29038=>"100100111",
  29039=>"010010000",
  29040=>"000001001",
  29041=>"001011110",
  29042=>"110111111",
  29043=>"101011100",
  29044=>"001111110",
  29045=>"100011011",
  29046=>"111011000",
  29047=>"001010101",
  29048=>"001101001",
  29049=>"010111011",
  29050=>"100101110",
  29051=>"111111010",
  29052=>"101000111",
  29053=>"111111011",
  29054=>"101000100",
  29055=>"111100011",
  29056=>"111110111",
  29057=>"010000100",
  29058=>"100010010",
  29059=>"010101100",
  29060=>"111111100",
  29061=>"000101001",
  29062=>"001101111",
  29063=>"001100111",
  29064=>"010011001",
  29065=>"111010110",
  29066=>"010101111",
  29067=>"011101111",
  29068=>"001000010",
  29069=>"011000100",
  29070=>"010001011",
  29071=>"100010111",
  29072=>"010110100",
  29073=>"010100111",
  29074=>"110101000",
  29075=>"001111010",
  29076=>"001101011",
  29077=>"000000010",
  29078=>"101000100",
  29079=>"000111001",
  29080=>"000011110",
  29081=>"100000111",
  29082=>"101101100",
  29083=>"011111011",
  29084=>"000000011",
  29085=>"011011110",
  29086=>"111010111",
  29087=>"111000000",
  29088=>"100100001",
  29089=>"000110010",
  29090=>"000010010",
  29091=>"001000001",
  29092=>"110100001",
  29093=>"100110100",
  29094=>"101011011",
  29095=>"000000101",
  29096=>"111100110",
  29097=>"010110011",
  29098=>"001001101",
  29099=>"000000011",
  29100=>"000110000",
  29101=>"111000101",
  29102=>"000000000",
  29103=>"101010110",
  29104=>"001010010",
  29105=>"111101100",
  29106=>"001000000",
  29107=>"100010100",
  29108=>"100001111",
  29109=>"111110101",
  29110=>"111010010",
  29111=>"110010011",
  29112=>"110101101",
  29113=>"011111001",
  29114=>"111000000",
  29115=>"101001100",
  29116=>"011101110",
  29117=>"101100001",
  29118=>"001010001",
  29119=>"001011011",
  29120=>"100101110",
  29121=>"010101001",
  29122=>"111000110",
  29123=>"101100000",
  29124=>"111111000",
  29125=>"010100100",
  29126=>"001000111",
  29127=>"100000101",
  29128=>"011001010",
  29129=>"011111011",
  29130=>"101000101",
  29131=>"000110100",
  29132=>"001111000",
  29133=>"011010101",
  29134=>"011100111",
  29135=>"100100100",
  29136=>"111111100",
  29137=>"000100110",
  29138=>"110111000",
  29139=>"000101010",
  29140=>"000100001",
  29141=>"111100001",
  29142=>"111000000",
  29143=>"101000111",
  29144=>"000101000",
  29145=>"101101001",
  29146=>"010001011",
  29147=>"101111100",
  29148=>"111000110",
  29149=>"111000111",
  29150=>"110011000",
  29151=>"011100111",
  29152=>"001111001",
  29153=>"010000000",
  29154=>"011011101",
  29155=>"111001111",
  29156=>"111001101",
  29157=>"110011101",
  29158=>"000001111",
  29159=>"111000011",
  29160=>"000010100",
  29161=>"101111110",
  29162=>"000011100",
  29163=>"001010000",
  29164=>"101101011",
  29165=>"100011000",
  29166=>"111001000",
  29167=>"011111011",
  29168=>"011011111",
  29169=>"111011111",
  29170=>"011100010",
  29171=>"110011111",
  29172=>"110001000",
  29173=>"001100101",
  29174=>"000110111",
  29175=>"000001010",
  29176=>"011111110",
  29177=>"100010100",
  29178=>"001110010",
  29179=>"001001100",
  29180=>"010111100",
  29181=>"001111101",
  29182=>"101001000",
  29183=>"111011001",
  29184=>"110100111",
  29185=>"100000100",
  29186=>"110100101",
  29187=>"001010011",
  29188=>"101001010",
  29189=>"110101010",
  29190=>"000111111",
  29191=>"010011110",
  29192=>"111110010",
  29193=>"011011110",
  29194=>"001011110",
  29195=>"111101000",
  29196=>"010011111",
  29197=>"111111010",
  29198=>"111001110",
  29199=>"100001010",
  29200=>"111010101",
  29201=>"000100011",
  29202=>"100101001",
  29203=>"100100101",
  29204=>"100000001",
  29205=>"010100000",
  29206=>"101100000",
  29207=>"011011000",
  29208=>"111011010",
  29209=>"101001110",
  29210=>"001010111",
  29211=>"010001101",
  29212=>"110001111",
  29213=>"110111010",
  29214=>"001011010",
  29215=>"011110011",
  29216=>"011000111",
  29217=>"000101100",
  29218=>"000011010",
  29219=>"001010110",
  29220=>"001111001",
  29221=>"010101001",
  29222=>"100111100",
  29223=>"001000101",
  29224=>"010000010",
  29225=>"100001101",
  29226=>"110101111",
  29227=>"011000000",
  29228=>"000001111",
  29229=>"011011010",
  29230=>"101011011",
  29231=>"110000101",
  29232=>"101111011",
  29233=>"100100011",
  29234=>"010110101",
  29235=>"000001000",
  29236=>"000101111",
  29237=>"000000001",
  29238=>"101011100",
  29239=>"111001000",
  29240=>"110100100",
  29241=>"001001001",
  29242=>"101111111",
  29243=>"001001110",
  29244=>"010111111",
  29245=>"110010010",
  29246=>"111000010",
  29247=>"110011001",
  29248=>"001011001",
  29249=>"000010000",
  29250=>"100000000",
  29251=>"011000110",
  29252=>"110010101",
  29253=>"111000000",
  29254=>"011000000",
  29255=>"101111110",
  29256=>"000101100",
  29257=>"101011001",
  29258=>"110010101",
  29259=>"101100101",
  29260=>"011110110",
  29261=>"001011110",
  29262=>"111111111",
  29263=>"110110100",
  29264=>"110110110",
  29265=>"010111101",
  29266=>"111100001",
  29267=>"110100100",
  29268=>"000010001",
  29269=>"111100011",
  29270=>"001010011",
  29271=>"000100011",
  29272=>"000101101",
  29273=>"001111101",
  29274=>"000111000",
  29275=>"000011011",
  29276=>"101010000",
  29277=>"000000000",
  29278=>"011111111",
  29279=>"100111111",
  29280=>"011001100",
  29281=>"011011101",
  29282=>"100010110",
  29283=>"100101111",
  29284=>"101011110",
  29285=>"101001110",
  29286=>"111000110",
  29287=>"011010011",
  29288=>"100000001",
  29289=>"010110101",
  29290=>"011101101",
  29291=>"000111000",
  29292=>"010101011",
  29293=>"100110010",
  29294=>"011110000",
  29295=>"000011101",
  29296=>"011110001",
  29297=>"001110000",
  29298=>"110111110",
  29299=>"000000001",
  29300=>"011011010",
  29301=>"101000101",
  29302=>"111101110",
  29303=>"101101111",
  29304=>"001111000",
  29305=>"011110111",
  29306=>"100000000",
  29307=>"011001111",
  29308=>"011010010",
  29309=>"111001110",
  29310=>"010110010",
  29311=>"001100010",
  29312=>"100101110",
  29313=>"101110100",
  29314=>"110111100",
  29315=>"111100001",
  29316=>"110001111",
  29317=>"001000000",
  29318=>"100111100",
  29319=>"000101001",
  29320=>"100101000",
  29321=>"111101000",
  29322=>"000001010",
  29323=>"111111000",
  29324=>"000000100",
  29325=>"101101111",
  29326=>"111000100",
  29327=>"110100011",
  29328=>"011111110",
  29329=>"001001000",
  29330=>"111100000",
  29331=>"101111101",
  29332=>"111100100",
  29333=>"010001101",
  29334=>"101010111",
  29335=>"000111100",
  29336=>"111010000",
  29337=>"010001010",
  29338=>"011011011",
  29339=>"001001101",
  29340=>"111001101",
  29341=>"011010000",
  29342=>"000100000",
  29343=>"011010110",
  29344=>"001000100",
  29345=>"110100110",
  29346=>"101111110",
  29347=>"011101010",
  29348=>"101101101",
  29349=>"000001000",
  29350=>"000100100",
  29351=>"001110011",
  29352=>"010110010",
  29353=>"001011100",
  29354=>"101011011",
  29355=>"100001001",
  29356=>"110110000",
  29357=>"001111000",
  29358=>"101110000",
  29359=>"011101100",
  29360=>"011001110",
  29361=>"110111110",
  29362=>"111010100",
  29363=>"000000010",
  29364=>"110101001",
  29365=>"110011111",
  29366=>"111000111",
  29367=>"010100100",
  29368=>"110110110",
  29369=>"010101100",
  29370=>"011101010",
  29371=>"000101010",
  29372=>"111001101",
  29373=>"100100100",
  29374=>"101110001",
  29375=>"000011110",
  29376=>"101101101",
  29377=>"101110000",
  29378=>"001111010",
  29379=>"111110101",
  29380=>"011101000",
  29381=>"011000011",
  29382=>"011110111",
  29383=>"111001110",
  29384=>"000110010",
  29385=>"111001110",
  29386=>"101111111",
  29387=>"010001010",
  29388=>"000000000",
  29389=>"010010000",
  29390=>"110010110",
  29391=>"000111101",
  29392=>"100010101",
  29393=>"011101001",
  29394=>"010000101",
  29395=>"000101111",
  29396=>"011110100",
  29397=>"000110100",
  29398=>"010011011",
  29399=>"001101001",
  29400=>"011110010",
  29401=>"011111101",
  29402=>"010110001",
  29403=>"111001101",
  29404=>"110001011",
  29405=>"011010010",
  29406=>"001001101",
  29407=>"101000000",
  29408=>"110100111",
  29409=>"001111111",
  29410=>"011000111",
  29411=>"111110000",
  29412=>"000001101",
  29413=>"110000100",
  29414=>"011100100",
  29415=>"001011001",
  29416=>"100101010",
  29417=>"110111011",
  29418=>"110111001",
  29419=>"101101110",
  29420=>"100110110",
  29421=>"100111110",
  29422=>"011110000",
  29423=>"100010010",
  29424=>"010100100",
  29425=>"011101010",
  29426=>"100111101",
  29427=>"000010101",
  29428=>"111111111",
  29429=>"001110011",
  29430=>"010111000",
  29431=>"111010000",
  29432=>"111110000",
  29433=>"101101100",
  29434=>"010110010",
  29435=>"011110101",
  29436=>"110011000",
  29437=>"110000101",
  29438=>"000100010",
  29439=>"000001110",
  29440=>"010000111",
  29441=>"101101011",
  29442=>"100101110",
  29443=>"111110111",
  29444=>"001001010",
  29445=>"100010011",
  29446=>"001010101",
  29447=>"000011111",
  29448=>"011101001",
  29449=>"110101000",
  29450=>"000001100",
  29451=>"000011010",
  29452=>"001011101",
  29453=>"001101000",
  29454=>"001110100",
  29455=>"010100101",
  29456=>"011110000",
  29457=>"111010101",
  29458=>"000011001",
  29459=>"110011010",
  29460=>"101011010",
  29461=>"011101010",
  29462=>"101101111",
  29463=>"000101001",
  29464=>"111111110",
  29465=>"110011001",
  29466=>"111000100",
  29467=>"011000000",
  29468=>"100010111",
  29469=>"110110110",
  29470=>"001110111",
  29471=>"001111001",
  29472=>"001010001",
  29473=>"111000100",
  29474=>"111101111",
  29475=>"010000110",
  29476=>"111111111",
  29477=>"100001111",
  29478=>"111101101",
  29479=>"110110111",
  29480=>"011111011",
  29481=>"101100000",
  29482=>"001101000",
  29483=>"010010111",
  29484=>"010000011",
  29485=>"001100000",
  29486=>"100011001",
  29487=>"110101101",
  29488=>"010010111",
  29489=>"100001111",
  29490=>"011111111",
  29491=>"000000010",
  29492=>"010010111",
  29493=>"101100101",
  29494=>"011100111",
  29495=>"010110111",
  29496=>"000000011",
  29497=>"110110010",
  29498=>"000011111",
  29499=>"100011101",
  29500=>"101110001",
  29501=>"010011011",
  29502=>"001100011",
  29503=>"001110100",
  29504=>"011001100",
  29505=>"001000000",
  29506=>"111111110",
  29507=>"101000111",
  29508=>"101110011",
  29509=>"010101100",
  29510=>"010010011",
  29511=>"000101010",
  29512=>"101011001",
  29513=>"111101110",
  29514=>"011000010",
  29515=>"100010011",
  29516=>"100000010",
  29517=>"100111110",
  29518=>"001100101",
  29519=>"001100110",
  29520=>"110010010",
  29521=>"011010000",
  29522=>"101000000",
  29523=>"001001001",
  29524=>"111100101",
  29525=>"100101000",
  29526=>"000100111",
  29527=>"001101000",
  29528=>"110001101",
  29529=>"110111001",
  29530=>"010101101",
  29531=>"110101110",
  29532=>"110000110",
  29533=>"111000101",
  29534=>"010001011",
  29535=>"101101111",
  29536=>"111011011",
  29537=>"101110011",
  29538=>"000111000",
  29539=>"001001100",
  29540=>"000110110",
  29541=>"011110011",
  29542=>"101100100",
  29543=>"001100101",
  29544=>"010000110",
  29545=>"110010011",
  29546=>"001110010",
  29547=>"010010110",
  29548=>"110000000",
  29549=>"011101110",
  29550=>"010001100",
  29551=>"000111001",
  29552=>"101110110",
  29553=>"011001110",
  29554=>"111111010",
  29555=>"000111000",
  29556=>"011100111",
  29557=>"101111011",
  29558=>"100000100",
  29559=>"000010011",
  29560=>"101111011",
  29561=>"111010010",
  29562=>"111111011",
  29563=>"010111001",
  29564=>"000001010",
  29565=>"000111111",
  29566=>"111111110",
  29567=>"010111101",
  29568=>"100000001",
  29569=>"101011000",
  29570=>"110110010",
  29571=>"100111010",
  29572=>"000100010",
  29573=>"001111011",
  29574=>"010001000",
  29575=>"101101001",
  29576=>"100110001",
  29577=>"011010001",
  29578=>"001011000",
  29579=>"000111111",
  29580=>"101000111",
  29581=>"101011010",
  29582=>"111000110",
  29583=>"000010010",
  29584=>"010011100",
  29585=>"101001000",
  29586=>"101001111",
  29587=>"010000111",
  29588=>"001000000",
  29589=>"001001101",
  29590=>"100100011",
  29591=>"000000010",
  29592=>"010010001",
  29593=>"110000111",
  29594=>"111010001",
  29595=>"000101111",
  29596=>"011011000",
  29597=>"011110001",
  29598=>"111010000",
  29599=>"010000011",
  29600=>"110001010",
  29601=>"101100101",
  29602=>"111011000",
  29603=>"001001010",
  29604=>"000111111",
  29605=>"001010001",
  29606=>"111010000",
  29607=>"101001000",
  29608=>"110100110",
  29609=>"010111111",
  29610=>"101111001",
  29611=>"001101100",
  29612=>"110001111",
  29613=>"011001101",
  29614=>"111010001",
  29615=>"001100100",
  29616=>"010000100",
  29617=>"110000100",
  29618=>"011111001",
  29619=>"010001001",
  29620=>"000111001",
  29621=>"000110001",
  29622=>"110110101",
  29623=>"100110101",
  29624=>"001101100",
  29625=>"101100001",
  29626=>"100011000",
  29627=>"000000100",
  29628=>"100101001",
  29629=>"000010100",
  29630=>"100001000",
  29631=>"110101001",
  29632=>"101110110",
  29633=>"000001101",
  29634=>"011011000",
  29635=>"010000000",
  29636=>"001100000",
  29637=>"001000001",
  29638=>"110000000",
  29639=>"100011010",
  29640=>"001100000",
  29641=>"111011110",
  29642=>"111011111",
  29643=>"110101111",
  29644=>"111000011",
  29645=>"011000000",
  29646=>"000001000",
  29647=>"010010101",
  29648=>"100101011",
  29649=>"100011000",
  29650=>"001001101",
  29651=>"001100011",
  29652=>"100001110",
  29653=>"011011000",
  29654=>"101111001",
  29655=>"001000111",
  29656=>"011101000",
  29657=>"001011001",
  29658=>"000001010",
  29659=>"001011000",
  29660=>"100010101",
  29661=>"100000010",
  29662=>"010010000",
  29663=>"111110110",
  29664=>"100011100",
  29665=>"100000011",
  29666=>"110011010",
  29667=>"001000101",
  29668=>"100000000",
  29669=>"111100110",
  29670=>"011101010",
  29671=>"011000010",
  29672=>"111110010",
  29673=>"000001110",
  29674=>"000110111",
  29675=>"111110110",
  29676=>"100000010",
  29677=>"000010101",
  29678=>"110000000",
  29679=>"011010010",
  29680=>"100000010",
  29681=>"101100001",
  29682=>"001011001",
  29683=>"010101000",
  29684=>"110011111",
  29685=>"010111100",
  29686=>"001110101",
  29687=>"111111111",
  29688=>"101001111",
  29689=>"101111000",
  29690=>"101000110",
  29691=>"001001110",
  29692=>"011110011",
  29693=>"000011011",
  29694=>"011100111",
  29695=>"100110100",
  29696=>"111110011",
  29697=>"111101100",
  29698=>"010010110",
  29699=>"111101100",
  29700=>"111101001",
  29701=>"011001001",
  29702=>"110001100",
  29703=>"000101110",
  29704=>"000000000",
  29705=>"111111110",
  29706=>"010011111",
  29707=>"101111011",
  29708=>"110010101",
  29709=>"111000111",
  29710=>"001001110",
  29711=>"111000000",
  29712=>"100010100",
  29713=>"110101001",
  29714=>"000000011",
  29715=>"000000000",
  29716=>"101110111",
  29717=>"111001010",
  29718=>"100000010",
  29719=>"111001100",
  29720=>"100001000",
  29721=>"000011001",
  29722=>"110010110",
  29723=>"100000101",
  29724=>"110111100",
  29725=>"011011110",
  29726=>"011011101",
  29727=>"110000110",
  29728=>"011111100",
  29729=>"000010101",
  29730=>"111111001",
  29731=>"001011011",
  29732=>"101111010",
  29733=>"011110100",
  29734=>"100111101",
  29735=>"001111101",
  29736=>"001110011",
  29737=>"110100110",
  29738=>"000100001",
  29739=>"010101001",
  29740=>"100101101",
  29741=>"101001100",
  29742=>"101110101",
  29743=>"111010001",
  29744=>"001000111",
  29745=>"101010101",
  29746=>"110001011",
  29747=>"111011110",
  29748=>"110100000",
  29749=>"001111111",
  29750=>"100001011",
  29751=>"010011100",
  29752=>"101001011",
  29753=>"010010100",
  29754=>"100001111",
  29755=>"101101101",
  29756=>"111111001",
  29757=>"100011001",
  29758=>"101110010",
  29759=>"101100001",
  29760=>"110010111",
  29761=>"010010000",
  29762=>"100101000",
  29763=>"000000001",
  29764=>"001001001",
  29765=>"010101000",
  29766=>"010000011",
  29767=>"100110011",
  29768=>"000101011",
  29769=>"101101100",
  29770=>"010000001",
  29771=>"111000000",
  29772=>"001100010",
  29773=>"110100111",
  29774=>"000000100",
  29775=>"100000010",
  29776=>"010000111",
  29777=>"111101101",
  29778=>"010110000",
  29779=>"101000111",
  29780=>"001101001",
  29781=>"001011001",
  29782=>"111110111",
  29783=>"000100000",
  29784=>"010101101",
  29785=>"110001010",
  29786=>"001100001",
  29787=>"110100010",
  29788=>"001010101",
  29789=>"101101100",
  29790=>"101000000",
  29791=>"010111001",
  29792=>"101001100",
  29793=>"111101110",
  29794=>"110011001",
  29795=>"111110010",
  29796=>"110110110",
  29797=>"111111010",
  29798=>"000001110",
  29799=>"110011110",
  29800=>"101001001",
  29801=>"101011000",
  29802=>"011110101",
  29803=>"010100111",
  29804=>"110011100",
  29805=>"101111110",
  29806=>"101110001",
  29807=>"111111010",
  29808=>"110001100",
  29809=>"110011110",
  29810=>"101011010",
  29811=>"110110011",
  29812=>"110001001",
  29813=>"110010101",
  29814=>"100010111",
  29815=>"100100100",
  29816=>"011111010",
  29817=>"110011001",
  29818=>"011111000",
  29819=>"100010011",
  29820=>"001111111",
  29821=>"001011100",
  29822=>"111111011",
  29823=>"010001011",
  29824=>"010101100",
  29825=>"000110111",
  29826=>"111000101",
  29827=>"110100111",
  29828=>"100100010",
  29829=>"111011101",
  29830=>"000111101",
  29831=>"001111100",
  29832=>"000011001",
  29833=>"111001001",
  29834=>"100000011",
  29835=>"110110110",
  29836=>"110110010",
  29837=>"001010010",
  29838=>"001010111",
  29839=>"111111100",
  29840=>"111011000",
  29841=>"000110010",
  29842=>"011001110",
  29843=>"011111001",
  29844=>"100111111",
  29845=>"100100110",
  29846=>"111001000",
  29847=>"000111000",
  29848=>"100100011",
  29849=>"010011001",
  29850=>"101100001",
  29851=>"000000010",
  29852=>"100010110",
  29853=>"110110110",
  29854=>"110101101",
  29855=>"110001111",
  29856=>"110100110",
  29857=>"111000111",
  29858=>"110010110",
  29859=>"101000101",
  29860=>"011010101",
  29861=>"010000001",
  29862=>"111101001",
  29863=>"110110011",
  29864=>"010100101",
  29865=>"001100010",
  29866=>"100100111",
  29867=>"111101100",
  29868=>"010001000",
  29869=>"001100010",
  29870=>"000000001",
  29871=>"100001110",
  29872=>"110111110",
  29873=>"001100110",
  29874=>"010110001",
  29875=>"110101001",
  29876=>"011011011",
  29877=>"001011111",
  29878=>"011111001",
  29879=>"110001101",
  29880=>"000001100",
  29881=>"111101000",
  29882=>"101100100",
  29883=>"100001011",
  29884=>"101001100",
  29885=>"111100010",
  29886=>"111100001",
  29887=>"110101101",
  29888=>"100111110",
  29889=>"100001101",
  29890=>"001111110",
  29891=>"111101101",
  29892=>"011010010",
  29893=>"010001011",
  29894=>"010100011",
  29895=>"001101111",
  29896=>"101100000",
  29897=>"010101110",
  29898=>"110010010",
  29899=>"001111010",
  29900=>"100000000",
  29901=>"011111111",
  29902=>"100100110",
  29903=>"100110011",
  29904=>"101001110",
  29905=>"101111110",
  29906=>"001111011",
  29907=>"010011011",
  29908=>"111100100",
  29909=>"101101100",
  29910=>"101011100",
  29911=>"001010110",
  29912=>"011001000",
  29913=>"100111000",
  29914=>"101101011",
  29915=>"011110101",
  29916=>"001001111",
  29917=>"100010110",
  29918=>"101001010",
  29919=>"100111011",
  29920=>"011100011",
  29921=>"001011011",
  29922=>"101110011",
  29923=>"101101000",
  29924=>"001010111",
  29925=>"100111111",
  29926=>"000001001",
  29927=>"110111110",
  29928=>"110010101",
  29929=>"110011001",
  29930=>"100101110",
  29931=>"010010011",
  29932=>"110101101",
  29933=>"111000000",
  29934=>"100101110",
  29935=>"001101101",
  29936=>"100011000",
  29937=>"000010001",
  29938=>"001000000",
  29939=>"110111100",
  29940=>"100101000",
  29941=>"110100101",
  29942=>"011111000",
  29943=>"000101100",
  29944=>"111101011",
  29945=>"000100111",
  29946=>"000001011",
  29947=>"010001001",
  29948=>"001100010",
  29949=>"100000101",
  29950=>"101101111",
  29951=>"011111011",
  29952=>"101110000",
  29953=>"000011000",
  29954=>"111001011",
  29955=>"110100100",
  29956=>"111011100",
  29957=>"001010000",
  29958=>"100001100",
  29959=>"110100110",
  29960=>"010011111",
  29961=>"011011101",
  29962=>"010000001",
  29963=>"001000001",
  29964=>"011010101",
  29965=>"111011000",
  29966=>"010010001",
  29967=>"010111001",
  29968=>"001011101",
  29969=>"101111101",
  29970=>"101001100",
  29971=>"111000000",
  29972=>"010111011",
  29973=>"001110001",
  29974=>"110001011",
  29975=>"011001100",
  29976=>"000100101",
  29977=>"110000011",
  29978=>"111110111",
  29979=>"000110111",
  29980=>"010011010",
  29981=>"101000110",
  29982=>"100011111",
  29983=>"111111111",
  29984=>"111100000",
  29985=>"000011100",
  29986=>"101010010",
  29987=>"001001110",
  29988=>"100000010",
  29989=>"101001001",
  29990=>"010001001",
  29991=>"011011010",
  29992=>"001000000",
  29993=>"101110100",
  29994=>"110111011",
  29995=>"011011000",
  29996=>"000101000",
  29997=>"101010010",
  29998=>"010111000",
  29999=>"011001010",
  30000=>"100000000",
  30001=>"110111001",
  30002=>"110001111",
  30003=>"110101010",
  30004=>"011100001",
  30005=>"000010010",
  30006=>"000111010",
  30007=>"110011100",
  30008=>"100101100",
  30009=>"110111011",
  30010=>"110010011",
  30011=>"010111111",
  30012=>"010100110",
  30013=>"111000110",
  30014=>"010111000",
  30015=>"110101110",
  30016=>"001000101",
  30017=>"001000000",
  30018=>"000001110",
  30019=>"011110011",
  30020=>"100010011",
  30021=>"101101011",
  30022=>"001010101",
  30023=>"011110001",
  30024=>"010101100",
  30025=>"001000001",
  30026=>"000000000",
  30027=>"000111011",
  30028=>"001010010",
  30029=>"011000000",
  30030=>"101011001",
  30031=>"010110101",
  30032=>"101001010",
  30033=>"001100001",
  30034=>"010110010",
  30035=>"010010001",
  30036=>"100101111",
  30037=>"100101101",
  30038=>"001000010",
  30039=>"110111111",
  30040=>"001011000",
  30041=>"101001110",
  30042=>"000110001",
  30043=>"101110010",
  30044=>"000101010",
  30045=>"011111111",
  30046=>"111100111",
  30047=>"100011100",
  30048=>"111100110",
  30049=>"001101101",
  30050=>"101100001",
  30051=>"111100101",
  30052=>"010011010",
  30053=>"111111101",
  30054=>"100101000",
  30055=>"010101111",
  30056=>"010001101",
  30057=>"100101100",
  30058=>"100010000",
  30059=>"101101010",
  30060=>"111011100",
  30061=>"100101000",
  30062=>"111101110",
  30063=>"010011001",
  30064=>"110000001",
  30065=>"110001101",
  30066=>"001101111",
  30067=>"111111101",
  30068=>"000100111",
  30069=>"101110000",
  30070=>"000000010",
  30071=>"100000101",
  30072=>"100010001",
  30073=>"010101100",
  30074=>"011010101",
  30075=>"110110001",
  30076=>"000010101",
  30077=>"100101110",
  30078=>"000010010",
  30079=>"110101111",
  30080=>"100110001",
  30081=>"000000110",
  30082=>"111101111",
  30083=>"000001111",
  30084=>"101000010",
  30085=>"101101111",
  30086=>"110101110",
  30087=>"101010001",
  30088=>"010001001",
  30089=>"110000110",
  30090=>"010001001",
  30091=>"111010001",
  30092=>"001001000",
  30093=>"111001011",
  30094=>"110001100",
  30095=>"111100010",
  30096=>"001001000",
  30097=>"111110011",
  30098=>"100000011",
  30099=>"101000010",
  30100=>"011011100",
  30101=>"000001101",
  30102=>"001100001",
  30103=>"000100110",
  30104=>"001010101",
  30105=>"101100010",
  30106=>"001111011",
  30107=>"001010001",
  30108=>"001111000",
  30109=>"100101100",
  30110=>"101110100",
  30111=>"110011111",
  30112=>"110100100",
  30113=>"001100001",
  30114=>"110101000",
  30115=>"000010011",
  30116=>"111101000",
  30117=>"101100101",
  30118=>"001110111",
  30119=>"101110100",
  30120=>"010110000",
  30121=>"001011100",
  30122=>"100110001",
  30123=>"110000011",
  30124=>"000010110",
  30125=>"011111111",
  30126=>"101001100",
  30127=>"111100001",
  30128=>"111101011",
  30129=>"000110100",
  30130=>"100100100",
  30131=>"100110100",
  30132=>"000110010",
  30133=>"011111010",
  30134=>"000100000",
  30135=>"001110110",
  30136=>"011001110",
  30137=>"110101010",
  30138=>"110010010",
  30139=>"001000011",
  30140=>"000000110",
  30141=>"001011100",
  30142=>"000001110",
  30143=>"101000110",
  30144=>"110011100",
  30145=>"100011010",
  30146=>"101001110",
  30147=>"000101001",
  30148=>"000010111",
  30149=>"011010010",
  30150=>"011100111",
  30151=>"011101110",
  30152=>"100101011",
  30153=>"011101111",
  30154=>"101011111",
  30155=>"111110100",
  30156=>"111111101",
  30157=>"011001100",
  30158=>"000111010",
  30159=>"011110110",
  30160=>"010000001",
  30161=>"101111101",
  30162=>"000110001",
  30163=>"000100010",
  30164=>"011000111",
  30165=>"011101101",
  30166=>"100100111",
  30167=>"011001000",
  30168=>"011010100",
  30169=>"110001000",
  30170=>"101001111",
  30171=>"101111111",
  30172=>"111110011",
  30173=>"000010000",
  30174=>"111000111",
  30175=>"001111110",
  30176=>"011000001",
  30177=>"001011000",
  30178=>"000010001",
  30179=>"001000011",
  30180=>"011110100",
  30181=>"110001011",
  30182=>"110010101",
  30183=>"000101001",
  30184=>"100101001",
  30185=>"000010101",
  30186=>"010110101",
  30187=>"111100100",
  30188=>"111001011",
  30189=>"011010000",
  30190=>"101001010",
  30191=>"001110001",
  30192=>"001111000",
  30193=>"101000000",
  30194=>"100011110",
  30195=>"011010001",
  30196=>"110000111",
  30197=>"111011000",
  30198=>"011101100",
  30199=>"110111101",
  30200=>"000100111",
  30201=>"001101000",
  30202=>"010100101",
  30203=>"110001111",
  30204=>"011001010",
  30205=>"100100000",
  30206=>"111111111",
  30207=>"101111011",
  30208=>"110101011",
  30209=>"000010101",
  30210=>"101011011",
  30211=>"110010100",
  30212=>"010110100",
  30213=>"010000111",
  30214=>"001011100",
  30215=>"111001011",
  30216=>"101100110",
  30217=>"111100101",
  30218=>"011101110",
  30219=>"011001101",
  30220=>"001000000",
  30221=>"001011010",
  30222=>"101001100",
  30223=>"110100000",
  30224=>"011001001",
  30225=>"110111111",
  30226=>"011001011",
  30227=>"000000111",
  30228=>"111000000",
  30229=>"011110011",
  30230=>"000001111",
  30231=>"100000011",
  30232=>"111111000",
  30233=>"001001111",
  30234=>"001001011",
  30235=>"111010100",
  30236=>"011001010",
  30237=>"011110100",
  30238=>"101111110",
  30239=>"111101100",
  30240=>"011011011",
  30241=>"001100110",
  30242=>"010000000",
  30243=>"001000110",
  30244=>"111111001",
  30245=>"101000011",
  30246=>"001001001",
  30247=>"000111101",
  30248=>"010000001",
  30249=>"110100011",
  30250=>"110100101",
  30251=>"111000111",
  30252=>"110000000",
  30253=>"000000101",
  30254=>"111111100",
  30255=>"110101011",
  30256=>"000100000",
  30257=>"010111101",
  30258=>"011110111",
  30259=>"011000000",
  30260=>"100100100",
  30261=>"111010110",
  30262=>"011111111",
  30263=>"010000101",
  30264=>"101011001",
  30265=>"101100000",
  30266=>"001001010",
  30267=>"001101101",
  30268=>"011001010",
  30269=>"111001001",
  30270=>"000111011",
  30271=>"101010001",
  30272=>"001010101",
  30273=>"111010000",
  30274=>"100011001",
  30275=>"101101111",
  30276=>"100001011",
  30277=>"111000010",
  30278=>"100010111",
  30279=>"101011100",
  30280=>"001000001",
  30281=>"001010100",
  30282=>"011100001",
  30283=>"011000010",
  30284=>"011011101",
  30285=>"010110111",
  30286=>"011011000",
  30287=>"000110000",
  30288=>"110011011",
  30289=>"110011011",
  30290=>"011000101",
  30291=>"101100001",
  30292=>"010100011",
  30293=>"110100100",
  30294=>"101111111",
  30295=>"000000000",
  30296=>"001101110",
  30297=>"000101001",
  30298=>"010000001",
  30299=>"110110111",
  30300=>"111110001",
  30301=>"111011110",
  30302=>"111000001",
  30303=>"010001001",
  30304=>"111010000",
  30305=>"110001011",
  30306=>"111111110",
  30307=>"100010011",
  30308=>"111111010",
  30309=>"101101110",
  30310=>"010001111",
  30311=>"110100011",
  30312=>"011011000",
  30313=>"111101000",
  30314=>"001101110",
  30315=>"101000110",
  30316=>"100010111",
  30317=>"100101011",
  30318=>"101000010",
  30319=>"001101111",
  30320=>"000111001",
  30321=>"101101010",
  30322=>"010001111",
  30323=>"011100110",
  30324=>"000011100",
  30325=>"110101000",
  30326=>"011001111",
  30327=>"001001000",
  30328=>"101001010",
  30329=>"000000000",
  30330=>"111101001",
  30331=>"100111101",
  30332=>"001000101",
  30333=>"011001001",
  30334=>"000101010",
  30335=>"101101011",
  30336=>"011011001",
  30337=>"101101000",
  30338=>"001000001",
  30339=>"000101001",
  30340=>"001101010",
  30341=>"100011110",
  30342=>"100001101",
  30343=>"000110000",
  30344=>"000101100",
  30345=>"100001001",
  30346=>"000010000",
  30347=>"101000111",
  30348=>"001100000",
  30349=>"111000101",
  30350=>"010010001",
  30351=>"010101100",
  30352=>"100110101",
  30353=>"111101011",
  30354=>"011010011",
  30355=>"001011011",
  30356=>"110111100",
  30357=>"101010110",
  30358=>"101010101",
  30359=>"101010001",
  30360=>"000010010",
  30361=>"000101100",
  30362=>"100011100",
  30363=>"011110100",
  30364=>"001010101",
  30365=>"001110000",
  30366=>"010001010",
  30367=>"011100111",
  30368=>"110000000",
  30369=>"100100000",
  30370=>"001001011",
  30371=>"001001111",
  30372=>"000001010",
  30373=>"000000011",
  30374=>"000001110",
  30375=>"010010111",
  30376=>"110101010",
  30377=>"100010011",
  30378=>"001000100",
  30379=>"011100111",
  30380=>"111000100",
  30381=>"011001101",
  30382=>"000001111",
  30383=>"010001111",
  30384=>"010010100",
  30385=>"111010100",
  30386=>"000101111",
  30387=>"111001111",
  30388=>"101001101",
  30389=>"010100101",
  30390=>"101011101",
  30391=>"011010011",
  30392=>"011111100",
  30393=>"011011011",
  30394=>"001111110",
  30395=>"000101101",
  30396=>"101101100",
  30397=>"101000001",
  30398=>"001101110",
  30399=>"110000001",
  30400=>"110000111",
  30401=>"100101011",
  30402=>"111011011",
  30403=>"001100001",
  30404=>"011011011",
  30405=>"101100101",
  30406=>"101011010",
  30407=>"011011001",
  30408=>"101100100",
  30409=>"010000111",
  30410=>"110100000",
  30411=>"110111100",
  30412=>"100111110",
  30413=>"010000100",
  30414=>"001101101",
  30415=>"011000101",
  30416=>"101000001",
  30417=>"011100000",
  30418=>"111010101",
  30419=>"100110001",
  30420=>"000100000",
  30421=>"111101000",
  30422=>"100110110",
  30423=>"111011101",
  30424=>"101000010",
  30425=>"100100110",
  30426=>"101001000",
  30427=>"101101011",
  30428=>"011001000",
  30429=>"111010000",
  30430=>"100000010",
  30431=>"100000111",
  30432=>"100101101",
  30433=>"101010010",
  30434=>"100010010",
  30435=>"010100000",
  30436=>"100100000",
  30437=>"100010011",
  30438=>"001101000",
  30439=>"000100010",
  30440=>"100100001",
  30441=>"001011011",
  30442=>"011000010",
  30443=>"100111011",
  30444=>"011100011",
  30445=>"101101101",
  30446=>"111000001",
  30447=>"001101001",
  30448=>"010111001",
  30449=>"111111110",
  30450=>"100101011",
  30451=>"101110000",
  30452=>"110110011",
  30453=>"101101011",
  30454=>"011110100",
  30455=>"001110000",
  30456=>"011000100",
  30457=>"010011111",
  30458=>"101111001",
  30459=>"100111101",
  30460=>"110001001",
  30461=>"011111111",
  30462=>"010101101",
  30463=>"011011111",
  30464=>"100100011",
  30465=>"100101100",
  30466=>"100010000",
  30467=>"100110010",
  30468=>"011101111",
  30469=>"111100001",
  30470=>"110110100",
  30471=>"000100000",
  30472=>"100111101",
  30473=>"110001100",
  30474=>"010101011",
  30475=>"111011000",
  30476=>"001100001",
  30477=>"111101011",
  30478=>"001110110",
  30479=>"010101111",
  30480=>"100110010",
  30481=>"001001000",
  30482=>"101011011",
  30483=>"111110111",
  30484=>"001101011",
  30485=>"001100100",
  30486=>"110111101",
  30487=>"101100011",
  30488=>"101101001",
  30489=>"100011000",
  30490=>"100111100",
  30491=>"001100000",
  30492=>"001001001",
  30493=>"000110010",
  30494=>"100100101",
  30495=>"100100111",
  30496=>"101110111",
  30497=>"100110111",
  30498=>"111001111",
  30499=>"110000011",
  30500=>"001111011",
  30501=>"110100000",
  30502=>"110110111",
  30503=>"010111110",
  30504=>"010101001",
  30505=>"000101101",
  30506=>"001100000",
  30507=>"011011011",
  30508=>"011011100",
  30509=>"011101000",
  30510=>"100100111",
  30511=>"000101111",
  30512=>"001011011",
  30513=>"110100011",
  30514=>"100111110",
  30515=>"101000111",
  30516=>"010011000",
  30517=>"110100100",
  30518=>"100010001",
  30519=>"000111100",
  30520=>"111111111",
  30521=>"000000000",
  30522=>"100100101",
  30523=>"100101110",
  30524=>"000010001",
  30525=>"101001001",
  30526=>"000101101",
  30527=>"111101000",
  30528=>"011101001",
  30529=>"010100000",
  30530=>"000010010",
  30531=>"000100010",
  30532=>"100101100",
  30533=>"010011100",
  30534=>"001100001",
  30535=>"100001010",
  30536=>"010011001",
  30537=>"101001100",
  30538=>"010010000",
  30539=>"000011001",
  30540=>"100001000",
  30541=>"100110011",
  30542=>"001000110",
  30543=>"110011100",
  30544=>"000000100",
  30545=>"100000000",
  30546=>"111100010",
  30547=>"101010000",
  30548=>"011101100",
  30549=>"100100010",
  30550=>"010110010",
  30551=>"000000011",
  30552=>"001001111",
  30553=>"110000011",
  30554=>"101011100",
  30555=>"101110100",
  30556=>"011111111",
  30557=>"011011110",
  30558=>"101000101",
  30559=>"101001010",
  30560=>"111111101",
  30561=>"111110111",
  30562=>"110010010",
  30563=>"010011011",
  30564=>"001111110",
  30565=>"100111101",
  30566=>"110010000",
  30567=>"111111010",
  30568=>"110000010",
  30569=>"010100100",
  30570=>"101100011",
  30571=>"011010110",
  30572=>"000001100",
  30573=>"000001000",
  30574=>"100100100",
  30575=>"111010110",
  30576=>"011010111",
  30577=>"010000001",
  30578=>"101011000",
  30579=>"010001101",
  30580=>"000010001",
  30581=>"010110000",
  30582=>"100110000",
  30583=>"110010110",
  30584=>"101101100",
  30585=>"000001000",
  30586=>"100100000",
  30587=>"101100001",
  30588=>"011010000",
  30589=>"011101101",
  30590=>"000000011",
  30591=>"101011111",
  30592=>"101011001",
  30593=>"001101101",
  30594=>"111001001",
  30595=>"100101110",
  30596=>"001101111",
  30597=>"111010001",
  30598=>"000101010",
  30599=>"001101111",
  30600=>"100010100",
  30601=>"100101101",
  30602=>"111100101",
  30603=>"011010111",
  30604=>"110110011",
  30605=>"010000101",
  30606=>"111011000",
  30607=>"000001101",
  30608=>"000010001",
  30609=>"000011111",
  30610=>"110100110",
  30611=>"111111011",
  30612=>"010010010",
  30613=>"000110000",
  30614=>"101010001",
  30615=>"000000001",
  30616=>"010010101",
  30617=>"110100111",
  30618=>"000001001",
  30619=>"110001000",
  30620=>"101010010",
  30621=>"011011110",
  30622=>"101010100",
  30623=>"001100011",
  30624=>"111000010",
  30625=>"010101010",
  30626=>"111000010",
  30627=>"001010101",
  30628=>"000010100",
  30629=>"000010110",
  30630=>"101101001",
  30631=>"101000110",
  30632=>"110000100",
  30633=>"010010010",
  30634=>"000100011",
  30635=>"011000010",
  30636=>"011101101",
  30637=>"111110011",
  30638=>"101100011",
  30639=>"011110101",
  30640=>"000011011",
  30641=>"100010101",
  30642=>"000111001",
  30643=>"000100010",
  30644=>"110101101",
  30645=>"001100100",
  30646=>"111011011",
  30647=>"011010100",
  30648=>"011111010",
  30649=>"110000010",
  30650=>"111111010",
  30651=>"000100011",
  30652=>"100110100",
  30653=>"011000001",
  30654=>"110101010",
  30655=>"000000111",
  30656=>"111010100",
  30657=>"101011011",
  30658=>"100001001",
  30659=>"001100100",
  30660=>"000110000",
  30661=>"100100001",
  30662=>"110111111",
  30663=>"010100111",
  30664=>"110110000",
  30665=>"110011000",
  30666=>"000110100",
  30667=>"100110111",
  30668=>"010100001",
  30669=>"111010111",
  30670=>"101100111",
  30671=>"010110011",
  30672=>"011011110",
  30673=>"001100111",
  30674=>"110111011",
  30675=>"011101001",
  30676=>"001101101",
  30677=>"101011011",
  30678=>"010010011",
  30679=>"101000111",
  30680=>"110000010",
  30681=>"101000010",
  30682=>"011010011",
  30683=>"100001010",
  30684=>"001011100",
  30685=>"001100111",
  30686=>"110001000",
  30687=>"011011101",
  30688=>"101100001",
  30689=>"010111001",
  30690=>"110110100",
  30691=>"101011000",
  30692=>"100000010",
  30693=>"000100110",
  30694=>"010100010",
  30695=>"111101011",
  30696=>"100101101",
  30697=>"011100000",
  30698=>"101101010",
  30699=>"101111001",
  30700=>"101111000",
  30701=>"000100100",
  30702=>"011011000",
  30703=>"100101110",
  30704=>"111110011",
  30705=>"101001111",
  30706=>"010010100",
  30707=>"001111010",
  30708=>"010110111",
  30709=>"001111010",
  30710=>"011101111",
  30711=>"010101110",
  30712=>"101110001",
  30713=>"111110011",
  30714=>"000100100",
  30715=>"110011111",
  30716=>"101011011",
  30717=>"100000111",
  30718=>"011111111",
  30719=>"011100110",
  30720=>"001111101",
  30721=>"011101110",
  30722=>"101011100",
  30723=>"000000011",
  30724=>"110111110",
  30725=>"011101110",
  30726=>"101011011",
  30727=>"111110100",
  30728=>"101101111",
  30729=>"100001101",
  30730=>"011010000",
  30731=>"001111101",
  30732=>"000101101",
  30733=>"011000100",
  30734=>"110101011",
  30735=>"101100001",
  30736=>"100010010",
  30737=>"111101101",
  30738=>"000001010",
  30739=>"111111011",
  30740=>"000110101",
  30741=>"001010000",
  30742=>"000100111",
  30743=>"000001000",
  30744=>"001000001",
  30745=>"000101111",
  30746=>"001111001",
  30747=>"010100101",
  30748=>"110100101",
  30749=>"000001110",
  30750=>"000000011",
  30751=>"001000001",
  30752=>"011000100",
  30753=>"001100000",
  30754=>"010110110",
  30755=>"000000011",
  30756=>"011010011",
  30757=>"011111011",
  30758=>"001111111",
  30759=>"010111110",
  30760=>"101000100",
  30761=>"111110101",
  30762=>"101101001",
  30763=>"011011011",
  30764=>"001000011",
  30765=>"011010010",
  30766=>"010110001",
  30767=>"100111101",
  30768=>"001010010",
  30769=>"001100000",
  30770=>"010001000",
  30771=>"111111100",
  30772=>"011010110",
  30773=>"011001000",
  30774=>"010011110",
  30775=>"111111111",
  30776=>"110000000",
  30777=>"000001111",
  30778=>"100001101",
  30779=>"111011101",
  30780=>"101110101",
  30781=>"110011110",
  30782=>"110000110",
  30783=>"000000110",
  30784=>"000000101",
  30785=>"001110010",
  30786=>"000111111",
  30787=>"010000110",
  30788=>"000100101",
  30789=>"111000010",
  30790=>"100110000",
  30791=>"001000101",
  30792=>"011110100",
  30793=>"001111111",
  30794=>"111101111",
  30795=>"111001100",
  30796=>"101101110",
  30797=>"000000010",
  30798=>"100101100",
  30799=>"011011110",
  30800=>"011100010",
  30801=>"000100000",
  30802=>"111000101",
  30803=>"110100100",
  30804=>"101010000",
  30805=>"100000100",
  30806=>"010100000",
  30807=>"110001111",
  30808=>"110010110",
  30809=>"110010111",
  30810=>"010110001",
  30811=>"110110101",
  30812=>"011010001",
  30813=>"111011010",
  30814=>"000001101",
  30815=>"110101011",
  30816=>"101000000",
  30817=>"011000001",
  30818=>"110110110",
  30819=>"011011100",
  30820=>"000110000",
  30821=>"011101010",
  30822=>"010000000",
  30823=>"101111010",
  30824=>"001110011",
  30825=>"100010000",
  30826=>"111011100",
  30827=>"101010101",
  30828=>"001100111",
  30829=>"100000000",
  30830=>"110111000",
  30831=>"011101111",
  30832=>"000101101",
  30833=>"111001111",
  30834=>"000000101",
  30835=>"111111111",
  30836=>"101001011",
  30837=>"101101111",
  30838=>"011011101",
  30839=>"100111010",
  30840=>"111011001",
  30841=>"100010111",
  30842=>"101001010",
  30843=>"010000010",
  30844=>"110110011",
  30845=>"111011111",
  30846=>"101100011",
  30847=>"010000101",
  30848=>"001011100",
  30849=>"110010101",
  30850=>"110000110",
  30851=>"000001011",
  30852=>"101001001",
  30853=>"111001111",
  30854=>"100110000",
  30855=>"001100100",
  30856=>"111001001",
  30857=>"000001000",
  30858=>"101100101",
  30859=>"101010001",
  30860=>"100011101",
  30861=>"001100101",
  30862=>"111010011",
  30863=>"110110101",
  30864=>"011100111",
  30865=>"100101111",
  30866=>"000000010",
  30867=>"100111100",
  30868=>"000110101",
  30869=>"110101010",
  30870=>"000000111",
  30871=>"110010010",
  30872=>"011110101",
  30873=>"001110110",
  30874=>"000001001",
  30875=>"110010101",
  30876=>"000010011",
  30877=>"000110010",
  30878=>"001101001",
  30879=>"010001001",
  30880=>"100010001",
  30881=>"111011010",
  30882=>"110110010",
  30883=>"111100100",
  30884=>"011101100",
  30885=>"000100100",
  30886=>"110011101",
  30887=>"011010011",
  30888=>"100001010",
  30889=>"111110111",
  30890=>"111001001",
  30891=>"110111011",
  30892=>"001110000",
  30893=>"111111101",
  30894=>"000101110",
  30895=>"010010100",
  30896=>"011000001",
  30897=>"101000000",
  30898=>"010101101",
  30899=>"000000101",
  30900=>"110001111",
  30901=>"001001111",
  30902=>"010110011",
  30903=>"011001001",
  30904=>"100000011",
  30905=>"011100100",
  30906=>"000100000",
  30907=>"111110000",
  30908=>"000001010",
  30909=>"010011001",
  30910=>"010010100",
  30911=>"110110100",
  30912=>"000011101",
  30913=>"010100010",
  30914=>"111100100",
  30915=>"010001111",
  30916=>"111111111",
  30917=>"001000110",
  30918=>"101111000",
  30919=>"001000011",
  30920=>"010110101",
  30921=>"100010011",
  30922=>"001000000",
  30923=>"010001111",
  30924=>"010110011",
  30925=>"001000011",
  30926=>"111111001",
  30927=>"100101110",
  30928=>"100100111",
  30929=>"111010110",
  30930=>"111010110",
  30931=>"100001101",
  30932=>"101011100",
  30933=>"010011001",
  30934=>"100011001",
  30935=>"100100110",
  30936=>"000000010",
  30937=>"000001001",
  30938=>"010000100",
  30939=>"101000011",
  30940=>"101001101",
  30941=>"010111000",
  30942=>"001101100",
  30943=>"011110111",
  30944=>"000001000",
  30945=>"111010110",
  30946=>"100100101",
  30947=>"010100011",
  30948=>"111010000",
  30949=>"000111110",
  30950=>"000110001",
  30951=>"101001111",
  30952=>"110001010",
  30953=>"101100001",
  30954=>"000001011",
  30955=>"111010111",
  30956=>"000110111",
  30957=>"010001001",
  30958=>"100100110",
  30959=>"000110000",
  30960=>"001001111",
  30961=>"011000101",
  30962=>"011000000",
  30963=>"001011010",
  30964=>"111110001",
  30965=>"011101110",
  30966=>"000010100",
  30967=>"000001110",
  30968=>"001010100",
  30969=>"100100011",
  30970=>"000000000",
  30971=>"000000000",
  30972=>"000001101",
  30973=>"101101110",
  30974=>"001101010",
  30975=>"111001110",
  30976=>"010010101",
  30977=>"101010100",
  30978=>"110010111",
  30979=>"111111000",
  30980=>"010011110",
  30981=>"100100000",
  30982=>"100011010",
  30983=>"011001101",
  30984=>"001000000",
  30985=>"010001111",
  30986=>"111101101",
  30987=>"001000110",
  30988=>"110000111",
  30989=>"111010000",
  30990=>"101011010",
  30991=>"001001111",
  30992=>"011010001",
  30993=>"000100110",
  30994=>"101110111",
  30995=>"101101010",
  30996=>"101001101",
  30997=>"010000000",
  30998=>"100010001",
  30999=>"110101011",
  31000=>"001011001",
  31001=>"000110001",
  31002=>"010000100",
  31003=>"010101100",
  31004=>"000011001",
  31005=>"100111111",
  31006=>"001101101",
  31007=>"100100010",
  31008=>"001110000",
  31009=>"010000010",
  31010=>"011101000",
  31011=>"011110010",
  31012=>"000100110",
  31013=>"010010110",
  31014=>"101111101",
  31015=>"001011101",
  31016=>"100000000",
  31017=>"001101001",
  31018=>"000101100",
  31019=>"011111100",
  31020=>"111100101",
  31021=>"000000101",
  31022=>"011101010",
  31023=>"011110011",
  31024=>"000100001",
  31025=>"100101001",
  31026=>"011010100",
  31027=>"011000000",
  31028=>"001001010",
  31029=>"001011111",
  31030=>"001001001",
  31031=>"100011010",
  31032=>"000000000",
  31033=>"010101010",
  31034=>"010001010",
  31035=>"110101110",
  31036=>"010101011",
  31037=>"000100000",
  31038=>"110000110",
  31039=>"000111101",
  31040=>"011001010",
  31041=>"001111100",
  31042=>"011100110",
  31043=>"110000000",
  31044=>"001111111",
  31045=>"101011000",
  31046=>"000011001",
  31047=>"111010111",
  31048=>"110010101",
  31049=>"100110100",
  31050=>"101010011",
  31051=>"011001001",
  31052=>"101010101",
  31053=>"011000101",
  31054=>"001111101",
  31055=>"000010001",
  31056=>"001101100",
  31057=>"101111101",
  31058=>"011000000",
  31059=>"010010011",
  31060=>"101110011",
  31061=>"001111111",
  31062=>"110101000",
  31063=>"111001001",
  31064=>"000110000",
  31065=>"000100100",
  31066=>"101100000",
  31067=>"000111100",
  31068=>"011110100",
  31069=>"111011010",
  31070=>"000101000",
  31071=>"110001011",
  31072=>"010111001",
  31073=>"101111100",
  31074=>"100101100",
  31075=>"100001111",
  31076=>"101011000",
  31077=>"000110010",
  31078=>"011000010",
  31079=>"001110101",
  31080=>"110110011",
  31081=>"111010101",
  31082=>"011011011",
  31083=>"110101011",
  31084=>"000101001",
  31085=>"011010000",
  31086=>"101010010",
  31087=>"011100110",
  31088=>"100000000",
  31089=>"100011100",
  31090=>"000111000",
  31091=>"100100001",
  31092=>"010100100",
  31093=>"100111100",
  31094=>"111100000",
  31095=>"001011100",
  31096=>"001111100",
  31097=>"101100101",
  31098=>"001110011",
  31099=>"100010100",
  31100=>"101010010",
  31101=>"111111101",
  31102=>"001100000",
  31103=>"101001100",
  31104=>"100011111",
  31105=>"011101000",
  31106=>"100001111",
  31107=>"011100101",
  31108=>"100000110",
  31109=>"100001100",
  31110=>"011100100",
  31111=>"000010101",
  31112=>"001100011",
  31113=>"111001100",
  31114=>"000100101",
  31115=>"000010011",
  31116=>"110111010",
  31117=>"000010000",
  31118=>"010011111",
  31119=>"011100110",
  31120=>"101100101",
  31121=>"101001111",
  31122=>"000100000",
  31123=>"110010000",
  31124=>"000001000",
  31125=>"100100010",
  31126=>"011111110",
  31127=>"011001001",
  31128=>"101001011",
  31129=>"101001110",
  31130=>"100011000",
  31131=>"000001110",
  31132=>"010000110",
  31133=>"000101001",
  31134=>"100011110",
  31135=>"001101000",
  31136=>"011101101",
  31137=>"101000100",
  31138=>"100101110",
  31139=>"001100001",
  31140=>"000111101",
  31141=>"110001001",
  31142=>"111001011",
  31143=>"100101110",
  31144=>"000001000",
  31145=>"010110110",
  31146=>"010000000",
  31147=>"010001001",
  31148=>"000111101",
  31149=>"110000001",
  31150=>"111101101",
  31151=>"000011000",
  31152=>"010111101",
  31153=>"010100110",
  31154=>"110000101",
  31155=>"001111111",
  31156=>"101100010",
  31157=>"010100010",
  31158=>"001001111",
  31159=>"101010110",
  31160=>"110001100",
  31161=>"101000011",
  31162=>"011001001",
  31163=>"000010101",
  31164=>"111110111",
  31165=>"001010101",
  31166=>"000000110",
  31167=>"010100000",
  31168=>"110101000",
  31169=>"100111000",
  31170=>"010001010",
  31171=>"111001010",
  31172=>"101111111",
  31173=>"111101011",
  31174=>"111010111",
  31175=>"000000000",
  31176=>"011001111",
  31177=>"110010011",
  31178=>"000000101",
  31179=>"011010011",
  31180=>"110100111",
  31181=>"111011110",
  31182=>"101000100",
  31183=>"000101011",
  31184=>"100100010",
  31185=>"011111100",
  31186=>"100000001",
  31187=>"100101001",
  31188=>"100101101",
  31189=>"011111110",
  31190=>"010111010",
  31191=>"100110111",
  31192=>"110001011",
  31193=>"011011010",
  31194=>"011011001",
  31195=>"001011001",
  31196=>"101001101",
  31197=>"010011011",
  31198=>"010001010",
  31199=>"110101010",
  31200=>"000010100",
  31201=>"010000111",
  31202=>"010110000",
  31203=>"011010100",
  31204=>"010000000",
  31205=>"010101111",
  31206=>"100010111",
  31207=>"001001001",
  31208=>"111001001",
  31209=>"011100000",
  31210=>"011110100",
  31211=>"111111000",
  31212=>"001011010",
  31213=>"000110111",
  31214=>"011101110",
  31215=>"001111000",
  31216=>"111101010",
  31217=>"000011010",
  31218=>"100010011",
  31219=>"110111111",
  31220=>"001101111",
  31221=>"010000110",
  31222=>"110110111",
  31223=>"100111001",
  31224=>"010100101",
  31225=>"011111100",
  31226=>"101100011",
  31227=>"100110101",
  31228=>"001111110",
  31229=>"011101001",
  31230=>"101111001",
  31231=>"011100111",
  31232=>"101000010",
  31233=>"001000110",
  31234=>"100001010",
  31235=>"001001110",
  31236=>"001110110",
  31237=>"111111001",
  31238=>"000111100",
  31239=>"001000011",
  31240=>"101000011",
  31241=>"001100001",
  31242=>"010100010",
  31243=>"000001101",
  31244=>"101101000",
  31245=>"110110000",
  31246=>"010111001",
  31247=>"110110101",
  31248=>"001100011",
  31249=>"000110111",
  31250=>"011111111",
  31251=>"011110010",
  31252=>"011100111",
  31253=>"011111010",
  31254=>"010111001",
  31255=>"110110110",
  31256=>"110111001",
  31257=>"110011111",
  31258=>"000110111",
  31259=>"010000101",
  31260=>"100011101",
  31261=>"111001101",
  31262=>"100001110",
  31263=>"101111111",
  31264=>"100101100",
  31265=>"001011010",
  31266=>"001101111",
  31267=>"100011111",
  31268=>"110000100",
  31269=>"111100100",
  31270=>"000001000",
  31271=>"101010111",
  31272=>"010010010",
  31273=>"000011100",
  31274=>"001110011",
  31275=>"111111111",
  31276=>"100001111",
  31277=>"101100111",
  31278=>"101100010",
  31279=>"010100110",
  31280=>"000000001",
  31281=>"010011001",
  31282=>"000110101",
  31283=>"011110111",
  31284=>"101011000",
  31285=>"001010011",
  31286=>"010011100",
  31287=>"010110101",
  31288=>"111000110",
  31289=>"011000101",
  31290=>"010101111",
  31291=>"000000001",
  31292=>"001000101",
  31293=>"011011001",
  31294=>"011110000",
  31295=>"111110000",
  31296=>"100000000",
  31297=>"110010000",
  31298=>"000101111",
  31299=>"101111000",
  31300=>"101001000",
  31301=>"111111101",
  31302=>"110000000",
  31303=>"001001100",
  31304=>"110010010",
  31305=>"101000101",
  31306=>"110111101",
  31307=>"001010001",
  31308=>"001000110",
  31309=>"011010010",
  31310=>"011101111",
  31311=>"100011100",
  31312=>"101000110",
  31313=>"010110011",
  31314=>"110000100",
  31315=>"100100101",
  31316=>"100110100",
  31317=>"111110000",
  31318=>"010010010",
  31319=>"101101101",
  31320=>"111111101",
  31321=>"111110010",
  31322=>"101101010",
  31323=>"101000000",
  31324=>"011110001",
  31325=>"000111001",
  31326=>"000101110",
  31327=>"000000001",
  31328=>"000101011",
  31329=>"000101010",
  31330=>"110010000",
  31331=>"100001001",
  31332=>"101001101",
  31333=>"001000000",
  31334=>"100001010",
  31335=>"011001100",
  31336=>"000010110",
  31337=>"000101101",
  31338=>"111110111",
  31339=>"111111110",
  31340=>"100010111",
  31341=>"000011100",
  31342=>"000011101",
  31343=>"011111110",
  31344=>"111111100",
  31345=>"000000000",
  31346=>"111000110",
  31347=>"001000010",
  31348=>"100011000",
  31349=>"111111001",
  31350=>"010000011",
  31351=>"100011101",
  31352=>"001110000",
  31353=>"011110101",
  31354=>"000100100",
  31355=>"010111101",
  31356=>"110001111",
  31357=>"110001010",
  31358=>"000110111",
  31359=>"101001001",
  31360=>"011111101",
  31361=>"100101010",
  31362=>"010101101",
  31363=>"100000101",
  31364=>"101010000",
  31365=>"000011101",
  31366=>"000010001",
  31367=>"101111110",
  31368=>"101000000",
  31369=>"111110000",
  31370=>"000100100",
  31371=>"011000000",
  31372=>"011000010",
  31373=>"010101111",
  31374=>"010011100",
  31375=>"101001011",
  31376=>"011110100",
  31377=>"100101101",
  31378=>"111011100",
  31379=>"001010000",
  31380=>"101000011",
  31381=>"011111011",
  31382=>"011000000",
  31383=>"100101111",
  31384=>"011100110",
  31385=>"010110111",
  31386=>"011000000",
  31387=>"111011111",
  31388=>"001000110",
  31389=>"111010100",
  31390=>"000010011",
  31391=>"111101111",
  31392=>"001100000",
  31393=>"000100011",
  31394=>"111011101",
  31395=>"111001010",
  31396=>"100110101",
  31397=>"010000001",
  31398=>"110111001",
  31399=>"000011111",
  31400=>"000111111",
  31401=>"100110110",
  31402=>"010001100",
  31403=>"100001000",
  31404=>"010100100",
  31405=>"001001111",
  31406=>"100111110",
  31407=>"111111110",
  31408=>"011011101",
  31409=>"000000101",
  31410=>"001110100",
  31411=>"001100010",
  31412=>"001011001",
  31413=>"100010010",
  31414=>"000111001",
  31415=>"100111101",
  31416=>"011001011",
  31417=>"110100001",
  31418=>"111101101",
  31419=>"110111011",
  31420=>"000111110",
  31421=>"110011000",
  31422=>"000101111",
  31423=>"010010100",
  31424=>"000010101",
  31425=>"111111101",
  31426=>"110001101",
  31427=>"001111101",
  31428=>"000011000",
  31429=>"010110001",
  31430=>"110000000",
  31431=>"001001000",
  31432=>"110110010",
  31433=>"010110101",
  31434=>"011100001",
  31435=>"101001010",
  31436=>"100010001",
  31437=>"000011001",
  31438=>"010100101",
  31439=>"110111010",
  31440=>"101011000",
  31441=>"010000011",
  31442=>"110000111",
  31443=>"000001100",
  31444=>"000010000",
  31445=>"101100110",
  31446=>"100100001",
  31447=>"110100111",
  31448=>"000100111",
  31449=>"011110000",
  31450=>"000000111",
  31451=>"110110110",
  31452=>"100100111",
  31453=>"110111101",
  31454=>"111100000",
  31455=>"010011100",
  31456=>"101000010",
  31457=>"000100110",
  31458=>"011001110",
  31459=>"101010100",
  31460=>"010101101",
  31461=>"111111101",
  31462=>"010000011",
  31463=>"001111110",
  31464=>"000101001",
  31465=>"011111100",
  31466=>"111110110",
  31467=>"100100001",
  31468=>"000100101",
  31469=>"100101111",
  31470=>"100001001",
  31471=>"001010011",
  31472=>"001011111",
  31473=>"100011000",
  31474=>"100001000",
  31475=>"111010111",
  31476=>"100011101",
  31477=>"000011100",
  31478=>"000100000",
  31479=>"001100010",
  31480=>"111010001",
  31481=>"100111001",
  31482=>"100110101",
  31483=>"000110000",
  31484=>"001001010",
  31485=>"001011000",
  31486=>"101101011",
  31487=>"011000111",
  31488=>"010110111",
  31489=>"100010101",
  31490=>"101010011",
  31491=>"000001001",
  31492=>"101101001",
  31493=>"101000101",
  31494=>"000111010",
  31495=>"101100000",
  31496=>"111000111",
  31497=>"101100001",
  31498=>"101000111",
  31499=>"000101111",
  31500=>"100010011",
  31501=>"001000100",
  31502=>"000100100",
  31503=>"001001111",
  31504=>"110101101",
  31505=>"111100111",
  31506=>"001110001",
  31507=>"010110100",
  31508=>"010110100",
  31509=>"000111101",
  31510=>"100110001",
  31511=>"000000101",
  31512=>"000001001",
  31513=>"000101000",
  31514=>"101001010",
  31515=>"111100110",
  31516=>"111010111",
  31517=>"110000111",
  31518=>"100000101",
  31519=>"110011110",
  31520=>"110000001",
  31521=>"010011110",
  31522=>"000100011",
  31523=>"111000000",
  31524=>"110101010",
  31525=>"000011110",
  31526=>"110110101",
  31527=>"101111011",
  31528=>"110101011",
  31529=>"111111000",
  31530=>"011111101",
  31531=>"000000010",
  31532=>"011111010",
  31533=>"000000111",
  31534=>"001111011",
  31535=>"011101111",
  31536=>"010001111",
  31537=>"001101000",
  31538=>"110100100",
  31539=>"011101100",
  31540=>"111011110",
  31541=>"111010000",
  31542=>"101100111",
  31543=>"001000100",
  31544=>"111111010",
  31545=>"000101111",
  31546=>"101010101",
  31547=>"001011100",
  31548=>"011101001",
  31549=>"011000101",
  31550=>"000000010",
  31551=>"111000011",
  31552=>"001100101",
  31553=>"101100011",
  31554=>"010010000",
  31555=>"000000101",
  31556=>"111111101",
  31557=>"100011100",
  31558=>"000011101",
  31559=>"011110110",
  31560=>"101010100",
  31561=>"000101111",
  31562=>"010101011",
  31563=>"110110110",
  31564=>"100110011",
  31565=>"000000000",
  31566=>"010001010",
  31567=>"101011111",
  31568=>"111111010",
  31569=>"010001101",
  31570=>"011110110",
  31571=>"011011101",
  31572=>"000000111",
  31573=>"010101001",
  31574=>"111010001",
  31575=>"111101110",
  31576=>"110101101",
  31577=>"111101011",
  31578=>"111111010",
  31579=>"000001010",
  31580=>"110101100",
  31581=>"111101101",
  31582=>"000111101",
  31583=>"001100011",
  31584=>"011011100",
  31585=>"111101111",
  31586=>"101110000",
  31587=>"010011010",
  31588=>"110111110",
  31589=>"101010010",
  31590=>"001100101",
  31591=>"011000000",
  31592=>"101110100",
  31593=>"100110100",
  31594=>"111100011",
  31595=>"101111001",
  31596=>"001111010",
  31597=>"100011100",
  31598=>"110010100",
  31599=>"111001010",
  31600=>"010101111",
  31601=>"100000101",
  31602=>"001010000",
  31603=>"110110010",
  31604=>"111010100",
  31605=>"100011001",
  31606=>"110011000",
  31607=>"101101101",
  31608=>"100111011",
  31609=>"111100110",
  31610=>"010101101",
  31611=>"010100110",
  31612=>"101111110",
  31613=>"001001011",
  31614=>"001100101",
  31615=>"011001101",
  31616=>"100100001",
  31617=>"001101100",
  31618=>"000000111",
  31619=>"111001010",
  31620=>"100101000",
  31621=>"001111110",
  31622=>"101000010",
  31623=>"100101110",
  31624=>"011111001",
  31625=>"010001110",
  31626=>"011110110",
  31627=>"100100010",
  31628=>"001011110",
  31629=>"111111000",
  31630=>"111100010",
  31631=>"100010100",
  31632=>"010010001",
  31633=>"101011000",
  31634=>"011110000",
  31635=>"101001110",
  31636=>"110111010",
  31637=>"000001000",
  31638=>"111011100",
  31639=>"011011110",
  31640=>"111101000",
  31641=>"011000111",
  31642=>"101101100",
  31643=>"001011011",
  31644=>"010111010",
  31645=>"111111111",
  31646=>"010110100",
  31647=>"000110101",
  31648=>"100100101",
  31649=>"100111011",
  31650=>"101110001",
  31651=>"001000000",
  31652=>"111011010",
  31653=>"011111101",
  31654=>"001000011",
  31655=>"001111000",
  31656=>"100011010",
  31657=>"101111111",
  31658=>"011110101",
  31659=>"111000010",
  31660=>"011110001",
  31661=>"101100100",
  31662=>"011010011",
  31663=>"110111101",
  31664=>"101111000",
  31665=>"100011111",
  31666=>"110001001",
  31667=>"011100000",
  31668=>"001001010",
  31669=>"001101100",
  31670=>"101000001",
  31671=>"011010111",
  31672=>"000101000",
  31673=>"111110111",
  31674=>"111110000",
  31675=>"001011010",
  31676=>"001001000",
  31677=>"011111011",
  31678=>"010111100",
  31679=>"111010000",
  31680=>"110010111",
  31681=>"111111110",
  31682=>"000100110",
  31683=>"000001101",
  31684=>"110000001",
  31685=>"010000101",
  31686=>"110111001",
  31687=>"010110001",
  31688=>"001000111",
  31689=>"111111110",
  31690=>"000010100",
  31691=>"111010111",
  31692=>"000100001",
  31693=>"101000111",
  31694=>"011010110",
  31695=>"010101101",
  31696=>"110100111",
  31697=>"111101001",
  31698=>"101101100",
  31699=>"110011000",
  31700=>"111011011",
  31701=>"110100011",
  31702=>"010000000",
  31703=>"011101011",
  31704=>"011101101",
  31705=>"111111100",
  31706=>"001011001",
  31707=>"010010110",
  31708=>"011000010",
  31709=>"010011101",
  31710=>"010110001",
  31711=>"011000000",
  31712=>"111010101",
  31713=>"011011010",
  31714=>"000000101",
  31715=>"100000100",
  31716=>"110100101",
  31717=>"000001000",
  31718=>"101110001",
  31719=>"001111101",
  31720=>"100101111",
  31721=>"100000110",
  31722=>"011101101",
  31723=>"110110110",
  31724=>"111001101",
  31725=>"001010101",
  31726=>"101011011",
  31727=>"111110100",
  31728=>"101000011",
  31729=>"100101001",
  31730=>"110001100",
  31731=>"110100111",
  31732=>"100111000",
  31733=>"111000100",
  31734=>"111110001",
  31735=>"000001110",
  31736=>"100110011",
  31737=>"111001100",
  31738=>"001000100",
  31739=>"001100001",
  31740=>"000110000",
  31741=>"010100001",
  31742=>"011001001",
  31743=>"000001111",
  31744=>"100000000",
  31745=>"110110001",
  31746=>"110000101",
  31747=>"000001111",
  31748=>"100000110",
  31749=>"001010010",
  31750=>"101010111",
  31751=>"110110111",
  31752=>"110000101",
  31753=>"101010101",
  31754=>"001010101",
  31755=>"111011011",
  31756=>"110101111",
  31757=>"101001011",
  31758=>"011001000",
  31759=>"110111010",
  31760=>"101110101",
  31761=>"000111010",
  31762=>"010010100",
  31763=>"100100110",
  31764=>"100001100",
  31765=>"100100110",
  31766=>"001000111",
  31767=>"100000100",
  31768=>"001111010",
  31769=>"000111001",
  31770=>"110000110",
  31771=>"000011011",
  31772=>"010011011",
  31773=>"101011000",
  31774=>"001000110",
  31775=>"111011100",
  31776=>"101000110",
  31777=>"100010001",
  31778=>"000110000",
  31779=>"110000011",
  31780=>"010010101",
  31781=>"001011101",
  31782=>"001101100",
  31783=>"110010100",
  31784=>"010110100",
  31785=>"000100000",
  31786=>"010101011",
  31787=>"011010110",
  31788=>"100000110",
  31789=>"101111111",
  31790=>"011000001",
  31791=>"010100011",
  31792=>"110101111",
  31793=>"001101111",
  31794=>"000110011",
  31795=>"111000111",
  31796=>"110111011",
  31797=>"001001100",
  31798=>"110001101",
  31799=>"000110000",
  31800=>"101110101",
  31801=>"010101111",
  31802=>"000011101",
  31803=>"100010010",
  31804=>"010000101",
  31805=>"100011011",
  31806=>"100000110",
  31807=>"111101011",
  31808=>"000010010",
  31809=>"000011000",
  31810=>"111101001",
  31811=>"000001000",
  31812=>"100010000",
  31813=>"110111000",
  31814=>"001000011",
  31815=>"001110110",
  31816=>"001111110",
  31817=>"101001100",
  31818=>"111010001",
  31819=>"010100110",
  31820=>"001001000",
  31821=>"101110100",
  31822=>"111100000",
  31823=>"010000011",
  31824=>"010100000",
  31825=>"000110000",
  31826=>"000100110",
  31827=>"011000001",
  31828=>"000010111",
  31829=>"011100010",
  31830=>"010110110",
  31831=>"001111100",
  31832=>"011000011",
  31833=>"111101001",
  31834=>"000110110",
  31835=>"010110010",
  31836=>"000100111",
  31837=>"000000100",
  31838=>"111011001",
  31839=>"110011011",
  31840=>"000000000",
  31841=>"100010111",
  31842=>"000101001",
  31843=>"001011111",
  31844=>"100000000",
  31845=>"101111111",
  31846=>"100000010",
  31847=>"100101011",
  31848=>"000111001",
  31849=>"110100111",
  31850=>"010111110",
  31851=>"000000010",
  31852=>"011010111",
  31853=>"111010100",
  31854=>"101101000",
  31855=>"111011111",
  31856=>"110011101",
  31857=>"000011001",
  31858=>"111011111",
  31859=>"101011110",
  31860=>"010010110",
  31861=>"100110101",
  31862=>"111110110",
  31863=>"000001111",
  31864=>"000000110",
  31865=>"000010111",
  31866=>"011011010",
  31867=>"001000101",
  31868=>"011100100",
  31869=>"001001101",
  31870=>"011010001",
  31871=>"101000111",
  31872=>"011001000",
  31873=>"000000000",
  31874=>"001001011",
  31875=>"001011011",
  31876=>"000000001",
  31877=>"011000111",
  31878=>"000001100",
  31879=>"101001110",
  31880=>"001001100",
  31881=>"011000100",
  31882=>"000011000",
  31883=>"111101110",
  31884=>"100110001",
  31885=>"111110000",
  31886=>"010000111",
  31887=>"111011011",
  31888=>"001111000",
  31889=>"111101011",
  31890=>"010110111",
  31891=>"111111101",
  31892=>"111011011",
  31893=>"101110101",
  31894=>"101010101",
  31895=>"000000111",
  31896=>"110001110",
  31897=>"000101110",
  31898=>"100010101",
  31899=>"001001010",
  31900=>"101100101",
  31901=>"110000110",
  31902=>"001000000",
  31903=>"111110011",
  31904=>"110010001",
  31905=>"100001010",
  31906=>"000110000",
  31907=>"110110000",
  31908=>"111011101",
  31909=>"111011011",
  31910=>"000010001",
  31911=>"100111001",
  31912=>"011010110",
  31913=>"101001011",
  31914=>"010010111",
  31915=>"100001101",
  31916=>"001010000",
  31917=>"100110100",
  31918=>"011000000",
  31919=>"001001011",
  31920=>"011011100",
  31921=>"000100000",
  31922=>"100001111",
  31923=>"111101100",
  31924=>"001011101",
  31925=>"010001000",
  31926=>"110100100",
  31927=>"010001000",
  31928=>"000001111",
  31929=>"000001110",
  31930=>"100110110",
  31931=>"011010001",
  31932=>"111111001",
  31933=>"111101011",
  31934=>"010101000",
  31935=>"011110001",
  31936=>"101000101",
  31937=>"000110100",
  31938=>"001001100",
  31939=>"100101100",
  31940=>"010001010",
  31941=>"110101001",
  31942=>"110011101",
  31943=>"001000100",
  31944=>"111100010",
  31945=>"011110000",
  31946=>"110000000",
  31947=>"110011010",
  31948=>"111101011",
  31949=>"000111010",
  31950=>"001000111",
  31951=>"110010111",
  31952=>"111001010",
  31953=>"010111001",
  31954=>"000101111",
  31955=>"000111000",
  31956=>"011001010",
  31957=>"000010000",
  31958=>"000100000",
  31959=>"110010100",
  31960=>"101110001",
  31961=>"011000011",
  31962=>"100000000",
  31963=>"111100100",
  31964=>"100000000",
  31965=>"010010010",
  31966=>"101110101",
  31967=>"110111001",
  31968=>"101110000",
  31969=>"011110101",
  31970=>"010110011",
  31971=>"011100000",
  31972=>"110111100",
  31973=>"001001000",
  31974=>"000011111",
  31975=>"010011001",
  31976=>"001110001",
  31977=>"111110011",
  31978=>"110110011",
  31979=>"001000010",
  31980=>"001110001",
  31981=>"000000111",
  31982=>"110010011",
  31983=>"011101010",
  31984=>"001010110",
  31985=>"110101011",
  31986=>"100010101",
  31987=>"110100110",
  31988=>"000101101",
  31989=>"111000100",
  31990=>"011111000",
  31991=>"101010110",
  31992=>"001001011",
  31993=>"101110101",
  31994=>"011001010",
  31995=>"001100111",
  31996=>"010101100",
  31997=>"010010101",
  31998=>"000101110",
  31999=>"000110100",
  32000=>"101110010",
  32001=>"000110011",
  32002=>"101011101",
  32003=>"111011110",
  32004=>"001010000",
  32005=>"101000011",
  32006=>"000010010",
  32007=>"011010011",
  32008=>"001101111",
  32009=>"000111100",
  32010=>"010010000",
  32011=>"100011011",
  32012=>"000001101",
  32013=>"000101001",
  32014=>"001110001",
  32015=>"000011110",
  32016=>"111001111",
  32017=>"101010010",
  32018=>"000000111",
  32019=>"111001111",
  32020=>"101111001",
  32021=>"000110100",
  32022=>"000101100",
  32023=>"001100010",
  32024=>"111010100",
  32025=>"100001101",
  32026=>"111100100",
  32027=>"011001100",
  32028=>"101101011",
  32029=>"101110011",
  32030=>"110111111",
  32031=>"011110010",
  32032=>"110000000",
  32033=>"111111001",
  32034=>"111111100",
  32035=>"101010000",
  32036=>"111100101",
  32037=>"001000001",
  32038=>"000000000",
  32039=>"111110111",
  32040=>"001010011",
  32041=>"110001110",
  32042=>"100110001",
  32043=>"110100011",
  32044=>"011101011",
  32045=>"000000100",
  32046=>"011111000",
  32047=>"000110001",
  32048=>"101100001",
  32049=>"001001000",
  32050=>"101100111",
  32051=>"100000111",
  32052=>"000100011",
  32053=>"011110110",
  32054=>"100111101",
  32055=>"101101101",
  32056=>"101101001",
  32057=>"110010100",
  32058=>"010010101",
  32059=>"101110001",
  32060=>"111111110",
  32061=>"010001000",
  32062=>"001111001",
  32063=>"000110111",
  32064=>"011110001",
  32065=>"110110111",
  32066=>"000010011",
  32067=>"011011111",
  32068=>"110111011",
  32069=>"111100101",
  32070=>"111100000",
  32071=>"111011100",
  32072=>"011011100",
  32073=>"110110000",
  32074=>"000100110",
  32075=>"110000101",
  32076=>"110100101",
  32077=>"000001100",
  32078=>"000001101",
  32079=>"001011110",
  32080=>"111110010",
  32081=>"110101100",
  32082=>"101100111",
  32083=>"000111000",
  32084=>"100100000",
  32085=>"101011000",
  32086=>"011000001",
  32087=>"000111000",
  32088=>"010100010",
  32089=>"011111111",
  32090=>"101110111",
  32091=>"110011000",
  32092=>"111110000",
  32093=>"110101111",
  32094=>"000011001",
  32095=>"000001001",
  32096=>"110001111",
  32097=>"001011001",
  32098=>"011011001",
  32099=>"001010011",
  32100=>"100101111",
  32101=>"001000000",
  32102=>"110010000",
  32103=>"100101010",
  32104=>"101011010",
  32105=>"000100010",
  32106=>"010000000",
  32107=>"111101011",
  32108=>"000011011",
  32109=>"111111111",
  32110=>"000000111",
  32111=>"001000110",
  32112=>"000000101",
  32113=>"111000100",
  32114=>"010100101",
  32115=>"110100100",
  32116=>"001010101",
  32117=>"111000111",
  32118=>"000110011",
  32119=>"011011111",
  32120=>"111110111",
  32121=>"010110000",
  32122=>"111011101",
  32123=>"010000100",
  32124=>"111110101",
  32125=>"111100100",
  32126=>"000010001",
  32127=>"000100111",
  32128=>"000011110",
  32129=>"011101101",
  32130=>"111111110",
  32131=>"001010010",
  32132=>"010101010",
  32133=>"100011001",
  32134=>"101110110",
  32135=>"001001001",
  32136=>"001111100",
  32137=>"101010011",
  32138=>"011010001",
  32139=>"111101000",
  32140=>"100010010",
  32141=>"000101101",
  32142=>"100010011",
  32143=>"111010001",
  32144=>"101001101",
  32145=>"000000001",
  32146=>"010000010",
  32147=>"100101011",
  32148=>"111100011",
  32149=>"000001001",
  32150=>"110100011",
  32151=>"110011101",
  32152=>"010110110",
  32153=>"001100001",
  32154=>"001111110",
  32155=>"111000011",
  32156=>"001101100",
  32157=>"000011110",
  32158=>"010100010",
  32159=>"111010110",
  32160=>"000101000",
  32161=>"100011100",
  32162=>"010101011",
  32163=>"000010111",
  32164=>"110010101",
  32165=>"001100011",
  32166=>"100000110",
  32167=>"110100110",
  32168=>"101111001",
  32169=>"111001000",
  32170=>"001111001",
  32171=>"101101011",
  32172=>"000110000",
  32173=>"000000101",
  32174=>"110011101",
  32175=>"001010001",
  32176=>"000100011",
  32177=>"001000000",
  32178=>"010101011",
  32179=>"101110111",
  32180=>"111111010",
  32181=>"000000100",
  32182=>"000100001",
  32183=>"100101000",
  32184=>"110010100",
  32185=>"100110010",
  32186=>"001011100",
  32187=>"011110110",
  32188=>"100010111",
  32189=>"111001000",
  32190=>"111001111",
  32191=>"110110011",
  32192=>"001000111",
  32193=>"110010110",
  32194=>"100111110",
  32195=>"010001110",
  32196=>"011000000",
  32197=>"111000101",
  32198=>"001111100",
  32199=>"100110111",
  32200=>"100011101",
  32201=>"101110110",
  32202=>"010100110",
  32203=>"100100110",
  32204=>"000101101",
  32205=>"011000111",
  32206=>"011110101",
  32207=>"010011111",
  32208=>"111111001",
  32209=>"011111011",
  32210=>"111011111",
  32211=>"011010011",
  32212=>"111101110",
  32213=>"001010001",
  32214=>"111101001",
  32215=>"001001011",
  32216=>"111101101",
  32217=>"000001100",
  32218=>"100011101",
  32219=>"101100010",
  32220=>"111010110",
  32221=>"011111111",
  32222=>"001001111",
  32223=>"111010100",
  32224=>"010000001",
  32225=>"111100000",
  32226=>"000111001",
  32227=>"001101011",
  32228=>"011011000",
  32229=>"011011000",
  32230=>"001100000",
  32231=>"100111101",
  32232=>"000101010",
  32233=>"111010001",
  32234=>"000000000",
  32235=>"111111110",
  32236=>"011001011",
  32237=>"010011010",
  32238=>"100100000",
  32239=>"110011001",
  32240=>"000011011",
  32241=>"010101111",
  32242=>"100100001",
  32243=>"100011000",
  32244=>"011011111",
  32245=>"011101001",
  32246=>"000000000",
  32247=>"100111110",
  32248=>"100010110",
  32249=>"111001000",
  32250=>"000101000",
  32251=>"000001001",
  32252=>"000010100",
  32253=>"110100000",
  32254=>"011111000",
  32255=>"101100110",
  32256=>"001010001",
  32257=>"001010000",
  32258=>"000000011",
  32259=>"100101000",
  32260=>"101100110",
  32261=>"011010001",
  32262=>"110000101",
  32263=>"111100000",
  32264=>"111101101",
  32265=>"010111000",
  32266=>"111000011",
  32267=>"001001000",
  32268=>"001111000",
  32269=>"010100001",
  32270=>"111000000",
  32271=>"101001111",
  32272=>"001010100",
  32273=>"100010001",
  32274=>"101100011",
  32275=>"111000010",
  32276=>"010100010",
  32277=>"000001010",
  32278=>"110111100",
  32279=>"000001000",
  32280=>"100111001",
  32281=>"010010011",
  32282=>"011101010",
  32283=>"100011111",
  32284=>"110011101",
  32285=>"000110000",
  32286=>"011010011",
  32287=>"011000000",
  32288=>"111001110",
  32289=>"000001001",
  32290=>"010000000",
  32291=>"000000111",
  32292=>"010010100",
  32293=>"100000100",
  32294=>"101110001",
  32295=>"011000110",
  32296=>"000110001",
  32297=>"111000000",
  32298=>"000000111",
  32299=>"000010000",
  32300=>"010101100",
  32301=>"000000110",
  32302=>"101000000",
  32303=>"100111011",
  32304=>"100110011",
  32305=>"011001010",
  32306=>"101100100",
  32307=>"101100100",
  32308=>"101100000",
  32309=>"010000110",
  32310=>"011001111",
  32311=>"001000000",
  32312=>"001000111",
  32313=>"010100000",
  32314=>"000001110",
  32315=>"110001010",
  32316=>"111010100",
  32317=>"110111011",
  32318=>"111110110",
  32319=>"110110010",
  32320=>"001000000",
  32321=>"111101000",
  32322=>"101011011",
  32323=>"100010100",
  32324=>"111100111",
  32325=>"011111011",
  32326=>"100100101",
  32327=>"011110111",
  32328=>"100111011",
  32329=>"101111011",
  32330=>"101100011",
  32331=>"000101011",
  32332=>"001101001",
  32333=>"100001001",
  32334=>"101101000",
  32335=>"001101000",
  32336=>"000100111",
  32337=>"101101011",
  32338=>"001001100",
  32339=>"100001100",
  32340=>"100010001",
  32341=>"000111110",
  32342=>"110110011",
  32343=>"110110100",
  32344=>"001110001",
  32345=>"001011010",
  32346=>"100101100",
  32347=>"110111101",
  32348=>"001101011",
  32349=>"000000111",
  32350=>"111101001",
  32351=>"111000001",
  32352=>"000101100",
  32353=>"000101001",
  32354=>"100011011",
  32355=>"111001110",
  32356=>"111111001",
  32357=>"101100110",
  32358=>"000001010",
  32359=>"000100011",
  32360=>"010111100",
  32361=>"110100111",
  32362=>"111011101",
  32363=>"011101110",
  32364=>"011111101",
  32365=>"101110011",
  32366=>"000010101",
  32367=>"100101010",
  32368=>"001001100",
  32369=>"111101011",
  32370=>"110100001",
  32371=>"111011110",
  32372=>"001111000",
  32373=>"001010010",
  32374=>"010010110",
  32375=>"111111000",
  32376=>"110111111",
  32377=>"001100010",
  32378=>"000011011",
  32379=>"110011111",
  32380=>"001001010",
  32381=>"100000000",
  32382=>"000111010",
  32383=>"001110101",
  32384=>"111001011",
  32385=>"110001101",
  32386=>"000000101",
  32387=>"010101011",
  32388=>"000100110",
  32389=>"100011010",
  32390=>"110010111",
  32391=>"111100001",
  32392=>"000100000",
  32393=>"000100000",
  32394=>"101001101",
  32395=>"000000000",
  32396=>"001110110",
  32397=>"001011111",
  32398=>"111000101",
  32399=>"001000010",
  32400=>"011111011",
  32401=>"010000010",
  32402=>"001101101",
  32403=>"101111101",
  32404=>"000110011",
  32405=>"010110000",
  32406=>"101111100",
  32407=>"011011100",
  32408=>"110101010",
  32409=>"110010111",
  32410=>"110000001",
  32411=>"110110100",
  32412=>"001111001",
  32413=>"011000010",
  32414=>"110100010",
  32415=>"011001001",
  32416=>"001000111",
  32417=>"000011111",
  32418=>"101111101",
  32419=>"011111110",
  32420=>"011111011",
  32421=>"000100101",
  32422=>"010110100",
  32423=>"001000101",
  32424=>"001001000",
  32425=>"101101100",
  32426=>"011001111",
  32427=>"011100101",
  32428=>"011001000",
  32429=>"011110101",
  32430=>"011001000",
  32431=>"111111000",
  32432=>"000111001",
  32433=>"010011001",
  32434=>"111110011",
  32435=>"101110001",
  32436=>"010100011",
  32437=>"010111100",
  32438=>"010111010",
  32439=>"111010000",
  32440=>"000100101",
  32441=>"000110011",
  32442=>"001011000",
  32443=>"011101111",
  32444=>"000110010",
  32445=>"001001011",
  32446=>"100011110",
  32447=>"010111011",
  32448=>"101011101",
  32449=>"100101111",
  32450=>"101000000",
  32451=>"010101010",
  32452=>"010110000",
  32453=>"001100000",
  32454=>"110010110",
  32455=>"000011010",
  32456=>"111011010",
  32457=>"000101001",
  32458=>"000001100",
  32459=>"011111100",
  32460=>"100110010",
  32461=>"001100001",
  32462=>"010000110",
  32463=>"000011000",
  32464=>"001010100",
  32465=>"010000100",
  32466=>"100110100",
  32467=>"000001011",
  32468=>"110100011",
  32469=>"101010110",
  32470=>"100110000",
  32471=>"011111010",
  32472=>"111010011",
  32473=>"111000100",
  32474=>"111110101",
  32475=>"101010110",
  32476=>"100111011",
  32477=>"000000000",
  32478=>"000111111",
  32479=>"010010001",
  32480=>"111001010",
  32481=>"010100011",
  32482=>"111010000",
  32483=>"010010101",
  32484=>"100110001",
  32485=>"000011101",
  32486=>"011011101",
  32487=>"111110111",
  32488=>"010101000",
  32489=>"011101101",
  32490=>"111111101",
  32491=>"110110101",
  32492=>"001010110",
  32493=>"110000001",
  32494=>"110001101",
  32495=>"011001111",
  32496=>"001010100",
  32497=>"100101000",
  32498=>"101100101",
  32499=>"110010100",
  32500=>"111110010",
  32501=>"011110001",
  32502=>"111011000",
  32503=>"101010010",
  32504=>"010001010",
  32505=>"110101001",
  32506=>"010110111",
  32507=>"011111111",
  32508=>"010100100",
  32509=>"111100111",
  32510=>"010110101",
  32511=>"010100001",
  32512=>"000111010",
  32513=>"110011100",
  32514=>"101111000",
  32515=>"100010111",
  32516=>"010001100",
  32517=>"010110111",
  32518=>"011100010",
  32519=>"101011010",
  32520=>"000110110",
  32521=>"001001010",
  32522=>"001110110",
  32523=>"011110001",
  32524=>"000001010",
  32525=>"111001111",
  32526=>"000010000",
  32527=>"101111010",
  32528=>"011011110",
  32529=>"111000100",
  32530=>"001111001",
  32531=>"110111111",
  32532=>"010010000",
  32533=>"101101011",
  32534=>"100111100",
  32535=>"100001010",
  32536=>"001101101",
  32537=>"000000001",
  32538=>"110000011",
  32539=>"100010100",
  32540=>"001101000",
  32541=>"110010011",
  32542=>"010010011",
  32543=>"110010101",
  32544=>"000010111",
  32545=>"100011011",
  32546=>"100010110",
  32547=>"110101010",
  32548=>"000100101",
  32549=>"001001100",
  32550=>"100100010",
  32551=>"001000010",
  32552=>"111111001",
  32553=>"011111110",
  32554=>"000100111",
  32555=>"101010111",
  32556=>"111011111",
  32557=>"111101111",
  32558=>"000110010",
  32559=>"011100110",
  32560=>"000001101",
  32561=>"101000011",
  32562=>"011100001",
  32563=>"110000000",
  32564=>"001110001",
  32565=>"010110100",
  32566=>"000000011",
  32567=>"000101101",
  32568=>"111010010",
  32569=>"101000001",
  32570=>"001111011",
  32571=>"101001101",
  32572=>"010101011",
  32573=>"000100101",
  32574=>"011100100",
  32575=>"010111101",
  32576=>"111110111",
  32577=>"100100010",
  32578=>"111111001",
  32579=>"000101011",
  32580=>"000001011",
  32581=>"101010101",
  32582=>"111101110",
  32583=>"000011111",
  32584=>"001111101",
  32585=>"110101011",
  32586=>"001011101",
  32587=>"010101011",
  32588=>"001100101",
  32589=>"111110000",
  32590=>"010110110",
  32591=>"001111000",
  32592=>"100110100",
  32593=>"001010110",
  32594=>"001001001",
  32595=>"111110110",
  32596=>"101100110",
  32597=>"000000000",
  32598=>"000100000",
  32599=>"111110010",
  32600=>"010111010",
  32601=>"100011001",
  32602=>"011000101",
  32603=>"001100011",
  32604=>"101011111",
  32605=>"000010011",
  32606=>"111110010",
  32607=>"001010001",
  32608=>"111100001",
  32609=>"000101011",
  32610=>"010111111",
  32611=>"011011011",
  32612=>"000101001",
  32613=>"000000011",
  32614=>"100100010",
  32615=>"111100101",
  32616=>"001011101",
  32617=>"011110000",
  32618=>"111111011",
  32619=>"011111101",
  32620=>"010100101",
  32621=>"001100111",
  32622=>"000010000",
  32623=>"100100110",
  32624=>"000100001",
  32625=>"111101100",
  32626=>"001001001",
  32627=>"001101011",
  32628=>"101101111",
  32629=>"110011101",
  32630=>"111110000",
  32631=>"010101010",
  32632=>"011010010",
  32633=>"010001011",
  32634=>"001001000",
  32635=>"010111010",
  32636=>"000001010",
  32637=>"000000111",
  32638=>"010010101",
  32639=>"111010110",
  32640=>"001110110",
  32641=>"110101011",
  32642=>"001000100",
  32643=>"010011000",
  32644=>"001100010",
  32645=>"110011010",
  32646=>"001111001",
  32647=>"001111100",
  32648=>"101001110",
  32649=>"010100101",
  32650=>"100011111",
  32651=>"101010100",
  32652=>"111111010",
  32653=>"101000001",
  32654=>"101111001",
  32655=>"000001000",
  32656=>"100010010",
  32657=>"111011101",
  32658=>"000111000",
  32659=>"001100111",
  32660=>"011111111",
  32661=>"011110101",
  32662=>"001100000",
  32663=>"101101000",
  32664=>"110010011",
  32665=>"000010110",
  32666=>"001101000",
  32667=>"110110000",
  32668=>"011101000",
  32669=>"001100100",
  32670=>"111100000",
  32671=>"110111111",
  32672=>"001100101",
  32673=>"011111111",
  32674=>"001111110",
  32675=>"111000001",
  32676=>"000010100",
  32677=>"011111100",
  32678=>"101110110",
  32679=>"111001111",
  32680=>"111000101",
  32681=>"100000101",
  32682=>"011011001",
  32683=>"000100110",
  32684=>"110110010",
  32685=>"000010111",
  32686=>"001010001",
  32687=>"000110111",
  32688=>"111000111",
  32689=>"101100101",
  32690=>"111010101",
  32691=>"101101000",
  32692=>"001010110",
  32693=>"100111101",
  32694=>"010010000",
  32695=>"011001001",
  32696=>"000000010",
  32697=>"001111000",
  32698=>"011111101",
  32699=>"000001001",
  32700=>"101100001",
  32701=>"100010111",
  32702=>"111010111",
  32703=>"001000101",
  32704=>"101100000",
  32705=>"001010010",
  32706=>"000110111",
  32707=>"011100101",
  32708=>"100110111",
  32709=>"001000001",
  32710=>"101001010",
  32711=>"101001001",
  32712=>"010000000",
  32713=>"000000100",
  32714=>"110001101",
  32715=>"110000111",
  32716=>"010001001",
  32717=>"000111011",
  32718=>"110000011",
  32719=>"100100100",
  32720=>"111011010",
  32721=>"110101010",
  32722=>"101111100",
  32723=>"101000000",
  32724=>"110001000",
  32725=>"100111101",
  32726=>"001100001",
  32727=>"110100111",
  32728=>"110110011",
  32729=>"100000101",
  32730=>"110101000",
  32731=>"011111100",
  32732=>"001011100",
  32733=>"110111001",
  32734=>"000111111",
  32735=>"010000100",
  32736=>"110110010",
  32737=>"101110100",
  32738=>"100101111",
  32739=>"100001111",
  32740=>"010111111",
  32741=>"001001000",
  32742=>"001000000",
  32743=>"010100111",
  32744=>"000011001",
  32745=>"001001010",
  32746=>"111110011",
  32747=>"000011001",
  32748=>"100100000",
  32749=>"010001101",
  32750=>"010011111",
  32751=>"111110110",
  32752=>"011101011",
  32753=>"101110000",
  32754=>"111111001",
  32755=>"010100000",
  32756=>"100101010",
  32757=>"011110100",
  32758=>"010111000",
  32759=>"010000110",
  32760=>"100010110",
  32761=>"000011101",
  32762=>"110111100",
  32763=>"000000110",
  32764=>"001010001",
  32765=>"010011011",
  32766=>"101100111",
  32767=>"011010010",
  32768=>"000010011",
  32769=>"010111101",
  32770=>"101101011",
  32771=>"111100101",
  32772=>"010010101",
  32773=>"000000010",
  32774=>"001111011",
  32775=>"111010101",
  32776=>"010101101",
  32777=>"010011100",
  32778=>"110111100",
  32779=>"110101111",
  32780=>"010011001",
  32781=>"001111101",
  32782=>"011111101",
  32783=>"101110011",
  32784=>"011101110",
  32785=>"100010000",
  32786=>"000000111",
  32787=>"111011101",
  32788=>"110111001",
  32789=>"100111001",
  32790=>"110010101",
  32791=>"110000000",
  32792=>"000001101",
  32793=>"001011010",
  32794=>"110100100",
  32795=>"010001110",
  32796=>"100001010",
  32797=>"100010000",
  32798=>"101110010",
  32799=>"011101111",
  32800=>"010100011",
  32801=>"001111000",
  32802=>"011111101",
  32803=>"100001000",
  32804=>"011010111",
  32805=>"111101101",
  32806=>"001110101",
  32807=>"100101101",
  32808=>"010100111",
  32809=>"000110101",
  32810=>"101100100",
  32811=>"100001101",
  32812=>"000100000",
  32813=>"001011010",
  32814=>"110100100",
  32815=>"111011011",
  32816=>"111111111",
  32817=>"110101001",
  32818=>"001011001",
  32819=>"000000010",
  32820=>"111111011",
  32821=>"111110000",
  32822=>"100111110",
  32823=>"101111111",
  32824=>"111010100",
  32825=>"001111100",
  32826=>"001011011",
  32827=>"001000100",
  32828=>"101000000",
  32829=>"001110001",
  32830=>"011010101",
  32831=>"100011011",
  32832=>"110011000",
  32833=>"010100100",
  32834=>"100001110",
  32835=>"011000001",
  32836=>"100101001",
  32837=>"010010010",
  32838=>"000001001",
  32839=>"010000001",
  32840=>"100110110",
  32841=>"100001010",
  32842=>"010101001",
  32843=>"000000011",
  32844=>"101100010",
  32845=>"000000000",
  32846=>"001010000",
  32847=>"110011000",
  32848=>"000010011",
  32849=>"000010010",
  32850=>"001111100",
  32851=>"000110101",
  32852=>"001010001",
  32853=>"101001100",
  32854=>"111100000",
  32855=>"010000001",
  32856=>"000000111",
  32857=>"100011100",
  32858=>"110110110",
  32859=>"110101101",
  32860=>"000010010",
  32861=>"001000011",
  32862=>"000110100",
  32863=>"000000011",
  32864=>"110010100",
  32865=>"010100010",
  32866=>"000111000",
  32867=>"101101001",
  32868=>"001101101",
  32869=>"001010110",
  32870=>"110111111",
  32871=>"001010111",
  32872=>"110101000",
  32873=>"000011001",
  32874=>"100001101",
  32875=>"011101011",
  32876=>"100000011",
  32877=>"111010001",
  32878=>"011001000",
  32879=>"100100111",
  32880=>"101111001",
  32881=>"110101000",
  32882=>"100100011",
  32883=>"010000000",
  32884=>"010111101",
  32885=>"100100000",
  32886=>"101001011",
  32887=>"001100100",
  32888=>"100101111",
  32889=>"000110010",
  32890=>"000110011",
  32891=>"101110000",
  32892=>"100100101",
  32893=>"101000001",
  32894=>"100001000",
  32895=>"011111111",
  32896=>"100101100",
  32897=>"000001010",
  32898=>"001010000",
  32899=>"000101001",
  32900=>"100101000",
  32901=>"110010101",
  32902=>"011011111",
  32903=>"011011111",
  32904=>"111010110",
  32905=>"110111001",
  32906=>"110010000",
  32907=>"111001011",
  32908=>"000100110",
  32909=>"110001011",
  32910=>"001100111",
  32911=>"001001111",
  32912=>"111100001",
  32913=>"001111100",
  32914=>"011000100",
  32915=>"110100011",
  32916=>"111110011",
  32917=>"010001000",
  32918=>"000110001",
  32919=>"010100101",
  32920=>"001010010",
  32921=>"011000001",
  32922=>"100000001",
  32923=>"101110011",
  32924=>"010010101",
  32925=>"111100111",
  32926=>"111000011",
  32927=>"010101111",
  32928=>"101100000",
  32929=>"011000001",
  32930=>"111111010",
  32931=>"111110001",
  32932=>"111001100",
  32933=>"000011100",
  32934=>"001001010",
  32935=>"010100110",
  32936=>"100000011",
  32937=>"100011101",
  32938=>"101011110",
  32939=>"111111010",
  32940=>"110111110",
  32941=>"010001001",
  32942=>"110100000",
  32943=>"001101110",
  32944=>"100101010",
  32945=>"111010010",
  32946=>"100011011",
  32947=>"110001011",
  32948=>"111101011",
  32949=>"010011011",
  32950=>"111100110",
  32951=>"001011000",
  32952=>"100001110",
  32953=>"111010111",
  32954=>"100010000",
  32955=>"101001000",
  32956=>"111100010",
  32957=>"100000000",
  32958=>"100101001",
  32959=>"011001100",
  32960=>"111101010",
  32961=>"100111010",
  32962=>"101000011",
  32963=>"010000001",
  32964=>"001011010",
  32965=>"010111001",
  32966=>"111110010",
  32967=>"010010100",
  32968=>"110000011",
  32969=>"101100001",
  32970=>"111101111",
  32971=>"011100100",
  32972=>"100101000",
  32973=>"100011000",
  32974=>"100000010",
  32975=>"011111010",
  32976=>"101010001",
  32977=>"000000111",
  32978=>"010000100",
  32979=>"001101001",
  32980=>"000000111",
  32981=>"110010100",
  32982=>"001010000",
  32983=>"011011000",
  32984=>"110010110",
  32985=>"110010101",
  32986=>"110100001",
  32987=>"000111000",
  32988=>"000101001",
  32989=>"000001011",
  32990=>"100100100",
  32991=>"100111101",
  32992=>"111011110",
  32993=>"000010010",
  32994=>"001111110",
  32995=>"000001101",
  32996=>"110010000",
  32997=>"000111101",
  32998=>"000001111",
  32999=>"111000000",
  33000=>"010111010",
  33001=>"101101111",
  33002=>"010100101",
  33003=>"000011011",
  33004=>"110011001",
  33005=>"110000110",
  33006=>"101011101",
  33007=>"000100001",
  33008=>"101101011",
  33009=>"001101100",
  33010=>"010101101",
  33011=>"101100100",
  33012=>"101110001",
  33013=>"111001011",
  33014=>"010100101",
  33015=>"011001111",
  33016=>"001011111",
  33017=>"111111010",
  33018=>"010110001",
  33019=>"111101101",
  33020=>"101001111",
  33021=>"000001001",
  33022=>"011110011",
  33023=>"110001111",
  33024=>"101101100",
  33025=>"110011001",
  33026=>"101101101",
  33027=>"100111001",
  33028=>"101011100",
  33029=>"100000011",
  33030=>"110001010",
  33031=>"111111000",
  33032=>"111101110",
  33033=>"001011010",
  33034=>"010110011",
  33035=>"101001001",
  33036=>"001011101",
  33037=>"110111101",
  33038=>"100101110",
  33039=>"001010011",
  33040=>"110001111",
  33041=>"101001111",
  33042=>"001111011",
  33043=>"000101101",
  33044=>"010101001",
  33045=>"001000001",
  33046=>"000010000",
  33047=>"111101010",
  33048=>"101111110",
  33049=>"101011011",
  33050=>"110011100",
  33051=>"101100011",
  33052=>"011001101",
  33053=>"010010010",
  33054=>"010111001",
  33055=>"001000110",
  33056=>"100000001",
  33057=>"111110001",
  33058=>"111100000",
  33059=>"100101011",
  33060=>"111011011",
  33061=>"011110101",
  33062=>"101010111",
  33063=>"001111101",
  33064=>"100010010",
  33065=>"000111101",
  33066=>"000100100",
  33067=>"000011000",
  33068=>"101111001",
  33069=>"100000110",
  33070=>"000011110",
  33071=>"101101000",
  33072=>"001101110",
  33073=>"100010000",
  33074=>"100010111",
  33075=>"101000100",
  33076=>"101100110",
  33077=>"010111011",
  33078=>"010011010",
  33079=>"010111011",
  33080=>"111100110",
  33081=>"110010111",
  33082=>"001000010",
  33083=>"101110101",
  33084=>"101010000",
  33085=>"011000110",
  33086=>"010010000",
  33087=>"010111001",
  33088=>"001010011",
  33089=>"000101110",
  33090=>"111111001",
  33091=>"001101010",
  33092=>"010010111",
  33093=>"101010111",
  33094=>"101001110",
  33095=>"101001011",
  33096=>"110101100",
  33097=>"000100100",
  33098=>"100101000",
  33099=>"010011010",
  33100=>"101001101",
  33101=>"100001001",
  33102=>"010000001",
  33103=>"000001110",
  33104=>"100110101",
  33105=>"000001010",
  33106=>"010011100",
  33107=>"111111101",
  33108=>"010000001",
  33109=>"111100000",
  33110=>"100110101",
  33111=>"011101100",
  33112=>"001001100",
  33113=>"000001100",
  33114=>"110010000",
  33115=>"111001111",
  33116=>"100101011",
  33117=>"100000011",
  33118=>"001101100",
  33119=>"010101001",
  33120=>"001001001",
  33121=>"010111101",
  33122=>"001000100",
  33123=>"000011111",
  33124=>"111100000",
  33125=>"111001010",
  33126=>"010001101",
  33127=>"001110110",
  33128=>"110000110",
  33129=>"110000100",
  33130=>"111011000",
  33131=>"011001100",
  33132=>"110001100",
  33133=>"100010011",
  33134=>"000110101",
  33135=>"010111111",
  33136=>"001000111",
  33137=>"011100011",
  33138=>"011101000",
  33139=>"001100000",
  33140=>"101101110",
  33141=>"110011111",
  33142=>"000000111",
  33143=>"001011001",
  33144=>"011001101",
  33145=>"000010011",
  33146=>"111111101",
  33147=>"001011100",
  33148=>"111001100",
  33149=>"010111001",
  33150=>"011110100",
  33151=>"000010100",
  33152=>"010110100",
  33153=>"111001111",
  33154=>"001001111",
  33155=>"101110010",
  33156=>"011101111",
  33157=>"001111110",
  33158=>"111010001",
  33159=>"101100101",
  33160=>"011010111",
  33161=>"000010001",
  33162=>"001011110",
  33163=>"000110000",
  33164=>"001110100",
  33165=>"000011101",
  33166=>"110001011",
  33167=>"100100001",
  33168=>"110100110",
  33169=>"110010010",
  33170=>"010100010",
  33171=>"001010111",
  33172=>"101110111",
  33173=>"000001001",
  33174=>"000111110",
  33175=>"001111111",
  33176=>"110011101",
  33177=>"100111010",
  33178=>"000101100",
  33179=>"011010011",
  33180=>"011010000",
  33181=>"010000011",
  33182=>"000111010",
  33183=>"110110101",
  33184=>"110011011",
  33185=>"111001011",
  33186=>"001011000",
  33187=>"111011011",
  33188=>"010111011",
  33189=>"010011101",
  33190=>"110001111",
  33191=>"010100011",
  33192=>"111110100",
  33193=>"111010111",
  33194=>"010110111",
  33195=>"110011111",
  33196=>"011101010",
  33197=>"000011101",
  33198=>"110000010",
  33199=>"010111110",
  33200=>"111011110",
  33201=>"100100010",
  33202=>"001100100",
  33203=>"000010011",
  33204=>"010010101",
  33205=>"000010000",
  33206=>"001001010",
  33207=>"000111010",
  33208=>"111011011",
  33209=>"000100000",
  33210=>"000010011",
  33211=>"001111111",
  33212=>"101000000",
  33213=>"111011001",
  33214=>"111101001",
  33215=>"011100111",
  33216=>"000011111",
  33217=>"101001101",
  33218=>"110111010",
  33219=>"100100011",
  33220=>"110011000",
  33221=>"001010110",
  33222=>"010010011",
  33223=>"000000000",
  33224=>"011111000",
  33225=>"101011110",
  33226=>"011000011",
  33227=>"001000110",
  33228=>"000000001",
  33229=>"101100111",
  33230=>"110100100",
  33231=>"100001011",
  33232=>"110100100",
  33233=>"110011111",
  33234=>"100000101",
  33235=>"111001010",
  33236=>"110010010",
  33237=>"111101010",
  33238=>"110001010",
  33239=>"110111010",
  33240=>"010011101",
  33241=>"111101101",
  33242=>"100000011",
  33243=>"001001000",
  33244=>"101110110",
  33245=>"111011011",
  33246=>"110010001",
  33247=>"110111011",
  33248=>"110011110",
  33249=>"011101011",
  33250=>"111000110",
  33251=>"001101100",
  33252=>"100111100",
  33253=>"100011001",
  33254=>"111110100",
  33255=>"001110100",
  33256=>"100001011",
  33257=>"101100101",
  33258=>"010110011",
  33259=>"111110011",
  33260=>"101100000",
  33261=>"110011011",
  33262=>"110000011",
  33263=>"001000011",
  33264=>"011001100",
  33265=>"011101001",
  33266=>"011000000",
  33267=>"000100010",
  33268=>"100011110",
  33269=>"101010000",
  33270=>"000111000",
  33271=>"011010110",
  33272=>"110100011",
  33273=>"000011110",
  33274=>"000001011",
  33275=>"100110100",
  33276=>"010010010",
  33277=>"100010001",
  33278=>"000100000",
  33279=>"001100100",
  33280=>"011100010",
  33281=>"010100111",
  33282=>"111100110",
  33283=>"101110111",
  33284=>"010001010",
  33285=>"011101111",
  33286=>"100001101",
  33287=>"001101111",
  33288=>"101100001",
  33289=>"010111011",
  33290=>"010110001",
  33291=>"100110010",
  33292=>"101011010",
  33293=>"010010011",
  33294=>"000000110",
  33295=>"000011010",
  33296=>"101010110",
  33297=>"111111011",
  33298=>"100000000",
  33299=>"001001100",
  33300=>"011001001",
  33301=>"000001100",
  33302=>"101101101",
  33303=>"100101111",
  33304=>"011000001",
  33305=>"010000010",
  33306=>"111101100",
  33307=>"101011001",
  33308=>"111011101",
  33309=>"101000111",
  33310=>"100100000",
  33311=>"000010011",
  33312=>"110101100",
  33313=>"101000010",
  33314=>"111011001",
  33315=>"000001111",
  33316=>"100111001",
  33317=>"010100001",
  33318=>"111110110",
  33319=>"000110000",
  33320=>"110010101",
  33321=>"110100100",
  33322=>"111111110",
  33323=>"010010110",
  33324=>"111101100",
  33325=>"100000100",
  33326=>"111001100",
  33327=>"000100111",
  33328=>"111111011",
  33329=>"111101101",
  33330=>"000010110",
  33331=>"001000011",
  33332=>"100001011",
  33333=>"000011001",
  33334=>"110101100",
  33335=>"010001111",
  33336=>"000001111",
  33337=>"101010100",
  33338=>"100100111",
  33339=>"010100011",
  33340=>"100010000",
  33341=>"000011010",
  33342=>"100110111",
  33343=>"010101011",
  33344=>"110100011",
  33345=>"100101011",
  33346=>"100110011",
  33347=>"111000001",
  33348=>"111101101",
  33349=>"101000101",
  33350=>"000010001",
  33351=>"011110000",
  33352=>"011010101",
  33353=>"101101001",
  33354=>"001101100",
  33355=>"110010110",
  33356=>"010110000",
  33357=>"000001100",
  33358=>"010110010",
  33359=>"110101010",
  33360=>"101100011",
  33361=>"101011110",
  33362=>"001101001",
  33363=>"001101011",
  33364=>"001000100",
  33365=>"001100110",
  33366=>"101000100",
  33367=>"110100000",
  33368=>"001110110",
  33369=>"100010101",
  33370=>"101010001",
  33371=>"001100111",
  33372=>"110001011",
  33373=>"010100100",
  33374=>"011110010",
  33375=>"101111111",
  33376=>"010001100",
  33377=>"011010111",
  33378=>"001011000",
  33379=>"000110000",
  33380=>"110110110",
  33381=>"111111101",
  33382=>"011000100",
  33383=>"111111011",
  33384=>"000000100",
  33385=>"000000001",
  33386=>"110111000",
  33387=>"001101010",
  33388=>"110101010",
  33389=>"100101010",
  33390=>"100001100",
  33391=>"100101110",
  33392=>"100110110",
  33393=>"100000110",
  33394=>"110101011",
  33395=>"111101011",
  33396=>"111110000",
  33397=>"011000101",
  33398=>"111101101",
  33399=>"001111010",
  33400=>"101101111",
  33401=>"011100101",
  33402=>"111111011",
  33403=>"010111111",
  33404=>"000111010",
  33405=>"100001011",
  33406=>"000100101",
  33407=>"110101010",
  33408=>"010000110",
  33409=>"000000101",
  33410=>"111010111",
  33411=>"111010100",
  33412=>"111001100",
  33413=>"011111110",
  33414=>"001101001",
  33415=>"011100000",
  33416=>"010010100",
  33417=>"001111101",
  33418=>"110010011",
  33419=>"111010100",
  33420=>"111000111",
  33421=>"100111101",
  33422=>"100110000",
  33423=>"100110111",
  33424=>"110101001",
  33425=>"101001110",
  33426=>"010010101",
  33427=>"111010111",
  33428=>"011110000",
  33429=>"011011010",
  33430=>"001101101",
  33431=>"110000010",
  33432=>"110111111",
  33433=>"010000010",
  33434=>"101011100",
  33435=>"000110101",
  33436=>"111111001",
  33437=>"000001000",
  33438=>"000010111",
  33439=>"110101000",
  33440=>"101000101",
  33441=>"110001001",
  33442=>"101100111",
  33443=>"011110100",
  33444=>"000010010",
  33445=>"111011101",
  33446=>"011100111",
  33447=>"100100110",
  33448=>"110110000",
  33449=>"011010011",
  33450=>"110101111",
  33451=>"101000000",
  33452=>"110000001",
  33453=>"100110011",
  33454=>"000010011",
  33455=>"100000000",
  33456=>"010001000",
  33457=>"100101110",
  33458=>"100101101",
  33459=>"100011101",
  33460=>"011110001",
  33461=>"001011111",
  33462=>"000100100",
  33463=>"000000001",
  33464=>"011001101",
  33465=>"010001000",
  33466=>"101011001",
  33467=>"000010010",
  33468=>"011110001",
  33469=>"011011110",
  33470=>"100011111",
  33471=>"111010111",
  33472=>"010101101",
  33473=>"000110111",
  33474=>"100001100",
  33475=>"111101101",
  33476=>"110110110",
  33477=>"101001001",
  33478=>"011011000",
  33479=>"001010110",
  33480=>"101001100",
  33481=>"010010001",
  33482=>"010011110",
  33483=>"101000100",
  33484=>"111100000",
  33485=>"000001111",
  33486=>"101101101",
  33487=>"100111110",
  33488=>"010011100",
  33489=>"111001010",
  33490=>"001001001",
  33491=>"010010110",
  33492=>"110110001",
  33493=>"011100010",
  33494=>"010100011",
  33495=>"001100110",
  33496=>"110111001",
  33497=>"000011101",
  33498=>"110000000",
  33499=>"001101101",
  33500=>"101101000",
  33501=>"000100011",
  33502=>"010011001",
  33503=>"000011100",
  33504=>"011000101",
  33505=>"000100001",
  33506=>"011100001",
  33507=>"100010001",
  33508=>"011001000",
  33509=>"101001011",
  33510=>"000010010",
  33511=>"010010111",
  33512=>"110001110",
  33513=>"100110110",
  33514=>"010010111",
  33515=>"110001001",
  33516=>"100111111",
  33517=>"110010001",
  33518=>"110111101",
  33519=>"101000000",
  33520=>"110110000",
  33521=>"000010000",
  33522=>"100000011",
  33523=>"111111101",
  33524=>"011010011",
  33525=>"101111101",
  33526=>"001100110",
  33527=>"111110110",
  33528=>"100000110",
  33529=>"110101000",
  33530=>"010101101",
  33531=>"110111001",
  33532=>"001000010",
  33533=>"010110110",
  33534=>"100010010",
  33535=>"011000100",
  33536=>"011101010",
  33537=>"001011111",
  33538=>"101101111",
  33539=>"100011001",
  33540=>"101010001",
  33541=>"001000110",
  33542=>"100000001",
  33543=>"001000000",
  33544=>"001011110",
  33545=>"011100101",
  33546=>"011000100",
  33547=>"011010111",
  33548=>"000111100",
  33549=>"000100000",
  33550=>"001110011",
  33551=>"011011110",
  33552=>"001000111",
  33553=>"010101010",
  33554=>"110101100",
  33555=>"011001111",
  33556=>"010010111",
  33557=>"000001011",
  33558=>"001101011",
  33559=>"011100110",
  33560=>"100000111",
  33561=>"101010001",
  33562=>"010010110",
  33563=>"001111110",
  33564=>"011101010",
  33565=>"001100001",
  33566=>"100111111",
  33567=>"001010011",
  33568=>"011001000",
  33569=>"011000000",
  33570=>"111010010",
  33571=>"101100011",
  33572=>"011010010",
  33573=>"000001010",
  33574=>"011001011",
  33575=>"100101111",
  33576=>"101010100",
  33577=>"100011100",
  33578=>"000111011",
  33579=>"001101100",
  33580=>"110001010",
  33581=>"000000110",
  33582=>"011110010",
  33583=>"010011111",
  33584=>"000001010",
  33585=>"101100100",
  33586=>"100111000",
  33587=>"010000111",
  33588=>"010011101",
  33589=>"011100100",
  33590=>"010001001",
  33591=>"101000100",
  33592=>"000100101",
  33593=>"001011000",
  33594=>"001101001",
  33595=>"100100000",
  33596=>"110100100",
  33597=>"110010111",
  33598=>"101110101",
  33599=>"111110110",
  33600=>"111111010",
  33601=>"010110001",
  33602=>"001100011",
  33603=>"011110110",
  33604=>"011010110",
  33605=>"111000011",
  33606=>"110000101",
  33607=>"010011001",
  33608=>"111110011",
  33609=>"100000100",
  33610=>"100010100",
  33611=>"000010111",
  33612=>"001110000",
  33613=>"111110001",
  33614=>"111110001",
  33615=>"000001100",
  33616=>"111100100",
  33617=>"110101001",
  33618=>"000010011",
  33619=>"111101111",
  33620=>"010111000",
  33621=>"010111010",
  33622=>"001110101",
  33623=>"010010001",
  33624=>"110110000",
  33625=>"100111110",
  33626=>"001111111",
  33627=>"110011110",
  33628=>"101011011",
  33629=>"101010001",
  33630=>"111011001",
  33631=>"110001000",
  33632=>"110011000",
  33633=>"000010010",
  33634=>"100001100",
  33635=>"111111010",
  33636=>"110000110",
  33637=>"110000010",
  33638=>"011010011",
  33639=>"111000111",
  33640=>"000100100",
  33641=>"011111000",
  33642=>"110101010",
  33643=>"110100010",
  33644=>"111110101",
  33645=>"011010111",
  33646=>"011110100",
  33647=>"010110110",
  33648=>"100000000",
  33649=>"111001110",
  33650=>"111000110",
  33651=>"001100010",
  33652=>"100100110",
  33653=>"001111001",
  33654=>"001001000",
  33655=>"011101000",
  33656=>"001000010",
  33657=>"010001111",
  33658=>"110100010",
  33659=>"001111010",
  33660=>"001000111",
  33661=>"000110000",
  33662=>"110110111",
  33663=>"010010001",
  33664=>"110010001",
  33665=>"010101101",
  33666=>"110000111",
  33667=>"000100001",
  33668=>"111110101",
  33669=>"111110001",
  33670=>"011001010",
  33671=>"111011101",
  33672=>"100010101",
  33673=>"010111010",
  33674=>"111001110",
  33675=>"110101001",
  33676=>"010011000",
  33677=>"111011010",
  33678=>"000101000",
  33679=>"100010010",
  33680=>"111010000",
  33681=>"101001000",
  33682=>"000010100",
  33683=>"111001001",
  33684=>"111110011",
  33685=>"101101101",
  33686=>"001000001",
  33687=>"100010001",
  33688=>"011100011",
  33689=>"010000111",
  33690=>"111110100",
  33691=>"101110001",
  33692=>"100110010",
  33693=>"110001011",
  33694=>"111111100",
  33695=>"001000000",
  33696=>"100010011",
  33697=>"000100011",
  33698=>"010001101",
  33699=>"111111111",
  33700=>"011101110",
  33701=>"000110101",
  33702=>"101101011",
  33703=>"010000100",
  33704=>"100111101",
  33705=>"011011010",
  33706=>"001001100",
  33707=>"100011101",
  33708=>"000101001",
  33709=>"010000000",
  33710=>"010010111",
  33711=>"100011010",
  33712=>"000110000",
  33713=>"010110100",
  33714=>"001011000",
  33715=>"010010010",
  33716=>"011100100",
  33717=>"111101101",
  33718=>"101010000",
  33719=>"000110000",
  33720=>"100000110",
  33721=>"000111001",
  33722=>"100000000",
  33723=>"010100111",
  33724=>"010111111",
  33725=>"100011011",
  33726=>"101001010",
  33727=>"111000110",
  33728=>"011101001",
  33729=>"101111110",
  33730=>"101011011",
  33731=>"111101001",
  33732=>"000000100",
  33733=>"010001010",
  33734=>"011110001",
  33735=>"000000101",
  33736=>"000000010",
  33737=>"010010011",
  33738=>"110110101",
  33739=>"110100101",
  33740=>"100001101",
  33741=>"111101000",
  33742=>"100010000",
  33743=>"011001000",
  33744=>"010110110",
  33745=>"110110111",
  33746=>"011000100",
  33747=>"110110111",
  33748=>"000000001",
  33749=>"100010001",
  33750=>"110110001",
  33751=>"000001101",
  33752=>"011001111",
  33753=>"011010000",
  33754=>"110010110",
  33755=>"011011111",
  33756=>"111111101",
  33757=>"001001111",
  33758=>"000111111",
  33759=>"110010111",
  33760=>"110111111",
  33761=>"110011010",
  33762=>"010101001",
  33763=>"001010011",
  33764=>"110100000",
  33765=>"011111100",
  33766=>"000010100",
  33767=>"100100010",
  33768=>"101000010",
  33769=>"111000000",
  33770=>"100000010",
  33771=>"010001111",
  33772=>"101100100",
  33773=>"001000000",
  33774=>"110000100",
  33775=>"001110010",
  33776=>"100011010",
  33777=>"000100000",
  33778=>"011111011",
  33779=>"111111110",
  33780=>"110110010",
  33781=>"101101101",
  33782=>"000000111",
  33783=>"111000100",
  33784=>"001001010",
  33785=>"100001101",
  33786=>"101000101",
  33787=>"001110110",
  33788=>"000100010",
  33789=>"010011111",
  33790=>"000101100",
  33791=>"010100000",
  33792=>"001010010",
  33793=>"010010010",
  33794=>"100000000",
  33795=>"000101110",
  33796=>"001100000",
  33797=>"001001110",
  33798=>"100011101",
  33799=>"111001110",
  33800=>"110001100",
  33801=>"100000000",
  33802=>"101101101",
  33803=>"111111111",
  33804=>"011100111",
  33805=>"110111111",
  33806=>"011001110",
  33807=>"011100101",
  33808=>"010110100",
  33809=>"100001101",
  33810=>"101010100",
  33811=>"000100110",
  33812=>"110000010",
  33813=>"101110001",
  33814=>"010110111",
  33815=>"100110110",
  33816=>"001011111",
  33817=>"000010000",
  33818=>"110111000",
  33819=>"010110110",
  33820=>"011000101",
  33821=>"110111000",
  33822=>"100010111",
  33823=>"011000000",
  33824=>"011001000",
  33825=>"000011101",
  33826=>"010110000",
  33827=>"100000111",
  33828=>"001000110",
  33829=>"110111111",
  33830=>"100111000",
  33831=>"110100000",
  33832=>"010011100",
  33833=>"000111011",
  33834=>"101101110",
  33835=>"110100010",
  33836=>"000000000",
  33837=>"100000000",
  33838=>"001001100",
  33839=>"011010101",
  33840=>"001000000",
  33841=>"111101110",
  33842=>"111110010",
  33843=>"000000100",
  33844=>"011001000",
  33845=>"001000011",
  33846=>"000010111",
  33847=>"010000100",
  33848=>"000011011",
  33849=>"011101001",
  33850=>"100100010",
  33851=>"111100010",
  33852=>"000010110",
  33853=>"101010100",
  33854=>"101011101",
  33855=>"100010110",
  33856=>"000010000",
  33857=>"000110110",
  33858=>"010001000",
  33859=>"000000010",
  33860=>"100110011",
  33861=>"001010100",
  33862=>"101010011",
  33863=>"000101010",
  33864=>"010100010",
  33865=>"100001101",
  33866=>"000111011",
  33867=>"111011001",
  33868=>"010111011",
  33869=>"011110000",
  33870=>"111100001",
  33871=>"010000011",
  33872=>"001100100",
  33873=>"000001101",
  33874=>"110011111",
  33875=>"101110001",
  33876=>"001100011",
  33877=>"101101110",
  33878=>"111111101",
  33879=>"101000111",
  33880=>"110011001",
  33881=>"101010001",
  33882=>"001110010",
  33883=>"110010001",
  33884=>"100100000",
  33885=>"100011111",
  33886=>"011101111",
  33887=>"111110100",
  33888=>"011001100",
  33889=>"000001010",
  33890=>"101101011",
  33891=>"001110011",
  33892=>"000010101",
  33893=>"100100110",
  33894=>"000110111",
  33895=>"001110110",
  33896=>"010101000",
  33897=>"111000001",
  33898=>"101001000",
  33899=>"010101010",
  33900=>"011000001",
  33901=>"010000110",
  33902=>"111100111",
  33903=>"101001110",
  33904=>"000000011",
  33905=>"111000100",
  33906=>"110110000",
  33907=>"110100111",
  33908=>"101010110",
  33909=>"101001010",
  33910=>"000010111",
  33911=>"001111111",
  33912=>"111101010",
  33913=>"000010100",
  33914=>"000100010",
  33915=>"001100011",
  33916=>"110001010",
  33917=>"111101000",
  33918=>"010010011",
  33919=>"110010010",
  33920=>"100000011",
  33921=>"111011011",
  33922=>"010000111",
  33923=>"111011000",
  33924=>"101000000",
  33925=>"101011111",
  33926=>"100100101",
  33927=>"000010000",
  33928=>"101001011",
  33929=>"011010110",
  33930=>"110100111",
  33931=>"001100001",
  33932=>"000110001",
  33933=>"110110100",
  33934=>"101001111",
  33935=>"000101000",
  33936=>"000100011",
  33937=>"010000001",
  33938=>"111111010",
  33939=>"000101011",
  33940=>"111100111",
  33941=>"010011111",
  33942=>"010101111",
  33943=>"000010100",
  33944=>"100011110",
  33945=>"110001011",
  33946=>"101011111",
  33947=>"100001010",
  33948=>"000101111",
  33949=>"010011100",
  33950=>"110111001",
  33951=>"111010000",
  33952=>"101010110",
  33953=>"110001111",
  33954=>"101010000",
  33955=>"011010001",
  33956=>"111111100",
  33957=>"010000011",
  33958=>"111001010",
  33959=>"011001110",
  33960=>"000010100",
  33961=>"100000100",
  33962=>"110001000",
  33963=>"111110000",
  33964=>"110000011",
  33965=>"101001011",
  33966=>"111100110",
  33967=>"011011010",
  33968=>"000011111",
  33969=>"110010011",
  33970=>"000111111",
  33971=>"011001000",
  33972=>"100010100",
  33973=>"000011101",
  33974=>"011011001",
  33975=>"100010000",
  33976=>"001011000",
  33977=>"001011000",
  33978=>"100101101",
  33979=>"010101000",
  33980=>"011111011",
  33981=>"001110000",
  33982=>"100101100",
  33983=>"010100011",
  33984=>"101111101",
  33985=>"101101010",
  33986=>"000010100",
  33987=>"111100001",
  33988=>"000110010",
  33989=>"001110110",
  33990=>"011011001",
  33991=>"110010010",
  33992=>"000100101",
  33993=>"001000101",
  33994=>"100011000",
  33995=>"111010011",
  33996=>"101011111",
  33997=>"111100111",
  33998=>"000100100",
  33999=>"110001111",
  34000=>"011110100",
  34001=>"011010011",
  34002=>"001010011",
  34003=>"101110010",
  34004=>"000101110",
  34005=>"011101101",
  34006=>"110001100",
  34007=>"101110011",
  34008=>"110010001",
  34009=>"011101011",
  34010=>"101110110",
  34011=>"011100001",
  34012=>"001011001",
  34013=>"100101011",
  34014=>"011010010",
  34015=>"110000011",
  34016=>"000101111",
  34017=>"101110010",
  34018=>"111101010",
  34019=>"101100001",
  34020=>"101011000",
  34021=>"001110000",
  34022=>"110111110",
  34023=>"011110000",
  34024=>"101001010",
  34025=>"011110010",
  34026=>"001011100",
  34027=>"000100011",
  34028=>"101111000",
  34029=>"110010001",
  34030=>"110000111",
  34031=>"001001110",
  34032=>"111110010",
  34033=>"110000100",
  34034=>"100100010",
  34035=>"110101000",
  34036=>"101111000",
  34037=>"011010101",
  34038=>"011100100",
  34039=>"100001000",
  34040=>"100110000",
  34041=>"101100000",
  34042=>"001001100",
  34043=>"000011110",
  34044=>"111101000",
  34045=>"001000110",
  34046=>"100000010",
  34047=>"111100111",
  34048=>"001111010",
  34049=>"000101100",
  34050=>"100011111",
  34051=>"001110100",
  34052=>"110001010",
  34053=>"110010000",
  34054=>"011110111",
  34055=>"100000000",
  34056=>"000000001",
  34057=>"101111100",
  34058=>"111010110",
  34059=>"100101011",
  34060=>"001100101",
  34061=>"010011010",
  34062=>"100010010",
  34063=>"011100101",
  34064=>"011111100",
  34065=>"110011010",
  34066=>"100111111",
  34067=>"001100100",
  34068=>"101111010",
  34069=>"101011100",
  34070=>"001101000",
  34071=>"100010110",
  34072=>"000010001",
  34073=>"000111011",
  34074=>"010011010",
  34075=>"110100010",
  34076=>"000011000",
  34077=>"101100000",
  34078=>"110111100",
  34079=>"000010111",
  34080=>"001000101",
  34081=>"001110110",
  34082=>"101110110",
  34083=>"011010001",
  34084=>"011100010",
  34085=>"100111010",
  34086=>"110111000",
  34087=>"100100101",
  34088=>"000001101",
  34089=>"000100010",
  34090=>"000100001",
  34091=>"011110011",
  34092=>"100101010",
  34093=>"000000101",
  34094=>"110001101",
  34095=>"101001111",
  34096=>"000110100",
  34097=>"001010000",
  34098=>"001001100",
  34099=>"011100111",
  34100=>"010010010",
  34101=>"000001111",
  34102=>"001101001",
  34103=>"101100100",
  34104=>"000010101",
  34105=>"010000000",
  34106=>"110110101",
  34107=>"101010010",
  34108=>"110100101",
  34109=>"001011001",
  34110=>"011100101",
  34111=>"011010100",
  34112=>"101011010",
  34113=>"111000011",
  34114=>"010011101",
  34115=>"001100001",
  34116=>"101000111",
  34117=>"001110110",
  34118=>"110011011",
  34119=>"011110111",
  34120=>"110110111",
  34121=>"100110100",
  34122=>"001101100",
  34123=>"100001111",
  34124=>"100011111",
  34125=>"011011010",
  34126=>"110011010",
  34127=>"100110011",
  34128=>"101110110",
  34129=>"110111110",
  34130=>"110010000",
  34131=>"001000100",
  34132=>"000010001",
  34133=>"001100110",
  34134=>"010001000",
  34135=>"000111101",
  34136=>"000111000",
  34137=>"101101011",
  34138=>"010111110",
  34139=>"100000101",
  34140=>"110011101",
  34141=>"110000001",
  34142=>"010101010",
  34143=>"011010110",
  34144=>"001010001",
  34145=>"010001100",
  34146=>"011100010",
  34147=>"101010110",
  34148=>"000011001",
  34149=>"010000011",
  34150=>"100101101",
  34151=>"111100001",
  34152=>"111101100",
  34153=>"001000110",
  34154=>"110100011",
  34155=>"011011011",
  34156=>"010001001",
  34157=>"011111100",
  34158=>"001011101",
  34159=>"011110111",
  34160=>"001001100",
  34161=>"101001111",
  34162=>"111110000",
  34163=>"111000010",
  34164=>"010110111",
  34165=>"111010000",
  34166=>"110100010",
  34167=>"100010011",
  34168=>"111010011",
  34169=>"001011100",
  34170=>"110010101",
  34171=>"100000111",
  34172=>"111101011",
  34173=>"101111101",
  34174=>"001010000",
  34175=>"111111101",
  34176=>"000100110",
  34177=>"010010100",
  34178=>"100110101",
  34179=>"010010000",
  34180=>"000010111",
  34181=>"000001000",
  34182=>"100110111",
  34183=>"010110100",
  34184=>"001110111",
  34185=>"110100100",
  34186=>"101101010",
  34187=>"110110101",
  34188=>"001010001",
  34189=>"001100100",
  34190=>"000001100",
  34191=>"110101000",
  34192=>"111100010",
  34193=>"000000101",
  34194=>"111111100",
  34195=>"011111010",
  34196=>"110111010",
  34197=>"100110110",
  34198=>"000100101",
  34199=>"100111101",
  34200=>"110111000",
  34201=>"100111011",
  34202=>"011000101",
  34203=>"110000101",
  34204=>"010100100",
  34205=>"000100100",
  34206=>"111111001",
  34207=>"010001010",
  34208=>"000001001",
  34209=>"011011010",
  34210=>"101001100",
  34211=>"111001110",
  34212=>"011010000",
  34213=>"000000011",
  34214=>"000011001",
  34215=>"001011110",
  34216=>"011110110",
  34217=>"000011000",
  34218=>"001111110",
  34219=>"010001111",
  34220=>"010100101",
  34221=>"010000011",
  34222=>"000000000",
  34223=>"000000000",
  34224=>"101001100",
  34225=>"111110001",
  34226=>"111011110",
  34227=>"000111111",
  34228=>"101100010",
  34229=>"000101001",
  34230=>"001000110",
  34231=>"111011011",
  34232=>"101101111",
  34233=>"100100111",
  34234=>"101100010",
  34235=>"011101001",
  34236=>"111011000",
  34237=>"101010011",
  34238=>"010011110",
  34239=>"000010100",
  34240=>"111101101",
  34241=>"000010010",
  34242=>"010000110",
  34243=>"100111010",
  34244=>"011001000",
  34245=>"110010000",
  34246=>"111000000",
  34247=>"010000000",
  34248=>"111110011",
  34249=>"000101100",
  34250=>"001000011",
  34251=>"001101010",
  34252=>"000101111",
  34253=>"011110110",
  34254=>"000110111",
  34255=>"110001111",
  34256=>"111010000",
  34257=>"000111110",
  34258=>"011110111",
  34259=>"000010111",
  34260=>"000111111",
  34261=>"010111001",
  34262=>"010111001",
  34263=>"000000101",
  34264=>"111110101",
  34265=>"001010110",
  34266=>"111101100",
  34267=>"000100000",
  34268=>"010001100",
  34269=>"011101010",
  34270=>"011011010",
  34271=>"011101000",
  34272=>"001110111",
  34273=>"001100000",
  34274=>"001011010",
  34275=>"101001110",
  34276=>"010110001",
  34277=>"001010001",
  34278=>"111101011",
  34279=>"001100000",
  34280=>"110111100",
  34281=>"111010101",
  34282=>"000011010",
  34283=>"111100000",
  34284=>"111000111",
  34285=>"011100010",
  34286=>"000111110",
  34287=>"110110001",
  34288=>"000110100",
  34289=>"011100111",
  34290=>"100100000",
  34291=>"001101000",
  34292=>"010101110",
  34293=>"001001100",
  34294=>"000100101",
  34295=>"000110100",
  34296=>"110100011",
  34297=>"011111010",
  34298=>"000001000",
  34299=>"101100110",
  34300=>"000010010",
  34301=>"011001010",
  34302=>"111000010",
  34303=>"010000110",
  34304=>"111111001",
  34305=>"001101111",
  34306=>"111010001",
  34307=>"110101111",
  34308=>"101010100",
  34309=>"100001001",
  34310=>"101010110",
  34311=>"110000010",
  34312=>"001001111",
  34313=>"000110100",
  34314=>"100111110",
  34315=>"010001010",
  34316=>"011111011",
  34317=>"001101101",
  34318=>"010000010",
  34319=>"001001100",
  34320=>"100011000",
  34321=>"100010101",
  34322=>"100101111",
  34323=>"111111001",
  34324=>"101010101",
  34325=>"110100001",
  34326=>"110001101",
  34327=>"101001001",
  34328=>"011011010",
  34329=>"000000001",
  34330=>"001011011",
  34331=>"110001101",
  34332=>"000001110",
  34333=>"000100010",
  34334=>"011101111",
  34335=>"111101011",
  34336=>"010000011",
  34337=>"100100100",
  34338=>"011010111",
  34339=>"110010010",
  34340=>"100000101",
  34341=>"101001111",
  34342=>"000101011",
  34343=>"010111100",
  34344=>"010101000",
  34345=>"110011011",
  34346=>"110000100",
  34347=>"111100111",
  34348=>"110000000",
  34349=>"101101010",
  34350=>"100100000",
  34351=>"010001101",
  34352=>"101100111",
  34353=>"110101001",
  34354=>"001000101",
  34355=>"010110111",
  34356=>"010100111",
  34357=>"010000110",
  34358=>"010000000",
  34359=>"110001111",
  34360=>"111001001",
  34361=>"100010110",
  34362=>"111011001",
  34363=>"010100100",
  34364=>"111110000",
  34365=>"111011111",
  34366=>"011010011",
  34367=>"010110101",
  34368=>"000001001",
  34369=>"000110010",
  34370=>"100010001",
  34371=>"010001001",
  34372=>"010010001",
  34373=>"111011110",
  34374=>"100101111",
  34375=>"001111110",
  34376=>"000001100",
  34377=>"111111001",
  34378=>"111011010",
  34379=>"110011001",
  34380=>"000110001",
  34381=>"000000111",
  34382=>"110010100",
  34383=>"000010001",
  34384=>"010010001",
  34385=>"111000010",
  34386=>"000001010",
  34387=>"101111001",
  34388=>"001001100",
  34389=>"000111111",
  34390=>"000111111",
  34391=>"111101111",
  34392=>"001011010",
  34393=>"000111010",
  34394=>"110000011",
  34395=>"100011001",
  34396=>"100000100",
  34397=>"000000001",
  34398=>"100111011",
  34399=>"100101100",
  34400=>"010000011",
  34401=>"011000100",
  34402=>"101010111",
  34403=>"001111100",
  34404=>"011001101",
  34405=>"001110010",
  34406=>"111010000",
  34407=>"001000000",
  34408=>"000101010",
  34409=>"000110001",
  34410=>"100110111",
  34411=>"110000111",
  34412=>"000111011",
  34413=>"011011010",
  34414=>"001011001",
  34415=>"111111001",
  34416=>"110000101",
  34417=>"101011111",
  34418=>"001011100",
  34419=>"101010100",
  34420=>"111010011",
  34421=>"001001010",
  34422=>"000000011",
  34423=>"111110010",
  34424=>"001000011",
  34425=>"010010001",
  34426=>"111011000",
  34427=>"010000111",
  34428=>"011110110",
  34429=>"000000001",
  34430=>"010010000",
  34431=>"110100000",
  34432=>"101110000",
  34433=>"111111110",
  34434=>"000100001",
  34435=>"011000011",
  34436=>"001110001",
  34437=>"110111111",
  34438=>"000100111",
  34439=>"010010001",
  34440=>"110011101",
  34441=>"001001100",
  34442=>"111111100",
  34443=>"011011010",
  34444=>"001110101",
  34445=>"010001001",
  34446=>"100000010",
  34447=>"010110011",
  34448=>"011111000",
  34449=>"011000011",
  34450=>"010011001",
  34451=>"111101111",
  34452=>"000101110",
  34453=>"100101111",
  34454=>"110011101",
  34455=>"111011000",
  34456=>"000000111",
  34457=>"100110101",
  34458=>"111101010",
  34459=>"101110110",
  34460=>"011010001",
  34461=>"101111011",
  34462=>"101001000",
  34463=>"000010101",
  34464=>"111110110",
  34465=>"001101010",
  34466=>"101011111",
  34467=>"110010011",
  34468=>"001110000",
  34469=>"101001111",
  34470=>"101011000",
  34471=>"111000100",
  34472=>"110011111",
  34473=>"010001000",
  34474=>"101100101",
  34475=>"100100001",
  34476=>"111010110",
  34477=>"010100100",
  34478=>"011011010",
  34479=>"111000111",
  34480=>"000100001",
  34481=>"010100011",
  34482=>"010000001",
  34483=>"011111001",
  34484=>"101111111",
  34485=>"010010100",
  34486=>"011000001",
  34487=>"111010111",
  34488=>"010010110",
  34489=>"101111000",
  34490=>"101101100",
  34491=>"100011101",
  34492=>"010101001",
  34493=>"011111111",
  34494=>"000100100",
  34495=>"101010001",
  34496=>"010111011",
  34497=>"001000100",
  34498=>"000110001",
  34499=>"111101110",
  34500=>"001111110",
  34501=>"000011111",
  34502=>"111010000",
  34503=>"100010111",
  34504=>"000101000",
  34505=>"101010000",
  34506=>"011111111",
  34507=>"001000111",
  34508=>"000001011",
  34509=>"111101110",
  34510=>"001110101",
  34511=>"111111100",
  34512=>"001111111",
  34513=>"100010011",
  34514=>"101001110",
  34515=>"001000000",
  34516=>"001100011",
  34517=>"010000111",
  34518=>"101010011",
  34519=>"001000010",
  34520=>"001100101",
  34521=>"010100010",
  34522=>"111010000",
  34523=>"100100010",
  34524=>"100101011",
  34525=>"110100101",
  34526=>"011100110",
  34527=>"010101101",
  34528=>"111110111",
  34529=>"011010101",
  34530=>"010010011",
  34531=>"001010000",
  34532=>"101001000",
  34533=>"111010110",
  34534=>"111110010",
  34535=>"011101110",
  34536=>"010111001",
  34537=>"111101111",
  34538=>"001010100",
  34539=>"010001010",
  34540=>"001010111",
  34541=>"000110111",
  34542=>"101011001",
  34543=>"001101011",
  34544=>"110110101",
  34545=>"001111101",
  34546=>"101110001",
  34547=>"010101110",
  34548=>"011011011",
  34549=>"011100111",
  34550=>"110101110",
  34551=>"010111101",
  34552=>"011110110",
  34553=>"011111011",
  34554=>"010000001",
  34555=>"010010110",
  34556=>"010011100",
  34557=>"011111011",
  34558=>"001010010",
  34559=>"110011010",
  34560=>"011001010",
  34561=>"100111110",
  34562=>"000101101",
  34563=>"110000001",
  34564=>"101001010",
  34565=>"000000000",
  34566=>"011110010",
  34567=>"101100100",
  34568=>"110010011",
  34569=>"101101101",
  34570=>"000101111",
  34571=>"111001010",
  34572=>"010000001",
  34573=>"101001100",
  34574=>"111011010",
  34575=>"101101010",
  34576=>"011111000",
  34577=>"000111100",
  34578=>"000000001",
  34579=>"101111000",
  34580=>"011011000",
  34581=>"111011110",
  34582=>"000011111",
  34583=>"000101111",
  34584=>"000110001",
  34585=>"000010110",
  34586=>"101111111",
  34587=>"000000010",
  34588=>"000011011",
  34589=>"000001001",
  34590=>"000111111",
  34591=>"111100000",
  34592=>"100010001",
  34593=>"111111010",
  34594=>"101101100",
  34595=>"100011001",
  34596=>"000111101",
  34597=>"000000010",
  34598=>"110101011",
  34599=>"001001010",
  34600=>"001100111",
  34601=>"010000100",
  34602=>"011101100",
  34603=>"111010111",
  34604=>"011100010",
  34605=>"001111111",
  34606=>"000101101",
  34607=>"101000011",
  34608=>"010111111",
  34609=>"001110100",
  34610=>"100100000",
  34611=>"010100010",
  34612=>"001101000",
  34613=>"100011110",
  34614=>"001000101",
  34615=>"100101000",
  34616=>"010010110",
  34617=>"111101000",
  34618=>"100000001",
  34619=>"001001010",
  34620=>"110101101",
  34621=>"010011100",
  34622=>"100001010",
  34623=>"111010111",
  34624=>"100010101",
  34625=>"010011000",
  34626=>"111111110",
  34627=>"011110001",
  34628=>"010000001",
  34629=>"010011101",
  34630=>"101110100",
  34631=>"101110111",
  34632=>"101110011",
  34633=>"010101000",
  34634=>"111111101",
  34635=>"010111010",
  34636=>"110011100",
  34637=>"010001100",
  34638=>"100010101",
  34639=>"010101100",
  34640=>"011100111",
  34641=>"110101000",
  34642=>"000000001",
  34643=>"111011011",
  34644=>"011100100",
  34645=>"001111010",
  34646=>"101001110",
  34647=>"010000011",
  34648=>"110000100",
  34649=>"110010110",
  34650=>"111100000",
  34651=>"000010010",
  34652=>"011011101",
  34653=>"101011101",
  34654=>"000010110",
  34655=>"000000111",
  34656=>"110110101",
  34657=>"110100100",
  34658=>"001111111",
  34659=>"111111100",
  34660=>"100100100",
  34661=>"001000011",
  34662=>"101011111",
  34663=>"000100111",
  34664=>"010010000",
  34665=>"110001001",
  34666=>"100100000",
  34667=>"001101111",
  34668=>"001110000",
  34669=>"101011111",
  34670=>"101101101",
  34671=>"101001000",
  34672=>"000111100",
  34673=>"011001100",
  34674=>"010000111",
  34675=>"001111011",
  34676=>"101101101",
  34677=>"011101110",
  34678=>"001110000",
  34679=>"011100000",
  34680=>"001010100",
  34681=>"111001111",
  34682=>"001010000",
  34683=>"100000000",
  34684=>"100010100",
  34685=>"110011100",
  34686=>"000011110",
  34687=>"110000010",
  34688=>"111010110",
  34689=>"000001001",
  34690=>"101110001",
  34691=>"000001110",
  34692=>"011000110",
  34693=>"011111011",
  34694=>"001110110",
  34695=>"000000010",
  34696=>"110111111",
  34697=>"000011011",
  34698=>"010101111",
  34699=>"110000001",
  34700=>"011001111",
  34701=>"010110010",
  34702=>"011111000",
  34703=>"001011111",
  34704=>"100111111",
  34705=>"011011010",
  34706=>"000101100",
  34707=>"000010000",
  34708=>"001000100",
  34709=>"110111100",
  34710=>"100010000",
  34711=>"101101000",
  34712=>"101010011",
  34713=>"001011011",
  34714=>"000110000",
  34715=>"100111110",
  34716=>"001101000",
  34717=>"010101011",
  34718=>"010101000",
  34719=>"001101011",
  34720=>"000011111",
  34721=>"111110001",
  34722=>"110000111",
  34723=>"011010001",
  34724=>"100001001",
  34725=>"101000101",
  34726=>"000110111",
  34727=>"110110011",
  34728=>"011110010",
  34729=>"110011010",
  34730=>"111101111",
  34731=>"011110111",
  34732=>"101010101",
  34733=>"110101111",
  34734=>"111011000",
  34735=>"110000010",
  34736=>"110001100",
  34737=>"111110011",
  34738=>"100010111",
  34739=>"000010100",
  34740=>"111110011",
  34741=>"111111010",
  34742=>"110110010",
  34743=>"010000011",
  34744=>"001001110",
  34745=>"010101100",
  34746=>"000101111",
  34747=>"011001100",
  34748=>"011111101",
  34749=>"100100100",
  34750=>"110000101",
  34751=>"101101100",
  34752=>"000111111",
  34753=>"110000100",
  34754=>"101101111",
  34755=>"010000110",
  34756=>"011111111",
  34757=>"001101011",
  34758=>"101101111",
  34759=>"010010101",
  34760=>"000011010",
  34761=>"100100111",
  34762=>"100101011",
  34763=>"001100010",
  34764=>"011010010",
  34765=>"110000000",
  34766=>"101101101",
  34767=>"110110100",
  34768=>"000111111",
  34769=>"001001010",
  34770=>"011010111",
  34771=>"000000000",
  34772=>"011000010",
  34773=>"001001100",
  34774=>"100100010",
  34775=>"100101110",
  34776=>"001010000",
  34777=>"100000011",
  34778=>"110100001",
  34779=>"111000000",
  34780=>"101101011",
  34781=>"111010000",
  34782=>"110110010",
  34783=>"111000100",
  34784=>"101111001",
  34785=>"010101000",
  34786=>"110110010",
  34787=>"010101110",
  34788=>"000010111",
  34789=>"000010111",
  34790=>"101010111",
  34791=>"101001100",
  34792=>"001110010",
  34793=>"011110110",
  34794=>"011000101",
  34795=>"101101100",
  34796=>"001011001",
  34797=>"001000000",
  34798=>"001001001",
  34799=>"001100111",
  34800=>"100110100",
  34801=>"101001100",
  34802=>"000011000",
  34803=>"101001010",
  34804=>"011100000",
  34805=>"101110111",
  34806=>"000110010",
  34807=>"000011001",
  34808=>"010100010",
  34809=>"100000111",
  34810=>"001100001",
  34811=>"100110000",
  34812=>"000111101",
  34813=>"100111100",
  34814=>"100001111",
  34815=>"100010001",
  34816=>"010011110",
  34817=>"111001110",
  34818=>"110000001",
  34819=>"000010000",
  34820=>"111010010",
  34821=>"010101101",
  34822=>"010010000",
  34823=>"010000001",
  34824=>"101110101",
  34825=>"001000010",
  34826=>"111100011",
  34827=>"010000111",
  34828=>"010000100",
  34829=>"011100001",
  34830=>"000101010",
  34831=>"110011010",
  34832=>"011000111",
  34833=>"011101110",
  34834=>"101111110",
  34835=>"100010100",
  34836=>"110011100",
  34837=>"111000001",
  34838=>"101011001",
  34839=>"110101000",
  34840=>"000001010",
  34841=>"000100000",
  34842=>"010100100",
  34843=>"000000000",
  34844=>"001110101",
  34845=>"010011110",
  34846=>"110111110",
  34847=>"011100111",
  34848=>"010111001",
  34849=>"111100001",
  34850=>"111001111",
  34851=>"011110010",
  34852=>"010010101",
  34853=>"011111111",
  34854=>"011111010",
  34855=>"101001110",
  34856=>"001100100",
  34857=>"111111010",
  34858=>"100000100",
  34859=>"011000111",
  34860=>"000010000",
  34861=>"000100110",
  34862=>"001111111",
  34863=>"101010100",
  34864=>"011111100",
  34865=>"101000101",
  34866=>"101000101",
  34867=>"101100001",
  34868=>"001000100",
  34869=>"001100000",
  34870=>"001011010",
  34871=>"001011001",
  34872=>"110010101",
  34873=>"100010110",
  34874=>"101110101",
  34875=>"000011010",
  34876=>"010111010",
  34877=>"000000011",
  34878=>"001010000",
  34879=>"110011001",
  34880=>"011110100",
  34881=>"000101001",
  34882=>"111000011",
  34883=>"001110000",
  34884=>"101001001",
  34885=>"100100110",
  34886=>"110110010",
  34887=>"100101001",
  34888=>"011001000",
  34889=>"111011000",
  34890=>"110001101",
  34891=>"001100000",
  34892=>"011000001",
  34893=>"111110111",
  34894=>"001001000",
  34895=>"001110111",
  34896=>"110000000",
  34897=>"101000101",
  34898=>"110000110",
  34899=>"111011110",
  34900=>"000000001",
  34901=>"111110110",
  34902=>"010001000",
  34903=>"110001001",
  34904=>"100111110",
  34905=>"111010010",
  34906=>"000100010",
  34907=>"101001101",
  34908=>"000001010",
  34909=>"000101010",
  34910=>"111011100",
  34911=>"100001000",
  34912=>"000110010",
  34913=>"011101011",
  34914=>"011010000",
  34915=>"000101011",
  34916=>"001011000",
  34917=>"001101000",
  34918=>"111001111",
  34919=>"101111011",
  34920=>"100010101",
  34921=>"110101010",
  34922=>"111100111",
  34923=>"101101100",
  34924=>"000111100",
  34925=>"111100001",
  34926=>"111011101",
  34927=>"000000010",
  34928=>"000000011",
  34929=>"100111010",
  34930=>"111000010",
  34931=>"000001011",
  34932=>"101001000",
  34933=>"010101100",
  34934=>"101011001",
  34935=>"010111001",
  34936=>"111011101",
  34937=>"011000000",
  34938=>"011010001",
  34939=>"011110111",
  34940=>"001101011",
  34941=>"100100001",
  34942=>"101101010",
  34943=>"101011000",
  34944=>"010000100",
  34945=>"011101011",
  34946=>"000010101",
  34947=>"100101110",
  34948=>"100010101",
  34949=>"001001101",
  34950=>"101110110",
  34951=>"010000010",
  34952=>"100011011",
  34953=>"110110111",
  34954=>"101010101",
  34955=>"011000110",
  34956=>"011011100",
  34957=>"110110000",
  34958=>"110100000",
  34959=>"001101110",
  34960=>"000001010",
  34961=>"111001111",
  34962=>"100011001",
  34963=>"010111000",
  34964=>"000000001",
  34965=>"001100001",
  34966=>"100100011",
  34967=>"110111101",
  34968=>"101011000",
  34969=>"010011011",
  34970=>"101010001",
  34971=>"101110001",
  34972=>"100111111",
  34973=>"000010101",
  34974=>"110010010",
  34975=>"111101111",
  34976=>"110001001",
  34977=>"101111100",
  34978=>"011001100",
  34979=>"100000110",
  34980=>"101011000",
  34981=>"011110101",
  34982=>"000100101",
  34983=>"101001110",
  34984=>"000111101",
  34985=>"110000010",
  34986=>"101100000",
  34987=>"100100000",
  34988=>"010110110",
  34989=>"011110011",
  34990=>"111010011",
  34991=>"011011100",
  34992=>"101010100",
  34993=>"011101000",
  34994=>"011000101",
  34995=>"000100000",
  34996=>"000000010",
  34997=>"100011111",
  34998=>"111110100",
  34999=>"001001110",
  35000=>"101000100",
  35001=>"100010111",
  35002=>"000000111",
  35003=>"111101101",
  35004=>"001010110",
  35005=>"111111101",
  35006=>"000101110",
  35007=>"001110110",
  35008=>"101101111",
  35009=>"010011011",
  35010=>"001111101",
  35011=>"010011011",
  35012=>"100111111",
  35013=>"100011111",
  35014=>"101001001",
  35015=>"100000000",
  35016=>"010100010",
  35017=>"111001001",
  35018=>"000101010",
  35019=>"110000001",
  35020=>"010001101",
  35021=>"110101111",
  35022=>"010110111",
  35023=>"111000110",
  35024=>"011001101",
  35025=>"101111100",
  35026=>"000101010",
  35027=>"101001010",
  35028=>"110100111",
  35029=>"110111001",
  35030=>"110000000",
  35031=>"111110100",
  35032=>"100110100",
  35033=>"010010111",
  35034=>"111000011",
  35035=>"010110000",
  35036=>"001110000",
  35037=>"000001100",
  35038=>"100110011",
  35039=>"001100011",
  35040=>"110100100",
  35041=>"100001010",
  35042=>"100011001",
  35043=>"101001001",
  35044=>"010111001",
  35045=>"011101100",
  35046=>"000011110",
  35047=>"000010101",
  35048=>"010001011",
  35049=>"001110011",
  35050=>"011001001",
  35051=>"100111011",
  35052=>"111110101",
  35053=>"011011101",
  35054=>"110000101",
  35055=>"010000000",
  35056=>"001000110",
  35057=>"001000110",
  35058=>"000110001",
  35059=>"111011010",
  35060=>"111000111",
  35061=>"111001101",
  35062=>"111010000",
  35063=>"100011011",
  35064=>"111111010",
  35065=>"111000010",
  35066=>"110010010",
  35067=>"101100001",
  35068=>"001000101",
  35069=>"010010111",
  35070=>"111011110",
  35071=>"110110101",
  35072=>"100101110",
  35073=>"111110011",
  35074=>"100100010",
  35075=>"110010001",
  35076=>"001111010",
  35077=>"011011111",
  35078=>"011010011",
  35079=>"111001111",
  35080=>"110000111",
  35081=>"001011010",
  35082=>"101011001",
  35083=>"101101101",
  35084=>"011001111",
  35085=>"101110111",
  35086=>"010011001",
  35087=>"101111011",
  35088=>"010100111",
  35089=>"101111111",
  35090=>"101000110",
  35091=>"001100001",
  35092=>"110100011",
  35093=>"011101001",
  35094=>"001011010",
  35095=>"010111110",
  35096=>"000111000",
  35097=>"111100001",
  35098=>"010100111",
  35099=>"111011000",
  35100=>"000110001",
  35101=>"011100011",
  35102=>"000001110",
  35103=>"110110001",
  35104=>"101000000",
  35105=>"111011111",
  35106=>"111010000",
  35107=>"001010011",
  35108=>"100011010",
  35109=>"000000100",
  35110=>"101011111",
  35111=>"010000010",
  35112=>"110000100",
  35113=>"111010111",
  35114=>"111110001",
  35115=>"101110010",
  35116=>"011001110",
  35117=>"110010000",
  35118=>"001000001",
  35119=>"101111110",
  35120=>"010111111",
  35121=>"010111101",
  35122=>"100011110",
  35123=>"100100000",
  35124=>"111100101",
  35125=>"011110001",
  35126=>"011111110",
  35127=>"010010111",
  35128=>"001101101",
  35129=>"000110101",
  35130=>"111010100",
  35131=>"111111110",
  35132=>"111010111",
  35133=>"001001111",
  35134=>"001111000",
  35135=>"001000001",
  35136=>"010101111",
  35137=>"001100010",
  35138=>"111110000",
  35139=>"101111010",
  35140=>"000001110",
  35141=>"101111111",
  35142=>"000110110",
  35143=>"110101111",
  35144=>"111111110",
  35145=>"010001011",
  35146=>"100110000",
  35147=>"101011010",
  35148=>"100011100",
  35149=>"001010111",
  35150=>"011011101",
  35151=>"100101101",
  35152=>"111100100",
  35153=>"100100001",
  35154=>"101010100",
  35155=>"111010000",
  35156=>"001001110",
  35157=>"100111000",
  35158=>"100111000",
  35159=>"000101101",
  35160=>"111111111",
  35161=>"001100100",
  35162=>"110110011",
  35163=>"001111000",
  35164=>"010111111",
  35165=>"011000010",
  35166=>"101001001",
  35167=>"110001000",
  35168=>"010101100",
  35169=>"011010111",
  35170=>"011011111",
  35171=>"101001001",
  35172=>"010010010",
  35173=>"010100111",
  35174=>"001011000",
  35175=>"000001010",
  35176=>"011000110",
  35177=>"100100000",
  35178=>"010011010",
  35179=>"001100011",
  35180=>"001110100",
  35181=>"111011110",
  35182=>"001010011",
  35183=>"011101001",
  35184=>"010111010",
  35185=>"100001011",
  35186=>"000000101",
  35187=>"100000111",
  35188=>"001101111",
  35189=>"110010111",
  35190=>"111000110",
  35191=>"010001110",
  35192=>"101100011",
  35193=>"011001010",
  35194=>"111011111",
  35195=>"000001000",
  35196=>"000011010",
  35197=>"101010101",
  35198=>"111111100",
  35199=>"000010011",
  35200=>"101000100",
  35201=>"000011101",
  35202=>"100000000",
  35203=>"001000000",
  35204=>"000000110",
  35205=>"111110110",
  35206=>"001011010",
  35207=>"111101111",
  35208=>"010110100",
  35209=>"011000101",
  35210=>"110110101",
  35211=>"100110000",
  35212=>"000100000",
  35213=>"001010000",
  35214=>"000100001",
  35215=>"100110001",
  35216=>"110001100",
  35217=>"011010110",
  35218=>"001111111",
  35219=>"011010011",
  35220=>"110011001",
  35221=>"011011011",
  35222=>"010000000",
  35223=>"111010010",
  35224=>"001101011",
  35225=>"000100101",
  35226=>"111001111",
  35227=>"001000101",
  35228=>"111011111",
  35229=>"001110010",
  35230=>"110110011",
  35231=>"101001000",
  35232=>"001101001",
  35233=>"111001010",
  35234=>"101110100",
  35235=>"011000011",
  35236=>"001101101",
  35237=>"010001001",
  35238=>"000000011",
  35239=>"011100010",
  35240=>"110000110",
  35241=>"100000101",
  35242=>"101100010",
  35243=>"000011000",
  35244=>"100110000",
  35245=>"010011101",
  35246=>"101011011",
  35247=>"010110100",
  35248=>"111101110",
  35249=>"110011011",
  35250=>"000110101",
  35251=>"011011001",
  35252=>"011100111",
  35253=>"011011111",
  35254=>"111011001",
  35255=>"101111100",
  35256=>"001110010",
  35257=>"100001011",
  35258=>"011110111",
  35259=>"100000001",
  35260=>"101010000",
  35261=>"001111111",
  35262=>"101000010",
  35263=>"101110101",
  35264=>"111000011",
  35265=>"100001001",
  35266=>"010110110",
  35267=>"111101001",
  35268=>"011000010",
  35269=>"001101010",
  35270=>"101000100",
  35271=>"110101010",
  35272=>"010110010",
  35273=>"110100100",
  35274=>"000101010",
  35275=>"111101111",
  35276=>"010011011",
  35277=>"110011011",
  35278=>"010011001",
  35279=>"001101110",
  35280=>"111110110",
  35281=>"101001110",
  35282=>"011001100",
  35283=>"111101101",
  35284=>"011101000",
  35285=>"011010110",
  35286=>"110000001",
  35287=>"100001010",
  35288=>"100000110",
  35289=>"100000100",
  35290=>"001001010",
  35291=>"111010111",
  35292=>"010001000",
  35293=>"101101111",
  35294=>"010110010",
  35295=>"111010010",
  35296=>"101000101",
  35297=>"011000111",
  35298=>"100110101",
  35299=>"001100100",
  35300=>"100011010",
  35301=>"101100001",
  35302=>"010100111",
  35303=>"100000001",
  35304=>"001001000",
  35305=>"010010010",
  35306=>"100011011",
  35307=>"110101011",
  35308=>"111100100",
  35309=>"110001010",
  35310=>"101011001",
  35311=>"001001110",
  35312=>"001110110",
  35313=>"001011001",
  35314=>"111100011",
  35315=>"000000110",
  35316=>"000011001",
  35317=>"000010100",
  35318=>"001111000",
  35319=>"100001110",
  35320=>"100110110",
  35321=>"011011111",
  35322=>"111001000",
  35323=>"011010111",
  35324=>"100011010",
  35325=>"101100111",
  35326=>"100111101",
  35327=>"110010111",
  35328=>"010001000",
  35329=>"100111011",
  35330=>"000101010",
  35331=>"001101100",
  35332=>"011101101",
  35333=>"100111110",
  35334=>"011111100",
  35335=>"111100011",
  35336=>"011100111",
  35337=>"111110110",
  35338=>"000010101",
  35339=>"010110000",
  35340=>"010001001",
  35341=>"100111000",
  35342=>"101010100",
  35343=>"101110011",
  35344=>"011100001",
  35345=>"101110001",
  35346=>"100101001",
  35347=>"001010100",
  35348=>"000001001",
  35349=>"101000111",
  35350=>"101110010",
  35351=>"000101010",
  35352=>"101111011",
  35353=>"110111110",
  35354=>"011000110",
  35355=>"111110001",
  35356=>"111100011",
  35357=>"010100000",
  35358=>"001101110",
  35359=>"101101010",
  35360=>"111001111",
  35361=>"101010010",
  35362=>"111100010",
  35363=>"101011101",
  35364=>"011110110",
  35365=>"111100100",
  35366=>"010010010",
  35367=>"010000011",
  35368=>"001001010",
  35369=>"010110001",
  35370=>"000110001",
  35371=>"101000010",
  35372=>"111101010",
  35373=>"101010100",
  35374=>"111001101",
  35375=>"111000100",
  35376=>"010101010",
  35377=>"101010101",
  35378=>"100001101",
  35379=>"000101000",
  35380=>"111010110",
  35381=>"000110011",
  35382=>"011111110",
  35383=>"111110111",
  35384=>"101000000",
  35385=>"100110101",
  35386=>"011110001",
  35387=>"010010011",
  35388=>"100001010",
  35389=>"000000101",
  35390=>"100110101",
  35391=>"101100100",
  35392=>"110101111",
  35393=>"011000011",
  35394=>"000000101",
  35395=>"111001110",
  35396=>"101110111",
  35397=>"001110111",
  35398=>"001101111",
  35399=>"101100111",
  35400=>"011010111",
  35401=>"111010111",
  35402=>"110111011",
  35403=>"001111110",
  35404=>"101011011",
  35405=>"010000100",
  35406=>"101000101",
  35407=>"010111100",
  35408=>"000111111",
  35409=>"110001001",
  35410=>"000100001",
  35411=>"111010011",
  35412=>"000101000",
  35413=>"100110100",
  35414=>"110100011",
  35415=>"101011001",
  35416=>"111100111",
  35417=>"011000111",
  35418=>"111111010",
  35419=>"001011010",
  35420=>"001110101",
  35421=>"101100011",
  35422=>"101000010",
  35423=>"011010011",
  35424=>"100001011",
  35425=>"010010010",
  35426=>"100110100",
  35427=>"111101011",
  35428=>"101111101",
  35429=>"001001101",
  35430=>"111110111",
  35431=>"111010111",
  35432=>"011000001",
  35433=>"001111010",
  35434=>"111001001",
  35435=>"011011000",
  35436=>"111111001",
  35437=>"110000000",
  35438=>"010001001",
  35439=>"011010100",
  35440=>"101000101",
  35441=>"110011000",
  35442=>"011110000",
  35443=>"110010101",
  35444=>"110011111",
  35445=>"000010100",
  35446=>"110110111",
  35447=>"111111101",
  35448=>"110101000",
  35449=>"111111101",
  35450=>"110011001",
  35451=>"111001101",
  35452=>"000101110",
  35453=>"101001000",
  35454=>"011011110",
  35455=>"100111110",
  35456=>"011100110",
  35457=>"001111110",
  35458=>"001000100",
  35459=>"100111010",
  35460=>"101011100",
  35461=>"011010000",
  35462=>"101011001",
  35463=>"010000000",
  35464=>"000110010",
  35465=>"001011111",
  35466=>"101000111",
  35467=>"001001110",
  35468=>"100000010",
  35469=>"010110000",
  35470=>"110010001",
  35471=>"111001001",
  35472=>"010010010",
  35473=>"100110000",
  35474=>"000001100",
  35475=>"100001001",
  35476=>"110000000",
  35477=>"111101101",
  35478=>"001111010",
  35479=>"001101001",
  35480=>"110001101",
  35481=>"011000101",
  35482=>"100101100",
  35483=>"001000000",
  35484=>"000110111",
  35485=>"110010100",
  35486=>"001010110",
  35487=>"100111001",
  35488=>"010010000",
  35489=>"100001000",
  35490=>"000001111",
  35491=>"110001111",
  35492=>"101001110",
  35493=>"001100111",
  35494=>"001101001",
  35495=>"101000010",
  35496=>"000010001",
  35497=>"110101001",
  35498=>"100101111",
  35499=>"110001001",
  35500=>"100001100",
  35501=>"100000110",
  35502=>"011011111",
  35503=>"101101111",
  35504=>"000001011",
  35505=>"101110011",
  35506=>"100111011",
  35507=>"100101011",
  35508=>"100000101",
  35509=>"001101010",
  35510=>"000110001",
  35511=>"011101000",
  35512=>"100100000",
  35513=>"110110010",
  35514=>"011010010",
  35515=>"000000001",
  35516=>"111010001",
  35517=>"101010011",
  35518=>"100000011",
  35519=>"100101101",
  35520=>"110111000",
  35521=>"101001000",
  35522=>"110100101",
  35523=>"011001101",
  35524=>"011001000",
  35525=>"011001101",
  35526=>"011110111",
  35527=>"110010111",
  35528=>"111000111",
  35529=>"101001110",
  35530=>"000000000",
  35531=>"100000000",
  35532=>"001111110",
  35533=>"010010001",
  35534=>"100000000",
  35535=>"001011110",
  35536=>"110101111",
  35537=>"001000000",
  35538=>"101011110",
  35539=>"111101010",
  35540=>"111100000",
  35541=>"111001110",
  35542=>"000001010",
  35543=>"110011000",
  35544=>"000101111",
  35545=>"101010010",
  35546=>"000010101",
  35547=>"000101110",
  35548=>"111100001",
  35549=>"001011001",
  35550=>"111010010",
  35551=>"011011001",
  35552=>"000011001",
  35553=>"010001000",
  35554=>"011110111",
  35555=>"111101111",
  35556=>"011010010",
  35557=>"011001100",
  35558=>"000010010",
  35559=>"010111000",
  35560=>"101010111",
  35561=>"110010010",
  35562=>"001010000",
  35563=>"110011000",
  35564=>"000011001",
  35565=>"100101101",
  35566=>"011011100",
  35567=>"001000010",
  35568=>"000011011",
  35569=>"110011000",
  35570=>"100000010",
  35571=>"111100110",
  35572=>"100011011",
  35573=>"110110001",
  35574=>"100110000",
  35575=>"101110001",
  35576=>"100101010",
  35577=>"010101111",
  35578=>"000101001",
  35579=>"101000100",
  35580=>"100000000",
  35581=>"010001110",
  35582=>"000010111",
  35583=>"101001000",
  35584=>"010000110",
  35585=>"100111000",
  35586=>"110010010",
  35587=>"001001010",
  35588=>"010011111",
  35589=>"111001011",
  35590=>"101101101",
  35591=>"000110011",
  35592=>"110101000",
  35593=>"101111010",
  35594=>"110101000",
  35595=>"001010001",
  35596=>"010011000",
  35597=>"000001011",
  35598=>"011001011",
  35599=>"100000011",
  35600=>"100001011",
  35601=>"101101010",
  35602=>"001011100",
  35603=>"111111100",
  35604=>"001001010",
  35605=>"110101101",
  35606=>"010010001",
  35607=>"101110100",
  35608=>"101001001",
  35609=>"010110001",
  35610=>"000000001",
  35611=>"010000001",
  35612=>"111101101",
  35613=>"101100100",
  35614=>"110111100",
  35615=>"000100111",
  35616=>"011001110",
  35617=>"111000011",
  35618=>"101000000",
  35619=>"111000101",
  35620=>"101000101",
  35621=>"000001110",
  35622=>"000110100",
  35623=>"101110111",
  35624=>"011110010",
  35625=>"101011001",
  35626=>"010110000",
  35627=>"000100101",
  35628=>"001011001",
  35629=>"000011010",
  35630=>"111100011",
  35631=>"001010111",
  35632=>"100001011",
  35633=>"110000001",
  35634=>"000011011",
  35635=>"110010011",
  35636=>"010110101",
  35637=>"011001110",
  35638=>"110010011",
  35639=>"000001110",
  35640=>"111010001",
  35641=>"111001101",
  35642=>"111100110",
  35643=>"110011001",
  35644=>"101100011",
  35645=>"010000000",
  35646=>"010010111",
  35647=>"001110101",
  35648=>"010111000",
  35649=>"000001000",
  35650=>"010010011",
  35651=>"100111101",
  35652=>"101110101",
  35653=>"101110110",
  35654=>"100101110",
  35655=>"101101111",
  35656=>"111001100",
  35657=>"010011000",
  35658=>"111000001",
  35659=>"010000111",
  35660=>"101011111",
  35661=>"100101000",
  35662=>"111000001",
  35663=>"000010101",
  35664=>"011010000",
  35665=>"011110001",
  35666=>"001001111",
  35667=>"101101000",
  35668=>"100000111",
  35669=>"001110111",
  35670=>"000001011",
  35671=>"111100001",
  35672=>"001101100",
  35673=>"100011101",
  35674=>"001000011",
  35675=>"000000101",
  35676=>"001001001",
  35677=>"000010011",
  35678=>"010000001",
  35679=>"001100111",
  35680=>"111010011",
  35681=>"110000101",
  35682=>"011001110",
  35683=>"111111000",
  35684=>"010111010",
  35685=>"111000000",
  35686=>"010101111",
  35687=>"110111100",
  35688=>"110110101",
  35689=>"011110000",
  35690=>"001010010",
  35691=>"011101000",
  35692=>"000001000",
  35693=>"111000111",
  35694=>"000011100",
  35695=>"101111010",
  35696=>"111111111",
  35697=>"101011011",
  35698=>"011000111",
  35699=>"111111101",
  35700=>"110111110",
  35701=>"000111100",
  35702=>"000010001",
  35703=>"110110100",
  35704=>"011101110",
  35705=>"101101110",
  35706=>"001100011",
  35707=>"010101111",
  35708=>"111100000",
  35709=>"101000000",
  35710=>"101000001",
  35711=>"111001011",
  35712=>"001000000",
  35713=>"110000011",
  35714=>"000011101",
  35715=>"001011000",
  35716=>"010001110",
  35717=>"000000011",
  35718=>"000100100",
  35719=>"110110000",
  35720=>"100001010",
  35721=>"010111110",
  35722=>"111101101",
  35723=>"101010011",
  35724=>"000010111",
  35725=>"101100111",
  35726=>"011101101",
  35727=>"010101111",
  35728=>"101100100",
  35729=>"110101001",
  35730=>"111101011",
  35731=>"110001010",
  35732=>"011000101",
  35733=>"000100111",
  35734=>"000011001",
  35735=>"101100000",
  35736=>"011100001",
  35737=>"111111111",
  35738=>"001111010",
  35739=>"101011011",
  35740=>"011110000",
  35741=>"000100000",
  35742=>"001101000",
  35743=>"101111001",
  35744=>"010100110",
  35745=>"000001011",
  35746=>"100010001",
  35747=>"000100100",
  35748=>"111000000",
  35749=>"000100110",
  35750=>"100001011",
  35751=>"010010011",
  35752=>"011100000",
  35753=>"000000000",
  35754=>"110101100",
  35755=>"011011101",
  35756=>"001110001",
  35757=>"010111001",
  35758=>"100111010",
  35759=>"010011001",
  35760=>"011110100",
  35761=>"110100100",
  35762=>"111100001",
  35763=>"000100000",
  35764=>"101110001",
  35765=>"110101111",
  35766=>"100110000",
  35767=>"011101101",
  35768=>"100101111",
  35769=>"101100101",
  35770=>"101010001",
  35771=>"100110111",
  35772=>"111100011",
  35773=>"011011101",
  35774=>"000000010",
  35775=>"101100010",
  35776=>"010101000",
  35777=>"000110111",
  35778=>"100001110",
  35779=>"111011010",
  35780=>"110101110",
  35781=>"010111011",
  35782=>"110010110",
  35783=>"001101001",
  35784=>"100000010",
  35785=>"000111000",
  35786=>"001011011",
  35787=>"110110011",
  35788=>"101101001",
  35789=>"100000100",
  35790=>"000010101",
  35791=>"111101000",
  35792=>"100001000",
  35793=>"110101011",
  35794=>"001000101",
  35795=>"011000000",
  35796=>"000000000",
  35797=>"110011010",
  35798=>"011010101",
  35799=>"111110001",
  35800=>"010011010",
  35801=>"010101001",
  35802=>"100001001",
  35803=>"000010111",
  35804=>"001100001",
  35805=>"010111111",
  35806=>"101011000",
  35807=>"111001010",
  35808=>"100111000",
  35809=>"100010100",
  35810=>"111100010",
  35811=>"110101011",
  35812=>"000110100",
  35813=>"110011100",
  35814=>"011110101",
  35815=>"011011000",
  35816=>"010010110",
  35817=>"111111100",
  35818=>"001110111",
  35819=>"011100010",
  35820=>"111011100",
  35821=>"101101000",
  35822=>"111001111",
  35823=>"001010001",
  35824=>"110010101",
  35825=>"011101001",
  35826=>"001000110",
  35827=>"110010111",
  35828=>"110100101",
  35829=>"011010001",
  35830=>"000011111",
  35831=>"101100111",
  35832=>"101011101",
  35833=>"111111110",
  35834=>"111000110",
  35835=>"100000100",
  35836=>"111111001",
  35837=>"010001010",
  35838=>"000100110",
  35839=>"011111001",
  35840=>"011011000",
  35841=>"000010110",
  35842=>"011101011",
  35843=>"100011010",
  35844=>"001101111",
  35845=>"100001010",
  35846=>"001110100",
  35847=>"100010100",
  35848=>"001001001",
  35849=>"111111011",
  35850=>"111000001",
  35851=>"001010011",
  35852=>"001010100",
  35853=>"100001000",
  35854=>"011001100",
  35855=>"011011101",
  35856=>"001110100",
  35857=>"000110010",
  35858=>"111101001",
  35859=>"001111001",
  35860=>"001111000",
  35861=>"010111011",
  35862=>"010111011",
  35863=>"010100110",
  35864=>"011100000",
  35865=>"011001111",
  35866=>"100101101",
  35867=>"010100010",
  35868=>"101001001",
  35869=>"111101111",
  35870=>"010001101",
  35871=>"111001111",
  35872=>"110111001",
  35873=>"100100011",
  35874=>"111101101",
  35875=>"101000011",
  35876=>"000110010",
  35877=>"110110111",
  35878=>"001100000",
  35879=>"010010000",
  35880=>"010110101",
  35881=>"000100100",
  35882=>"000111110",
  35883=>"011101111",
  35884=>"001010110",
  35885=>"010011110",
  35886=>"001101111",
  35887=>"110000010",
  35888=>"001001111",
  35889=>"000000001",
  35890=>"010101001",
  35891=>"010011000",
  35892=>"111110100",
  35893=>"011111010",
  35894=>"111110001",
  35895=>"101101111",
  35896=>"110010101",
  35897=>"110100100",
  35898=>"100100111",
  35899=>"011100011",
  35900=>"000001110",
  35901=>"000001001",
  35902=>"111001000",
  35903=>"001000110",
  35904=>"010001100",
  35905=>"110100111",
  35906=>"101010101",
  35907=>"011010111",
  35908=>"110101100",
  35909=>"011101111",
  35910=>"111110100",
  35911=>"111000111",
  35912=>"111111010",
  35913=>"001000110",
  35914=>"100100100",
  35915=>"011100111",
  35916=>"010001001",
  35917=>"101110000",
  35918=>"001000100",
  35919=>"011101000",
  35920=>"000110111",
  35921=>"100000111",
  35922=>"011011010",
  35923=>"110110010",
  35924=>"100000110",
  35925=>"111010110",
  35926=>"011010010",
  35927=>"010111100",
  35928=>"110001010",
  35929=>"100111011",
  35930=>"100110010",
  35931=>"000001110",
  35932=>"011010001",
  35933=>"111000101",
  35934=>"011010000",
  35935=>"010010001",
  35936=>"010000100",
  35937=>"101110011",
  35938=>"101101001",
  35939=>"011001000",
  35940=>"001101100",
  35941=>"101000010",
  35942=>"101000000",
  35943=>"011001001",
  35944=>"010000000",
  35945=>"111001111",
  35946=>"000001100",
  35947=>"100100101",
  35948=>"010101000",
  35949=>"001100010",
  35950=>"001000111",
  35951=>"111110110",
  35952=>"000000000",
  35953=>"001111111",
  35954=>"101100110",
  35955=>"111001100",
  35956=>"010010011",
  35957=>"110101111",
  35958=>"011011011",
  35959=>"111011001",
  35960=>"010101011",
  35961=>"110001000",
  35962=>"010010010",
  35963=>"110000101",
  35964=>"001011101",
  35965=>"100011011",
  35966=>"010000000",
  35967=>"000000110",
  35968=>"000010010",
  35969=>"111101001",
  35970=>"000110101",
  35971=>"000000010",
  35972=>"000010011",
  35973=>"101010000",
  35974=>"110110101",
  35975=>"011011001",
  35976=>"100011110",
  35977=>"000001101",
  35978=>"011101001",
  35979=>"001110011",
  35980=>"111110001",
  35981=>"101101101",
  35982=>"010010011",
  35983=>"010010110",
  35984=>"011011100",
  35985=>"100011011",
  35986=>"110010001",
  35987=>"111101101",
  35988=>"100110011",
  35989=>"101010100",
  35990=>"100010010",
  35991=>"000101110",
  35992=>"010011101",
  35993=>"111101101",
  35994=>"010011111",
  35995=>"100000000",
  35996=>"000110011",
  35997=>"011111010",
  35998=>"111000111",
  35999=>"100011000",
  36000=>"011110111",
  36001=>"011111111",
  36002=>"110101100",
  36003=>"010011011",
  36004=>"011011000",
  36005=>"000110111",
  36006=>"000110100",
  36007=>"101001010",
  36008=>"101000010",
  36009=>"111100110",
  36010=>"110010101",
  36011=>"111101100",
  36012=>"111101011",
  36013=>"110110111",
  36014=>"011000111",
  36015=>"110101000",
  36016=>"010111001",
  36017=>"000000100",
  36018=>"001010001",
  36019=>"011001010",
  36020=>"000110011",
  36021=>"110000101",
  36022=>"100000010",
  36023=>"000000101",
  36024=>"011111111",
  36025=>"011000110",
  36026=>"110000001",
  36027=>"110010001",
  36028=>"000101000",
  36029=>"111011111",
  36030=>"010101001",
  36031=>"010111000",
  36032=>"111110011",
  36033=>"011001000",
  36034=>"010111011",
  36035=>"101111000",
  36036=>"000001000",
  36037=>"101110000",
  36038=>"001100001",
  36039=>"000111110",
  36040=>"110001101",
  36041=>"001101001",
  36042=>"001100000",
  36043=>"001110011",
  36044=>"111010001",
  36045=>"111100101",
  36046=>"000110010",
  36047=>"010010100",
  36048=>"101000010",
  36049=>"000011111",
  36050=>"111001100",
  36051=>"000001101",
  36052=>"111011101",
  36053=>"110010001",
  36054=>"110010100",
  36055=>"111010101",
  36056=>"111000010",
  36057=>"110010001",
  36058=>"010101111",
  36059=>"011101001",
  36060=>"001011010",
  36061=>"000010011",
  36062=>"100011000",
  36063=>"101101001",
  36064=>"000010010",
  36065=>"011110001",
  36066=>"011011101",
  36067=>"110000110",
  36068=>"011001000",
  36069=>"001000111",
  36070=>"011011011",
  36071=>"100010101",
  36072=>"001110111",
  36073=>"000010110",
  36074=>"100110010",
  36075=>"010001000",
  36076=>"000001100",
  36077=>"100010110",
  36078=>"000001000",
  36079=>"100011001",
  36080=>"010111110",
  36081=>"001000101",
  36082=>"010001101",
  36083=>"111111101",
  36084=>"101111110",
  36085=>"101011100",
  36086=>"100111000",
  36087=>"101110110",
  36088=>"100100001",
  36089=>"110110000",
  36090=>"000101101",
  36091=>"010100010",
  36092=>"000011011",
  36093=>"010101011",
  36094=>"000001010",
  36095=>"101011111",
  36096=>"100110111",
  36097=>"010001001",
  36098=>"011001010",
  36099=>"011110001",
  36100=>"110010101",
  36101=>"001001010",
  36102=>"111010010",
  36103=>"010100010",
  36104=>"100010001",
  36105=>"100110101",
  36106=>"000000101",
  36107=>"100101001",
  36108=>"000001101",
  36109=>"111101000",
  36110=>"000011011",
  36111=>"001100010",
  36112=>"011110101",
  36113=>"111101101",
  36114=>"111011010",
  36115=>"110101101",
  36116=>"101000010",
  36117=>"010000111",
  36118=>"100010110",
  36119=>"001100111",
  36120=>"010010001",
  36121=>"011111010",
  36122=>"000110001",
  36123=>"100001011",
  36124=>"111011010",
  36125=>"110001000",
  36126=>"111001010",
  36127=>"011100000",
  36128=>"000111100",
  36129=>"101000101",
  36130=>"110110101",
  36131=>"011001011",
  36132=>"011100000",
  36133=>"000001010",
  36134=>"000010110",
  36135=>"100111000",
  36136=>"000000001",
  36137=>"011100001",
  36138=>"101001010",
  36139=>"010011100",
  36140=>"011011111",
  36141=>"110111010",
  36142=>"001001011",
  36143=>"101010110",
  36144=>"001000100",
  36145=>"100100101",
  36146=>"101000001",
  36147=>"001110101",
  36148=>"101010010",
  36149=>"000001010",
  36150=>"011011110",
  36151=>"010110010",
  36152=>"000101010",
  36153=>"011000000",
  36154=>"100101011",
  36155=>"101011000",
  36156=>"000000000",
  36157=>"111101101",
  36158=>"100101100",
  36159=>"010110111",
  36160=>"010011100",
  36161=>"100001000",
  36162=>"101111100",
  36163=>"000000011",
  36164=>"010000111",
  36165=>"011110001",
  36166=>"000000001",
  36167=>"100111100",
  36168=>"001100110",
  36169=>"100100010",
  36170=>"111010111",
  36171=>"001000100",
  36172=>"000111110",
  36173=>"011000101",
  36174=>"011010011",
  36175=>"111010010",
  36176=>"101111111",
  36177=>"011001100",
  36178=>"100101001",
  36179=>"000101101",
  36180=>"000100101",
  36181=>"001101111",
  36182=>"001010000",
  36183=>"111111010",
  36184=>"000001001",
  36185=>"011001101",
  36186=>"101001111",
  36187=>"010000001",
  36188=>"111101111",
  36189=>"110110111",
  36190=>"010100001",
  36191=>"100100101",
  36192=>"000011010",
  36193=>"111010011",
  36194=>"000010011",
  36195=>"001100100",
  36196=>"010001001",
  36197=>"110101101",
  36198=>"000110100",
  36199=>"111001111",
  36200=>"000101011",
  36201=>"001100101",
  36202=>"100000000",
  36203=>"111111101",
  36204=>"111101010",
  36205=>"101101111",
  36206=>"110111100",
  36207=>"000000010",
  36208=>"000000011",
  36209=>"111110100",
  36210=>"111100101",
  36211=>"011010000",
  36212=>"100111000",
  36213=>"101100111",
  36214=>"111110011",
  36215=>"000001110",
  36216=>"100111011",
  36217=>"100011100",
  36218=>"111110110",
  36219=>"001011111",
  36220=>"000110000",
  36221=>"101001011",
  36222=>"010111000",
  36223=>"011111011",
  36224=>"010110111",
  36225=>"010001001",
  36226=>"111110110",
  36227=>"110100101",
  36228=>"011111111",
  36229=>"010001101",
  36230=>"110110000",
  36231=>"100100001",
  36232=>"000101000",
  36233=>"000111011",
  36234=>"010101010",
  36235=>"111110110",
  36236=>"010101110",
  36237=>"010001010",
  36238=>"011000011",
  36239=>"011101011",
  36240=>"010100111",
  36241=>"110100000",
  36242=>"101111010",
  36243=>"101101101",
  36244=>"111111011",
  36245=>"000111100",
  36246=>"111011000",
  36247=>"100110001",
  36248=>"110110100",
  36249=>"000000000",
  36250=>"100111011",
  36251=>"011110000",
  36252=>"100100111",
  36253=>"111010111",
  36254=>"110111101",
  36255=>"011000000",
  36256=>"000101111",
  36257=>"100111110",
  36258=>"110000001",
  36259=>"011100101",
  36260=>"100011010",
  36261=>"011010000",
  36262=>"111001011",
  36263=>"010000010",
  36264=>"001011111",
  36265=>"001110000",
  36266=>"000001010",
  36267=>"000110110",
  36268=>"111111110",
  36269=>"100101101",
  36270=>"100010011",
  36271=>"101011100",
  36272=>"111001000",
  36273=>"110110110",
  36274=>"011111110",
  36275=>"100001000",
  36276=>"110010001",
  36277=>"101001110",
  36278=>"100101100",
  36279=>"100000011",
  36280=>"111001101",
  36281=>"001110100",
  36282=>"001000101",
  36283=>"100011100",
  36284=>"001010001",
  36285=>"010100010",
  36286=>"111010000",
  36287=>"000111110",
  36288=>"110000110",
  36289=>"000110101",
  36290=>"111110011",
  36291=>"101101011",
  36292=>"011101001",
  36293=>"011100100",
  36294=>"101000011",
  36295=>"110100011",
  36296=>"011011011",
  36297=>"101110100",
  36298=>"100001100",
  36299=>"001101111",
  36300=>"001001110",
  36301=>"000001000",
  36302=>"000001000",
  36303=>"011100101",
  36304=>"001101010",
  36305=>"010001110",
  36306=>"000000000",
  36307=>"011010000",
  36308=>"110101000",
  36309=>"001000000",
  36310=>"100010110",
  36311=>"111001011",
  36312=>"000101100",
  36313=>"110111111",
  36314=>"101100100",
  36315=>"110101110",
  36316=>"001110111",
  36317=>"100111111",
  36318=>"110000010",
  36319=>"010001111",
  36320=>"000010010",
  36321=>"100000100",
  36322=>"010110100",
  36323=>"111000101",
  36324=>"111001010",
  36325=>"010110001",
  36326=>"000010000",
  36327=>"000011110",
  36328=>"101111001",
  36329=>"011010010",
  36330=>"001001101",
  36331=>"100111000",
  36332=>"011010111",
  36333=>"011101100",
  36334=>"100010100",
  36335=>"001010010",
  36336=>"110110100",
  36337=>"101100001",
  36338=>"101101101",
  36339=>"000101111",
  36340=>"101010110",
  36341=>"100101000",
  36342=>"001100100",
  36343=>"010111110",
  36344=>"001101000",
  36345=>"111011000",
  36346=>"110101101",
  36347=>"010101110",
  36348=>"100111010",
  36349=>"111000000",
  36350=>"000110000",
  36351=>"100111001",
  36352=>"111010111",
  36353=>"011110011",
  36354=>"110010000",
  36355=>"001100100",
  36356=>"101101010",
  36357=>"010000101",
  36358=>"010101011",
  36359=>"000000011",
  36360=>"111010111",
  36361=>"001010000",
  36362=>"100111101",
  36363=>"001100001",
  36364=>"111100001",
  36365=>"101100011",
  36366=>"101100000",
  36367=>"101100000",
  36368=>"101110100",
  36369=>"110101100",
  36370=>"000001001",
  36371=>"110110101",
  36372=>"100001010",
  36373=>"000000111",
  36374=>"001011000",
  36375=>"001000100",
  36376=>"100110101",
  36377=>"111011011",
  36378=>"111000000",
  36379=>"000111111",
  36380=>"001011010",
  36381=>"100010100",
  36382=>"100100011",
  36383=>"001011011",
  36384=>"110010100",
  36385=>"111000100",
  36386=>"101100111",
  36387=>"011100010",
  36388=>"101000011",
  36389=>"001000000",
  36390=>"101111010",
  36391=>"000010100",
  36392=>"000110001",
  36393=>"111110110",
  36394=>"001111001",
  36395=>"100000000",
  36396=>"110100000",
  36397=>"000000001",
  36398=>"000101110",
  36399=>"000001010",
  36400=>"100001100",
  36401=>"100000101",
  36402=>"011001100",
  36403=>"110100001",
  36404=>"011001010",
  36405=>"100011000",
  36406=>"111000001",
  36407=>"001110001",
  36408=>"000001100",
  36409=>"111110111",
  36410=>"110011111",
  36411=>"001010110",
  36412=>"001110011",
  36413=>"010010010",
  36414=>"001011100",
  36415=>"110101111",
  36416=>"110100010",
  36417=>"001000101",
  36418=>"101010011",
  36419=>"011001101",
  36420=>"000000100",
  36421=>"001101101",
  36422=>"011000001",
  36423=>"100100001",
  36424=>"001100000",
  36425=>"010000011",
  36426=>"010100101",
  36427=>"000110110",
  36428=>"100110010",
  36429=>"111001110",
  36430=>"100000100",
  36431=>"101101000",
  36432=>"000100110",
  36433=>"011000001",
  36434=>"110110000",
  36435=>"010101011",
  36436=>"001000010",
  36437=>"011001100",
  36438=>"011001111",
  36439=>"110101101",
  36440=>"100000010",
  36441=>"000100100",
  36442=>"010010010",
  36443=>"100000000",
  36444=>"000100000",
  36445=>"010100101",
  36446=>"011111101",
  36447=>"110101100",
  36448=>"011001011",
  36449=>"010011100",
  36450=>"001010000",
  36451=>"100000100",
  36452=>"011000100",
  36453=>"101000010",
  36454=>"101111001",
  36455=>"000011101",
  36456=>"010100111",
  36457=>"010000100",
  36458=>"101001101",
  36459=>"001000000",
  36460=>"100011100",
  36461=>"001011011",
  36462=>"000110111",
  36463=>"000101100",
  36464=>"000100010",
  36465=>"001100011",
  36466=>"001100010",
  36467=>"101111010",
  36468=>"100100100",
  36469=>"001010100",
  36470=>"010001000",
  36471=>"010000101",
  36472=>"011100001",
  36473=>"100001010",
  36474=>"100000010",
  36475=>"001011101",
  36476=>"111111111",
  36477=>"101111000",
  36478=>"011101000",
  36479=>"111111110",
  36480=>"001001011",
  36481=>"110101111",
  36482=>"000110011",
  36483=>"001010000",
  36484=>"001111011",
  36485=>"100111101",
  36486=>"101110100",
  36487=>"100101000",
  36488=>"110001101",
  36489=>"010011010",
  36490=>"000111100",
  36491=>"011100011",
  36492=>"101011101",
  36493=>"000110000",
  36494=>"001101000",
  36495=>"100000011",
  36496=>"111100111",
  36497=>"001111000",
  36498=>"100101110",
  36499=>"111111101",
  36500=>"100001000",
  36501=>"010001101",
  36502=>"110010001",
  36503=>"000011000",
  36504=>"010011000",
  36505=>"001111000",
  36506=>"001011111",
  36507=>"011010111",
  36508=>"000011100",
  36509=>"000111001",
  36510=>"111000101",
  36511=>"111000011",
  36512=>"111110011",
  36513=>"010100000",
  36514=>"110011111",
  36515=>"100011001",
  36516=>"000011101",
  36517=>"010100011",
  36518=>"110010100",
  36519=>"100101010",
  36520=>"111101000",
  36521=>"001101000",
  36522=>"100001110",
  36523=>"111010011",
  36524=>"110110100",
  36525=>"111010100",
  36526=>"010000011",
  36527=>"011010010",
  36528=>"011101101",
  36529=>"111011110",
  36530=>"110110111",
  36531=>"110001000",
  36532=>"100111101",
  36533=>"111110101",
  36534=>"111111110",
  36535=>"110110100",
  36536=>"111001110",
  36537=>"110100011",
  36538=>"110101001",
  36539=>"001111010",
  36540=>"010111100",
  36541=>"000101000",
  36542=>"000110110",
  36543=>"000001110",
  36544=>"000011001",
  36545=>"011010111",
  36546=>"100101111",
  36547=>"100101010",
  36548=>"001000101",
  36549=>"010010100",
  36550=>"010101011",
  36551=>"000100001",
  36552=>"100001000",
  36553=>"000101001",
  36554=>"101010000",
  36555=>"111010011",
  36556=>"010000011",
  36557=>"100111001",
  36558=>"001101010",
  36559=>"101011011",
  36560=>"101001000",
  36561=>"011100101",
  36562=>"110101100",
  36563=>"110110110",
  36564=>"110000000",
  36565=>"110001001",
  36566=>"011100100",
  36567=>"110001010",
  36568=>"000100111",
  36569=>"100101010",
  36570=>"100101010",
  36571=>"101110001",
  36572=>"000110011",
  36573=>"100111000",
  36574=>"110100001",
  36575=>"111110000",
  36576=>"001001101",
  36577=>"100000001",
  36578=>"110001011",
  36579=>"011010011",
  36580=>"011010110",
  36581=>"110001100",
  36582=>"110110101",
  36583=>"110000001",
  36584=>"010000101",
  36585=>"110101101",
  36586=>"000101010",
  36587=>"110000111",
  36588=>"011101000",
  36589=>"100101111",
  36590=>"100111001",
  36591=>"010001000",
  36592=>"101001001",
  36593=>"001111000",
  36594=>"110110000",
  36595=>"001101101",
  36596=>"010011111",
  36597=>"110111001",
  36598=>"111011101",
  36599=>"010001111",
  36600=>"100010011",
  36601=>"000111011",
  36602=>"001101000",
  36603=>"101010100",
  36604=>"011010000",
  36605=>"111011111",
  36606=>"011100010",
  36607=>"010001100",
  36608=>"111101100",
  36609=>"001111110",
  36610=>"010000010",
  36611=>"001101010",
  36612=>"011110111",
  36613=>"011010111",
  36614=>"101011011",
  36615=>"111011111",
  36616=>"110101011",
  36617=>"001000111",
  36618=>"101101101",
  36619=>"010111000",
  36620=>"111100011",
  36621=>"011001111",
  36622=>"110011101",
  36623=>"100100101",
  36624=>"100111110",
  36625=>"111100010",
  36626=>"001011100",
  36627=>"110011110",
  36628=>"000111100",
  36629=>"011000111",
  36630=>"100110000",
  36631=>"101100001",
  36632=>"110010010",
  36633=>"011000000",
  36634=>"100110111",
  36635=>"101111110",
  36636=>"110001100",
  36637=>"110101001",
  36638=>"100101111",
  36639=>"010000000",
  36640=>"000001100",
  36641=>"010101000",
  36642=>"111000001",
  36643=>"110011101",
  36644=>"110111100",
  36645=>"111100111",
  36646=>"000111001",
  36647=>"111100011",
  36648=>"010100000",
  36649=>"101000000",
  36650=>"010111110",
  36651=>"110111100",
  36652=>"110001011",
  36653=>"000000001",
  36654=>"010010001",
  36655=>"010011000",
  36656=>"000100110",
  36657=>"001101010",
  36658=>"000010000",
  36659=>"110001010",
  36660=>"110010111",
  36661=>"111101000",
  36662=>"100000110",
  36663=>"010010010",
  36664=>"110101110",
  36665=>"000001101",
  36666=>"000010100",
  36667=>"110011001",
  36668=>"101010000",
  36669=>"100101000",
  36670=>"110110011",
  36671=>"110111111",
  36672=>"101101111",
  36673=>"100110011",
  36674=>"101011100",
  36675=>"010110000",
  36676=>"000111011",
  36677=>"000010100",
  36678=>"001101100",
  36679=>"011111011",
  36680=>"000101011",
  36681=>"100010001",
  36682=>"001011101",
  36683=>"101011110",
  36684=>"101000101",
  36685=>"010010000",
  36686=>"000011101",
  36687=>"010011001",
  36688=>"001000000",
  36689=>"100110010",
  36690=>"100000111",
  36691=>"000000100",
  36692=>"101000010",
  36693=>"101100111",
  36694=>"011101100",
  36695=>"000000001",
  36696=>"101100100",
  36697=>"101101011",
  36698=>"010010100",
  36699=>"110001011",
  36700=>"011001000",
  36701=>"111001011",
  36702=>"001110110",
  36703=>"000001000",
  36704=>"111011001",
  36705=>"011100111",
  36706=>"001001111",
  36707=>"110001011",
  36708=>"101100000",
  36709=>"100001011",
  36710=>"010010111",
  36711=>"000110011",
  36712=>"110000000",
  36713=>"100110111",
  36714=>"001101111",
  36715=>"110100100",
  36716=>"110011101",
  36717=>"001001010",
  36718=>"001100000",
  36719=>"011111100",
  36720=>"001101110",
  36721=>"010001011",
  36722=>"010101100",
  36723=>"101101100",
  36724=>"011111101",
  36725=>"001011011",
  36726=>"010000101",
  36727=>"110101101",
  36728=>"101110100",
  36729=>"001000101",
  36730=>"101110111",
  36731=>"011000001",
  36732=>"000010010",
  36733=>"111101000",
  36734=>"110001000",
  36735=>"000011111",
  36736=>"010101000",
  36737=>"010011010",
  36738=>"000011011",
  36739=>"110000111",
  36740=>"000100111",
  36741=>"101111010",
  36742=>"000101011",
  36743=>"101100111",
  36744=>"110101001",
  36745=>"000111111",
  36746=>"100101011",
  36747=>"011111001",
  36748=>"011101110",
  36749=>"100110100",
  36750=>"001111100",
  36751=>"000001000",
  36752=>"101110000",
  36753=>"101100101",
  36754=>"000001110",
  36755=>"010100110",
  36756=>"100010101",
  36757=>"010110000",
  36758=>"100011010",
  36759=>"100101001",
  36760=>"101001111",
  36761=>"001001011",
  36762=>"100001111",
  36763=>"100001010",
  36764=>"101110111",
  36765=>"000111011",
  36766=>"001101001",
  36767=>"101101111",
  36768=>"100110010",
  36769=>"100001001",
  36770=>"100101001",
  36771=>"011101110",
  36772=>"010000110",
  36773=>"110111111",
  36774=>"001100011",
  36775=>"000110001",
  36776=>"010110011",
  36777=>"010110101",
  36778=>"010111011",
  36779=>"011111100",
  36780=>"010111010",
  36781=>"100100101",
  36782=>"101001000",
  36783=>"101001110",
  36784=>"101000011",
  36785=>"111101011",
  36786=>"111011111",
  36787=>"001101101",
  36788=>"111010000",
  36789=>"011000011",
  36790=>"111000110",
  36791=>"111100000",
  36792=>"011010100",
  36793=>"000011010",
  36794=>"011100011",
  36795=>"000101010",
  36796=>"011111000",
  36797=>"000010101",
  36798=>"010001000",
  36799=>"001110000",
  36800=>"111010011",
  36801=>"110100000",
  36802=>"110111111",
  36803=>"101001110",
  36804=>"011110000",
  36805=>"001010111",
  36806=>"001101000",
  36807=>"000101000",
  36808=>"000000010",
  36809=>"001011101",
  36810=>"010100111",
  36811=>"111100000",
  36812=>"010110100",
  36813=>"010000100",
  36814=>"010101100",
  36815=>"101110010",
  36816=>"101000111",
  36817=>"000000101",
  36818=>"010001001",
  36819=>"000010101",
  36820=>"010100001",
  36821=>"111010101",
  36822=>"100000010",
  36823=>"010010111",
  36824=>"111101111",
  36825=>"110101100",
  36826=>"001011100",
  36827=>"010001000",
  36828=>"011010100",
  36829=>"111111101",
  36830=>"001000111",
  36831=>"000001010",
  36832=>"111000011",
  36833=>"000001011",
  36834=>"111100101",
  36835=>"011110001",
  36836=>"000000101",
  36837=>"011001001",
  36838=>"110010111",
  36839=>"110000100",
  36840=>"010001010",
  36841=>"011100100",
  36842=>"001111100",
  36843=>"100010001",
  36844=>"010110001",
  36845=>"110010101",
  36846=>"110001011",
  36847=>"100011101",
  36848=>"110000011",
  36849=>"001101110",
  36850=>"000010001",
  36851=>"010110001",
  36852=>"010000111",
  36853=>"100000000",
  36854=>"110110111",
  36855=>"100001111",
  36856=>"111000011",
  36857=>"111111100",
  36858=>"100110101",
  36859=>"001000001",
  36860=>"010001010",
  36861=>"101001001",
  36862=>"111000110",
  36863=>"000110110",
  36864=>"000000100",
  36865=>"010100111",
  36866=>"110010101",
  36867=>"110101000",
  36868=>"100110010",
  36869=>"000101100",
  36870=>"111111110",
  36871=>"011001101",
  36872=>"000001010",
  36873=>"010000001",
  36874=>"110000111",
  36875=>"111100100",
  36876=>"010010001",
  36877=>"111011110",
  36878=>"100000010",
  36879=>"011100111",
  36880=>"010101101",
  36881=>"001101110",
  36882=>"110101011",
  36883=>"111110100",
  36884=>"011001001",
  36885=>"100100010",
  36886=>"100111000",
  36887=>"001111011",
  36888=>"100101000",
  36889=>"000101011",
  36890=>"100010101",
  36891=>"001010010",
  36892=>"110001101",
  36893=>"001011001",
  36894=>"001001011",
  36895=>"010010010",
  36896=>"000111111",
  36897=>"101011100",
  36898=>"101100000",
  36899=>"001000011",
  36900=>"111111010",
  36901=>"000000001",
  36902=>"101111101",
  36903=>"101000100",
  36904=>"111111101",
  36905=>"010111010",
  36906=>"000101110",
  36907=>"001011000",
  36908=>"101101110",
  36909=>"011000100",
  36910=>"111101101",
  36911=>"010111011",
  36912=>"000010100",
  36913=>"000000100",
  36914=>"111011110",
  36915=>"110110101",
  36916=>"000001100",
  36917=>"100010100",
  36918=>"011011100",
  36919=>"001001111",
  36920=>"000100010",
  36921=>"000110000",
  36922=>"000001101",
  36923=>"011000111",
  36924=>"011000111",
  36925=>"011011111",
  36926=>"001011011",
  36927=>"001111001",
  36928=>"001011110",
  36929=>"001010001",
  36930=>"101101110",
  36931=>"001010010",
  36932=>"100001100",
  36933=>"011101011",
  36934=>"011001000",
  36935=>"010101101",
  36936=>"100001100",
  36937=>"010010100",
  36938=>"100001010",
  36939=>"011110111",
  36940=>"101010010",
  36941=>"110010011",
  36942=>"000110000",
  36943=>"001100001",
  36944=>"101001000",
  36945=>"011010101",
  36946=>"100000100",
  36947=>"011100000",
  36948=>"111100101",
  36949=>"011010010",
  36950=>"111010001",
  36951=>"010010110",
  36952=>"011111100",
  36953=>"111100010",
  36954=>"011010000",
  36955=>"100111001",
  36956=>"101000001",
  36957=>"101010110",
  36958=>"001111100",
  36959=>"111011001",
  36960=>"010111111",
  36961=>"001011100",
  36962=>"101000010",
  36963=>"101000100",
  36964=>"001000110",
  36965=>"001110111",
  36966=>"110001000",
  36967=>"010100100",
  36968=>"010011010",
  36969=>"011111010",
  36970=>"010100101",
  36971=>"000101111",
  36972=>"110100001",
  36973=>"001001101",
  36974=>"110001111",
  36975=>"011111001",
  36976=>"110010101",
  36977=>"011001011",
  36978=>"101011010",
  36979=>"001010010",
  36980=>"010000001",
  36981=>"111100001",
  36982=>"011111010",
  36983=>"010100000",
  36984=>"111101000",
  36985=>"110011000",
  36986=>"101011001",
  36987=>"010001111",
  36988=>"001011100",
  36989=>"001111101",
  36990=>"000000000",
  36991=>"101101111",
  36992=>"011110000",
  36993=>"010111011",
  36994=>"000110011",
  36995=>"000100111",
  36996=>"100101101",
  36997=>"101111110",
  36998=>"111100101",
  36999=>"010010000",
  37000=>"101011000",
  37001=>"100000010",
  37002=>"000010111",
  37003=>"111110000",
  37004=>"111001000",
  37005=>"001110101",
  37006=>"111000000",
  37007=>"010001000",
  37008=>"010011100",
  37009=>"110010111",
  37010=>"001011101",
  37011=>"101110011",
  37012=>"100101110",
  37013=>"100000110",
  37014=>"000011111",
  37015=>"010100100",
  37016=>"101000111",
  37017=>"001010001",
  37018=>"000001000",
  37019=>"100011001",
  37020=>"010011110",
  37021=>"000101110",
  37022=>"000000100",
  37023=>"111010100",
  37024=>"000100111",
  37025=>"111100010",
  37026=>"110000111",
  37027=>"000100111",
  37028=>"011000100",
  37029=>"100011101",
  37030=>"100101111",
  37031=>"011111010",
  37032=>"110110110",
  37033=>"100010101",
  37034=>"001001111",
  37035=>"011100101",
  37036=>"111101111",
  37037=>"000010110",
  37038=>"100011100",
  37039=>"100110111",
  37040=>"100000001",
  37041=>"001111110",
  37042=>"111110001",
  37043=>"100000010",
  37044=>"101011101",
  37045=>"011100101",
  37046=>"110110111",
  37047=>"001101101",
  37048=>"101011110",
  37049=>"001101101",
  37050=>"011111111",
  37051=>"100011000",
  37052=>"100001001",
  37053=>"000101010",
  37054=>"001000101",
  37055=>"101001010",
  37056=>"010100000",
  37057=>"110011001",
  37058=>"000110101",
  37059=>"110110010",
  37060=>"000001001",
  37061=>"010011011",
  37062=>"000001111",
  37063=>"011000100",
  37064=>"101000011",
  37065=>"110000100",
  37066=>"110010000",
  37067=>"000011110",
  37068=>"001100110",
  37069=>"000011101",
  37070=>"100000100",
  37071=>"001000010",
  37072=>"110110000",
  37073=>"010011101",
  37074=>"101110100",
  37075=>"010111100",
  37076=>"011000000",
  37077=>"011111110",
  37078=>"101011000",
  37079=>"001000001",
  37080=>"110110011",
  37081=>"001001111",
  37082=>"111110000",
  37083=>"100010111",
  37084=>"100101010",
  37085=>"010100110",
  37086=>"101111001",
  37087=>"001010111",
  37088=>"010001110",
  37089=>"001000011",
  37090=>"000110100",
  37091=>"011101101",
  37092=>"101100110",
  37093=>"110100011",
  37094=>"010110110",
  37095=>"000101100",
  37096=>"100100010",
  37097=>"010001011",
  37098=>"100111010",
  37099=>"100011011",
  37100=>"011011001",
  37101=>"011100001",
  37102=>"100100001",
  37103=>"000111101",
  37104=>"111111011",
  37105=>"011010010",
  37106=>"001100001",
  37107=>"101000000",
  37108=>"000110111",
  37109=>"011111010",
  37110=>"011111100",
  37111=>"000011110",
  37112=>"100111001",
  37113=>"001001000",
  37114=>"110101000",
  37115=>"111011001",
  37116=>"000011001",
  37117=>"100010000",
  37118=>"011110011",
  37119=>"001110010",
  37120=>"010010011",
  37121=>"011011110",
  37122=>"000100101",
  37123=>"010010010",
  37124=>"001000010",
  37125=>"001001100",
  37126=>"001110110",
  37127=>"101110000",
  37128=>"100111101",
  37129=>"000100011",
  37130=>"000011000",
  37131=>"000000000",
  37132=>"000010100",
  37133=>"100111000",
  37134=>"000100001",
  37135=>"000100111",
  37136=>"011110000",
  37137=>"100111001",
  37138=>"110010000",
  37139=>"000101100",
  37140=>"000110100",
  37141=>"111101101",
  37142=>"010010011",
  37143=>"011011010",
  37144=>"101101011",
  37145=>"010111001",
  37146=>"111000100",
  37147=>"110001111",
  37148=>"101000000",
  37149=>"000110001",
  37150=>"101010100",
  37151=>"110010000",
  37152=>"011110110",
  37153=>"010000011",
  37154=>"011000110",
  37155=>"010001111",
  37156=>"000001010",
  37157=>"110101000",
  37158=>"000001000",
  37159=>"001110110",
  37160=>"100011000",
  37161=>"001001110",
  37162=>"111100001",
  37163=>"000100100",
  37164=>"110011101",
  37165=>"110100001",
  37166=>"111011111",
  37167=>"010111111",
  37168=>"011011110",
  37169=>"100001111",
  37170=>"101110101",
  37171=>"011001000",
  37172=>"110000011",
  37173=>"010100001",
  37174=>"001011001",
  37175=>"000000101",
  37176=>"001110111",
  37177=>"010001011",
  37178=>"111101011",
  37179=>"110010110",
  37180=>"001111011",
  37181=>"100000011",
  37182=>"100110100",
  37183=>"001100000",
  37184=>"100100110",
  37185=>"000111110",
  37186=>"000010001",
  37187=>"011100110",
  37188=>"100000010",
  37189=>"101100000",
  37190=>"000101011",
  37191=>"110001011",
  37192=>"100110111",
  37193=>"100101001",
  37194=>"010010010",
  37195=>"110100000",
  37196=>"110011111",
  37197=>"010110101",
  37198=>"001001100",
  37199=>"100110101",
  37200=>"110010110",
  37201=>"110100001",
  37202=>"110110000",
  37203=>"001011010",
  37204=>"001101110",
  37205=>"000000000",
  37206=>"101111011",
  37207=>"101110100",
  37208=>"000011111",
  37209=>"001000011",
  37210=>"100111010",
  37211=>"001110001",
  37212=>"101001010",
  37213=>"000110101",
  37214=>"010110110",
  37215=>"000001111",
  37216=>"100010101",
  37217=>"010001011",
  37218=>"000011101",
  37219=>"000001110",
  37220=>"101101101",
  37221=>"100001011",
  37222=>"101111110",
  37223=>"100001110",
  37224=>"110010011",
  37225=>"000001111",
  37226=>"110001101",
  37227=>"001011000",
  37228=>"110011110",
  37229=>"111000010",
  37230=>"101101101",
  37231=>"011100010",
  37232=>"001010111",
  37233=>"001111010",
  37234=>"001100101",
  37235=>"100110100",
  37236=>"100100110",
  37237=>"001101011",
  37238=>"000011011",
  37239=>"101000001",
  37240=>"011011111",
  37241=>"111001101",
  37242=>"111001000",
  37243=>"000011111",
  37244=>"010011110",
  37245=>"110000010",
  37246=>"111000001",
  37247=>"001111010",
  37248=>"000000010",
  37249=>"010110110",
  37250=>"000000101",
  37251=>"000001100",
  37252=>"111011100",
  37253=>"111001100",
  37254=>"100000111",
  37255=>"111101011",
  37256=>"101101001",
  37257=>"110100110",
  37258=>"001110011",
  37259=>"110111001",
  37260=>"000010001",
  37261=>"000101011",
  37262=>"100000111",
  37263=>"000001010",
  37264=>"011111011",
  37265=>"111001111",
  37266=>"011101100",
  37267=>"011110010",
  37268=>"111111010",
  37269=>"100101001",
  37270=>"000011001",
  37271=>"100100110",
  37272=>"111111111",
  37273=>"100101111",
  37274=>"001010110",
  37275=>"000110101",
  37276=>"111101101",
  37277=>"011111010",
  37278=>"100100111",
  37279=>"111111100",
  37280=>"010000101",
  37281=>"000111011",
  37282=>"010000101",
  37283=>"000100100",
  37284=>"101011111",
  37285=>"111000111",
  37286=>"100110101",
  37287=>"100011101",
  37288=>"101101111",
  37289=>"111101101",
  37290=>"001000000",
  37291=>"000001100",
  37292=>"000001110",
  37293=>"010100111",
  37294=>"000011111",
  37295=>"101111000",
  37296=>"110101000",
  37297=>"101001001",
  37298=>"100011011",
  37299=>"011011000",
  37300=>"001011010",
  37301=>"001101001",
  37302=>"100101101",
  37303=>"101100010",
  37304=>"110010100",
  37305=>"111010110",
  37306=>"000010011",
  37307=>"010010010",
  37308=>"100111100",
  37309=>"111000101",
  37310=>"101000101",
  37311=>"010011001",
  37312=>"001101101",
  37313=>"101111000",
  37314=>"001001110",
  37315=>"101010111",
  37316=>"000000100",
  37317=>"111111101",
  37318=>"010101111",
  37319=>"110011001",
  37320=>"000011111",
  37321=>"001110001",
  37322=>"111010010",
  37323=>"000010000",
  37324=>"101001110",
  37325=>"111011000",
  37326=>"000110011",
  37327=>"010010010",
  37328=>"010100011",
  37329=>"011110001",
  37330=>"101111100",
  37331=>"100101010",
  37332=>"011011000",
  37333=>"110011010",
  37334=>"100100001",
  37335=>"100111001",
  37336=>"001011101",
  37337=>"001100001",
  37338=>"001010000",
  37339=>"010111101",
  37340=>"111100110",
  37341=>"110010011",
  37342=>"100000011",
  37343=>"000101011",
  37344=>"101001110",
  37345=>"101111010",
  37346=>"000001011",
  37347=>"000000110",
  37348=>"100010100",
  37349=>"110000001",
  37350=>"111011110",
  37351=>"111000001",
  37352=>"110110110",
  37353=>"010010100",
  37354=>"101111100",
  37355=>"011010111",
  37356=>"011100000",
  37357=>"010000001",
  37358=>"011001001",
  37359=>"111101011",
  37360=>"111100100",
  37361=>"011010010",
  37362=>"001110110",
  37363=>"010001111",
  37364=>"110000101",
  37365=>"001101001",
  37366=>"100100110",
  37367=>"110111011",
  37368=>"000111100",
  37369=>"101011110",
  37370=>"100001000",
  37371=>"101100000",
  37372=>"110101111",
  37373=>"010100101",
  37374=>"101100100",
  37375=>"100000101",
  37376=>"111000110",
  37377=>"111010111",
  37378=>"100011101",
  37379=>"011001001",
  37380=>"101110111",
  37381=>"110110100",
  37382=>"000000001",
  37383=>"100110000",
  37384=>"100000110",
  37385=>"000110011",
  37386=>"000010000",
  37387=>"110000000",
  37388=>"101111111",
  37389=>"001101001",
  37390=>"011011000",
  37391=>"010100011",
  37392=>"011001100",
  37393=>"100000010",
  37394=>"101000001",
  37395=>"111000000",
  37396=>"101001101",
  37397=>"010110011",
  37398=>"101010000",
  37399=>"110111011",
  37400=>"000001010",
  37401=>"100110000",
  37402=>"001000111",
  37403=>"010011001",
  37404=>"011011110",
  37405=>"011110010",
  37406=>"101110010",
  37407=>"111001011",
  37408=>"100000101",
  37409=>"111000111",
  37410=>"011011001",
  37411=>"100011101",
  37412=>"101100001",
  37413=>"000000111",
  37414=>"011000010",
  37415=>"100100110",
  37416=>"010110011",
  37417=>"111000001",
  37418=>"100101111",
  37419=>"001000101",
  37420=>"001110100",
  37421=>"011100100",
  37422=>"001000011",
  37423=>"010001010",
  37424=>"100000100",
  37425=>"110100111",
  37426=>"010000100",
  37427=>"101001101",
  37428=>"111111110",
  37429=>"010101000",
  37430=>"011111111",
  37431=>"111101111",
  37432=>"110110110",
  37433=>"111110001",
  37434=>"010110111",
  37435=>"111111000",
  37436=>"111100010",
  37437=>"000100000",
  37438=>"110000001",
  37439=>"100011101",
  37440=>"001001001",
  37441=>"111011111",
  37442=>"011010011",
  37443=>"110010101",
  37444=>"000000001",
  37445=>"000110111",
  37446=>"111110100",
  37447=>"011001010",
  37448=>"011011010",
  37449=>"000000011",
  37450=>"011101000",
  37451=>"001010110",
  37452=>"101010011",
  37453=>"010001001",
  37454=>"110111000",
  37455=>"100011010",
  37456=>"000100101",
  37457=>"111100100",
  37458=>"000000100",
  37459=>"001111100",
  37460=>"011110101",
  37461=>"001010010",
  37462=>"101110101",
  37463=>"101011100",
  37464=>"010100010",
  37465=>"101001000",
  37466=>"001010001",
  37467=>"001100101",
  37468=>"010011101",
  37469=>"000010010",
  37470=>"010000111",
  37471=>"111011110",
  37472=>"010001010",
  37473=>"011001001",
  37474=>"101110100",
  37475=>"001001101",
  37476=>"011010001",
  37477=>"111100000",
  37478=>"100100111",
  37479=>"001000100",
  37480=>"010110110",
  37481=>"001011111",
  37482=>"000011101",
  37483=>"001100000",
  37484=>"001101010",
  37485=>"001000000",
  37486=>"010100001",
  37487=>"100100001",
  37488=>"110011011",
  37489=>"101101100",
  37490=>"000100111",
  37491=>"000000100",
  37492=>"101101111",
  37493=>"011010000",
  37494=>"100110110",
  37495=>"000100010",
  37496=>"110011000",
  37497=>"011000101",
  37498=>"101111000",
  37499=>"101100010",
  37500=>"110001000",
  37501=>"001010111",
  37502=>"100000100",
  37503=>"001011101",
  37504=>"000000110",
  37505=>"010011011",
  37506=>"011110000",
  37507=>"010101101",
  37508=>"001100001",
  37509=>"100110100",
  37510=>"100000011",
  37511=>"100111110",
  37512=>"011010110",
  37513=>"010011010",
  37514=>"000111011",
  37515=>"011101011",
  37516=>"000001111",
  37517=>"010000110",
  37518=>"101000010",
  37519=>"000011000",
  37520=>"101001001",
  37521=>"111101010",
  37522=>"111001011",
  37523=>"101011000",
  37524=>"101100011",
  37525=>"000110011",
  37526=>"110011001",
  37527=>"101000100",
  37528=>"011100011",
  37529=>"100100110",
  37530=>"011011110",
  37531=>"110011000",
  37532=>"011101011",
  37533=>"100010101",
  37534=>"110011111",
  37535=>"111001000",
  37536=>"001000110",
  37537=>"110110010",
  37538=>"001101111",
  37539=>"011000001",
  37540=>"011110011",
  37541=>"011001010",
  37542=>"000011010",
  37543=>"000000000",
  37544=>"100000010",
  37545=>"000010010",
  37546=>"001011100",
  37547=>"101111100",
  37548=>"100000011",
  37549=>"101101010",
  37550=>"100101011",
  37551=>"010011010",
  37552=>"111111000",
  37553=>"111000100",
  37554=>"101100111",
  37555=>"001010011",
  37556=>"110111101",
  37557=>"111011110",
  37558=>"001000000",
  37559=>"111100100",
  37560=>"000100100",
  37561=>"000001011",
  37562=>"110111100",
  37563=>"011011111",
  37564=>"100110010",
  37565=>"100110001",
  37566=>"010111010",
  37567=>"000001000",
  37568=>"010101000",
  37569=>"101100110",
  37570=>"011101101",
  37571=>"001110101",
  37572=>"011100001",
  37573=>"110010100",
  37574=>"111001011",
  37575=>"110001000",
  37576=>"010101101",
  37577=>"110010110",
  37578=>"000010001",
  37579=>"001010101",
  37580=>"001011010",
  37581=>"010110111",
  37582=>"101000001",
  37583=>"000110010",
  37584=>"000000010",
  37585=>"110000010",
  37586=>"110100111",
  37587=>"100010001",
  37588=>"011101010",
  37589=>"100000110",
  37590=>"000001100",
  37591=>"001010010",
  37592=>"100011001",
  37593=>"110111001",
  37594=>"100011101",
  37595=>"001001101",
  37596=>"101010110",
  37597=>"010000010",
  37598=>"011001111",
  37599=>"110001000",
  37600=>"110110011",
  37601=>"001000100",
  37602=>"000011000",
  37603=>"100110100",
  37604=>"111110001",
  37605=>"100000100",
  37606=>"010010100",
  37607=>"011010000",
  37608=>"011011011",
  37609=>"101110011",
  37610=>"011111001",
  37611=>"100111000",
  37612=>"000000111",
  37613=>"111101111",
  37614=>"111010100",
  37615=>"110011010",
  37616=>"100000000",
  37617=>"100010001",
  37618=>"011011110",
  37619=>"110001101",
  37620=>"100010000",
  37621=>"000100111",
  37622=>"000111101",
  37623=>"010000110",
  37624=>"011001100",
  37625=>"110000010",
  37626=>"000000011",
  37627=>"110010111",
  37628=>"101001001",
  37629=>"011011000",
  37630=>"110001111",
  37631=>"101000000",
  37632=>"100101011",
  37633=>"000111100",
  37634=>"111110011",
  37635=>"010010110",
  37636=>"111000110",
  37637=>"010011000",
  37638=>"000010001",
  37639=>"110101110",
  37640=>"100111101",
  37641=>"100011001",
  37642=>"001000010",
  37643=>"000001010",
  37644=>"000001011",
  37645=>"001110010",
  37646=>"101000010",
  37647=>"100111110",
  37648=>"100000110",
  37649=>"101010110",
  37650=>"000001001",
  37651=>"001111110",
  37652=>"010010110",
  37653=>"111010000",
  37654=>"110001010",
  37655=>"110101111",
  37656=>"001011001",
  37657=>"001010100",
  37658=>"111100000",
  37659=>"100111011",
  37660=>"100011001",
  37661=>"110001111",
  37662=>"111000000",
  37663=>"100011111",
  37664=>"000000001",
  37665=>"111100101",
  37666=>"111011011",
  37667=>"000111101",
  37668=>"000000011",
  37669=>"100010111",
  37670=>"101100111",
  37671=>"010000111",
  37672=>"000001101",
  37673=>"111100011",
  37674=>"000011010",
  37675=>"110110000",
  37676=>"111100100",
  37677=>"001100011",
  37678=>"001001110",
  37679=>"110110111",
  37680=>"101111111",
  37681=>"111111110",
  37682=>"001000110",
  37683=>"000100111",
  37684=>"110000001",
  37685=>"010001001",
  37686=>"001110111",
  37687=>"000011110",
  37688=>"101011100",
  37689=>"000010101",
  37690=>"000000110",
  37691=>"000111010",
  37692=>"001010010",
  37693=>"110111000",
  37694=>"110100000",
  37695=>"000111010",
  37696=>"100111011",
  37697=>"001001000",
  37698=>"101111101",
  37699=>"000100010",
  37700=>"111000010",
  37701=>"011001101",
  37702=>"001011101",
  37703=>"100111111",
  37704=>"100000111",
  37705=>"101011010",
  37706=>"100101000",
  37707=>"000100001",
  37708=>"100010100",
  37709=>"100000011",
  37710=>"111000001",
  37711=>"000010000",
  37712=>"110111110",
  37713=>"001100101",
  37714=>"001010000",
  37715=>"100000010",
  37716=>"111111110",
  37717=>"110011001",
  37718=>"011010110",
  37719=>"010001101",
  37720=>"010100111",
  37721=>"110011000",
  37722=>"001011111",
  37723=>"001110011",
  37724=>"001010000",
  37725=>"000001011",
  37726=>"100011001",
  37727=>"010000110",
  37728=>"001001110",
  37729=>"011100011",
  37730=>"000101110",
  37731=>"001110001",
  37732=>"010101110",
  37733=>"101000101",
  37734=>"011001000",
  37735=>"111100110",
  37736=>"000010101",
  37737=>"111000001",
  37738=>"110101000",
  37739=>"001011011",
  37740=>"101001001",
  37741=>"100010111",
  37742=>"111100110",
  37743=>"011011001",
  37744=>"100011100",
  37745=>"010100100",
  37746=>"100100001",
  37747=>"000100010",
  37748=>"111011000",
  37749=>"110101011",
  37750=>"100000000",
  37751=>"001100011",
  37752=>"010001100",
  37753=>"000010010",
  37754=>"001110100",
  37755=>"010010011",
  37756=>"101110101",
  37757=>"011111011",
  37758=>"001010110",
  37759=>"010110101",
  37760=>"101100010",
  37761=>"001110111",
  37762=>"010001010",
  37763=>"110101010",
  37764=>"111110001",
  37765=>"100000010",
  37766=>"010111101",
  37767=>"001100110",
  37768=>"111101010",
  37769=>"001100010",
  37770=>"110100010",
  37771=>"111011100",
  37772=>"100010100",
  37773=>"001100010",
  37774=>"000001000",
  37775=>"100101100",
  37776=>"000111001",
  37777=>"101100110",
  37778=>"111010000",
  37779=>"010011110",
  37780=>"010001111",
  37781=>"110010011",
  37782=>"010001101",
  37783=>"000001100",
  37784=>"000101010",
  37785=>"010011011",
  37786=>"110010001",
  37787=>"000101101",
  37788=>"000111110",
  37789=>"100111001",
  37790=>"011001010",
  37791=>"100110110",
  37792=>"001000111",
  37793=>"010000111",
  37794=>"101001011",
  37795=>"101100110",
  37796=>"000110111",
  37797=>"010110010",
  37798=>"000100011",
  37799=>"001100110",
  37800=>"111011111",
  37801=>"011110110",
  37802=>"001010101",
  37803=>"001010000",
  37804=>"100101111",
  37805=>"110000001",
  37806=>"101001101",
  37807=>"000000000",
  37808=>"000110100",
  37809=>"110001010",
  37810=>"100101110",
  37811=>"000111111",
  37812=>"011000011",
  37813=>"111111010",
  37814=>"101100111",
  37815=>"011110101",
  37816=>"010100000",
  37817=>"011001100",
  37818=>"001110000",
  37819=>"011110011",
  37820=>"100101001",
  37821=>"000000000",
  37822=>"001111100",
  37823=>"010110101",
  37824=>"111100101",
  37825=>"001110011",
  37826=>"110011111",
  37827=>"101011001",
  37828=>"111100010",
  37829=>"011101100",
  37830=>"110001010",
  37831=>"100110000",
  37832=>"111111111",
  37833=>"010101110",
  37834=>"010110000",
  37835=>"100001101",
  37836=>"010001000",
  37837=>"101011000",
  37838=>"010101100",
  37839=>"010100011",
  37840=>"111101100",
  37841=>"000011101",
  37842=>"111101100",
  37843=>"001000000",
  37844=>"111000011",
  37845=>"011011001",
  37846=>"001001011",
  37847=>"111111011",
  37848=>"001111101",
  37849=>"001111101",
  37850=>"000001101",
  37851=>"111110111",
  37852=>"000000001",
  37853=>"111010010",
  37854=>"011101110",
  37855=>"100101110",
  37856=>"010111101",
  37857=>"001100001",
  37858=>"001010011",
  37859=>"111110010",
  37860=>"110111000",
  37861=>"000000110",
  37862=>"000101011",
  37863=>"000010101",
  37864=>"010001111",
  37865=>"111111101",
  37866=>"101001101",
  37867=>"110100110",
  37868=>"001110000",
  37869=>"000101010",
  37870=>"010010100",
  37871=>"011000000",
  37872=>"011110000",
  37873=>"110001000",
  37874=>"000010001",
  37875=>"100100000",
  37876=>"101001001",
  37877=>"010101011",
  37878=>"010011000",
  37879=>"111010111",
  37880=>"000000010",
  37881=>"011101100",
  37882=>"111111010",
  37883=>"110010101",
  37884=>"111110001",
  37885=>"000111111",
  37886=>"010111111",
  37887=>"010110001",
  37888=>"110011111",
  37889=>"001011010",
  37890=>"111011101",
  37891=>"100010000",
  37892=>"110000100",
  37893=>"001000011",
  37894=>"100101100",
  37895=>"000110100",
  37896=>"010101011",
  37897=>"110000110",
  37898=>"011111111",
  37899=>"110011010",
  37900=>"001111011",
  37901=>"111111110",
  37902=>"110101111",
  37903=>"100100111",
  37904=>"011000000",
  37905=>"100001010",
  37906=>"010000110",
  37907=>"010010101",
  37908=>"101000110",
  37909=>"101010010",
  37910=>"000011111",
  37911=>"001000010",
  37912=>"101111010",
  37913=>"110010100",
  37914=>"110110010",
  37915=>"101011100",
  37916=>"110111001",
  37917=>"110111100",
  37918=>"010010010",
  37919=>"100011001",
  37920=>"011101101",
  37921=>"111011100",
  37922=>"001000000",
  37923=>"011011111",
  37924=>"111111001",
  37925=>"111010010",
  37926=>"101111010",
  37927=>"110101111",
  37928=>"111011100",
  37929=>"100011100",
  37930=>"010001101",
  37931=>"101110010",
  37932=>"100001100",
  37933=>"011111100",
  37934=>"101101010",
  37935=>"000111000",
  37936=>"111000001",
  37937=>"100111001",
  37938=>"000000000",
  37939=>"000010101",
  37940=>"101111111",
  37941=>"001100100",
  37942=>"000000100",
  37943=>"101100110",
  37944=>"111011100",
  37945=>"011011011",
  37946=>"000111101",
  37947=>"010111010",
  37948=>"000000110",
  37949=>"000011100",
  37950=>"001110111",
  37951=>"111011000",
  37952=>"111010111",
  37953=>"001110100",
  37954=>"101100000",
  37955=>"000000000",
  37956=>"010001100",
  37957=>"010000001",
  37958=>"110110000",
  37959=>"001111010",
  37960=>"100110001",
  37961=>"110011111",
  37962=>"111010011",
  37963=>"110001001",
  37964=>"100011000",
  37965=>"001100100",
  37966=>"110111110",
  37967=>"100001001",
  37968=>"010111011",
  37969=>"110010001",
  37970=>"111110010",
  37971=>"101111100",
  37972=>"010001100",
  37973=>"100100001",
  37974=>"101000011",
  37975=>"110101000",
  37976=>"101010110",
  37977=>"100101110",
  37978=>"110111000",
  37979=>"110000110",
  37980=>"100101000",
  37981=>"011011010",
  37982=>"011110111",
  37983=>"001100000",
  37984=>"100111100",
  37985=>"011101000",
  37986=>"111011111",
  37987=>"011110011",
  37988=>"100111111",
  37989=>"010001010",
  37990=>"111010100",
  37991=>"001110101",
  37992=>"010010001",
  37993=>"100001100",
  37994=>"000001100",
  37995=>"100110010",
  37996=>"100001100",
  37997=>"100001100",
  37998=>"100111110",
  37999=>"010011111",
  38000=>"010000111",
  38001=>"111011101",
  38002=>"000000101",
  38003=>"011011111",
  38004=>"100111100",
  38005=>"001001011",
  38006=>"110110011",
  38007=>"100110100",
  38008=>"110111001",
  38009=>"100101111",
  38010=>"110011101",
  38011=>"000101011",
  38012=>"011110011",
  38013=>"100000110",
  38014=>"111111111",
  38015=>"111011000",
  38016=>"111000111",
  38017=>"011000111",
  38018=>"010000111",
  38019=>"111010111",
  38020=>"011010101",
  38021=>"010010101",
  38022=>"000110111",
  38023=>"011101101",
  38024=>"011100001",
  38025=>"000010001",
  38026=>"011110111",
  38027=>"111111110",
  38028=>"111110111",
  38029=>"100110001",
  38030=>"101010010",
  38031=>"001111100",
  38032=>"110100000",
  38033=>"001000001",
  38034=>"011010001",
  38035=>"110111000",
  38036=>"111111100",
  38037=>"100101100",
  38038=>"100111110",
  38039=>"101010010",
  38040=>"000010011",
  38041=>"101100011",
  38042=>"011111110",
  38043=>"111001001",
  38044=>"001100100",
  38045=>"100101001",
  38046=>"110010100",
  38047=>"100100011",
  38048=>"001111101",
  38049=>"101001001",
  38050=>"101100010",
  38051=>"101010101",
  38052=>"101000010",
  38053=>"101010010",
  38054=>"010110111",
  38055=>"100010000",
  38056=>"101110101",
  38057=>"111110110",
  38058=>"000010000",
  38059=>"110011010",
  38060=>"011000000",
  38061=>"111001001",
  38062=>"100101001",
  38063=>"000100000",
  38064=>"101111011",
  38065=>"101011010",
  38066=>"111001100",
  38067=>"001001100",
  38068=>"110100000",
  38069=>"110001111",
  38070=>"101111111",
  38071=>"111000110",
  38072=>"001100110",
  38073=>"100110111",
  38074=>"110101110",
  38075=>"111000101",
  38076=>"000111000",
  38077=>"010001001",
  38078=>"000001000",
  38079=>"110010111",
  38080=>"010101100",
  38081=>"001010010",
  38082=>"001000111",
  38083=>"100100010",
  38084=>"100000000",
  38085=>"000101011",
  38086=>"101101001",
  38087=>"001101100",
  38088=>"111000011",
  38089=>"101101010",
  38090=>"001111001",
  38091=>"010100010",
  38092=>"011010110",
  38093=>"111110011",
  38094=>"100010101",
  38095=>"101100110",
  38096=>"101001101",
  38097=>"000000110",
  38098=>"000100100",
  38099=>"011010000",
  38100=>"101100010",
  38101=>"110001011",
  38102=>"101111101",
  38103=>"101011110",
  38104=>"111011011",
  38105=>"101110110",
  38106=>"010110011",
  38107=>"000100000",
  38108=>"011101101",
  38109=>"110100011",
  38110=>"000011100",
  38111=>"100011110",
  38112=>"100011010",
  38113=>"111100101",
  38114=>"110111010",
  38115=>"100011111",
  38116=>"100100000",
  38117=>"100100011",
  38118=>"110010100",
  38119=>"010101111",
  38120=>"000011101",
  38121=>"100100000",
  38122=>"000101110",
  38123=>"011011011",
  38124=>"110111110",
  38125=>"111100010",
  38126=>"000011011",
  38127=>"111000101",
  38128=>"101010011",
  38129=>"000100100",
  38130=>"100000011",
  38131=>"010010110",
  38132=>"100000100",
  38133=>"111010001",
  38134=>"100011010",
  38135=>"010100111",
  38136=>"111111100",
  38137=>"001101101",
  38138=>"110010000",
  38139=>"111101001",
  38140=>"001101010",
  38141=>"010101000",
  38142=>"101011100",
  38143=>"101001101",
  38144=>"100111010",
  38145=>"101111011",
  38146=>"111111011",
  38147=>"111010111",
  38148=>"110111101",
  38149=>"100100010",
  38150=>"111111001",
  38151=>"110100001",
  38152=>"010111000",
  38153=>"101111101",
  38154=>"010010011",
  38155=>"001001110",
  38156=>"000110000",
  38157=>"000010111",
  38158=>"010100011",
  38159=>"001111100",
  38160=>"011010001",
  38161=>"110000111",
  38162=>"000011111",
  38163=>"010111110",
  38164=>"100010100",
  38165=>"001110010",
  38166=>"110111100",
  38167=>"000010101",
  38168=>"110010110",
  38169=>"010001111",
  38170=>"000110101",
  38171=>"111111110",
  38172=>"111110001",
  38173=>"100000111",
  38174=>"110101110",
  38175=>"111111101",
  38176=>"101001110",
  38177=>"100101110",
  38178=>"100001110",
  38179=>"010011111",
  38180=>"011100000",
  38181=>"110010011",
  38182=>"100010011",
  38183=>"001010101",
  38184=>"101001000",
  38185=>"101001101",
  38186=>"000010111",
  38187=>"111010001",
  38188=>"101110001",
  38189=>"001111101",
  38190=>"011100111",
  38191=>"011100100",
  38192=>"010110110",
  38193=>"000100001",
  38194=>"001011010",
  38195=>"001001001",
  38196=>"001110001",
  38197=>"111110011",
  38198=>"000000111",
  38199=>"100100101",
  38200=>"100101001",
  38201=>"111001011",
  38202=>"101101100",
  38203=>"011110001",
  38204=>"011101011",
  38205=>"110111001",
  38206=>"010101000",
  38207=>"100000111",
  38208=>"000100101",
  38209=>"000010010",
  38210=>"010100111",
  38211=>"110011111",
  38212=>"001010010",
  38213=>"101101110",
  38214=>"011100010",
  38215=>"100111110",
  38216=>"010010010",
  38217=>"101110101",
  38218=>"010110111",
  38219=>"001100111",
  38220=>"011000100",
  38221=>"000100011",
  38222=>"000001010",
  38223=>"111100111",
  38224=>"110110101",
  38225=>"000001110",
  38226=>"011011011",
  38227=>"001000110",
  38228=>"011010011",
  38229=>"110010111",
  38230=>"000011110",
  38231=>"110101101",
  38232=>"111010111",
  38233=>"101001111",
  38234=>"001001111",
  38235=>"110011000",
  38236=>"010001001",
  38237=>"001001011",
  38238=>"010000011",
  38239=>"111100011",
  38240=>"110110000",
  38241=>"110011110",
  38242=>"111111011",
  38243=>"010010010",
  38244=>"000100011",
  38245=>"011011010",
  38246=>"101111010",
  38247=>"001010111",
  38248=>"110000001",
  38249=>"000101010",
  38250=>"010001001",
  38251=>"100011010",
  38252=>"001010110",
  38253=>"000101101",
  38254=>"010100100",
  38255=>"111110110",
  38256=>"111001011",
  38257=>"100111001",
  38258=>"011100000",
  38259=>"110111111",
  38260=>"111010011",
  38261=>"010101110",
  38262=>"001111110",
  38263=>"111111001",
  38264=>"110011111",
  38265=>"110011100",
  38266=>"110100110",
  38267=>"101011010",
  38268=>"100111001",
  38269=>"110111110",
  38270=>"000110110",
  38271=>"101101111",
  38272=>"101101100",
  38273=>"001100100",
  38274=>"000010100",
  38275=>"100001011",
  38276=>"100010011",
  38277=>"000000000",
  38278=>"100000000",
  38279=>"001000001",
  38280=>"110111001",
  38281=>"100101101",
  38282=>"010101100",
  38283=>"111100000",
  38284=>"000110000",
  38285=>"001011111",
  38286=>"001110011",
  38287=>"111110000",
  38288=>"111000100",
  38289=>"010101010",
  38290=>"000100111",
  38291=>"110111101",
  38292=>"000001111",
  38293=>"011101011",
  38294=>"001101000",
  38295=>"011010000",
  38296=>"010101000",
  38297=>"110011111",
  38298=>"010101101",
  38299=>"100101001",
  38300=>"011000010",
  38301=>"100110100",
  38302=>"101111110",
  38303=>"110110011",
  38304=>"101011001",
  38305=>"010110111",
  38306=>"010000111",
  38307=>"101111010",
  38308=>"101111110",
  38309=>"100000101",
  38310=>"001111101",
  38311=>"001101111",
  38312=>"001101010",
  38313=>"111111011",
  38314=>"001010110",
  38315=>"000001101",
  38316=>"100000010",
  38317=>"101110111",
  38318=>"110110101",
  38319=>"010011111",
  38320=>"110110110",
  38321=>"110101001",
  38322=>"101101100",
  38323=>"100110111",
  38324=>"000100101",
  38325=>"000110100",
  38326=>"011011101",
  38327=>"100111000",
  38328=>"010001101",
  38329=>"010011111",
  38330=>"100111010",
  38331=>"111001010",
  38332=>"010001101",
  38333=>"110111101",
  38334=>"110010111",
  38335=>"101000110",
  38336=>"100110001",
  38337=>"100000000",
  38338=>"000110000",
  38339=>"101110111",
  38340=>"110110001",
  38341=>"001101011",
  38342=>"011110111",
  38343=>"101000111",
  38344=>"000010100",
  38345=>"100010000",
  38346=>"111100110",
  38347=>"000010011",
  38348=>"010111100",
  38349=>"010000010",
  38350=>"101110010",
  38351=>"110101110",
  38352=>"111110000",
  38353=>"010101110",
  38354=>"110110100",
  38355=>"110011110",
  38356=>"010101111",
  38357=>"010000000",
  38358=>"100110001",
  38359=>"000101010",
  38360=>"110011101",
  38361=>"110110110",
  38362=>"110000000",
  38363=>"101111101",
  38364=>"000001000",
  38365=>"011110100",
  38366=>"011101010",
  38367=>"000001010",
  38368=>"010111101",
  38369=>"111000100",
  38370=>"000111010",
  38371=>"101100010",
  38372=>"100010010",
  38373=>"000111010",
  38374=>"100010110",
  38375=>"000010001",
  38376=>"001110110",
  38377=>"111011011",
  38378=>"101011011",
  38379=>"100011001",
  38380=>"000111111",
  38381=>"000011001",
  38382=>"110001100",
  38383=>"010100010",
  38384=>"001110000",
  38385=>"100110101",
  38386=>"101000100",
  38387=>"101111101",
  38388=>"101101011",
  38389=>"010110111",
  38390=>"001110001",
  38391=>"011100100",
  38392=>"100100101",
  38393=>"000101111",
  38394=>"111101100",
  38395=>"110010100",
  38396=>"111101011",
  38397=>"010110100",
  38398=>"110010001",
  38399=>"110000100",
  38400=>"110011010",
  38401=>"101101010",
  38402=>"100100101",
  38403=>"100110001",
  38404=>"111000000",
  38405=>"110011111",
  38406=>"100100100",
  38407=>"100110001",
  38408=>"000001100",
  38409=>"111100110",
  38410=>"010010100",
  38411=>"110101001",
  38412=>"111111101",
  38413=>"001001010",
  38414=>"101001111",
  38415=>"000011110",
  38416=>"010010011",
  38417=>"100001010",
  38418=>"000100000",
  38419=>"001010100",
  38420=>"000011100",
  38421=>"111111100",
  38422=>"011011000",
  38423=>"110101101",
  38424=>"111110011",
  38425=>"110110000",
  38426=>"110000100",
  38427=>"001110001",
  38428=>"100101100",
  38429=>"011000000",
  38430=>"101110001",
  38431=>"110011101",
  38432=>"000100111",
  38433=>"101011010",
  38434=>"001011001",
  38435=>"010001010",
  38436=>"100100010",
  38437=>"001100101",
  38438=>"001000011",
  38439=>"010111111",
  38440=>"101111110",
  38441=>"100111110",
  38442=>"001101011",
  38443=>"000011110",
  38444=>"011111101",
  38445=>"110001001",
  38446=>"010110000",
  38447=>"110001110",
  38448=>"111001110",
  38449=>"010011101",
  38450=>"010101111",
  38451=>"111110111",
  38452=>"110101110",
  38453=>"110111100",
  38454=>"000011110",
  38455=>"110000010",
  38456=>"100101011",
  38457=>"000110000",
  38458=>"110011010",
  38459=>"101000000",
  38460=>"101000100",
  38461=>"111101010",
  38462=>"101111011",
  38463=>"010110101",
  38464=>"000000001",
  38465=>"000001001",
  38466=>"010000100",
  38467=>"110111011",
  38468=>"111111100",
  38469=>"110001000",
  38470=>"110001011",
  38471=>"110000000",
  38472=>"010100110",
  38473=>"010000001",
  38474=>"010000010",
  38475=>"001000011",
  38476=>"000010100",
  38477=>"000000101",
  38478=>"110001010",
  38479=>"110101110",
  38480=>"000011111",
  38481=>"100001100",
  38482=>"110000010",
  38483=>"011000001",
  38484=>"001000010",
  38485=>"001010001",
  38486=>"101101001",
  38487=>"100101011",
  38488=>"111101111",
  38489=>"101011011",
  38490=>"000000111",
  38491=>"010011101",
  38492=>"010000110",
  38493=>"011001010",
  38494=>"111010001",
  38495=>"010111000",
  38496=>"100010111",
  38497=>"100110100",
  38498=>"100001101",
  38499=>"110010010",
  38500=>"100000010",
  38501=>"000101110",
  38502=>"111100111",
  38503=>"000011101",
  38504=>"101101101",
  38505=>"101110001",
  38506=>"000101010",
  38507=>"101011110",
  38508=>"000000110",
  38509=>"011011111",
  38510=>"010001111",
  38511=>"110111001",
  38512=>"000100000",
  38513=>"101111010",
  38514=>"111001111",
  38515=>"111111000",
  38516=>"101100101",
  38517=>"011100111",
  38518=>"000000010",
  38519=>"100011100",
  38520=>"100110010",
  38521=>"001100100",
  38522=>"001000001",
  38523=>"100110000",
  38524=>"010111110",
  38525=>"100101111",
  38526=>"110010010",
  38527=>"110101010",
  38528=>"010010101",
  38529=>"000111101",
  38530=>"010010100",
  38531=>"011111100",
  38532=>"010111011",
  38533=>"110011110",
  38534=>"101111100",
  38535=>"000000001",
  38536=>"100101110",
  38537=>"100001110",
  38538=>"011101011",
  38539=>"011010110",
  38540=>"001110010",
  38541=>"110001111",
  38542=>"110000000",
  38543=>"011011011",
  38544=>"000000000",
  38545=>"000110010",
  38546=>"000001111",
  38547=>"100001111",
  38548=>"100110111",
  38549=>"101111100",
  38550=>"101010111",
  38551=>"111011010",
  38552=>"001010100",
  38553=>"010000000",
  38554=>"000011110",
  38555=>"100101010",
  38556=>"101110100",
  38557=>"111110110",
  38558=>"110100001",
  38559=>"111101101",
  38560=>"000110101",
  38561=>"100010010",
  38562=>"110011100",
  38563=>"100000001",
  38564=>"011011110",
  38565=>"000110011",
  38566=>"110000001",
  38567=>"011000000",
  38568=>"111111101",
  38569=>"110100100",
  38570=>"011100111",
  38571=>"010010000",
  38572=>"001100011",
  38573=>"010111000",
  38574=>"101001101",
  38575=>"111010000",
  38576=>"000111100",
  38577=>"111101111",
  38578=>"100111111",
  38579=>"110000000",
  38580=>"011000101",
  38581=>"101011010",
  38582=>"100100100",
  38583=>"111100000",
  38584=>"101100001",
  38585=>"110010010",
  38586=>"110000010",
  38587=>"001001111",
  38588=>"100100000",
  38589=>"111100100",
  38590=>"110110000",
  38591=>"010111001",
  38592=>"111111010",
  38593=>"110110110",
  38594=>"111110010",
  38595=>"010100111",
  38596=>"110100001",
  38597=>"100111000",
  38598=>"111101110",
  38599=>"111001100",
  38600=>"100111111",
  38601=>"000111111",
  38602=>"111101110",
  38603=>"000000110",
  38604=>"010110010",
  38605=>"010100100",
  38606=>"100111011",
  38607=>"111110111",
  38608=>"011011111",
  38609=>"110001100",
  38610=>"000111001",
  38611=>"010010010",
  38612=>"101011001",
  38613=>"001100101",
  38614=>"100011101",
  38615=>"000011011",
  38616=>"001100010",
  38617=>"000011000",
  38618=>"001000101",
  38619=>"111001000",
  38620=>"001011110",
  38621=>"011111100",
  38622=>"111000001",
  38623=>"010010001",
  38624=>"110100111",
  38625=>"011011000",
  38626=>"110011101",
  38627=>"101101100",
  38628=>"110110000",
  38629=>"011001001",
  38630=>"011000101",
  38631=>"011110000",
  38632=>"111110110",
  38633=>"100000100",
  38634=>"001101110",
  38635=>"001110001",
  38636=>"011111000",
  38637=>"001110010",
  38638=>"101110001",
  38639=>"001100000",
  38640=>"110110001",
  38641=>"100111110",
  38642=>"111110000",
  38643=>"011001100",
  38644=>"011101001",
  38645=>"010000110",
  38646=>"100110101",
  38647=>"011011111",
  38648=>"101101000",
  38649=>"000100001",
  38650=>"110001000",
  38651=>"100110110",
  38652=>"011010010",
  38653=>"111100110",
  38654=>"101001011",
  38655=>"000010100",
  38656=>"010111010",
  38657=>"110010010",
  38658=>"010100100",
  38659=>"100000011",
  38660=>"000011110",
  38661=>"101001000",
  38662=>"011110011",
  38663=>"001001011",
  38664=>"000100101",
  38665=>"011101100",
  38666=>"100100001",
  38667=>"110001100",
  38668=>"010101010",
  38669=>"000000111",
  38670=>"100000100",
  38671=>"101110100",
  38672=>"111100110",
  38673=>"000000010",
  38674=>"101011100",
  38675=>"001011011",
  38676=>"111001001",
  38677=>"010010010",
  38678=>"010010000",
  38679=>"010100000",
  38680=>"111100111",
  38681=>"011101110",
  38682=>"011111010",
  38683=>"001010100",
  38684=>"011111101",
  38685=>"001100101",
  38686=>"101101011",
  38687=>"000110000",
  38688=>"000000101",
  38689=>"111101010",
  38690=>"111001100",
  38691=>"111101010",
  38692=>"001010111",
  38693=>"100000001",
  38694=>"101101001",
  38695=>"000011111",
  38696=>"110011111",
  38697=>"000000111",
  38698=>"010011000",
  38699=>"111010011",
  38700=>"100111011",
  38701=>"111110010",
  38702=>"000100001",
  38703=>"100011001",
  38704=>"111001111",
  38705=>"010010000",
  38706=>"111000011",
  38707=>"101110011",
  38708=>"110011000",
  38709=>"011101010",
  38710=>"011111111",
  38711=>"010110001",
  38712=>"010111110",
  38713=>"001001101",
  38714=>"110011110",
  38715=>"111110100",
  38716=>"111000000",
  38717=>"111101111",
  38718=>"100000010",
  38719=>"011101001",
  38720=>"110011011",
  38721=>"111101111",
  38722=>"011001111",
  38723=>"100111101",
  38724=>"100000100",
  38725=>"100101011",
  38726=>"111101111",
  38727=>"110001111",
  38728=>"110011100",
  38729=>"001000101",
  38730=>"101010101",
  38731=>"110010110",
  38732=>"000000010",
  38733=>"001001100",
  38734=>"001110011",
  38735=>"011111000",
  38736=>"100111101",
  38737=>"000100001",
  38738=>"001010101",
  38739=>"111001101",
  38740=>"001001010",
  38741=>"100101100",
  38742=>"101011001",
  38743=>"010110101",
  38744=>"010000101",
  38745=>"111101111",
  38746=>"011000110",
  38747=>"111110011",
  38748=>"111100001",
  38749=>"111000001",
  38750=>"110011101",
  38751=>"100000100",
  38752=>"100110100",
  38753=>"010110100",
  38754=>"110100010",
  38755=>"010010100",
  38756=>"111001111",
  38757=>"101100011",
  38758=>"000101010",
  38759=>"010110010",
  38760=>"001010010",
  38761=>"110000100",
  38762=>"110101101",
  38763=>"010001101",
  38764=>"100010100",
  38765=>"111000001",
  38766=>"011100100",
  38767=>"101001001",
  38768=>"111111010",
  38769=>"000010100",
  38770=>"000110000",
  38771=>"001001010",
  38772=>"100011001",
  38773=>"001000010",
  38774=>"000001010",
  38775=>"011110011",
  38776=>"101001010",
  38777=>"100110010",
  38778=>"000001011",
  38779=>"011001100",
  38780=>"111010001",
  38781=>"001101111",
  38782=>"101100001",
  38783=>"001000001",
  38784=>"001010111",
  38785=>"101111110",
  38786=>"010000000",
  38787=>"111001000",
  38788=>"101110000",
  38789=>"001010111",
  38790=>"111111111",
  38791=>"101010000",
  38792=>"011010111",
  38793=>"001101111",
  38794=>"111011011",
  38795=>"000101111",
  38796=>"111110110",
  38797=>"011000111",
  38798=>"101101101",
  38799=>"111111001",
  38800=>"001100001",
  38801=>"010010100",
  38802=>"100100010",
  38803=>"010100100",
  38804=>"110110001",
  38805=>"000111011",
  38806=>"010110100",
  38807=>"111010110",
  38808=>"001011000",
  38809=>"101000010",
  38810=>"000110100",
  38811=>"110010011",
  38812=>"011101010",
  38813=>"110111010",
  38814=>"100000101",
  38815=>"110110101",
  38816=>"011010011",
  38817=>"011011111",
  38818=>"101000110",
  38819=>"001000010",
  38820=>"100101011",
  38821=>"100001011",
  38822=>"111001100",
  38823=>"101001001",
  38824=>"000111000",
  38825=>"001001111",
  38826=>"110111000",
  38827=>"110000000",
  38828=>"111110110",
  38829=>"110101010",
  38830=>"001001111",
  38831=>"110011000",
  38832=>"000010100",
  38833=>"110010000",
  38834=>"110101111",
  38835=>"110010010",
  38836=>"001100100",
  38837=>"000111110",
  38838=>"101010000",
  38839=>"000010111",
  38840=>"011011001",
  38841=>"000011001",
  38842=>"111010100",
  38843=>"111101010",
  38844=>"101111001",
  38845=>"111000001",
  38846=>"011111110",
  38847=>"001100000",
  38848=>"101100110",
  38849=>"100111100",
  38850=>"000110000",
  38851=>"111100010",
  38852=>"111101110",
  38853=>"011100111",
  38854=>"110001010",
  38855=>"100111001",
  38856=>"111110111",
  38857=>"100001001",
  38858=>"011001000",
  38859=>"101100010",
  38860=>"111001000",
  38861=>"001110001",
  38862=>"011110100",
  38863=>"110001101",
  38864=>"110111001",
  38865=>"010101110",
  38866=>"111110110",
  38867=>"101000001",
  38868=>"010010001",
  38869=>"110001101",
  38870=>"100011101",
  38871=>"101110010",
  38872=>"110010001",
  38873=>"101110000",
  38874=>"110111111",
  38875=>"010000100",
  38876=>"110000100",
  38877=>"111101111",
  38878=>"111011010",
  38879=>"111100011",
  38880=>"101110000",
  38881=>"110001000",
  38882=>"111100011",
  38883=>"100000000",
  38884=>"111101001",
  38885=>"101001101",
  38886=>"111101101",
  38887=>"010111111",
  38888=>"000111001",
  38889=>"111000110",
  38890=>"001010000",
  38891=>"110110110",
  38892=>"011011010",
  38893=>"000100010",
  38894=>"111011010",
  38895=>"111101010",
  38896=>"001000000",
  38897=>"110010110",
  38898=>"101011001",
  38899=>"101101111",
  38900=>"111011110",
  38901=>"111100011",
  38902=>"111011001",
  38903=>"000010101",
  38904=>"011001100",
  38905=>"111000111",
  38906=>"110100100",
  38907=>"001100101",
  38908=>"110001100",
  38909=>"001010010",
  38910=>"101011110",
  38911=>"010011011",
  38912=>"010000001",
  38913=>"111100000",
  38914=>"101001000",
  38915=>"011010000",
  38916=>"101100111",
  38917=>"011111010",
  38918=>"001000100",
  38919=>"011110010",
  38920=>"011111110",
  38921=>"100100000",
  38922=>"101111100",
  38923=>"100111100",
  38924=>"001101100",
  38925=>"110111101",
  38926=>"001111111",
  38927=>"110011101",
  38928=>"111010101",
  38929=>"110010100",
  38930=>"101010010",
  38931=>"011111110",
  38932=>"111110111",
  38933=>"100010100",
  38934=>"010111001",
  38935=>"111110111",
  38936=>"101100101",
  38937=>"100111101",
  38938=>"110100000",
  38939=>"111100100",
  38940=>"111101101",
  38941=>"100111001",
  38942=>"010101000",
  38943=>"010010000",
  38944=>"001101101",
  38945=>"101110101",
  38946=>"111111000",
  38947=>"011111010",
  38948=>"000101110",
  38949=>"011110010",
  38950=>"010001111",
  38951=>"100101011",
  38952=>"001111000",
  38953=>"011010101",
  38954=>"111011011",
  38955=>"000001010",
  38956=>"101001011",
  38957=>"110011111",
  38958=>"110010110",
  38959=>"110010011",
  38960=>"111110110",
  38961=>"111010010",
  38962=>"011101100",
  38963=>"100100001",
  38964=>"110100110",
  38965=>"010001110",
  38966=>"000100000",
  38967=>"000100011",
  38968=>"100100100",
  38969=>"100111000",
  38970=>"010111011",
  38971=>"100000101",
  38972=>"001010111",
  38973=>"100101001",
  38974=>"111000111",
  38975=>"101010000",
  38976=>"100000100",
  38977=>"000001000",
  38978=>"001010001",
  38979=>"100111100",
  38980=>"110001111",
  38981=>"111100011",
  38982=>"101111000",
  38983=>"100001000",
  38984=>"101101100",
  38985=>"011011101",
  38986=>"001000100",
  38987=>"111100011",
  38988=>"001000010",
  38989=>"110011010",
  38990=>"101000110",
  38991=>"000100100",
  38992=>"000001111",
  38993=>"101101001",
  38994=>"010001111",
  38995=>"010011001",
  38996=>"001110010",
  38997=>"110010100",
  38998=>"010001101",
  38999=>"011010101",
  39000=>"010011011",
  39001=>"110000000",
  39002=>"011110110",
  39003=>"111110001",
  39004=>"011001001",
  39005=>"011101101",
  39006=>"010010110",
  39007=>"011000011",
  39008=>"100100000",
  39009=>"010100100",
  39010=>"100000110",
  39011=>"011000001",
  39012=>"011110110",
  39013=>"011011010",
  39014=>"010111011",
  39015=>"111000110",
  39016=>"111001011",
  39017=>"001110100",
  39018=>"010001110",
  39019=>"011101101",
  39020=>"110111010",
  39021=>"011100111",
  39022=>"100111100",
  39023=>"001100010",
  39024=>"010100011",
  39025=>"110000100",
  39026=>"111110010",
  39027=>"111111001",
  39028=>"011000011",
  39029=>"111001101",
  39030=>"010010101",
  39031=>"010101000",
  39032=>"110011110",
  39033=>"010111001",
  39034=>"000100100",
  39035=>"111101001",
  39036=>"001010110",
  39037=>"111001100",
  39038=>"010011000",
  39039=>"011111010",
  39040=>"110000110",
  39041=>"010100010",
  39042=>"001000011",
  39043=>"001110001",
  39044=>"010100011",
  39045=>"100101000",
  39046=>"110101110",
  39047=>"000100100",
  39048=>"110000101",
  39049=>"111010000",
  39050=>"010110011",
  39051=>"000111010",
  39052=>"011111110",
  39053=>"100011111",
  39054=>"101101100",
  39055=>"100010011",
  39056=>"111101011",
  39057=>"001100011",
  39058=>"011000011",
  39059=>"101010010",
  39060=>"100100100",
  39061=>"010011110",
  39062=>"010001111",
  39063=>"110010101",
  39064=>"101000001",
  39065=>"101010010",
  39066=>"100001111",
  39067=>"101001100",
  39068=>"100101000",
  39069=>"011100000",
  39070=>"000111111",
  39071=>"011001111",
  39072=>"000111001",
  39073=>"110011110",
  39074=>"010101000",
  39075=>"010000000",
  39076=>"111111001",
  39077=>"100000000",
  39078=>"111010111",
  39079=>"100100101",
  39080=>"000100110",
  39081=>"000011011",
  39082=>"101011110",
  39083=>"100111110",
  39084=>"110111010",
  39085=>"000100000",
  39086=>"011100010",
  39087=>"101110011",
  39088=>"011110010",
  39089=>"000111110",
  39090=>"111001101",
  39091=>"010111111",
  39092=>"110101110",
  39093=>"000001000",
  39094=>"001100100",
  39095=>"010011000",
  39096=>"000111100",
  39097=>"001010101",
  39098=>"010001101",
  39099=>"111111001",
  39100=>"111010001",
  39101=>"001111100",
  39102=>"111100000",
  39103=>"000100000",
  39104=>"000011010",
  39105=>"010011100",
  39106=>"010000000",
  39107=>"011000110",
  39108=>"010111001",
  39109=>"101100001",
  39110=>"011111001",
  39111=>"100010011",
  39112=>"100000000",
  39113=>"011011101",
  39114=>"000010000",
  39115=>"001000011",
  39116=>"100111010",
  39117=>"001011011",
  39118=>"001001110",
  39119=>"101111110",
  39120=>"001111010",
  39121=>"001000111",
  39122=>"100100000",
  39123=>"000100011",
  39124=>"100101100",
  39125=>"101111110",
  39126=>"001001000",
  39127=>"110110011",
  39128=>"100001111",
  39129=>"100111100",
  39130=>"111110100",
  39131=>"001000101",
  39132=>"101010111",
  39133=>"001011110",
  39134=>"100001101",
  39135=>"001010100",
  39136=>"111101101",
  39137=>"111111110",
  39138=>"011100100",
  39139=>"010010000",
  39140=>"101111101",
  39141=>"101100001",
  39142=>"101101101",
  39143=>"111110111",
  39144=>"000100011",
  39145=>"111100000",
  39146=>"011100110",
  39147=>"100001011",
  39148=>"100000011",
  39149=>"001001011",
  39150=>"001001110",
  39151=>"110110111",
  39152=>"000000110",
  39153=>"001001000",
  39154=>"110011010",
  39155=>"010100000",
  39156=>"101011100",
  39157=>"100000001",
  39158=>"011111110",
  39159=>"010000010",
  39160=>"110111110",
  39161=>"001000110",
  39162=>"111101011",
  39163=>"101100001",
  39164=>"011101001",
  39165=>"101110100",
  39166=>"100000010",
  39167=>"001011101",
  39168=>"111011011",
  39169=>"110011011",
  39170=>"111000101",
  39171=>"000011100",
  39172=>"110001100",
  39173=>"011101110",
  39174=>"100001101",
  39175=>"100001001",
  39176=>"100100100",
  39177=>"101110010",
  39178=>"000100100",
  39179=>"101101000",
  39180=>"000010010",
  39181=>"011000110",
  39182=>"110011000",
  39183=>"001011101",
  39184=>"000001011",
  39185=>"001101010",
  39186=>"000101001",
  39187=>"001001110",
  39188=>"010101010",
  39189=>"101101000",
  39190=>"011111111",
  39191=>"001111001",
  39192=>"011001001",
  39193=>"010000100",
  39194=>"010001000",
  39195=>"101111110",
  39196=>"010000011",
  39197=>"001011110",
  39198=>"011111001",
  39199=>"010000110",
  39200=>"011100100",
  39201=>"101100011",
  39202=>"101111111",
  39203=>"101010010",
  39204=>"001101010",
  39205=>"100110011",
  39206=>"000101000",
  39207=>"111000110",
  39208=>"100000010",
  39209=>"101101110",
  39210=>"000110010",
  39211=>"111100110",
  39212=>"100100010",
  39213=>"010100010",
  39214=>"000010010",
  39215=>"100000001",
  39216=>"010101011",
  39217=>"101000111",
  39218=>"001110101",
  39219=>"000111100",
  39220=>"100101101",
  39221=>"100001011",
  39222=>"111010101",
  39223=>"000101101",
  39224=>"010000110",
  39225=>"010001111",
  39226=>"001100000",
  39227=>"110101100",
  39228=>"010100100",
  39229=>"101111100",
  39230=>"110010101",
  39231=>"001000011",
  39232=>"101110111",
  39233=>"001000101",
  39234=>"010100011",
  39235=>"010101101",
  39236=>"101110001",
  39237=>"100101100",
  39238=>"001100001",
  39239=>"100000111",
  39240=>"011110100",
  39241=>"110111111",
  39242=>"101001011",
  39243=>"111010010",
  39244=>"001100111",
  39245=>"100001010",
  39246=>"011010110",
  39247=>"111111101",
  39248=>"001000110",
  39249=>"110110010",
  39250=>"100101011",
  39251=>"000001011",
  39252=>"000001110",
  39253=>"000111111",
  39254=>"001000000",
  39255=>"010010011",
  39256=>"010100010",
  39257=>"000010111",
  39258=>"010110111",
  39259=>"001100000",
  39260=>"110000001",
  39261=>"101011100",
  39262=>"100111011",
  39263=>"110010010",
  39264=>"011001011",
  39265=>"101000111",
  39266=>"011000010",
  39267=>"101101000",
  39268=>"011110011",
  39269=>"010011111",
  39270=>"001011111",
  39271=>"110000011",
  39272=>"101000000",
  39273=>"010110101",
  39274=>"010001000",
  39275=>"000000101",
  39276=>"011000011",
  39277=>"111111100",
  39278=>"100011111",
  39279=>"000110101",
  39280=>"111110000",
  39281=>"100000100",
  39282=>"011011110",
  39283=>"101010101",
  39284=>"100000011",
  39285=>"101001100",
  39286=>"110110000",
  39287=>"011010101",
  39288=>"000100100",
  39289=>"101001000",
  39290=>"111101111",
  39291=>"110101111",
  39292=>"000000001",
  39293=>"010101001",
  39294=>"110000010",
  39295=>"011010000",
  39296=>"000010110",
  39297=>"101001101",
  39298=>"110010000",
  39299=>"001001101",
  39300=>"101010000",
  39301=>"011110000",
  39302=>"100101011",
  39303=>"001001111",
  39304=>"111001101",
  39305=>"001111110",
  39306=>"101101000",
  39307=>"100010000",
  39308=>"010111001",
  39309=>"111010000",
  39310=>"011011101",
  39311=>"001111111",
  39312=>"111000011",
  39313=>"010000000",
  39314=>"000011000",
  39315=>"111001010",
  39316=>"011011111",
  39317=>"010001000",
  39318=>"000010000",
  39319=>"000001000",
  39320=>"010000000",
  39321=>"010011100",
  39322=>"111011001",
  39323=>"011111111",
  39324=>"000001111",
  39325=>"101110010",
  39326=>"111101011",
  39327=>"001011100",
  39328=>"011101110",
  39329=>"001010100",
  39330=>"110101101",
  39331=>"110110010",
  39332=>"000010110",
  39333=>"111110111",
  39334=>"011101001",
  39335=>"110001101",
  39336=>"001100011",
  39337=>"100010111",
  39338=>"101000111",
  39339=>"111011101",
  39340=>"000111000",
  39341=>"010101111",
  39342=>"001000111",
  39343=>"000010100",
  39344=>"011110011",
  39345=>"110111000",
  39346=>"110101110",
  39347=>"001010001",
  39348=>"011010101",
  39349=>"111001010",
  39350=>"111000010",
  39351=>"111101000",
  39352=>"001010010",
  39353=>"110010011",
  39354=>"101000010",
  39355=>"101001111",
  39356=>"110010010",
  39357=>"101100111",
  39358=>"100100101",
  39359=>"010010101",
  39360=>"111001000",
  39361=>"111111111",
  39362=>"001111110",
  39363=>"000100101",
  39364=>"100010001",
  39365=>"110011000",
  39366=>"100000011",
  39367=>"010011011",
  39368=>"101011011",
  39369=>"100000001",
  39370=>"110100111",
  39371=>"110100000",
  39372=>"001000100",
  39373=>"101111001",
  39374=>"100101111",
  39375=>"001000010",
  39376=>"000110110",
  39377=>"000111101",
  39378=>"011010100",
  39379=>"101010001",
  39380=>"101001100",
  39381=>"010101001",
  39382=>"000101000",
  39383=>"011011100",
  39384=>"000110100",
  39385=>"111000101",
  39386=>"010011001",
  39387=>"010010110",
  39388=>"111111100",
  39389=>"000101111",
  39390=>"000000010",
  39391=>"110101000",
  39392=>"111011011",
  39393=>"100011110",
  39394=>"110100010",
  39395=>"000100100",
  39396=>"001001110",
  39397=>"000101000",
  39398=>"001000000",
  39399=>"011011100",
  39400=>"001101100",
  39401=>"111101110",
  39402=>"010001001",
  39403=>"110011111",
  39404=>"111011100",
  39405=>"000000110",
  39406=>"011010010",
  39407=>"010011110",
  39408=>"011111100",
  39409=>"011101100",
  39410=>"110010000",
  39411=>"011010000",
  39412=>"110000110",
  39413=>"101100010",
  39414=>"001000011",
  39415=>"110011111",
  39416=>"111110111",
  39417=>"011011101",
  39418=>"100100100",
  39419=>"110110011",
  39420=>"101000110",
  39421=>"000001100",
  39422=>"010010001",
  39423=>"000100100",
  39424=>"001011100",
  39425=>"110010001",
  39426=>"001000000",
  39427=>"011000110",
  39428=>"110011111",
  39429=>"111100000",
  39430=>"111011001",
  39431=>"000101100",
  39432=>"011011000",
  39433=>"111010010",
  39434=>"000001011",
  39435=>"001101100",
  39436=>"010110101",
  39437=>"001011100",
  39438=>"000011011",
  39439=>"100110011",
  39440=>"101101011",
  39441=>"011010010",
  39442=>"010110010",
  39443=>"001110101",
  39444=>"000000101",
  39445=>"001101100",
  39446=>"001001010",
  39447=>"101011110",
  39448=>"111101111",
  39449=>"100101111",
  39450=>"100100100",
  39451=>"010011111",
  39452=>"101111110",
  39453=>"110001101",
  39454=>"100010111",
  39455=>"011011000",
  39456=>"000011000",
  39457=>"000011010",
  39458=>"001000000",
  39459=>"100111101",
  39460=>"111100001",
  39461=>"011101100",
  39462=>"001100010",
  39463=>"110011011",
  39464=>"010001111",
  39465=>"110111110",
  39466=>"111110100",
  39467=>"101111101",
  39468=>"011000100",
  39469=>"111100000",
  39470=>"000110000",
  39471=>"001110101",
  39472=>"011000111",
  39473=>"000001010",
  39474=>"001110101",
  39475=>"001101001",
  39476=>"100010101",
  39477=>"011010001",
  39478=>"000101100",
  39479=>"111000101",
  39480=>"011111000",
  39481=>"100000101",
  39482=>"001010101",
  39483=>"111011001",
  39484=>"011000111",
  39485=>"100000010",
  39486=>"110010001",
  39487=>"110110111",
  39488=>"101101110",
  39489=>"011010111",
  39490=>"111110101",
  39491=>"011111110",
  39492=>"001011010",
  39493=>"101101110",
  39494=>"100110110",
  39495=>"111110101",
  39496=>"001110000",
  39497=>"011000000",
  39498=>"101111111",
  39499=>"101101011",
  39500=>"001110100",
  39501=>"001011100",
  39502=>"011011000",
  39503=>"110001100",
  39504=>"000100011",
  39505=>"101011001",
  39506=>"000010001",
  39507=>"111101111",
  39508=>"100011001",
  39509=>"000001111",
  39510=>"101011110",
  39511=>"110010100",
  39512=>"000101000",
  39513=>"010010000",
  39514=>"001011100",
  39515=>"110001100",
  39516=>"010100100",
  39517=>"010000000",
  39518=>"100011100",
  39519=>"000010110",
  39520=>"001101111",
  39521=>"000000001",
  39522=>"010000111",
  39523=>"110011110",
  39524=>"000110000",
  39525=>"011010000",
  39526=>"000001101",
  39527=>"110001000",
  39528=>"101000100",
  39529=>"011101101",
  39530=>"011011110",
  39531=>"010011010",
  39532=>"100110010",
  39533=>"110000111",
  39534=>"010000011",
  39535=>"111001110",
  39536=>"100110000",
  39537=>"111011101",
  39538=>"001100111",
  39539=>"011111011",
  39540=>"101110100",
  39541=>"011010111",
  39542=>"011011110",
  39543=>"111011011",
  39544=>"100010100",
  39545=>"010101001",
  39546=>"100111010",
  39547=>"010100000",
  39548=>"100010000",
  39549=>"011101101",
  39550=>"010100001",
  39551=>"010101010",
  39552=>"001000111",
  39553=>"110000001",
  39554=>"101000101",
  39555=>"100100101",
  39556=>"011100011",
  39557=>"001111000",
  39558=>"010001001",
  39559=>"101001000",
  39560=>"000000000",
  39561=>"011110111",
  39562=>"000010010",
  39563=>"010001100",
  39564=>"001000000",
  39565=>"100110100",
  39566=>"001011100",
  39567=>"111101000",
  39568=>"011111001",
  39569=>"001010000",
  39570=>"111111101",
  39571=>"001011111",
  39572=>"110001010",
  39573=>"011111011",
  39574=>"100000011",
  39575=>"111010101",
  39576=>"000101001",
  39577=>"110000011",
  39578=>"101110001",
  39579=>"110000111",
  39580=>"110111111",
  39581=>"001001111",
  39582=>"000110100",
  39583=>"000010011",
  39584=>"000111111",
  39585=>"001101001",
  39586=>"000100111",
  39587=>"111000011",
  39588=>"110110011",
  39589=>"110000101",
  39590=>"000111011",
  39591=>"011010010",
  39592=>"100111001",
  39593=>"100001010",
  39594=>"001011011",
  39595=>"000111101",
  39596=>"100110001",
  39597=>"111001001",
  39598=>"111101011",
  39599=>"001000101",
  39600=>"000000110",
  39601=>"111000101",
  39602=>"110110111",
  39603=>"111110010",
  39604=>"010111000",
  39605=>"111010010",
  39606=>"111001100",
  39607=>"110010010",
  39608=>"000001011",
  39609=>"101111111",
  39610=>"011110111",
  39611=>"100001110",
  39612=>"100011000",
  39613=>"111110101",
  39614=>"110110001",
  39615=>"111000111",
  39616=>"100111101",
  39617=>"101001111",
  39618=>"001010000",
  39619=>"010000000",
  39620=>"111001011",
  39621=>"001011001",
  39622=>"101111001",
  39623=>"110111000",
  39624=>"101100001",
  39625=>"001100101",
  39626=>"001011010",
  39627=>"010011000",
  39628=>"000001000",
  39629=>"010001101",
  39630=>"100010111",
  39631=>"111111001",
  39632=>"000011111",
  39633=>"000111101",
  39634=>"111100010",
  39635=>"101101100",
  39636=>"111110110",
  39637=>"100010111",
  39638=>"001111111",
  39639=>"110101001",
  39640=>"110001101",
  39641=>"000010000",
  39642=>"100001000",
  39643=>"011001111",
  39644=>"010011111",
  39645=>"111001010",
  39646=>"000111000",
  39647=>"100111011",
  39648=>"100001110",
  39649=>"110001001",
  39650=>"001101111",
  39651=>"100011001",
  39652=>"110110101",
  39653=>"001110000",
  39654=>"000001000",
  39655=>"001100000",
  39656=>"110100100",
  39657=>"111001100",
  39658=>"110010110",
  39659=>"100010011",
  39660=>"101001101",
  39661=>"110001000",
  39662=>"000100100",
  39663=>"001110110",
  39664=>"011110010",
  39665=>"111011001",
  39666=>"100110100",
  39667=>"110101110",
  39668=>"101010101",
  39669=>"110100101",
  39670=>"110010010",
  39671=>"000100010",
  39672=>"000001010",
  39673=>"100100111",
  39674=>"111001010",
  39675=>"011000111",
  39676=>"100101000",
  39677=>"011010111",
  39678=>"100000011",
  39679=>"000011100",
  39680=>"110110100",
  39681=>"000010101",
  39682=>"000111000",
  39683=>"010001101",
  39684=>"111110110",
  39685=>"000110000",
  39686=>"110000010",
  39687=>"011100000",
  39688=>"111100111",
  39689=>"010011100",
  39690=>"000001100",
  39691=>"010000010",
  39692=>"111111100",
  39693=>"100011100",
  39694=>"100001010",
  39695=>"100011001",
  39696=>"100001011",
  39697=>"010000011",
  39698=>"010001101",
  39699=>"000000101",
  39700=>"111011000",
  39701=>"110001110",
  39702=>"101010000",
  39703=>"100110010",
  39704=>"100000011",
  39705=>"000000100",
  39706=>"101011100",
  39707=>"000000111",
  39708=>"111000000",
  39709=>"100010110",
  39710=>"110111110",
  39711=>"100100010",
  39712=>"110111110",
  39713=>"011010110",
  39714=>"100000001",
  39715=>"000110101",
  39716=>"100101011",
  39717=>"110101010",
  39718=>"001011001",
  39719=>"111110011",
  39720=>"100000111",
  39721=>"101011100",
  39722=>"100011011",
  39723=>"101011110",
  39724=>"001100010",
  39725=>"110001111",
  39726=>"101111011",
  39727=>"110110111",
  39728=>"101100001",
  39729=>"111111010",
  39730=>"100011111",
  39731=>"001001100",
  39732=>"000110000",
  39733=>"100101011",
  39734=>"001101100",
  39735=>"100100000",
  39736=>"010101000",
  39737=>"101001100",
  39738=>"111101010",
  39739=>"010101011",
  39740=>"010000111",
  39741=>"110100000",
  39742=>"000000101",
  39743=>"100000101",
  39744=>"101000101",
  39745=>"111110001",
  39746=>"001011000",
  39747=>"010001000",
  39748=>"100000011",
  39749=>"010100101",
  39750=>"001000011",
  39751=>"010001111",
  39752=>"100100000",
  39753=>"001000011",
  39754=>"100100101",
  39755=>"001011010",
  39756=>"111101010",
  39757=>"110010100",
  39758=>"001111111",
  39759=>"100110110",
  39760=>"000111111",
  39761=>"000000000",
  39762=>"110110110",
  39763=>"010110110",
  39764=>"111111100",
  39765=>"101001010",
  39766=>"100100101",
  39767=>"001101010",
  39768=>"000001101",
  39769=>"111101001",
  39770=>"100101010",
  39771=>"111010100",
  39772=>"001010000",
  39773=>"010100111",
  39774=>"101100100",
  39775=>"100011011",
  39776=>"011111011",
  39777=>"101001011",
  39778=>"000000001",
  39779=>"111001001",
  39780=>"110111001",
  39781=>"001100010",
  39782=>"111011011",
  39783=>"100011111",
  39784=>"000000111",
  39785=>"111001011",
  39786=>"111111111",
  39787=>"100011001",
  39788=>"100100000",
  39789=>"000101011",
  39790=>"010001101",
  39791=>"111110110",
  39792=>"001110110",
  39793=>"101001011",
  39794=>"010010100",
  39795=>"001000010",
  39796=>"011001010",
  39797=>"001101000",
  39798=>"100110100",
  39799=>"000001100",
  39800=>"111111010",
  39801=>"001100111",
  39802=>"111011010",
  39803=>"011101001",
  39804=>"111111101",
  39805=>"111111010",
  39806=>"010011001",
  39807=>"110101101",
  39808=>"111110101",
  39809=>"011000010",
  39810=>"110101110",
  39811=>"110110001",
  39812=>"100101110",
  39813=>"010010111",
  39814=>"111101100",
  39815=>"100000100",
  39816=>"010111001",
  39817=>"110110000",
  39818=>"001101100",
  39819=>"000010000",
  39820=>"101000111",
  39821=>"110101111",
  39822=>"000111001",
  39823=>"111110110",
  39824=>"011001100",
  39825=>"001110100",
  39826=>"010101110",
  39827=>"011101101",
  39828=>"011000000",
  39829=>"111110110",
  39830=>"000001101",
  39831=>"000100110",
  39832=>"111011111",
  39833=>"101100100",
  39834=>"001101100",
  39835=>"011011100",
  39836=>"110010000",
  39837=>"011011000",
  39838=>"001010010",
  39839=>"010110100",
  39840=>"000110011",
  39841=>"010000011",
  39842=>"111001010",
  39843=>"110010101",
  39844=>"110110000",
  39845=>"101011111",
  39846=>"000100110",
  39847=>"100000101",
  39848=>"010100010",
  39849=>"110101010",
  39850=>"110101000",
  39851=>"101000000",
  39852=>"011010111",
  39853=>"100111010",
  39854=>"100101100",
  39855=>"010011101",
  39856=>"010101111",
  39857=>"111001101",
  39858=>"101001001",
  39859=>"001001100",
  39860=>"101111001",
  39861=>"000110100",
  39862=>"111111100",
  39863=>"011111001",
  39864=>"101010000",
  39865=>"100111000",
  39866=>"000100001",
  39867=>"001010011",
  39868=>"000000001",
  39869=>"010010110",
  39870=>"011011110",
  39871=>"011010001",
  39872=>"111111001",
  39873=>"100101000",
  39874=>"000101111",
  39875=>"100011010",
  39876=>"100111111",
  39877=>"110000011",
  39878=>"000000000",
  39879=>"110010100",
  39880=>"000010000",
  39881=>"100101011",
  39882=>"110000001",
  39883=>"100010010",
  39884=>"100111010",
  39885=>"000000000",
  39886=>"100101000",
  39887=>"001011101",
  39888=>"010101011",
  39889=>"001010000",
  39890=>"110111101",
  39891=>"101110100",
  39892=>"111010011",
  39893=>"110100001",
  39894=>"110000011",
  39895=>"001000000",
  39896=>"100010001",
  39897=>"011000011",
  39898=>"111010000",
  39899=>"111100011",
  39900=>"110010011",
  39901=>"100110000",
  39902=>"110110100",
  39903=>"101101010",
  39904=>"010100110",
  39905=>"011010101",
  39906=>"100011010",
  39907=>"001111101",
  39908=>"100001110",
  39909=>"101101111",
  39910=>"100101100",
  39911=>"011010111",
  39912=>"000001001",
  39913=>"101111111",
  39914=>"111010010",
  39915=>"110010101",
  39916=>"010000110",
  39917=>"110001101",
  39918=>"011100110",
  39919=>"001000010",
  39920=>"110001000",
  39921=>"111110101",
  39922=>"100000111",
  39923=>"101010011",
  39924=>"010010100",
  39925=>"001111101",
  39926=>"010110010",
  39927=>"100000010",
  39928=>"111101001",
  39929=>"101101111",
  39930=>"010111110",
  39931=>"000111010",
  39932=>"100110000",
  39933=>"111001110",
  39934=>"110101111",
  39935=>"110110100",
  39936=>"010000010",
  39937=>"110000110",
  39938=>"010100001",
  39939=>"110101111",
  39940=>"011111010",
  39941=>"000111110",
  39942=>"100100110",
  39943=>"101110001",
  39944=>"111000000",
  39945=>"011010110",
  39946=>"111000111",
  39947=>"001010110",
  39948=>"001111011",
  39949=>"110101100",
  39950=>"001101101",
  39951=>"101111101",
  39952=>"111001000",
  39953=>"000001011",
  39954=>"111000000",
  39955=>"101010111",
  39956=>"111101111",
  39957=>"011110100",
  39958=>"101010001",
  39959=>"101010111",
  39960=>"100001001",
  39961=>"011111011",
  39962=>"000010011",
  39963=>"011101011",
  39964=>"011101010",
  39965=>"010101010",
  39966=>"011011111",
  39967=>"011011000",
  39968=>"010000110",
  39969=>"111101000",
  39970=>"100101010",
  39971=>"100011100",
  39972=>"010111100",
  39973=>"000100101",
  39974=>"001000011",
  39975=>"011011001",
  39976=>"011000110",
  39977=>"000001000",
  39978=>"110011000",
  39979=>"001111101",
  39980=>"111000110",
  39981=>"000001100",
  39982=>"011101011",
  39983=>"100101001",
  39984=>"011101110",
  39985=>"111010010",
  39986=>"010111001",
  39987=>"110101011",
  39988=>"111010101",
  39989=>"000100010",
  39990=>"111011100",
  39991=>"001101101",
  39992=>"101101000",
  39993=>"111101100",
  39994=>"110111111",
  39995=>"111000111",
  39996=>"110101101",
  39997=>"100111111",
  39998=>"011001100",
  39999=>"111001111",
  40000=>"110010010",
  40001=>"101101001",
  40002=>"101101111",
  40003=>"001010010",
  40004=>"111110100",
  40005=>"010000111",
  40006=>"111101000",
  40007=>"101111011",
  40008=>"011100100",
  40009=>"001101010",
  40010=>"001111101",
  40011=>"010111100",
  40012=>"101001101",
  40013=>"111101110",
  40014=>"000100001",
  40015=>"010000011",
  40016=>"010000100",
  40017=>"001111011",
  40018=>"011010001",
  40019=>"110111000",
  40020=>"000011001",
  40021=>"011110010",
  40022=>"000001001",
  40023=>"110110001",
  40024=>"111100010",
  40025=>"111110000",
  40026=>"011110010",
  40027=>"011000000",
  40028=>"010101100",
  40029=>"101111010",
  40030=>"001110000",
  40031=>"000110001",
  40032=>"001000111",
  40033=>"001010010",
  40034=>"010000011",
  40035=>"001010001",
  40036=>"111111011",
  40037=>"000010101",
  40038=>"110000011",
  40039=>"111111001",
  40040=>"001101010",
  40041=>"001010100",
  40042=>"100001010",
  40043=>"110101010",
  40044=>"111100000",
  40045=>"100011000",
  40046=>"011111001",
  40047=>"111101111",
  40048=>"010000000",
  40049=>"011001010",
  40050=>"111111011",
  40051=>"111110010",
  40052=>"001111111",
  40053=>"010100001",
  40054=>"001100101",
  40055=>"101111011",
  40056=>"100000111",
  40057=>"101100000",
  40058=>"110011010",
  40059=>"111011000",
  40060=>"010000100",
  40061=>"110000110",
  40062=>"011111000",
  40063=>"000100101",
  40064=>"000101110",
  40065=>"101001100",
  40066=>"110101010",
  40067=>"110111111",
  40068=>"000010001",
  40069=>"110000100",
  40070=>"010010100",
  40071=>"011001111",
  40072=>"000001010",
  40073=>"001010101",
  40074=>"111101010",
  40075=>"100100001",
  40076=>"101111000",
  40077=>"110000001",
  40078=>"010010001",
  40079=>"101000100",
  40080=>"000001100",
  40081=>"111010101",
  40082=>"000111101",
  40083=>"010000010",
  40084=>"101101111",
  40085=>"101101111",
  40086=>"011011010",
  40087=>"111000010",
  40088=>"000011010",
  40089=>"101111110",
  40090=>"100110111",
  40091=>"111110100",
  40092=>"001100111",
  40093=>"001001111",
  40094=>"000100100",
  40095=>"110100101",
  40096=>"111101110",
  40097=>"001010111",
  40098=>"001011100",
  40099=>"011101101",
  40100=>"001100011",
  40101=>"100000101",
  40102=>"100001100",
  40103=>"011001110",
  40104=>"101110110",
  40105=>"111011010",
  40106=>"000110000",
  40107=>"010010010",
  40108=>"110110101",
  40109=>"100111000",
  40110=>"111010000",
  40111=>"111000000",
  40112=>"010011011",
  40113=>"000011101",
  40114=>"001000010",
  40115=>"111100000",
  40116=>"111010001",
  40117=>"101000101",
  40118=>"111001001",
  40119=>"101100110",
  40120=>"011111111",
  40121=>"000010111",
  40122=>"011001000",
  40123=>"101001000",
  40124=>"001101010",
  40125=>"001100111",
  40126=>"110100000",
  40127=>"011011110",
  40128=>"111100101",
  40129=>"100110110",
  40130=>"001001001",
  40131=>"100100111",
  40132=>"101001101",
  40133=>"000110011",
  40134=>"101000010",
  40135=>"010101111",
  40136=>"010110100",
  40137=>"100010110",
  40138=>"011000010",
  40139=>"100111001",
  40140=>"011101011",
  40141=>"110010111",
  40142=>"000001010",
  40143=>"010111101",
  40144=>"010000100",
  40145=>"110101010",
  40146=>"111111000",
  40147=>"001110110",
  40148=>"101000111",
  40149=>"010001101",
  40150=>"100100101",
  40151=>"111001101",
  40152=>"000011011",
  40153=>"010111010",
  40154=>"111111001",
  40155=>"110000101",
  40156=>"101000101",
  40157=>"010000011",
  40158=>"101111001",
  40159=>"110111011",
  40160=>"000001000",
  40161=>"001011010",
  40162=>"010100010",
  40163=>"011110110",
  40164=>"110100111",
  40165=>"010101010",
  40166=>"100110110",
  40167=>"011101000",
  40168=>"100110100",
  40169=>"100010000",
  40170=>"000000011",
  40171=>"011100111",
  40172=>"111111111",
  40173=>"110110110",
  40174=>"110001011",
  40175=>"011000000",
  40176=>"101011001",
  40177=>"010001110",
  40178=>"110011010",
  40179=>"111001011",
  40180=>"111000011",
  40181=>"000100000",
  40182=>"111011111",
  40183=>"010100010",
  40184=>"110101110",
  40185=>"111111000",
  40186=>"010001000",
  40187=>"010101110",
  40188=>"110100101",
  40189=>"000101000",
  40190=>"111111101",
  40191=>"111111110",
  40192=>"111111111",
  40193=>"110011110",
  40194=>"010100000",
  40195=>"111010011",
  40196=>"001000110",
  40197=>"000001100",
  40198=>"000000110",
  40199=>"111100110",
  40200=>"100001000",
  40201=>"100100010",
  40202=>"000000001",
  40203=>"010010010",
  40204=>"110110011",
  40205=>"010010101",
  40206=>"011011000",
  40207=>"100011011",
  40208=>"111001111",
  40209=>"111011000",
  40210=>"000100100",
  40211=>"110010010",
  40212=>"101010000",
  40213=>"100011010",
  40214=>"001000010",
  40215=>"111111011",
  40216=>"101100001",
  40217=>"001000000",
  40218=>"110001111",
  40219=>"100111011",
  40220=>"011010101",
  40221=>"101000101",
  40222=>"001110000",
  40223=>"110101010",
  40224=>"100000011",
  40225=>"101011111",
  40226=>"110110011",
  40227=>"100101000",
  40228=>"011000011",
  40229=>"000000010",
  40230=>"111000100",
  40231=>"001010010",
  40232=>"000001100",
  40233=>"111100111",
  40234=>"010010101",
  40235=>"011110010",
  40236=>"001010111",
  40237=>"001000010",
  40238=>"111100010",
  40239=>"111111011",
  40240=>"010011100",
  40241=>"000111001",
  40242=>"111000000",
  40243=>"000110110",
  40244=>"110101101",
  40245=>"110110110",
  40246=>"000001100",
  40247=>"010001000",
  40248=>"000010010",
  40249=>"101001101",
  40250=>"101101100",
  40251=>"000001001",
  40252=>"001011100",
  40253=>"110000011",
  40254=>"001010111",
  40255=>"100000000",
  40256=>"010100100",
  40257=>"011010000",
  40258=>"001110110",
  40259=>"110011010",
  40260=>"001110100",
  40261=>"001001111",
  40262=>"100000010",
  40263=>"000001111",
  40264=>"100101011",
  40265=>"000011000",
  40266=>"001010101",
  40267=>"100011101",
  40268=>"111110000",
  40269=>"000010110",
  40270=>"110010111",
  40271=>"011011100",
  40272=>"001000011",
  40273=>"101101110",
  40274=>"000101110",
  40275=>"010111010",
  40276=>"001010110",
  40277=>"101100001",
  40278=>"010110001",
  40279=>"001001001",
  40280=>"000100101",
  40281=>"100101000",
  40282=>"010010001",
  40283=>"000101011",
  40284=>"101100101",
  40285=>"000010100",
  40286=>"111011011",
  40287=>"011100111",
  40288=>"001010001",
  40289=>"100111010",
  40290=>"000000101",
  40291=>"001100111",
  40292=>"010000001",
  40293=>"101101110",
  40294=>"000010111",
  40295=>"000101110",
  40296=>"010110111",
  40297=>"000011110",
  40298=>"111110010",
  40299=>"111111010",
  40300=>"011000101",
  40301=>"001100110",
  40302=>"011011011",
  40303=>"110000010",
  40304=>"010010110",
  40305=>"100111111",
  40306=>"010110011",
  40307=>"110001001",
  40308=>"100011111",
  40309=>"001100100",
  40310=>"100010100",
  40311=>"101101011",
  40312=>"000001101",
  40313=>"011100110",
  40314=>"100011111",
  40315=>"010001000",
  40316=>"100110111",
  40317=>"100001001",
  40318=>"110100010",
  40319=>"101100010",
  40320=>"000000110",
  40321=>"001010011",
  40322=>"010100100",
  40323=>"100100001",
  40324=>"111101001",
  40325=>"110000100",
  40326=>"001000110",
  40327=>"000010110",
  40328=>"001000110",
  40329=>"011110101",
  40330=>"000000110",
  40331=>"000111011",
  40332=>"000110011",
  40333=>"001000000",
  40334=>"101010100",
  40335=>"010001100",
  40336=>"111001001",
  40337=>"000111111",
  40338=>"111011111",
  40339=>"100001110",
  40340=>"101000011",
  40341=>"001101110",
  40342=>"001101000",
  40343=>"011000101",
  40344=>"011101110",
  40345=>"001101001",
  40346=>"000101011",
  40347=>"000110010",
  40348=>"011001010",
  40349=>"000010001",
  40350=>"100110011",
  40351=>"000000001",
  40352=>"111111010",
  40353=>"011000110",
  40354=>"111100001",
  40355=>"111100001",
  40356=>"011010110",
  40357=>"011001011",
  40358=>"110000001",
  40359=>"111111110",
  40360=>"010101001",
  40361=>"111001100",
  40362=>"000000010",
  40363=>"000010100",
  40364=>"101100111",
  40365=>"001000100",
  40366=>"011010000",
  40367=>"000001001",
  40368=>"010110101",
  40369=>"010000000",
  40370=>"100110001",
  40371=>"000110011",
  40372=>"101101111",
  40373=>"100111010",
  40374=>"100100101",
  40375=>"000100111",
  40376=>"110011011",
  40377=>"101111011",
  40378=>"000001101",
  40379=>"011110010",
  40380=>"001001101",
  40381=>"100110101",
  40382=>"011111110",
  40383=>"100101111",
  40384=>"101010100",
  40385=>"010101111",
  40386=>"001101000",
  40387=>"110010000",
  40388=>"111111101",
  40389=>"111111011",
  40390=>"110111011",
  40391=>"001110011",
  40392=>"000001101",
  40393=>"000010010",
  40394=>"010011111",
  40395=>"110001001",
  40396=>"011100010",
  40397=>"000011111",
  40398=>"000111001",
  40399=>"111101101",
  40400=>"100010011",
  40401=>"010111011",
  40402=>"101101011",
  40403=>"101000001",
  40404=>"101100011",
  40405=>"010101111",
  40406=>"010001000",
  40407=>"100101000",
  40408=>"101101100",
  40409=>"110001000",
  40410=>"011010011",
  40411=>"101110101",
  40412=>"101100110",
  40413=>"101100100",
  40414=>"011101001",
  40415=>"101011111",
  40416=>"001101001",
  40417=>"101100010",
  40418=>"101111011",
  40419=>"111011000",
  40420=>"000110101",
  40421=>"111000000",
  40422=>"011101100",
  40423=>"011011101",
  40424=>"011110111",
  40425=>"101100110",
  40426=>"000100011",
  40427=>"100110111",
  40428=>"100110111",
  40429=>"011100010",
  40430=>"010111011",
  40431=>"010000000",
  40432=>"100101001",
  40433=>"111110100",
  40434=>"010000101",
  40435=>"000000101",
  40436=>"001000111",
  40437=>"011000111",
  40438=>"100100011",
  40439=>"111001101",
  40440=>"100000011",
  40441=>"101101100",
  40442=>"100001011",
  40443=>"110010101",
  40444=>"010111010",
  40445=>"010000010",
  40446=>"000100011",
  40447=>"100010110",
  40448=>"101101101",
  40449=>"111111111",
  40450=>"110101010",
  40451=>"010000010",
  40452=>"111100011",
  40453=>"000100010",
  40454=>"110001001",
  40455=>"111110010",
  40456=>"101010101",
  40457=>"111101110",
  40458=>"011001101",
  40459=>"010001010",
  40460=>"111110000",
  40461=>"011001101",
  40462=>"000101011",
  40463=>"110110000",
  40464=>"110111110",
  40465=>"011001110",
  40466=>"000010111",
  40467=>"100101001",
  40468=>"001000110",
  40469=>"100000010",
  40470=>"101010011",
  40471=>"000100101",
  40472=>"100000001",
  40473=>"000110110",
  40474=>"101000100",
  40475=>"011111111",
  40476=>"010100100",
  40477=>"101111110",
  40478=>"100000100",
  40479=>"111001110",
  40480=>"011111011",
  40481=>"110100011",
  40482=>"101101111",
  40483=>"011111010",
  40484=>"110001000",
  40485=>"101000000",
  40486=>"010001110",
  40487=>"011110001",
  40488=>"100100001",
  40489=>"110010010",
  40490=>"110000001",
  40491=>"110101110",
  40492=>"000011001",
  40493=>"111110011",
  40494=>"001000000",
  40495=>"110000010",
  40496=>"011100101",
  40497=>"001101110",
  40498=>"010110110",
  40499=>"001011110",
  40500=>"111101010",
  40501=>"100001000",
  40502=>"011111100",
  40503=>"000100111",
  40504=>"110011010",
  40505=>"010001111",
  40506=>"101101011",
  40507=>"011110111",
  40508=>"111100100",
  40509=>"110111001",
  40510=>"011001110",
  40511=>"110100011",
  40512=>"011000100",
  40513=>"011000000",
  40514=>"100101101",
  40515=>"100001001",
  40516=>"011000111",
  40517=>"011110101",
  40518=>"011101110",
  40519=>"000100111",
  40520=>"100111101",
  40521=>"101000101",
  40522=>"000110111",
  40523=>"000000011",
  40524=>"000100110",
  40525=>"001001110",
  40526=>"111000100",
  40527=>"000110010",
  40528=>"111010100",
  40529=>"011100010",
  40530=>"110111110",
  40531=>"010101100",
  40532=>"100100110",
  40533=>"000111111",
  40534=>"000111101",
  40535=>"001001100",
  40536=>"000110000",
  40537=>"111001011",
  40538=>"111011001",
  40539=>"100000011",
  40540=>"110110110",
  40541=>"000000000",
  40542=>"000100111",
  40543=>"011010000",
  40544=>"001111100",
  40545=>"000001000",
  40546=>"001001111",
  40547=>"010000010",
  40548=>"010110101",
  40549=>"111000101",
  40550=>"101000101",
  40551=>"110111001",
  40552=>"001000001",
  40553=>"001011100",
  40554=>"110001111",
  40555=>"101010010",
  40556=>"010100100",
  40557=>"001101010",
  40558=>"101111111",
  40559=>"110100000",
  40560=>"010101000",
  40561=>"100001100",
  40562=>"110000101",
  40563=>"101111110",
  40564=>"101101000",
  40565=>"000101100",
  40566=>"100010000",
  40567=>"111001101",
  40568=>"001100110",
  40569=>"111111011",
  40570=>"010111010",
  40571=>"100111101",
  40572=>"101111111",
  40573=>"000011100",
  40574=>"101000011",
  40575=>"101111111",
  40576=>"001110001",
  40577=>"001000000",
  40578=>"110000000",
  40579=>"001000010",
  40580=>"010101111",
  40581=>"101000011",
  40582=>"000000001",
  40583=>"011001101",
  40584=>"011011110",
  40585=>"010101100",
  40586=>"011110001",
  40587=>"010100101",
  40588=>"100100100",
  40589=>"001100001",
  40590=>"101101101",
  40591=>"011110000",
  40592=>"110100101",
  40593=>"011000101",
  40594=>"100000011",
  40595=>"001111110",
  40596=>"000000101",
  40597=>"100010010",
  40598=>"000100001",
  40599=>"001010110",
  40600=>"001111110",
  40601=>"001010011",
  40602=>"101110011",
  40603=>"010010110",
  40604=>"010010000",
  40605=>"000000000",
  40606=>"010110111",
  40607=>"101000000",
  40608=>"111101011",
  40609=>"110100000",
  40610=>"000001100",
  40611=>"111000011",
  40612=>"111111111",
  40613=>"111000111",
  40614=>"110101100",
  40615=>"001011100",
  40616=>"110011010",
  40617=>"011110100",
  40618=>"110110100",
  40619=>"111001000",
  40620=>"100101010",
  40621=>"000100111",
  40622=>"011001111",
  40623=>"100011011",
  40624=>"000101011",
  40625=>"010010101",
  40626=>"100110000",
  40627=>"110100111",
  40628=>"111000100",
  40629=>"001011111",
  40630=>"011010000",
  40631=>"000011100",
  40632=>"100100000",
  40633=>"101001110",
  40634=>"010001100",
  40635=>"011011000",
  40636=>"111011101",
  40637=>"001101111",
  40638=>"000000001",
  40639=>"110111111",
  40640=>"011011100",
  40641=>"101001111",
  40642=>"111111110",
  40643=>"011000100",
  40644=>"111111111",
  40645=>"001001110",
  40646=>"101111110",
  40647=>"110011100",
  40648=>"010001000",
  40649=>"111001111",
  40650=>"010110111",
  40651=>"000110111",
  40652=>"100101011",
  40653=>"001110100",
  40654=>"111100111",
  40655=>"011101000",
  40656=>"011101000",
  40657=>"100001110",
  40658=>"011111111",
  40659=>"100101101",
  40660=>"011100111",
  40661=>"101110100",
  40662=>"000010111",
  40663=>"000001110",
  40664=>"001100001",
  40665=>"101101011",
  40666=>"000110111",
  40667=>"110011110",
  40668=>"111101000",
  40669=>"000110001",
  40670=>"001100000",
  40671=>"101001110",
  40672=>"011100110",
  40673=>"111101000",
  40674=>"100101111",
  40675=>"001111001",
  40676=>"110110011",
  40677=>"101000101",
  40678=>"010001110",
  40679=>"101101100",
  40680=>"111000010",
  40681=>"100010000",
  40682=>"100110110",
  40683=>"011001010",
  40684=>"010110101",
  40685=>"010010001",
  40686=>"111000110",
  40687=>"010010010",
  40688=>"001011011",
  40689=>"101001101",
  40690=>"010000110",
  40691=>"111000100",
  40692=>"000011111",
  40693=>"010000100",
  40694=>"100110010",
  40695=>"011000011",
  40696=>"011001001",
  40697=>"100100000",
  40698=>"010100001",
  40699=>"010000010",
  40700=>"011100001",
  40701=>"101010101",
  40702=>"111001101",
  40703=>"010011000",
  40704=>"010100111",
  40705=>"010111101",
  40706=>"100100101",
  40707=>"110110010",
  40708=>"100111111",
  40709=>"010000111",
  40710=>"100101000",
  40711=>"111010000",
  40712=>"111000100",
  40713=>"001100110",
  40714=>"001010011",
  40715=>"010110000",
  40716=>"001100010",
  40717=>"001100011",
  40718=>"010000101",
  40719=>"110010110",
  40720=>"101010100",
  40721=>"011101000",
  40722=>"011011011",
  40723=>"001101100",
  40724=>"101010000",
  40725=>"100011110",
  40726=>"001000111",
  40727=>"110001110",
  40728=>"011110110",
  40729=>"110000001",
  40730=>"000110110",
  40731=>"010111000",
  40732=>"010110110",
  40733=>"110000110",
  40734=>"000011111",
  40735=>"011101001",
  40736=>"011010100",
  40737=>"100100010",
  40738=>"110111010",
  40739=>"001100010",
  40740=>"101000001",
  40741=>"100100111",
  40742=>"001101000",
  40743=>"010101001",
  40744=>"011010100",
  40745=>"101011010",
  40746=>"000001011",
  40747=>"000110111",
  40748=>"101010011",
  40749=>"011001011",
  40750=>"000100000",
  40751=>"010110000",
  40752=>"101101100",
  40753=>"011011100",
  40754=>"000010000",
  40755=>"100010011",
  40756=>"100101100",
  40757=>"111101010",
  40758=>"101001011",
  40759=>"110000000",
  40760=>"101011111",
  40761=>"000111111",
  40762=>"100011000",
  40763=>"011001110",
  40764=>"000000100",
  40765=>"010001001",
  40766=>"111001100",
  40767=>"011000011",
  40768=>"101101001",
  40769=>"110101001",
  40770=>"100101110",
  40771=>"111001001",
  40772=>"110101010",
  40773=>"101111110",
  40774=>"100000111",
  40775=>"010011100",
  40776=>"100111001",
  40777=>"100110010",
  40778=>"111001110",
  40779=>"001101011",
  40780=>"111001000",
  40781=>"100100100",
  40782=>"010000100",
  40783=>"100000101",
  40784=>"110111111",
  40785=>"000000011",
  40786=>"011110001",
  40787=>"001011000",
  40788=>"010101000",
  40789=>"101001111",
  40790=>"011101000",
  40791=>"011011110",
  40792=>"010000000",
  40793=>"100111000",
  40794=>"111010010",
  40795=>"101001011",
  40796=>"010110101",
  40797=>"000100010",
  40798=>"110110111",
  40799=>"000001011",
  40800=>"001010011",
  40801=>"000010010",
  40802=>"111100101",
  40803=>"000110101",
  40804=>"110110010",
  40805=>"000101101",
  40806=>"101010000",
  40807=>"100001111",
  40808=>"111011000",
  40809=>"111100001",
  40810=>"110110000",
  40811=>"000111000",
  40812=>"000000110",
  40813=>"110000101",
  40814=>"100111101",
  40815=>"000110011",
  40816=>"011111110",
  40817=>"100100111",
  40818=>"011000111",
  40819=>"001100001",
  40820=>"001010010",
  40821=>"101111101",
  40822=>"011111000",
  40823=>"010010010",
  40824=>"000101001",
  40825=>"010011111",
  40826=>"100000110",
  40827=>"010100101",
  40828=>"001010010",
  40829=>"010100011",
  40830=>"000111110",
  40831=>"110111010",
  40832=>"100001000",
  40833=>"000001110",
  40834=>"000100111",
  40835=>"001011010",
  40836=>"100011001",
  40837=>"110001011",
  40838=>"101101110",
  40839=>"110110111",
  40840=>"110111010",
  40841=>"101001000",
  40842=>"110101001",
  40843=>"000010011",
  40844=>"011011000",
  40845=>"000010110",
  40846=>"010111001",
  40847=>"000001011",
  40848=>"011000011",
  40849=>"001101001",
  40850=>"011000110",
  40851=>"110110000",
  40852=>"001011010",
  40853=>"101001011",
  40854=>"011101111",
  40855=>"101000100",
  40856=>"111001011",
  40857=>"111110000",
  40858=>"001101101",
  40859=>"100101101",
  40860=>"000001101",
  40861=>"011111010",
  40862=>"101101111",
  40863=>"010101011",
  40864=>"000001101",
  40865=>"111100001",
  40866=>"011101000",
  40867=>"101000111",
  40868=>"001010011",
  40869=>"101101101",
  40870=>"101010011",
  40871=>"000110100",
  40872=>"011010111",
  40873=>"111110110",
  40874=>"110001001",
  40875=>"110100100",
  40876=>"100011000",
  40877=>"011011111",
  40878=>"101010001",
  40879=>"100100000",
  40880=>"101011111",
  40881=>"011101000",
  40882=>"111011100",
  40883=>"001101111",
  40884=>"000001101",
  40885=>"010101010",
  40886=>"001010100",
  40887=>"011011100",
  40888=>"110101111",
  40889=>"110001100",
  40890=>"100010111",
  40891=>"111101111",
  40892=>"010010110",
  40893=>"001101100",
  40894=>"110011000",
  40895=>"001101010",
  40896=>"111110011",
  40897=>"111001110",
  40898=>"000000001",
  40899=>"011000001",
  40900=>"101100101",
  40901=>"011000011",
  40902=>"100001100",
  40903=>"010101101",
  40904=>"010111100",
  40905=>"001001001",
  40906=>"000100100",
  40907=>"000101101",
  40908=>"111100110",
  40909=>"001010111",
  40910=>"100110010",
  40911=>"110111110",
  40912=>"001100110",
  40913=>"100111100",
  40914=>"100000001",
  40915=>"010000011",
  40916=>"010111111",
  40917=>"101011110",
  40918=>"101001111",
  40919=>"110111110",
  40920=>"100001011",
  40921=>"101011101",
  40922=>"010110010",
  40923=>"001100001",
  40924=>"111010010",
  40925=>"110111010",
  40926=>"110110001",
  40927=>"000001011",
  40928=>"010010001",
  40929=>"011110111",
  40930=>"010001001",
  40931=>"000110011",
  40932=>"000001101",
  40933=>"000010011",
  40934=>"110111010",
  40935=>"010010101",
  40936=>"000000000",
  40937=>"101000010",
  40938=>"111100100",
  40939=>"001111011",
  40940=>"100111011",
  40941=>"000110010",
  40942=>"010010010",
  40943=>"010111010",
  40944=>"010010100",
  40945=>"101001010",
  40946=>"110010011",
  40947=>"110100011",
  40948=>"000100000",
  40949=>"000111111",
  40950=>"011111001",
  40951=>"000011111",
  40952=>"000000111",
  40953=>"110000010",
  40954=>"111000111",
  40955=>"110111111",
  40956=>"000100111",
  40957=>"100000111",
  40958=>"100100010",
  40959=>"111011110",
  40960=>"000010000",
  40961=>"111010110",
  40962=>"111100110",
  40963=>"010000000",
  40964=>"110000000",
  40965=>"001000001",
  40966=>"110110100",
  40967=>"010011110",
  40968=>"111101111",
  40969=>"011100000",
  40970=>"000000101",
  40971=>"101111010",
  40972=>"101100101",
  40973=>"000010100",
  40974=>"010110110",
  40975=>"110110101",
  40976=>"011110001",
  40977=>"011111011",
  40978=>"011000101",
  40979=>"110111111",
  40980=>"110100111",
  40981=>"000101010",
  40982=>"100100110",
  40983=>"001001111",
  40984=>"111100110",
  40985=>"000101010",
  40986=>"110101100",
  40987=>"101010001",
  40988=>"001111010",
  40989=>"001010110",
  40990=>"101110110",
  40991=>"000101001",
  40992=>"010010000",
  40993=>"101000011",
  40994=>"101111000",
  40995=>"110100010",
  40996=>"101010000",
  40997=>"101110001",
  40998=>"000010111",
  40999=>"110010101",
  41000=>"101000001",
  41001=>"011001111",
  41002=>"000100110",
  41003=>"100101111",
  41004=>"110001001",
  41005=>"110011100",
  41006=>"011010110",
  41007=>"011010100",
  41008=>"101010110",
  41009=>"100100100",
  41010=>"111100100",
  41011=>"010100010",
  41012=>"000000001",
  41013=>"010100000",
  41014=>"010010000",
  41015=>"110101111",
  41016=>"101011101",
  41017=>"000111001",
  41018=>"000110110",
  41019=>"111101110",
  41020=>"100101000",
  41021=>"100000100",
  41022=>"111111010",
  41023=>"101111010",
  41024=>"100000010",
  41025=>"100010110",
  41026=>"001110110",
  41027=>"011001111",
  41028=>"101010110",
  41029=>"101000011",
  41030=>"011110001",
  41031=>"010111010",
  41032=>"000001001",
  41033=>"001000110",
  41034=>"111010011",
  41035=>"011100100",
  41036=>"111011011",
  41037=>"011101110",
  41038=>"001001010",
  41039=>"011000010",
  41040=>"101110001",
  41041=>"111010011",
  41042=>"011010100",
  41043=>"101101110",
  41044=>"001000111",
  41045=>"011100110",
  41046=>"000111111",
  41047=>"111110100",
  41048=>"001001000",
  41049=>"101110110",
  41050=>"100011110",
  41051=>"001010011",
  41052=>"011111000",
  41053=>"110001001",
  41054=>"100011011",
  41055=>"000000111",
  41056=>"001001001",
  41057=>"011001110",
  41058=>"101010111",
  41059=>"000010101",
  41060=>"100101000",
  41061=>"110000011",
  41062=>"001110110",
  41063=>"110011111",
  41064=>"011000010",
  41065=>"111100010",
  41066=>"010000101",
  41067=>"110011100",
  41068=>"001011001",
  41069=>"111000011",
  41070=>"100111011",
  41071=>"111010010",
  41072=>"101000010",
  41073=>"000010110",
  41074=>"110001011",
  41075=>"111101010",
  41076=>"100010100",
  41077=>"100000010",
  41078=>"011001001",
  41079=>"101001111",
  41080=>"111011111",
  41081=>"100100111",
  41082=>"001000110",
  41083=>"101101101",
  41084=>"000100000",
  41085=>"110000000",
  41086=>"000100010",
  41087=>"000111000",
  41088=>"000100010",
  41089=>"011011000",
  41090=>"011100111",
  41091=>"100101000",
  41092=>"001001000",
  41093=>"101111101",
  41094=>"101001010",
  41095=>"100111011",
  41096=>"010010010",
  41097=>"110111001",
  41098=>"111101010",
  41099=>"001001011",
  41100=>"111010000",
  41101=>"100101000",
  41102=>"001010011",
  41103=>"001101011",
  41104=>"111110111",
  41105=>"110101100",
  41106=>"111010001",
  41107=>"110000010",
  41108=>"011000001",
  41109=>"100011001",
  41110=>"101011001",
  41111=>"101100010",
  41112=>"011110001",
  41113=>"101000011",
  41114=>"101100010",
  41115=>"000100100",
  41116=>"100101101",
  41117=>"110111101",
  41118=>"000010111",
  41119=>"011110001",
  41120=>"111100101",
  41121=>"110001010",
  41122=>"010100100",
  41123=>"011111100",
  41124=>"110100010",
  41125=>"110000010",
  41126=>"101111000",
  41127=>"000010000",
  41128=>"000100000",
  41129=>"101100111",
  41130=>"001100000",
  41131=>"100010101",
  41132=>"111100111",
  41133=>"011010101",
  41134=>"000010001",
  41135=>"110001100",
  41136=>"000101100",
  41137=>"101001011",
  41138=>"010001000",
  41139=>"101011011",
  41140=>"100011110",
  41141=>"001010011",
  41142=>"000000001",
  41143=>"100100001",
  41144=>"111100001",
  41145=>"101110110",
  41146=>"100001001",
  41147=>"101001011",
  41148=>"001001010",
  41149=>"000010101",
  41150=>"011100110",
  41151=>"011100100",
  41152=>"001101111",
  41153=>"000000101",
  41154=>"100101101",
  41155=>"111000110",
  41156=>"110100001",
  41157=>"011000010",
  41158=>"111010011",
  41159=>"011010001",
  41160=>"011011010",
  41161=>"000000101",
  41162=>"011100001",
  41163=>"011111111",
  41164=>"011011101",
  41165=>"111100110",
  41166=>"000001000",
  41167=>"000100100",
  41168=>"111010100",
  41169=>"000101110",
  41170=>"101011100",
  41171=>"100110001",
  41172=>"110110101",
  41173=>"110100111",
  41174=>"000111000",
  41175=>"111100011",
  41176=>"011001000",
  41177=>"011001010",
  41178=>"001111101",
  41179=>"111110001",
  41180=>"010100000",
  41181=>"010110111",
  41182=>"000011111",
  41183=>"111110000",
  41184=>"001111000",
  41185=>"100010010",
  41186=>"110011101",
  41187=>"000010001",
  41188=>"010101010",
  41189=>"111111101",
  41190=>"101000000",
  41191=>"111010111",
  41192=>"001110111",
  41193=>"101001100",
  41194=>"010010101",
  41195=>"001100111",
  41196=>"101100000",
  41197=>"001100010",
  41198=>"000000010",
  41199=>"011010000",
  41200=>"111011011",
  41201=>"011011100",
  41202=>"000000110",
  41203=>"100001001",
  41204=>"110110000",
  41205=>"010101010",
  41206=>"101001010",
  41207=>"010000011",
  41208=>"111101000",
  41209=>"111110010",
  41210=>"001000111",
  41211=>"010110000",
  41212=>"001011000",
  41213=>"010111000",
  41214=>"101101000",
  41215=>"111100110",
  41216=>"101000000",
  41217=>"011011000",
  41218=>"111000101",
  41219=>"010010111",
  41220=>"101000111",
  41221=>"110011000",
  41222=>"101000001",
  41223=>"111011001",
  41224=>"011010110",
  41225=>"110110010",
  41226=>"100010101",
  41227=>"111001000",
  41228=>"000001110",
  41229=>"001010100",
  41230=>"100111101",
  41231=>"110011100",
  41232=>"011101011",
  41233=>"100100000",
  41234=>"101100000",
  41235=>"111001101",
  41236=>"110111100",
  41237=>"101001011",
  41238=>"110100010",
  41239=>"110011000",
  41240=>"110011101",
  41241=>"101110101",
  41242=>"111001000",
  41243=>"011111010",
  41244=>"110101011",
  41245=>"111100100",
  41246=>"001111001",
  41247=>"110000101",
  41248=>"101100111",
  41249=>"100111100",
  41250=>"111010111",
  41251=>"000000001",
  41252=>"001011111",
  41253=>"010001111",
  41254=>"000010000",
  41255=>"100000110",
  41256=>"101000001",
  41257=>"000111011",
  41258=>"011110110",
  41259=>"010000010",
  41260=>"001110011",
  41261=>"101111000",
  41262=>"000001000",
  41263=>"010111111",
  41264=>"111101110",
  41265=>"000100101",
  41266=>"101010101",
  41267=>"100111010",
  41268=>"101000000",
  41269=>"111010000",
  41270=>"011001001",
  41271=>"000000000",
  41272=>"011011110",
  41273=>"111100001",
  41274=>"111000011",
  41275=>"110000001",
  41276=>"101001001",
  41277=>"100000010",
  41278=>"011111011",
  41279=>"010010011",
  41280=>"000010001",
  41281=>"111110101",
  41282=>"000010001",
  41283=>"111111011",
  41284=>"000111010",
  41285=>"000111000",
  41286=>"000001010",
  41287=>"010000000",
  41288=>"001110100",
  41289=>"000100010",
  41290=>"100000000",
  41291=>"101101110",
  41292=>"111110110",
  41293=>"110110111",
  41294=>"100100010",
  41295=>"111001100",
  41296=>"110001000",
  41297=>"111110110",
  41298=>"000111011",
  41299=>"101001000",
  41300=>"110010000",
  41301=>"010100111",
  41302=>"010010110",
  41303=>"101101000",
  41304=>"000010100",
  41305=>"001101100",
  41306=>"001111111",
  41307=>"010111001",
  41308=>"100000110",
  41309=>"111000101",
  41310=>"011000111",
  41311=>"100010010",
  41312=>"110101100",
  41313=>"110100010",
  41314=>"000011100",
  41315=>"001111111",
  41316=>"110000001",
  41317=>"010100100",
  41318=>"010101101",
  41319=>"001010011",
  41320=>"000110000",
  41321=>"101111111",
  41322=>"001011011",
  41323=>"001001010",
  41324=>"010000001",
  41325=>"100101010",
  41326=>"000010100",
  41327=>"111001111",
  41328=>"001010011",
  41329=>"110001001",
  41330=>"110011111",
  41331=>"000011010",
  41332=>"001011111",
  41333=>"001101000",
  41334=>"100111010",
  41335=>"001101110",
  41336=>"001000101",
  41337=>"000100000",
  41338=>"110110000",
  41339=>"101000000",
  41340=>"101010000",
  41341=>"110110011",
  41342=>"000100101",
  41343=>"000110001",
  41344=>"110111011",
  41345=>"011000110",
  41346=>"011101101",
  41347=>"110110010",
  41348=>"111101111",
  41349=>"101100111",
  41350=>"011011000",
  41351=>"000111110",
  41352=>"011001100",
  41353=>"101011101",
  41354=>"001100011",
  41355=>"101000111",
  41356=>"110111101",
  41357=>"111100100",
  41358=>"011100110",
  41359=>"011001111",
  41360=>"101111010",
  41361=>"100100111",
  41362=>"110011111",
  41363=>"111011101",
  41364=>"100000101",
  41365=>"001110001",
  41366=>"101110110",
  41367=>"110111010",
  41368=>"110010000",
  41369=>"000100110",
  41370=>"011011111",
  41371=>"010001110",
  41372=>"111010110",
  41373=>"100011110",
  41374=>"111100101",
  41375=>"000001101",
  41376=>"000101100",
  41377=>"111101001",
  41378=>"100001000",
  41379=>"101100100",
  41380=>"110100101",
  41381=>"010001001",
  41382=>"011001000",
  41383=>"010100001",
  41384=>"111100101",
  41385=>"011110101",
  41386=>"111001110",
  41387=>"110111010",
  41388=>"111010010",
  41389=>"000000110",
  41390=>"010000111",
  41391=>"101110000",
  41392=>"100111010",
  41393=>"001111110",
  41394=>"001100101",
  41395=>"101101100",
  41396=>"101110100",
  41397=>"001000000",
  41398=>"011110111",
  41399=>"110001100",
  41400=>"011010010",
  41401=>"001001001",
  41402=>"010000001",
  41403=>"010011000",
  41404=>"110110101",
  41405=>"101001010",
  41406=>"101100110",
  41407=>"100011010",
  41408=>"001001001",
  41409=>"000100001",
  41410=>"101111110",
  41411=>"000111001",
  41412=>"110111010",
  41413=>"011101101",
  41414=>"111000001",
  41415=>"000000000",
  41416=>"001011110",
  41417=>"110000111",
  41418=>"001000000",
  41419=>"111010000",
  41420=>"111011011",
  41421=>"000010111",
  41422=>"000110000",
  41423=>"000010011",
  41424=>"100011011",
  41425=>"010001111",
  41426=>"100100110",
  41427=>"010000111",
  41428=>"111111111",
  41429=>"000100000",
  41430=>"101100011",
  41431=>"010000001",
  41432=>"101000001",
  41433=>"111100000",
  41434=>"000101011",
  41435=>"111010000",
  41436=>"000000000",
  41437=>"111111000",
  41438=>"011101000",
  41439=>"011000111",
  41440=>"111000101",
  41441=>"000111101",
  41442=>"110010000",
  41443=>"010100001",
  41444=>"001010000",
  41445=>"010100110",
  41446=>"110001010",
  41447=>"110000000",
  41448=>"010000101",
  41449=>"101011001",
  41450=>"100110001",
  41451=>"101111000",
  41452=>"001101001",
  41453=>"100001000",
  41454=>"000000000",
  41455=>"000010001",
  41456=>"010101001",
  41457=>"001010000",
  41458=>"101110000",
  41459=>"110100110",
  41460=>"000001011",
  41461=>"001111101",
  41462=>"110111111",
  41463=>"101111000",
  41464=>"000010011",
  41465=>"010111100",
  41466=>"111101001",
  41467=>"000110111",
  41468=>"110010111",
  41469=>"100011100",
  41470=>"100110100",
  41471=>"111100000",
  41472=>"011011100",
  41473=>"001010000",
  41474=>"101100111",
  41475=>"100000111",
  41476=>"111101010",
  41477=>"001010111",
  41478=>"000100111",
  41479=>"100010100",
  41480=>"000100110",
  41481=>"101100000",
  41482=>"010111011",
  41483=>"001111100",
  41484=>"100011100",
  41485=>"111000001",
  41486=>"000000111",
  41487=>"010010110",
  41488=>"011110010",
  41489=>"011111001",
  41490=>"101001110",
  41491=>"000011100",
  41492=>"010110000",
  41493=>"101110100",
  41494=>"100100011",
  41495=>"110011011",
  41496=>"101001000",
  41497=>"010110111",
  41498=>"000001011",
  41499=>"000110011",
  41500=>"101000110",
  41501=>"101010011",
  41502=>"000101000",
  41503=>"100000011",
  41504=>"100110100",
  41505=>"110010101",
  41506=>"011100010",
  41507=>"001100000",
  41508=>"010110001",
  41509=>"100101101",
  41510=>"100101100",
  41511=>"110010001",
  41512=>"000000011",
  41513=>"101111110",
  41514=>"101101111",
  41515=>"011000000",
  41516=>"011010101",
  41517=>"101010100",
  41518=>"111011011",
  41519=>"010100111",
  41520=>"110100000",
  41521=>"101111110",
  41522=>"011001100",
  41523=>"010110011",
  41524=>"111111000",
  41525=>"010100111",
  41526=>"100000001",
  41527=>"110100001",
  41528=>"110000010",
  41529=>"110010011",
  41530=>"110111101",
  41531=>"010101011",
  41532=>"001111100",
  41533=>"001101100",
  41534=>"001000001",
  41535=>"011011000",
  41536=>"111110110",
  41537=>"011000010",
  41538=>"001000001",
  41539=>"011101000",
  41540=>"110111010",
  41541=>"111100100",
  41542=>"001000011",
  41543=>"101011001",
  41544=>"010100110",
  41545=>"001000100",
  41546=>"001001010",
  41547=>"110000110",
  41548=>"100001101",
  41549=>"000000101",
  41550=>"011100001",
  41551=>"011010010",
  41552=>"010111111",
  41553=>"010100111",
  41554=>"101111111",
  41555=>"100011101",
  41556=>"001000100",
  41557=>"101111101",
  41558=>"001100001",
  41559=>"001101011",
  41560=>"001000001",
  41561=>"010001100",
  41562=>"000101101",
  41563=>"100100111",
  41564=>"101100101",
  41565=>"100100001",
  41566=>"101111110",
  41567=>"110101011",
  41568=>"111001010",
  41569=>"100001111",
  41570=>"101010100",
  41571=>"100111100",
  41572=>"110101011",
  41573=>"101101011",
  41574=>"000110000",
  41575=>"000010110",
  41576=>"011101000",
  41577=>"011100110",
  41578=>"011101100",
  41579=>"110000111",
  41580=>"110111111",
  41581=>"000010100",
  41582=>"101001101",
  41583=>"110000100",
  41584=>"000100000",
  41585=>"000100000",
  41586=>"001011100",
  41587=>"011111110",
  41588=>"011100100",
  41589=>"000101101",
  41590=>"011001111",
  41591=>"110101111",
  41592=>"111111010",
  41593=>"001101110",
  41594=>"010111010",
  41595=>"100101101",
  41596=>"011000011",
  41597=>"011001000",
  41598=>"000110000",
  41599=>"101110110",
  41600=>"100101110",
  41601=>"010110100",
  41602=>"000111010",
  41603=>"010000100",
  41604=>"111101111",
  41605=>"000001110",
  41606=>"011000110",
  41607=>"000000010",
  41608=>"010101110",
  41609=>"010110111",
  41610=>"100001111",
  41611=>"001101011",
  41612=>"011000101",
  41613=>"011010110",
  41614=>"111011011",
  41615=>"100100101",
  41616=>"000101111",
  41617=>"111000110",
  41618=>"110011001",
  41619=>"100110101",
  41620=>"100001001",
  41621=>"010100111",
  41622=>"010010011",
  41623=>"000100000",
  41624=>"011000111",
  41625=>"111110110",
  41626=>"001111011",
  41627=>"010010100",
  41628=>"001010110",
  41629=>"011111010",
  41630=>"110101001",
  41631=>"011010011",
  41632=>"001010000",
  41633=>"001000101",
  41634=>"101000000",
  41635=>"010001111",
  41636=>"011110001",
  41637=>"111011110",
  41638=>"001111101",
  41639=>"100011001",
  41640=>"000111100",
  41641=>"010000001",
  41642=>"100010100",
  41643=>"000010111",
  41644=>"000000110",
  41645=>"011110001",
  41646=>"011100110",
  41647=>"001110001",
  41648=>"000101100",
  41649=>"000011111",
  41650=>"000001000",
  41651=>"001001110",
  41652=>"110011000",
  41653=>"101110010",
  41654=>"101011110",
  41655=>"100101010",
  41656=>"100000010",
  41657=>"000110001",
  41658=>"001010110",
  41659=>"011110101",
  41660=>"000100111",
  41661=>"011011111",
  41662=>"110000010",
  41663=>"010111010",
  41664=>"100011010",
  41665=>"111101011",
  41666=>"000110010",
  41667=>"111110011",
  41668=>"101111110",
  41669=>"111100000",
  41670=>"001001100",
  41671=>"000111111",
  41672=>"010011000",
  41673=>"110001000",
  41674=>"110010111",
  41675=>"000001101",
  41676=>"110101011",
  41677=>"010001010",
  41678=>"111011000",
  41679=>"010101001",
  41680=>"111101001",
  41681=>"111011111",
  41682=>"101101000",
  41683=>"011110111",
  41684=>"111101000",
  41685=>"000010111",
  41686=>"110101110",
  41687=>"001100101",
  41688=>"110111100",
  41689=>"010110010",
  41690=>"100001101",
  41691=>"011000000",
  41692=>"110000101",
  41693=>"100001001",
  41694=>"100001100",
  41695=>"111011101",
  41696=>"111011111",
  41697=>"101110110",
  41698=>"101001111",
  41699=>"001111010",
  41700=>"100000000",
  41701=>"101000101",
  41702=>"010011110",
  41703=>"111011111",
  41704=>"101010110",
  41705=>"010000110",
  41706=>"111001100",
  41707=>"111011111",
  41708=>"110000111",
  41709=>"000000000",
  41710=>"011110011",
  41711=>"111010110",
  41712=>"001110010",
  41713=>"010100001",
  41714=>"101100000",
  41715=>"111011110",
  41716=>"000010111",
  41717=>"101110110",
  41718=>"111110110",
  41719=>"111110111",
  41720=>"111001101",
  41721=>"011011010",
  41722=>"101111000",
  41723=>"111000101",
  41724=>"101101110",
  41725=>"101010001",
  41726=>"111110000",
  41727=>"101111110",
  41728=>"110000001",
  41729=>"000110111",
  41730=>"100011000",
  41731=>"011000000",
  41732=>"010101001",
  41733=>"010000000",
  41734=>"101010101",
  41735=>"011110011",
  41736=>"011101011",
  41737=>"101010010",
  41738=>"111010111",
  41739=>"001011011",
  41740=>"010100110",
  41741=>"010000110",
  41742=>"100111100",
  41743=>"001011100",
  41744=>"010100011",
  41745=>"001110110",
  41746=>"100001111",
  41747=>"101101100",
  41748=>"101011101",
  41749=>"000010011",
  41750=>"010100111",
  41751=>"111110111",
  41752=>"111001000",
  41753=>"101100001",
  41754=>"000010111",
  41755=>"111000000",
  41756=>"010110011",
  41757=>"111000000",
  41758=>"100100110",
  41759=>"011100100",
  41760=>"101000101",
  41761=>"011111011",
  41762=>"000101001",
  41763=>"110000111",
  41764=>"000101101",
  41765=>"000010101",
  41766=>"111101000",
  41767=>"111100111",
  41768=>"001110011",
  41769=>"001001000",
  41770=>"010100010",
  41771=>"110011010",
  41772=>"010101000",
  41773=>"000001010",
  41774=>"000000100",
  41775=>"010110001",
  41776=>"101000000",
  41777=>"100000000",
  41778=>"111001010",
  41779=>"010110011",
  41780=>"010010010",
  41781=>"101110001",
  41782=>"101110010",
  41783=>"101001000",
  41784=>"010110000",
  41785=>"110101011",
  41786=>"110100101",
  41787=>"010100110",
  41788=>"000110111",
  41789=>"101100111",
  41790=>"000000000",
  41791=>"101010100",
  41792=>"110001111",
  41793=>"011101000",
  41794=>"011011000",
  41795=>"010000101",
  41796=>"101100101",
  41797=>"011111001",
  41798=>"011011101",
  41799=>"100100011",
  41800=>"001010000",
  41801=>"110110100",
  41802=>"010001011",
  41803=>"100011100",
  41804=>"001011111",
  41805=>"101100101",
  41806=>"011000111",
  41807=>"010110100",
  41808=>"111001111",
  41809=>"011010011",
  41810=>"011100101",
  41811=>"011001111",
  41812=>"010010100",
  41813=>"001101000",
  41814=>"000000000",
  41815=>"010001011",
  41816=>"001101101",
  41817=>"100110011",
  41818=>"001111110",
  41819=>"001110110",
  41820=>"010001000",
  41821=>"110010010",
  41822=>"111000100",
  41823=>"101010101",
  41824=>"001100000",
  41825=>"000101100",
  41826=>"111111111",
  41827=>"111110010",
  41828=>"010100101",
  41829=>"111101001",
  41830=>"000100011",
  41831=>"111100001",
  41832=>"101011010",
  41833=>"100000010",
  41834=>"101111010",
  41835=>"010000000",
  41836=>"111000000",
  41837=>"010000100",
  41838=>"100111100",
  41839=>"001000010",
  41840=>"001010111",
  41841=>"011000100",
  41842=>"101001000",
  41843=>"111101000",
  41844=>"010011010",
  41845=>"000000100",
  41846=>"001110110",
  41847=>"100000010",
  41848=>"011101000",
  41849=>"101000111",
  41850=>"111101000",
  41851=>"000101100",
  41852=>"000100110",
  41853=>"011010000",
  41854=>"110010001",
  41855=>"000011101",
  41856=>"111111111",
  41857=>"001100001",
  41858=>"010010101",
  41859=>"111111100",
  41860=>"000000001",
  41861=>"110011011",
  41862=>"111010110",
  41863=>"110111110",
  41864=>"000111110",
  41865=>"100011110",
  41866=>"010001100",
  41867=>"000000110",
  41868=>"110000000",
  41869=>"001111010",
  41870=>"010111011",
  41871=>"101010011",
  41872=>"110000110",
  41873=>"001001110",
  41874=>"000100111",
  41875=>"001111000",
  41876=>"110110110",
  41877=>"001001101",
  41878=>"011101101",
  41879=>"001111111",
  41880=>"011001000",
  41881=>"000111111",
  41882=>"001111101",
  41883=>"000101110",
  41884=>"011111010",
  41885=>"100110010",
  41886=>"110100011",
  41887=>"010011111",
  41888=>"101001000",
  41889=>"111110100",
  41890=>"010111111",
  41891=>"010000000",
  41892=>"010101010",
  41893=>"111100011",
  41894=>"100000001",
  41895=>"100000001",
  41896=>"010100101",
  41897=>"000010000",
  41898=>"111111100",
  41899=>"011111111",
  41900=>"011101001",
  41901=>"001011111",
  41902=>"111110110",
  41903=>"001110100",
  41904=>"111010001",
  41905=>"011111000",
  41906=>"000100001",
  41907=>"000011000",
  41908=>"000100001",
  41909=>"000000110",
  41910=>"100111010",
  41911=>"110011011",
  41912=>"101100110",
  41913=>"010110001",
  41914=>"101000100",
  41915=>"110001111",
  41916=>"011000001",
  41917=>"100000111",
  41918=>"000101101",
  41919=>"011000000",
  41920=>"100010000",
  41921=>"000101101",
  41922=>"101101001",
  41923=>"000010000",
  41924=>"110100011",
  41925=>"100100011",
  41926=>"001000001",
  41927=>"110111010",
  41928=>"001000010",
  41929=>"101100000",
  41930=>"111101110",
  41931=>"111100001",
  41932=>"110011010",
  41933=>"000000011",
  41934=>"110100000",
  41935=>"011010010",
  41936=>"011011101",
  41937=>"001010001",
  41938=>"111001000",
  41939=>"111111101",
  41940=>"101000000",
  41941=>"101001101",
  41942=>"110000000",
  41943=>"101011111",
  41944=>"111111101",
  41945=>"011011011",
  41946=>"110110101",
  41947=>"000111011",
  41948=>"001101110",
  41949=>"010000011",
  41950=>"011010010",
  41951=>"000000010",
  41952=>"101011010",
  41953=>"001011011",
  41954=>"000100111",
  41955=>"010001111",
  41956=>"010000001",
  41957=>"111011000",
  41958=>"001111110",
  41959=>"101110010",
  41960=>"001000011",
  41961=>"110001011",
  41962=>"111100101",
  41963=>"100011111",
  41964=>"000100000",
  41965=>"101100011",
  41966=>"001000000",
  41967=>"011111010",
  41968=>"000011111",
  41969=>"111101110",
  41970=>"111100010",
  41971=>"001001110",
  41972=>"001101110",
  41973=>"011101000",
  41974=>"110010100",
  41975=>"010010110",
  41976=>"000111010",
  41977=>"010011001",
  41978=>"011101111",
  41979=>"011011001",
  41980=>"110110111",
  41981=>"101111110",
  41982=>"011110000",
  41983=>"000010101",
  41984=>"101100111",
  41985=>"111110110",
  41986=>"010101111",
  41987=>"011100100",
  41988=>"111110100",
  41989=>"111111001",
  41990=>"001100101",
  41991=>"111101100",
  41992=>"110010110",
  41993=>"111100010",
  41994=>"000100111",
  41995=>"001001100",
  41996=>"101001111",
  41997=>"111001111",
  41998=>"111110100",
  41999=>"001000000",
  42000=>"101101101",
  42001=>"001100000",
  42002=>"000101011",
  42003=>"101100110",
  42004=>"011111011",
  42005=>"110001110",
  42006=>"000110110",
  42007=>"111110000",
  42008=>"010010010",
  42009=>"010010010",
  42010=>"011110111",
  42011=>"001001010",
  42012=>"100101100",
  42013=>"011100111",
  42014=>"111011010",
  42015=>"101001001",
  42016=>"010110000",
  42017=>"110111000",
  42018=>"111101111",
  42019=>"000000110",
  42020=>"100101111",
  42021=>"111110011",
  42022=>"000100110",
  42023=>"010001011",
  42024=>"100110100",
  42025=>"101010111",
  42026=>"100000111",
  42027=>"000111010",
  42028=>"000000001",
  42029=>"010110001",
  42030=>"010111010",
  42031=>"110000110",
  42032=>"111111101",
  42033=>"111101011",
  42034=>"100000000",
  42035=>"111010000",
  42036=>"111110111",
  42037=>"010000010",
  42038=>"001111110",
  42039=>"001000011",
  42040=>"000110001",
  42041=>"001111010",
  42042=>"000000010",
  42043=>"000101011",
  42044=>"011000000",
  42045=>"011000100",
  42046=>"011001101",
  42047=>"100110011",
  42048=>"100100110",
  42049=>"000000001",
  42050=>"011010001",
  42051=>"010101000",
  42052=>"100111110",
  42053=>"110110011",
  42054=>"100101000",
  42055=>"011001101",
  42056=>"010010101",
  42057=>"011011101",
  42058=>"001000011",
  42059=>"101001100",
  42060=>"001001110",
  42061=>"110001111",
  42062=>"011110101",
  42063=>"011101010",
  42064=>"101001010",
  42065=>"001011100",
  42066=>"100010001",
  42067=>"010011010",
  42068=>"000000100",
  42069=>"010111001",
  42070=>"101001110",
  42071=>"000101001",
  42072=>"001111100",
  42073=>"110110101",
  42074=>"111011111",
  42075=>"001101110",
  42076=>"011011000",
  42077=>"100100101",
  42078=>"000101101",
  42079=>"100010011",
  42080=>"011010000",
  42081=>"011011010",
  42082=>"110000111",
  42083=>"101000000",
  42084=>"010100000",
  42085=>"011100100",
  42086=>"001110100",
  42087=>"001000111",
  42088=>"100001001",
  42089=>"110111110",
  42090=>"111100110",
  42091=>"001000000",
  42092=>"000000111",
  42093=>"001100000",
  42094=>"011010000",
  42095=>"000110000",
  42096=>"111111010",
  42097=>"000010000",
  42098=>"000110011",
  42099=>"011101111",
  42100=>"011110010",
  42101=>"010100010",
  42102=>"000000010",
  42103=>"110000011",
  42104=>"000010110",
  42105=>"011000110",
  42106=>"110010010",
  42107=>"000000100",
  42108=>"101001010",
  42109=>"001110001",
  42110=>"001110000",
  42111=>"101101000",
  42112=>"111100010",
  42113=>"100110000",
  42114=>"111110110",
  42115=>"101100010",
  42116=>"000000011",
  42117=>"000011000",
  42118=>"110100011",
  42119=>"101011000",
  42120=>"111000001",
  42121=>"000010100",
  42122=>"110110011",
  42123=>"011000010",
  42124=>"000000010",
  42125=>"001101100",
  42126=>"011111100",
  42127=>"011001000",
  42128=>"011010101",
  42129=>"101100000",
  42130=>"001111011",
  42131=>"111001111",
  42132=>"010111011",
  42133=>"001011000",
  42134=>"001010110",
  42135=>"111010100",
  42136=>"000010100",
  42137=>"111100111",
  42138=>"111000000",
  42139=>"010001001",
  42140=>"100011100",
  42141=>"101111101",
  42142=>"101001100",
  42143=>"000000010",
  42144=>"001011101",
  42145=>"011110110",
  42146=>"000001100",
  42147=>"011110001",
  42148=>"011111110",
  42149=>"111110010",
  42150=>"010011001",
  42151=>"111011001",
  42152=>"100111110",
  42153=>"100000010",
  42154=>"101010010",
  42155=>"111001101",
  42156=>"100011100",
  42157=>"111101100",
  42158=>"100101111",
  42159=>"000110010",
  42160=>"101000110",
  42161=>"101000000",
  42162=>"010001001",
  42163=>"111110010",
  42164=>"100001110",
  42165=>"010010111",
  42166=>"101110000",
  42167=>"001110000",
  42168=>"010010100",
  42169=>"100100111",
  42170=>"100010110",
  42171=>"001101000",
  42172=>"001011001",
  42173=>"011011011",
  42174=>"110011111",
  42175=>"110010000",
  42176=>"101111111",
  42177=>"000010110",
  42178=>"001101010",
  42179=>"011010001",
  42180=>"111011111",
  42181=>"000111101",
  42182=>"001100111",
  42183=>"110110011",
  42184=>"000111101",
  42185=>"010000100",
  42186=>"000111010",
  42187=>"100000010",
  42188=>"010010000",
  42189=>"111011011",
  42190=>"010000100",
  42191=>"000001101",
  42192=>"101000000",
  42193=>"111011100",
  42194=>"011111111",
  42195=>"001000111",
  42196=>"010000010",
  42197=>"111010101",
  42198=>"111000001",
  42199=>"100010110",
  42200=>"001010101",
  42201=>"011101110",
  42202=>"011101010",
  42203=>"010110000",
  42204=>"010011110",
  42205=>"111111010",
  42206=>"100011001",
  42207=>"011001101",
  42208=>"001110000",
  42209=>"001000000",
  42210=>"001010100",
  42211=>"111101010",
  42212=>"000101111",
  42213=>"101001100",
  42214=>"001110011",
  42215=>"100010001",
  42216=>"000110111",
  42217=>"010100011",
  42218=>"000110010",
  42219=>"001011011",
  42220=>"101011001",
  42221=>"111011110",
  42222=>"011101100",
  42223=>"011000010",
  42224=>"101010100",
  42225=>"001101001",
  42226=>"100011000",
  42227=>"001010001",
  42228=>"000010001",
  42229=>"101000001",
  42230=>"011000011",
  42231=>"011000001",
  42232=>"011000111",
  42233=>"100101110",
  42234=>"111111101",
  42235=>"100011010",
  42236=>"111001001",
  42237=>"011010100",
  42238=>"100111000",
  42239=>"000011010",
  42240=>"101101000",
  42241=>"001011100",
  42242=>"000111111",
  42243=>"110011100",
  42244=>"110101111",
  42245=>"000101010",
  42246=>"010111001",
  42247=>"000011100",
  42248=>"001001000",
  42249=>"110010001",
  42250=>"110110001",
  42251=>"011001000",
  42252=>"000000011",
  42253=>"100001101",
  42254=>"101110010",
  42255=>"010011100",
  42256=>"110000010",
  42257=>"011100101",
  42258=>"110011101",
  42259=>"111000011",
  42260=>"010000001",
  42261=>"110010011",
  42262=>"000001100",
  42263=>"000000101",
  42264=>"101100101",
  42265=>"111110010",
  42266=>"100110011",
  42267=>"111100100",
  42268=>"000011111",
  42269=>"101010000",
  42270=>"101100111",
  42271=>"000010000",
  42272=>"001101001",
  42273=>"110000000",
  42274=>"110101111",
  42275=>"111111110",
  42276=>"110101110",
  42277=>"000100100",
  42278=>"111010010",
  42279=>"001001010",
  42280=>"010001111",
  42281=>"111001111",
  42282=>"000001000",
  42283=>"111101001",
  42284=>"011011010",
  42285=>"010100111",
  42286=>"011001101",
  42287=>"000000001",
  42288=>"111111001",
  42289=>"010111000",
  42290=>"011100100",
  42291=>"111101101",
  42292=>"001101100",
  42293=>"000000000",
  42294=>"001001110",
  42295=>"101011100",
  42296=>"010001110",
  42297=>"001001111",
  42298=>"101100001",
  42299=>"011001110",
  42300=>"011110110",
  42301=>"111010110",
  42302=>"010100101",
  42303=>"101100100",
  42304=>"010111100",
  42305=>"001101000",
  42306=>"110000111",
  42307=>"110101101",
  42308=>"100000010",
  42309=>"011001111",
  42310=>"011010011",
  42311=>"001001001",
  42312=>"001110011",
  42313=>"110110010",
  42314=>"101010110",
  42315=>"001010010",
  42316=>"100111100",
  42317=>"110000001",
  42318=>"100111001",
  42319=>"101100110",
  42320=>"011110011",
  42321=>"001010011",
  42322=>"001110010",
  42323=>"001100011",
  42324=>"111001000",
  42325=>"010010110",
  42326=>"001000000",
  42327=>"110000101",
  42328=>"101011010",
  42329=>"110110101",
  42330=>"001111101",
  42331=>"000110011",
  42332=>"100010001",
  42333=>"001100000",
  42334=>"010001000",
  42335=>"100100001",
  42336=>"111011000",
  42337=>"110110100",
  42338=>"001101101",
  42339=>"000010100",
  42340=>"101110010",
  42341=>"000110010",
  42342=>"100101110",
  42343=>"001011011",
  42344=>"010101001",
  42345=>"001111010",
  42346=>"000100010",
  42347=>"001100000",
  42348=>"100010110",
  42349=>"101000011",
  42350=>"111111110",
  42351=>"010111101",
  42352=>"100010000",
  42353=>"000001111",
  42354=>"100111000",
  42355=>"010101011",
  42356=>"100011101",
  42357=>"001010011",
  42358=>"101001110",
  42359=>"001110000",
  42360=>"010000100",
  42361=>"000110110",
  42362=>"010110010",
  42363=>"011000001",
  42364=>"000000000",
  42365=>"111100110",
  42366=>"011001101",
  42367=>"010010000",
  42368=>"111101101",
  42369=>"010010000",
  42370=>"001001010",
  42371=>"111100101",
  42372=>"111101001",
  42373=>"011111010",
  42374=>"101010011",
  42375=>"100000010",
  42376=>"111000010",
  42377=>"100110000",
  42378=>"101100110",
  42379=>"111010100",
  42380=>"000110110",
  42381=>"000110000",
  42382=>"101000000",
  42383=>"100000100",
  42384=>"001010001",
  42385=>"000010101",
  42386=>"011110101",
  42387=>"011101100",
  42388=>"000011110",
  42389=>"000111101",
  42390=>"101011111",
  42391=>"100100000",
  42392=>"101000001",
  42393=>"010100111",
  42394=>"001010010",
  42395=>"010010101",
  42396=>"101110111",
  42397=>"000100000",
  42398=>"111111010",
  42399=>"010010000",
  42400=>"100101001",
  42401=>"110101011",
  42402=>"011010001",
  42403=>"000000011",
  42404=>"101111110",
  42405=>"100001011",
  42406=>"100101100",
  42407=>"101110000",
  42408=>"001011010",
  42409=>"101111000",
  42410=>"011111011",
  42411=>"000000011",
  42412=>"101011011",
  42413=>"101101111",
  42414=>"000100111",
  42415=>"010011010",
  42416=>"100010011",
  42417=>"011111111",
  42418=>"100111110",
  42419=>"111111001",
  42420=>"010011100",
  42421=>"101000011",
  42422=>"000101011",
  42423=>"101001100",
  42424=>"101011000",
  42425=>"001110000",
  42426=>"110110000",
  42427=>"001010000",
  42428=>"010011100",
  42429=>"111001000",
  42430=>"011011101",
  42431=>"100101000",
  42432=>"101000101",
  42433=>"111100101",
  42434=>"011010010",
  42435=>"111111011",
  42436=>"010101001",
  42437=>"001001001",
  42438=>"000100011",
  42439=>"000000000",
  42440=>"110000010",
  42441=>"100101101",
  42442=>"011011110",
  42443=>"101011100",
  42444=>"111111100",
  42445=>"101000001",
  42446=>"101011001",
  42447=>"110010101",
  42448=>"101010100",
  42449=>"101101111",
  42450=>"111110110",
  42451=>"110111000",
  42452=>"111111100",
  42453=>"010100110",
  42454=>"011000101",
  42455=>"010100011",
  42456=>"000000100",
  42457=>"110011010",
  42458=>"110110101",
  42459=>"010100000",
  42460=>"001010100",
  42461=>"010101010",
  42462=>"011110100",
  42463=>"011110001",
  42464=>"011100010",
  42465=>"011010111",
  42466=>"010011001",
  42467=>"010110100",
  42468=>"111010101",
  42469=>"010000111",
  42470=>"010100010",
  42471=>"011000000",
  42472=>"010110000",
  42473=>"011100110",
  42474=>"011100011",
  42475=>"100101010",
  42476=>"010110010",
  42477=>"101011100",
  42478=>"111101100",
  42479=>"001011101",
  42480=>"111001111",
  42481=>"110011100",
  42482=>"110111100",
  42483=>"111010111",
  42484=>"011000001",
  42485=>"001000000",
  42486=>"010110011",
  42487=>"100110001",
  42488=>"100001001",
  42489=>"111111000",
  42490=>"011100011",
  42491=>"001110001",
  42492=>"101011011",
  42493=>"111010101",
  42494=>"011101101",
  42495=>"001111101",
  42496=>"000111110",
  42497=>"011111011",
  42498=>"010000100",
  42499=>"110001000",
  42500=>"110011000",
  42501=>"111100001",
  42502=>"001011101",
  42503=>"001001011",
  42504=>"001001000",
  42505=>"111011000",
  42506=>"011100100",
  42507=>"111011000",
  42508=>"101110001",
  42509=>"110111010",
  42510=>"011000101",
  42511=>"001000100",
  42512=>"000001010",
  42513=>"101000111",
  42514=>"101111111",
  42515=>"010010001",
  42516=>"000100001",
  42517=>"111010001",
  42518=>"100101111",
  42519=>"010001101",
  42520=>"010010001",
  42521=>"000000110",
  42522=>"011101000",
  42523=>"010000010",
  42524=>"011101111",
  42525=>"011101111",
  42526=>"101101010",
  42527=>"110110011",
  42528=>"000011101",
  42529=>"101010000",
  42530=>"001110110",
  42531=>"101000000",
  42532=>"101111100",
  42533=>"101010001",
  42534=>"010000000",
  42535=>"111010010",
  42536=>"100001100",
  42537=>"001011100",
  42538=>"111010111",
  42539=>"110011001",
  42540=>"001100001",
  42541=>"010011110",
  42542=>"100000101",
  42543=>"000000101",
  42544=>"111111110",
  42545=>"111100001",
  42546=>"010000001",
  42547=>"101001110",
  42548=>"010101100",
  42549=>"000101010",
  42550=>"101111010",
  42551=>"111001001",
  42552=>"111110111",
  42553=>"110011100",
  42554=>"110110110",
  42555=>"000100101",
  42556=>"000100000",
  42557=>"001100110",
  42558=>"000000101",
  42559=>"001011101",
  42560=>"000100010",
  42561=>"110111000",
  42562=>"100101000",
  42563=>"011000010",
  42564=>"110000000",
  42565=>"010111101",
  42566=>"010110110",
  42567=>"101001100",
  42568=>"001000111",
  42569=>"010010000",
  42570=>"000110100",
  42571=>"011011100",
  42572=>"010011010",
  42573=>"101110100",
  42574=>"010100000",
  42575=>"010011010",
  42576=>"001011111",
  42577=>"111111101",
  42578=>"110111001",
  42579=>"110011001",
  42580=>"110001001",
  42581=>"111010111",
  42582=>"011110000",
  42583=>"001100011",
  42584=>"111000000",
  42585=>"010101101",
  42586=>"111010110",
  42587=>"001101000",
  42588=>"011010001",
  42589=>"100001101",
  42590=>"100001011",
  42591=>"101001111",
  42592=>"000010001",
  42593=>"001101101",
  42594=>"101001010",
  42595=>"010100000",
  42596=>"011111101",
  42597=>"000111000",
  42598=>"111111101",
  42599=>"000111011",
  42600=>"101100100",
  42601=>"000001001",
  42602=>"101110001",
  42603=>"111101100",
  42604=>"101111000",
  42605=>"001101000",
  42606=>"000011100",
  42607=>"101111110",
  42608=>"110011001",
  42609=>"001011111",
  42610=>"100011000",
  42611=>"011011100",
  42612=>"010001010",
  42613=>"100100000",
  42614=>"111011011",
  42615=>"101011111",
  42616=>"010011000",
  42617=>"110011001",
  42618=>"000101101",
  42619=>"000110001",
  42620=>"010010011",
  42621=>"001000110",
  42622=>"011011111",
  42623=>"101100111",
  42624=>"111101011",
  42625=>"101110011",
  42626=>"011101001",
  42627=>"100100101",
  42628=>"011000111",
  42629=>"111110011",
  42630=>"100101000",
  42631=>"110111011",
  42632=>"001001100",
  42633=>"100101001",
  42634=>"001001000",
  42635=>"000110111",
  42636=>"001100001",
  42637=>"101100111",
  42638=>"011101101",
  42639=>"010010011",
  42640=>"010100101",
  42641=>"100000001",
  42642=>"010100010",
  42643=>"110000111",
  42644=>"001101010",
  42645=>"100101001",
  42646=>"000110100",
  42647=>"011110011",
  42648=>"101101010",
  42649=>"111101111",
  42650=>"111011011",
  42651=>"101010001",
  42652=>"010000111",
  42653=>"000000001",
  42654=>"100110000",
  42655=>"110111010",
  42656=>"111100111",
  42657=>"011100000",
  42658=>"111100111",
  42659=>"101101110",
  42660=>"111000000",
  42661=>"111010110",
  42662=>"000100101",
  42663=>"010011100",
  42664=>"111000010",
  42665=>"011010010",
  42666=>"011111100",
  42667=>"101000111",
  42668=>"011000001",
  42669=>"011110110",
  42670=>"110001100",
  42671=>"011001001",
  42672=>"010100000",
  42673=>"111100011",
  42674=>"101111101",
  42675=>"000001001",
  42676=>"010001000",
  42677=>"001111011",
  42678=>"111100101",
  42679=>"111011000",
  42680=>"010010110",
  42681=>"101101011",
  42682=>"101010000",
  42683=>"011010100",
  42684=>"101100110",
  42685=>"101010000",
  42686=>"110010110",
  42687=>"011001001",
  42688=>"001111111",
  42689=>"010111010",
  42690=>"000001011",
  42691=>"100110001",
  42692=>"000100111",
  42693=>"111101110",
  42694=>"110011000",
  42695=>"110111010",
  42696=>"111111100",
  42697=>"101011101",
  42698=>"011101011",
  42699=>"111000011",
  42700=>"010110111",
  42701=>"001110101",
  42702=>"000110001",
  42703=>"011000101",
  42704=>"100111110",
  42705=>"101000111",
  42706=>"000010101",
  42707=>"011000110",
  42708=>"101101110",
  42709=>"100010100",
  42710=>"010100110",
  42711=>"100011111",
  42712=>"111011001",
  42713=>"100011000",
  42714=>"101101001",
  42715=>"101101101",
  42716=>"110101110",
  42717=>"111000000",
  42718=>"100000001",
  42719=>"101110011",
  42720=>"110000100",
  42721=>"101010001",
  42722=>"001101111",
  42723=>"100110110",
  42724=>"101001110",
  42725=>"000101111",
  42726=>"101001101",
  42727=>"100000101",
  42728=>"000110010",
  42729=>"100111001",
  42730=>"011111010",
  42731=>"011101010",
  42732=>"011101110",
  42733=>"001100110",
  42734=>"111101001",
  42735=>"100001110",
  42736=>"110010110",
  42737=>"010001000",
  42738=>"100000000",
  42739=>"001100100",
  42740=>"100001001",
  42741=>"000010001",
  42742=>"111000110",
  42743=>"011011011",
  42744=>"101100110",
  42745=>"010101110",
  42746=>"010011011",
  42747=>"100000011",
  42748=>"010000001",
  42749=>"111100100",
  42750=>"110000010",
  42751=>"110000110",
  42752=>"000000110",
  42753=>"111000100",
  42754=>"111101110",
  42755=>"011011110",
  42756=>"110011111",
  42757=>"001000001",
  42758=>"001100001",
  42759=>"101100101",
  42760=>"011011001",
  42761=>"111100010",
  42762=>"011011101",
  42763=>"000010110",
  42764=>"100010100",
  42765=>"101011111",
  42766=>"110100101",
  42767=>"010011111",
  42768=>"110000110",
  42769=>"000001001",
  42770=>"001001100",
  42771=>"010111110",
  42772=>"001101111",
  42773=>"110100100",
  42774=>"010100100",
  42775=>"001000000",
  42776=>"111100010",
  42777=>"100000100",
  42778=>"010001110",
  42779=>"000011001",
  42780=>"101111000",
  42781=>"011111011",
  42782=>"011011001",
  42783=>"011110101",
  42784=>"101011111",
  42785=>"010010101",
  42786=>"000001000",
  42787=>"000100110",
  42788=>"001101011",
  42789=>"001110110",
  42790=>"011001110",
  42791=>"010100101",
  42792=>"110011001",
  42793=>"000110110",
  42794=>"010100110",
  42795=>"010100010",
  42796=>"110001111",
  42797=>"111010010",
  42798=>"000101000",
  42799=>"001000110",
  42800=>"000001011",
  42801=>"010000001",
  42802=>"010011100",
  42803=>"001000111",
  42804=>"100011010",
  42805=>"000000011",
  42806=>"110110111",
  42807=>"101111011",
  42808=>"010101010",
  42809=>"010011011",
  42810=>"000100010",
  42811=>"010110000",
  42812=>"010011101",
  42813=>"001001010",
  42814=>"010011111",
  42815=>"010111101",
  42816=>"111000000",
  42817=>"111101111",
  42818=>"110011001",
  42819=>"001011101",
  42820=>"000000010",
  42821=>"010101100",
  42822=>"110001001",
  42823=>"000001010",
  42824=>"100001011",
  42825=>"100000110",
  42826=>"100000001",
  42827=>"000000010",
  42828=>"001010100",
  42829=>"110000000",
  42830=>"100000011",
  42831=>"000110110",
  42832=>"100000000",
  42833=>"110000100",
  42834=>"110001010",
  42835=>"111010101",
  42836=>"110010010",
  42837=>"101011011",
  42838=>"101111100",
  42839=>"010010011",
  42840=>"111111101",
  42841=>"000000001",
  42842=>"101001000",
  42843=>"010101000",
  42844=>"010101100",
  42845=>"010110111",
  42846=>"100111010",
  42847=>"000100010",
  42848=>"010011001",
  42849=>"100010011",
  42850=>"000111110",
  42851=>"011100001",
  42852=>"010101001",
  42853=>"111111010",
  42854=>"001001111",
  42855=>"001010011",
  42856=>"111111001",
  42857=>"000110001",
  42858=>"000101000",
  42859=>"110010001",
  42860=>"110111111",
  42861=>"001101010",
  42862=>"000001100",
  42863=>"111111101",
  42864=>"111001010",
  42865=>"101100000",
  42866=>"000010001",
  42867=>"011011111",
  42868=>"101111111",
  42869=>"100001110",
  42870=>"101011010",
  42871=>"010100100",
  42872=>"100110001",
  42873=>"111001000",
  42874=>"110111010",
  42875=>"000000110",
  42876=>"110011000",
  42877=>"101010011",
  42878=>"110001010",
  42879=>"101101001",
  42880=>"011011111",
  42881=>"110110010",
  42882=>"100110110",
  42883=>"111010100",
  42884=>"110001101",
  42885=>"100000000",
  42886=>"010111111",
  42887=>"110010011",
  42888=>"111101000",
  42889=>"010100001",
  42890=>"011110011",
  42891=>"001010111",
  42892=>"110100100",
  42893=>"110110001",
  42894=>"111110011",
  42895=>"111101100",
  42896=>"000001111",
  42897=>"111101011",
  42898=>"001010111",
  42899=>"111001111",
  42900=>"000110010",
  42901=>"000000100",
  42902=>"001001010",
  42903=>"110101110",
  42904=>"100010010",
  42905=>"011111000",
  42906=>"001000111",
  42907=>"110101010",
  42908=>"010001111",
  42909=>"111110100",
  42910=>"000111011",
  42911=>"110101000",
  42912=>"100011101",
  42913=>"000000101",
  42914=>"100011010",
  42915=>"011001101",
  42916=>"001000000",
  42917=>"001101000",
  42918=>"000010001",
  42919=>"111001011",
  42920=>"010001011",
  42921=>"000100010",
  42922=>"010110101",
  42923=>"110011111",
  42924=>"101011000",
  42925=>"010011110",
  42926=>"111000111",
  42927=>"111111010",
  42928=>"011101111",
  42929=>"000101010",
  42930=>"101111011",
  42931=>"101100111",
  42932=>"000011011",
  42933=>"001001010",
  42934=>"100110011",
  42935=>"111000100",
  42936=>"011001110",
  42937=>"100111111",
  42938=>"101011001",
  42939=>"011001011",
  42940=>"010100110",
  42941=>"110000111",
  42942=>"101011000",
  42943=>"001100001",
  42944=>"111101111",
  42945=>"000101100",
  42946=>"110111110",
  42947=>"010010101",
  42948=>"000010011",
  42949=>"001001101",
  42950=>"010000101",
  42951=>"110111101",
  42952=>"010110111",
  42953=>"101011100",
  42954=>"011110001",
  42955=>"000111100",
  42956=>"000111101",
  42957=>"100100101",
  42958=>"000010100",
  42959=>"110001100",
  42960=>"101011110",
  42961=>"100011110",
  42962=>"001001111",
  42963=>"101011101",
  42964=>"110000010",
  42965=>"001110011",
  42966=>"111001000",
  42967=>"000100000",
  42968=>"010111110",
  42969=>"010110101",
  42970=>"111111001",
  42971=>"110000100",
  42972=>"001101000",
  42973=>"111011111",
  42974=>"000011101",
  42975=>"101101010",
  42976=>"101011010",
  42977=>"000111000",
  42978=>"111100011",
  42979=>"000100000",
  42980=>"011010111",
  42981=>"010011001",
  42982=>"001100010",
  42983=>"010110000",
  42984=>"110001001",
  42985=>"011010100",
  42986=>"100111101",
  42987=>"111101011",
  42988=>"000101000",
  42989=>"101011111",
  42990=>"011000100",
  42991=>"001001000",
  42992=>"011001010",
  42993=>"000111000",
  42994=>"111100101",
  42995=>"111100011",
  42996=>"110011001",
  42997=>"011101000",
  42998=>"001110100",
  42999=>"111000100",
  43000=>"110010011",
  43001=>"011011111",
  43002=>"001001011",
  43003=>"110100010",
  43004=>"111010000",
  43005=>"011110100",
  43006=>"000001010",
  43007=>"101110000",
  43008=>"111100110",
  43009=>"100011011",
  43010=>"011001111",
  43011=>"000100011",
  43012=>"100101000",
  43013=>"111011010",
  43014=>"010010011",
  43015=>"010101001",
  43016=>"000011001",
  43017=>"010010000",
  43018=>"000010111",
  43019=>"011011001",
  43020=>"000101011",
  43021=>"101111010",
  43022=>"100011011",
  43023=>"100100001",
  43024=>"111101100",
  43025=>"100001000",
  43026=>"100100101",
  43027=>"000000100",
  43028=>"111111111",
  43029=>"000111010",
  43030=>"101101110",
  43031=>"110001010",
  43032=>"101111010",
  43033=>"011001110",
  43034=>"100101101",
  43035=>"101111110",
  43036=>"001100010",
  43037=>"010101100",
  43038=>"100010110",
  43039=>"000110000",
  43040=>"110001000",
  43041=>"100010010",
  43042=>"101110011",
  43043=>"000101100",
  43044=>"110100010",
  43045=>"101110010",
  43046=>"110000010",
  43047=>"000000111",
  43048=>"000111001",
  43049=>"110000010",
  43050=>"101110100",
  43051=>"000010111",
  43052=>"000000101",
  43053=>"111001100",
  43054=>"011001100",
  43055=>"110110000",
  43056=>"101010000",
  43057=>"011101011",
  43058=>"101111110",
  43059=>"011101011",
  43060=>"011101011",
  43061=>"000110110",
  43062=>"111001110",
  43063=>"101111011",
  43064=>"001001101",
  43065=>"001100100",
  43066=>"000010000",
  43067=>"110100001",
  43068=>"010100010",
  43069=>"001101111",
  43070=>"000001100",
  43071=>"000110011",
  43072=>"000010101",
  43073=>"000011000",
  43074=>"010010111",
  43075=>"111001010",
  43076=>"111001110",
  43077=>"011100110",
  43078=>"000101101",
  43079=>"000111000",
  43080=>"011101011",
  43081=>"110110111",
  43082=>"110010110",
  43083=>"000110011",
  43084=>"010110010",
  43085=>"100101110",
  43086=>"110001110",
  43087=>"001101000",
  43088=>"111100110",
  43089=>"111101010",
  43090=>"101100100",
  43091=>"010100011",
  43092=>"110111011",
  43093=>"010001000",
  43094=>"000000000",
  43095=>"001000110",
  43096=>"111000111",
  43097=>"010010101",
  43098=>"111010100",
  43099=>"001001011",
  43100=>"100010110",
  43101=>"001000010",
  43102=>"011011000",
  43103=>"110100011",
  43104=>"111111010",
  43105=>"101100010",
  43106=>"011000100",
  43107=>"111111100",
  43108=>"010100001",
  43109=>"000111000",
  43110=>"111111111",
  43111=>"011110101",
  43112=>"011100101",
  43113=>"110000100",
  43114=>"111000010",
  43115=>"011110001",
  43116=>"101000011",
  43117=>"101101100",
  43118=>"000101111",
  43119=>"001001000",
  43120=>"100001011",
  43121=>"000010000",
  43122=>"100011111",
  43123=>"111100111",
  43124=>"110111100",
  43125=>"011001000",
  43126=>"101010010",
  43127=>"110001111",
  43128=>"010011000",
  43129=>"000000010",
  43130=>"010101110",
  43131=>"111001101",
  43132=>"111110111",
  43133=>"010100100",
  43134=>"111111101",
  43135=>"010101000",
  43136=>"001111110",
  43137=>"010001000",
  43138=>"111010000",
  43139=>"101000000",
  43140=>"101001000",
  43141=>"000000100",
  43142=>"011010110",
  43143=>"000010010",
  43144=>"101100110",
  43145=>"111111010",
  43146=>"010110000",
  43147=>"000110111",
  43148=>"101001010",
  43149=>"000110001",
  43150=>"010010010",
  43151=>"111010110",
  43152=>"111110001",
  43153=>"000011011",
  43154=>"000110011",
  43155=>"111011110",
  43156=>"110011100",
  43157=>"000111001",
  43158=>"010011100",
  43159=>"111110000",
  43160=>"000101011",
  43161=>"101001111",
  43162=>"011011110",
  43163=>"001001101",
  43164=>"101111110",
  43165=>"110111000",
  43166=>"001010110",
  43167=>"111111000",
  43168=>"010111111",
  43169=>"101000010",
  43170=>"011101000",
  43171=>"111110100",
  43172=>"010111101",
  43173=>"100010100",
  43174=>"001111001",
  43175=>"011010110",
  43176=>"010001100",
  43177=>"100001110",
  43178=>"111001110",
  43179=>"010000101",
  43180=>"011111010",
  43181=>"001111010",
  43182=>"111001011",
  43183=>"101011000",
  43184=>"000001001",
  43185=>"011010010",
  43186=>"101110011",
  43187=>"010001101",
  43188=>"101000111",
  43189=>"110010000",
  43190=>"001000111",
  43191=>"110000101",
  43192=>"010110001",
  43193=>"001000011",
  43194=>"100001100",
  43195=>"000110000",
  43196=>"000111100",
  43197=>"001000010",
  43198=>"011111100",
  43199=>"011010111",
  43200=>"010001010",
  43201=>"010101111",
  43202=>"011110101",
  43203=>"000100000",
  43204=>"011001010",
  43205=>"001011011",
  43206=>"100100111",
  43207=>"010111000",
  43208=>"010010000",
  43209=>"111110101",
  43210=>"100001011",
  43211=>"001110010",
  43212=>"101001110",
  43213=>"001011010",
  43214=>"001010100",
  43215=>"010011011",
  43216=>"010100000",
  43217=>"010000100",
  43218=>"100000110",
  43219=>"010111001",
  43220=>"000101100",
  43221=>"010001010",
  43222=>"101111110",
  43223=>"111101100",
  43224=>"111100001",
  43225=>"110101110",
  43226=>"011101000",
  43227=>"010110010",
  43228=>"101010111",
  43229=>"010000011",
  43230=>"001001110",
  43231=>"100100110",
  43232=>"101000110",
  43233=>"100000011",
  43234=>"101010010",
  43235=>"000100011",
  43236=>"110000011",
  43237=>"101111001",
  43238=>"001111100",
  43239=>"011111011",
  43240=>"001111101",
  43241=>"111000100",
  43242=>"101100110",
  43243=>"011001001",
  43244=>"000110101",
  43245=>"101111111",
  43246=>"011011100",
  43247=>"100001100",
  43248=>"001101011",
  43249=>"010111111",
  43250=>"101101010",
  43251=>"101101001",
  43252=>"001100101",
  43253=>"100011101",
  43254=>"101001010",
  43255=>"110100101",
  43256=>"000010100",
  43257=>"100011101",
  43258=>"001100101",
  43259=>"110000100",
  43260=>"000011110",
  43261=>"011001100",
  43262=>"000110001",
  43263=>"111100011",
  43264=>"111000001",
  43265=>"100000101",
  43266=>"100110010",
  43267=>"010010101",
  43268=>"000101000",
  43269=>"111011001",
  43270=>"010100000",
  43271=>"111111011",
  43272=>"110000100",
  43273=>"000001111",
  43274=>"001011110",
  43275=>"000010110",
  43276=>"101110010",
  43277=>"100000011",
  43278=>"001111101",
  43279=>"010010111",
  43280=>"011110111",
  43281=>"111100010",
  43282=>"010111111",
  43283=>"010000011",
  43284=>"000010000",
  43285=>"010011000",
  43286=>"010000101",
  43287=>"000110101",
  43288=>"000101100",
  43289=>"111100000",
  43290=>"111100011",
  43291=>"011001000",
  43292=>"001111000",
  43293=>"110000101",
  43294=>"101111010",
  43295=>"000000001",
  43296=>"000100001",
  43297=>"111010101",
  43298=>"111101110",
  43299=>"100101110",
  43300=>"010100101",
  43301=>"100111001",
  43302=>"010100001",
  43303=>"001001011",
  43304=>"100000101",
  43305=>"111101010",
  43306=>"100100010",
  43307=>"000111100",
  43308=>"100111000",
  43309=>"111100001",
  43310=>"010110001",
  43311=>"000000110",
  43312=>"010010000",
  43313=>"111000011",
  43314=>"100101111",
  43315=>"100110101",
  43316=>"110000010",
  43317=>"000011111",
  43318=>"000110110",
  43319=>"000100000",
  43320=>"110110010",
  43321=>"101101101",
  43322=>"001100100",
  43323=>"111101101",
  43324=>"100000110",
  43325=>"011111110",
  43326=>"101100010",
  43327=>"000001001",
  43328=>"001100000",
  43329=>"011111100",
  43330=>"111011110",
  43331=>"100101001",
  43332=>"010010111",
  43333=>"100101011",
  43334=>"001111000",
  43335=>"100111111",
  43336=>"010001000",
  43337=>"001110000",
  43338=>"000001010",
  43339=>"000100011",
  43340=>"111010110",
  43341=>"001000100",
  43342=>"110101000",
  43343=>"101101101",
  43344=>"101001011",
  43345=>"100000000",
  43346=>"001011001",
  43347=>"010110001",
  43348=>"100101001",
  43349=>"111101111",
  43350=>"010001101",
  43351=>"111111101",
  43352=>"000010010",
  43353=>"001111011",
  43354=>"011101010",
  43355=>"010001011",
  43356=>"111000111",
  43357=>"101100111",
  43358=>"100010111",
  43359=>"010000110",
  43360=>"100110000",
  43361=>"011010000",
  43362=>"000001010",
  43363=>"010111101",
  43364=>"110001101",
  43365=>"010101100",
  43366=>"111101010",
  43367=>"010000010",
  43368=>"000100000",
  43369=>"111110001",
  43370=>"110001100",
  43371=>"101101000",
  43372=>"101111110",
  43373=>"111110110",
  43374=>"101101000",
  43375=>"000111010",
  43376=>"001100001",
  43377=>"001011011",
  43378=>"001110100",
  43379=>"111100000",
  43380=>"100111011",
  43381=>"001011001",
  43382=>"100001100",
  43383=>"010011111",
  43384=>"101011011",
  43385=>"100100100",
  43386=>"101001100",
  43387=>"011000010",
  43388=>"010011001",
  43389=>"101111011",
  43390=>"100111110",
  43391=>"111111000",
  43392=>"101011000",
  43393=>"010001001",
  43394=>"100001011",
  43395=>"111000110",
  43396=>"101000000",
  43397=>"000100000",
  43398=>"011111111",
  43399=>"111001000",
  43400=>"000110001",
  43401=>"010110001",
  43402=>"001010100",
  43403=>"111100001",
  43404=>"100111000",
  43405=>"001001101",
  43406=>"001010011",
  43407=>"010000001",
  43408=>"000110010",
  43409=>"011111101",
  43410=>"100111110",
  43411=>"000001010",
  43412=>"101000010",
  43413=>"100111100",
  43414=>"100100001",
  43415=>"111001000",
  43416=>"000000110",
  43417=>"010000001",
  43418=>"111111011",
  43419=>"011001010",
  43420=>"010000101",
  43421=>"111100111",
  43422=>"011011111",
  43423=>"000100100",
  43424=>"111010110",
  43425=>"011100001",
  43426=>"011110100",
  43427=>"001110000",
  43428=>"101101001",
  43429=>"101100000",
  43430=>"010111000",
  43431=>"111111100",
  43432=>"010101100",
  43433=>"101010110",
  43434=>"001111110",
  43435=>"100111100",
  43436=>"110111011",
  43437=>"010010110",
  43438=>"010001110",
  43439=>"110010010",
  43440=>"010111001",
  43441=>"111000010",
  43442=>"110001100",
  43443=>"011011001",
  43444=>"011011110",
  43445=>"110011010",
  43446=>"000100011",
  43447=>"001100111",
  43448=>"000001111",
  43449=>"010001110",
  43450=>"101100110",
  43451=>"100011101",
  43452=>"110010000",
  43453=>"101111111",
  43454=>"101001000",
  43455=>"101110110",
  43456=>"100101111",
  43457=>"011001001",
  43458=>"110010000",
  43459=>"001100100",
  43460=>"010101011",
  43461=>"010110100",
  43462=>"001011011",
  43463=>"001001110",
  43464=>"011000110",
  43465=>"010010100",
  43466=>"101011111",
  43467=>"001011010",
  43468=>"111101011",
  43469=>"111101011",
  43470=>"001100011",
  43471=>"110011101",
  43472=>"100111101",
  43473=>"111010001",
  43474=>"010110011",
  43475=>"011100111",
  43476=>"111100000",
  43477=>"100110101",
  43478=>"111000010",
  43479=>"000101111",
  43480=>"010101010",
  43481=>"011010110",
  43482=>"100101100",
  43483=>"011001110",
  43484=>"000011111",
  43485=>"000010111",
  43486=>"011001010",
  43487=>"010010111",
  43488=>"000101010",
  43489=>"110111000",
  43490=>"000010000",
  43491=>"011100000",
  43492=>"100001010",
  43493=>"101000001",
  43494=>"101010111",
  43495=>"111000111",
  43496=>"001101110",
  43497=>"110111011",
  43498=>"111111000",
  43499=>"111000101",
  43500=>"110101011",
  43501=>"000100111",
  43502=>"001111001",
  43503=>"001110111",
  43504=>"111001110",
  43505=>"001100111",
  43506=>"010110001",
  43507=>"111110110",
  43508=>"100100101",
  43509=>"111010010",
  43510=>"100000101",
  43511=>"000001110",
  43512=>"000110000",
  43513=>"110100010",
  43514=>"011110000",
  43515=>"100000110",
  43516=>"001001010",
  43517=>"110000000",
  43518=>"000000101",
  43519=>"011011001",
  43520=>"011111111",
  43521=>"011001110",
  43522=>"000100010",
  43523=>"000010101",
  43524=>"000100100",
  43525=>"101100011",
  43526=>"111111011",
  43527=>"011010110",
  43528=>"111001011",
  43529=>"011000110",
  43530=>"111000101",
  43531=>"101000111",
  43532=>"110101000",
  43533=>"111001001",
  43534=>"100000001",
  43535=>"001101011",
  43536=>"001011110",
  43537=>"101011011",
  43538=>"100011111",
  43539=>"000110110",
  43540=>"111110001",
  43541=>"001001000",
  43542=>"101101100",
  43543=>"000011010",
  43544=>"001011110",
  43545=>"000110101",
  43546=>"001011111",
  43547=>"001111010",
  43548=>"001011001",
  43549=>"100001110",
  43550=>"100110000",
  43551=>"001010010",
  43552=>"000110011",
  43553=>"111001001",
  43554=>"000000001",
  43555=>"101100001",
  43556=>"111111011",
  43557=>"010101010",
  43558=>"100101010",
  43559=>"001000011",
  43560=>"110001110",
  43561=>"010110001",
  43562=>"111001110",
  43563=>"011111001",
  43564=>"011001011",
  43565=>"110011110",
  43566=>"001111100",
  43567=>"011011111",
  43568=>"000000001",
  43569=>"000011011",
  43570=>"101010100",
  43571=>"010000100",
  43572=>"101001111",
  43573=>"110011001",
  43574=>"001001001",
  43575=>"100011001",
  43576=>"011110111",
  43577=>"011101010",
  43578=>"001001111",
  43579=>"011001100",
  43580=>"100110110",
  43581=>"100111100",
  43582=>"111001001",
  43583=>"111010000",
  43584=>"001110010",
  43585=>"101111101",
  43586=>"000000111",
  43587=>"010001010",
  43588=>"111111100",
  43589=>"010001000",
  43590=>"000000101",
  43591=>"000000010",
  43592=>"111000001",
  43593=>"010001110",
  43594=>"000100000",
  43595=>"111100001",
  43596=>"110000001",
  43597=>"100111101",
  43598=>"000001110",
  43599=>"111001111",
  43600=>"101010011",
  43601=>"011100000",
  43602=>"000011100",
  43603=>"000110110",
  43604=>"101111100",
  43605=>"010010111",
  43606=>"011101111",
  43607=>"010001000",
  43608=>"001000000",
  43609=>"100010000",
  43610=>"001100010",
  43611=>"100000001",
  43612=>"110000011",
  43613=>"010010001",
  43614=>"101101011",
  43615=>"110111111",
  43616=>"110000010",
  43617=>"111011011",
  43618=>"111111010",
  43619=>"001110001",
  43620=>"110100111",
  43621=>"010010111",
  43622=>"001000010",
  43623=>"000000110",
  43624=>"100010100",
  43625=>"010100111",
  43626=>"010011110",
  43627=>"101001111",
  43628=>"001101100",
  43629=>"101001110",
  43630=>"101000110",
  43631=>"101011000",
  43632=>"100100111",
  43633=>"000001000",
  43634=>"011100010",
  43635=>"011000100",
  43636=>"010100000",
  43637=>"100110100",
  43638=>"011011000",
  43639=>"010100110",
  43640=>"010011111",
  43641=>"100001011",
  43642=>"111111011",
  43643=>"111111000",
  43644=>"001100111",
  43645=>"110001001",
  43646=>"011010110",
  43647=>"100001000",
  43648=>"001100001",
  43649=>"001110110",
  43650=>"110000001",
  43651=>"001010000",
  43652=>"111010011",
  43653=>"000101100",
  43654=>"111110001",
  43655=>"100111010",
  43656=>"110000110",
  43657=>"111000101",
  43658=>"111001100",
  43659=>"010110100",
  43660=>"010011110",
  43661=>"101000001",
  43662=>"011101101",
  43663=>"101001011",
  43664=>"100001111",
  43665=>"110010001",
  43666=>"001111110",
  43667=>"001111000",
  43668=>"101000010",
  43669=>"101011111",
  43670=>"101101001",
  43671=>"001011100",
  43672=>"000111100",
  43673=>"111011000",
  43674=>"011011001",
  43675=>"100010110",
  43676=>"010000011",
  43677=>"000101011",
  43678=>"001001000",
  43679=>"111010100",
  43680=>"110110111",
  43681=>"110000100",
  43682=>"111111110",
  43683=>"001000010",
  43684=>"101001100",
  43685=>"100000001",
  43686=>"100001111",
  43687=>"111100100",
  43688=>"111110001",
  43689=>"000111000",
  43690=>"010000011",
  43691=>"001101010",
  43692=>"111100010",
  43693=>"100000000",
  43694=>"101111010",
  43695=>"011101011",
  43696=>"001011010",
  43697=>"101001110",
  43698=>"011111110",
  43699=>"110000110",
  43700=>"100000100",
  43701=>"111101111",
  43702=>"010100100",
  43703=>"100001001",
  43704=>"001111101",
  43705=>"101000110",
  43706=>"011110110",
  43707=>"011101111",
  43708=>"000001111",
  43709=>"001100101",
  43710=>"110000010",
  43711=>"011110110",
  43712=>"111000111",
  43713=>"011111011",
  43714=>"001100000",
  43715=>"100011110",
  43716=>"010111010",
  43717=>"100100011",
  43718=>"101101100",
  43719=>"100000010",
  43720=>"101001110",
  43721=>"000111101",
  43722=>"000100001",
  43723=>"100101100",
  43724=>"110110011",
  43725=>"000010010",
  43726=>"110011111",
  43727=>"111001001",
  43728=>"010011000",
  43729=>"110000111",
  43730=>"111011011",
  43731=>"110100111",
  43732=>"000101111",
  43733=>"101000001",
  43734=>"110110001",
  43735=>"001011011",
  43736=>"000110100",
  43737=>"101100000",
  43738=>"101011110",
  43739=>"000001100",
  43740=>"010111110",
  43741=>"010011110",
  43742=>"000011011",
  43743=>"010100010",
  43744=>"101111010",
  43745=>"111001100",
  43746=>"010010000",
  43747=>"000101000",
  43748=>"010001000",
  43749=>"110101101",
  43750=>"101010000",
  43751=>"111111010",
  43752=>"101010111",
  43753=>"000101100",
  43754=>"101001100",
  43755=>"100110010",
  43756=>"101110010",
  43757=>"011000110",
  43758=>"110100010",
  43759=>"010101000",
  43760=>"111010001",
  43761=>"011100100",
  43762=>"011111100",
  43763=>"010110110",
  43764=>"010000111",
  43765=>"111000010",
  43766=>"111001000",
  43767=>"111101101",
  43768=>"101110010",
  43769=>"110111010",
  43770=>"000000010",
  43771=>"111111100",
  43772=>"110000100",
  43773=>"110110101",
  43774=>"001101001",
  43775=>"111000111",
  43776=>"110111111",
  43777=>"001010100",
  43778=>"000111000",
  43779=>"000000000",
  43780=>"011100101",
  43781=>"101000110",
  43782=>"000110011",
  43783=>"010101000",
  43784=>"111011001",
  43785=>"011100001",
  43786=>"000010010",
  43787=>"000110001",
  43788=>"010001110",
  43789=>"011000111",
  43790=>"111001110",
  43791=>"100101101",
  43792=>"101100111",
  43793=>"000001101",
  43794=>"011101101",
  43795=>"100110011",
  43796=>"000110000",
  43797=>"101100001",
  43798=>"001011001",
  43799=>"000010010",
  43800=>"110110011",
  43801=>"100000111",
  43802=>"000000100",
  43803=>"110001000",
  43804=>"110110110",
  43805=>"101111100",
  43806=>"011110111",
  43807=>"101010001",
  43808=>"011100110",
  43809=>"110100011",
  43810=>"001111111",
  43811=>"001111101",
  43812=>"011101011",
  43813=>"010001111",
  43814=>"001101000",
  43815=>"000110100",
  43816=>"000110111",
  43817=>"100001100",
  43818=>"001000011",
  43819=>"000111001",
  43820=>"111011110",
  43821=>"001011011",
  43822=>"101010111",
  43823=>"001011110",
  43824=>"000110110",
  43825=>"010110000",
  43826=>"110010110",
  43827=>"001100100",
  43828=>"011001011",
  43829=>"100011011",
  43830=>"010010001",
  43831=>"110010000",
  43832=>"110001110",
  43833=>"110000011",
  43834=>"100111100",
  43835=>"101000111",
  43836=>"000101101",
  43837=>"010100100",
  43838=>"011101000",
  43839=>"101000110",
  43840=>"011011100",
  43841=>"001110011",
  43842=>"001101010",
  43843=>"110010101",
  43844=>"100001101",
  43845=>"010001110",
  43846=>"100011010",
  43847=>"011011010",
  43848=>"001101011",
  43849=>"100010010",
  43850=>"101111010",
  43851=>"001101010",
  43852=>"111111101",
  43853=>"011001010",
  43854=>"101001111",
  43855=>"101000110",
  43856=>"110011111",
  43857=>"001101100",
  43858=>"101100000",
  43859=>"111100111",
  43860=>"001001110",
  43861=>"111110100",
  43862=>"111100110",
  43863=>"101110101",
  43864=>"110110011",
  43865=>"001101100",
  43866=>"111011011",
  43867=>"010100000",
  43868=>"001110000",
  43869=>"011010010",
  43870=>"111101000",
  43871=>"000111111",
  43872=>"011101010",
  43873=>"010101100",
  43874=>"000101111",
  43875=>"100010101",
  43876=>"110100101",
  43877=>"111100010",
  43878=>"010001000",
  43879=>"100011100",
  43880=>"110001001",
  43881=>"011000101",
  43882=>"010000110",
  43883=>"100110101",
  43884=>"000010100",
  43885=>"011101100",
  43886=>"010110110",
  43887=>"000011010",
  43888=>"111001011",
  43889=>"011001010",
  43890=>"110010010",
  43891=>"111001100",
  43892=>"000101110",
  43893=>"001101001",
  43894=>"111100100",
  43895=>"100101100",
  43896=>"111010011",
  43897=>"111010010",
  43898=>"011001000",
  43899=>"000001001",
  43900=>"000001111",
  43901=>"111010001",
  43902=>"111010011",
  43903=>"011110110",
  43904=>"100101011",
  43905=>"011010011",
  43906=>"010000011",
  43907=>"010111101",
  43908=>"110000001",
  43909=>"100100010",
  43910=>"110111001",
  43911=>"101110011",
  43912=>"001111100",
  43913=>"010000001",
  43914=>"000100101",
  43915=>"001100001",
  43916=>"100000010",
  43917=>"001010011",
  43918=>"111011000",
  43919=>"011011111",
  43920=>"011000000",
  43921=>"011111100",
  43922=>"001100011",
  43923=>"100000010",
  43924=>"011011010",
  43925=>"100010111",
  43926=>"011101010",
  43927=>"010100000",
  43928=>"011000110",
  43929=>"001000101",
  43930=>"111100011",
  43931=>"101111110",
  43932=>"101100001",
  43933=>"000100010",
  43934=>"100010001",
  43935=>"111100101",
  43936=>"001101010",
  43937=>"000010010",
  43938=>"100110011",
  43939=>"000010010",
  43940=>"000010000",
  43941=>"110100000",
  43942=>"011100111",
  43943=>"010001011",
  43944=>"101010011",
  43945=>"111101001",
  43946=>"110110001",
  43947=>"110010111",
  43948=>"100010010",
  43949=>"100100010",
  43950=>"010110001",
  43951=>"011011011",
  43952=>"101011111",
  43953=>"111011101",
  43954=>"100000001",
  43955=>"101111101",
  43956=>"011010111",
  43957=>"110100011",
  43958=>"110110010",
  43959=>"010100001",
  43960=>"111100101",
  43961=>"010000111",
  43962=>"000000111",
  43963=>"101101010",
  43964=>"110010110",
  43965=>"100100010",
  43966=>"010001111",
  43967=>"001010110",
  43968=>"100001010",
  43969=>"110101001",
  43970=>"011101111",
  43971=>"011001001",
  43972=>"111011001",
  43973=>"110101000",
  43974=>"001101111",
  43975=>"010010011",
  43976=>"011010000",
  43977=>"011001000",
  43978=>"111100001",
  43979=>"001111100",
  43980=>"001101010",
  43981=>"000001100",
  43982=>"000011111",
  43983=>"001111100",
  43984=>"100110001",
  43985=>"011001101",
  43986=>"001110011",
  43987=>"100011011",
  43988=>"111011011",
  43989=>"010100111",
  43990=>"100101000",
  43991=>"110001111",
  43992=>"000001010",
  43993=>"000100010",
  43994=>"111111001",
  43995=>"111001101",
  43996=>"111111111",
  43997=>"011101000",
  43998=>"100100111",
  43999=>"010001101",
  44000=>"000000011",
  44001=>"100001100",
  44002=>"010111010",
  44003=>"100010101",
  44004=>"011000110",
  44005=>"100010011",
  44006=>"111010000",
  44007=>"111000100",
  44008=>"100011110",
  44009=>"100101000",
  44010=>"101010101",
  44011=>"000000000",
  44012=>"100000000",
  44013=>"110001101",
  44014=>"010010010",
  44015=>"111111110",
  44016=>"010111001",
  44017=>"000110011",
  44018=>"010000101",
  44019=>"100101100",
  44020=>"101101101",
  44021=>"000000001",
  44022=>"011111000",
  44023=>"110010111",
  44024=>"001010100",
  44025=>"000111010",
  44026=>"011000010",
  44027=>"111010111",
  44028=>"111010101",
  44029=>"110000101",
  44030=>"010001100",
  44031=>"100100011",
  44032=>"110000000",
  44033=>"001100101",
  44034=>"101000111",
  44035=>"100111100",
  44036=>"001011001",
  44037=>"100011000",
  44038=>"010000110",
  44039=>"110110000",
  44040=>"111100001",
  44041=>"010001000",
  44042=>"110101010",
  44043=>"100011011",
  44044=>"000001001",
  44045=>"111011011",
  44046=>"001111101",
  44047=>"000001001",
  44048=>"100001101",
  44049=>"000000101",
  44050=>"100100000",
  44051=>"100001100",
  44052=>"001111111",
  44053=>"011011000",
  44054=>"111111001",
  44055=>"100110011",
  44056=>"011101111",
  44057=>"011110010",
  44058=>"110111101",
  44059=>"001001001",
  44060=>"110001011",
  44061=>"010111110",
  44062=>"110110101",
  44063=>"101011000",
  44064=>"101011001",
  44065=>"100000100",
  44066=>"110100001",
  44067=>"010000001",
  44068=>"010011101",
  44069=>"011011001",
  44070=>"010000001",
  44071=>"110001100",
  44072=>"000100001",
  44073=>"000011011",
  44074=>"100100100",
  44075=>"111000110",
  44076=>"111010011",
  44077=>"011001100",
  44078=>"100011001",
  44079=>"111111110",
  44080=>"001011100",
  44081=>"010111111",
  44082=>"111000001",
  44083=>"111100100",
  44084=>"000000100",
  44085=>"110000111",
  44086=>"010001101",
  44087=>"110011000",
  44088=>"000111000",
  44089=>"001000000",
  44090=>"001100100",
  44091=>"100010010",
  44092=>"110100111",
  44093=>"011100000",
  44094=>"100100000",
  44095=>"001101101",
  44096=>"000100100",
  44097=>"010111110",
  44098=>"000000010",
  44099=>"101111000",
  44100=>"111101011",
  44101=>"011111001",
  44102=>"010101001",
  44103=>"001111111",
  44104=>"101001000",
  44105=>"101000111",
  44106=>"001101110",
  44107=>"001101100",
  44108=>"010100001",
  44109=>"010100011",
  44110=>"111000000",
  44111=>"101000001",
  44112=>"101101001",
  44113=>"011000111",
  44114=>"010111110",
  44115=>"000100111",
  44116=>"110001011",
  44117=>"011010010",
  44118=>"101010000",
  44119=>"100010101",
  44120=>"111010111",
  44121=>"001011000",
  44122=>"001101010",
  44123=>"000001101",
  44124=>"000001100",
  44125=>"000111111",
  44126=>"010011110",
  44127=>"110011110",
  44128=>"000100011",
  44129=>"011100011",
  44130=>"011111001",
  44131=>"011001101",
  44132=>"101101000",
  44133=>"011010101",
  44134=>"001001010",
  44135=>"000011101",
  44136=>"011011001",
  44137=>"101010011",
  44138=>"000110001",
  44139=>"011110000",
  44140=>"001101011",
  44141=>"110101000",
  44142=>"001110101",
  44143=>"000101011",
  44144=>"000100000",
  44145=>"011110010",
  44146=>"111011000",
  44147=>"011110010",
  44148=>"001100100",
  44149=>"010000000",
  44150=>"011110010",
  44151=>"011100100",
  44152=>"010100110",
  44153=>"000000011",
  44154=>"011011011",
  44155=>"001111000",
  44156=>"001001110",
  44157=>"110001011",
  44158=>"100111010",
  44159=>"111101100",
  44160=>"011101011",
  44161=>"101001101",
  44162=>"111010101",
  44163=>"101011001",
  44164=>"101000010",
  44165=>"001010110",
  44166=>"011001110",
  44167=>"010001001",
  44168=>"110100000",
  44169=>"101010110",
  44170=>"011000110",
  44171=>"000010010",
  44172=>"101100000",
  44173=>"011001110",
  44174=>"001011110",
  44175=>"000011001",
  44176=>"010100100",
  44177=>"011100010",
  44178=>"001100011",
  44179=>"111000010",
  44180=>"011110100",
  44181=>"000010001",
  44182=>"000001111",
  44183=>"111100100",
  44184=>"000000011",
  44185=>"110001110",
  44186=>"110000010",
  44187=>"111111001",
  44188=>"000000111",
  44189=>"000110000",
  44190=>"000111011",
  44191=>"111101000",
  44192=>"010000110",
  44193=>"110001010",
  44194=>"100011000",
  44195=>"111000011",
  44196=>"110100010",
  44197=>"010010000",
  44198=>"011011111",
  44199=>"001011110",
  44200=>"111101111",
  44201=>"000001110",
  44202=>"010000101",
  44203=>"110001100",
  44204=>"100010011",
  44205=>"010000010",
  44206=>"011111110",
  44207=>"111000011",
  44208=>"010110001",
  44209=>"010001010",
  44210=>"101100111",
  44211=>"110000100",
  44212=>"010110010",
  44213=>"010111011",
  44214=>"100000001",
  44215=>"111100011",
  44216=>"001101110",
  44217=>"011010001",
  44218=>"111001001",
  44219=>"101001000",
  44220=>"101001000",
  44221=>"011001100",
  44222=>"100101000",
  44223=>"011011111",
  44224=>"100011111",
  44225=>"011101011",
  44226=>"110111000",
  44227=>"100111110",
  44228=>"111100000",
  44229=>"010001001",
  44230=>"010100011",
  44231=>"111000001",
  44232=>"010010000",
  44233=>"011010011",
  44234=>"010010011",
  44235=>"010100001",
  44236=>"010111010",
  44237=>"000110011",
  44238=>"011001100",
  44239=>"011010000",
  44240=>"110010011",
  44241=>"001011100",
  44242=>"000101001",
  44243=>"100111010",
  44244=>"001000110",
  44245=>"100110010",
  44246=>"100110110",
  44247=>"111101100",
  44248=>"010001111",
  44249=>"111111001",
  44250=>"100010111",
  44251=>"111100000",
  44252=>"010110101",
  44253=>"010011101",
  44254=>"011010101",
  44255=>"100011001",
  44256=>"001001100",
  44257=>"110000001",
  44258=>"101010001",
  44259=>"000010101",
  44260=>"010001110",
  44261=>"010101110",
  44262=>"001010000",
  44263=>"110000000",
  44264=>"100101000",
  44265=>"101000000",
  44266=>"010110000",
  44267=>"001110000",
  44268=>"000001011",
  44269=>"010100010",
  44270=>"101001110",
  44271=>"011010000",
  44272=>"010110010",
  44273=>"100110011",
  44274=>"110001110",
  44275=>"001100000",
  44276=>"000010000",
  44277=>"110000000",
  44278=>"001101001",
  44279=>"101010110",
  44280=>"100101000",
  44281=>"010111011",
  44282=>"100100111",
  44283=>"001000000",
  44284=>"101101011",
  44285=>"000011001",
  44286=>"100111111",
  44287=>"101011000",
  44288=>"111100111",
  44289=>"000111010",
  44290=>"101110001",
  44291=>"000001011",
  44292=>"000110100",
  44293=>"001101101",
  44294=>"100011101",
  44295=>"101011110",
  44296=>"010110001",
  44297=>"001010010",
  44298=>"000111100",
  44299=>"010101011",
  44300=>"011111101",
  44301=>"000000100",
  44302=>"011001111",
  44303=>"000111111",
  44304=>"111000001",
  44305=>"010011001",
  44306=>"100010001",
  44307=>"100110100",
  44308=>"101110100",
  44309=>"101111010",
  44310=>"011011100",
  44311=>"101000111",
  44312=>"111101100",
  44313=>"100110111",
  44314=>"010111011",
  44315=>"111000011",
  44316=>"101110111",
  44317=>"001000110",
  44318=>"101011011",
  44319=>"011010110",
  44320=>"101110001",
  44321=>"000010001",
  44322=>"101111111",
  44323=>"110010101",
  44324=>"011100001",
  44325=>"110110011",
  44326=>"001010001",
  44327=>"001001001",
  44328=>"000010001",
  44329=>"010010110",
  44330=>"000000011",
  44331=>"111101001",
  44332=>"010101011",
  44333=>"101001100",
  44334=>"000100100",
  44335=>"001000000",
  44336=>"000101100",
  44337=>"010100111",
  44338=>"101011101",
  44339=>"000110110",
  44340=>"001010111",
  44341=>"000101011",
  44342=>"001110101",
  44343=>"010101000",
  44344=>"100001100",
  44345=>"101010011",
  44346=>"011010100",
  44347=>"111010001",
  44348=>"011000111",
  44349=>"100101010",
  44350=>"011001000",
  44351=>"010110101",
  44352=>"111111110",
  44353=>"101010001",
  44354=>"110011111",
  44355=>"011111101",
  44356=>"001011111",
  44357=>"011110100",
  44358=>"100101110",
  44359=>"000000010",
  44360=>"010011011",
  44361=>"100000010",
  44362=>"010101110",
  44363=>"001000000",
  44364=>"110001001",
  44365=>"111010000",
  44366=>"001010000",
  44367=>"110001010",
  44368=>"011110110",
  44369=>"001000011",
  44370=>"101100111",
  44371=>"110110011",
  44372=>"000100011",
  44373=>"101111111",
  44374=>"000110110",
  44375=>"100101000",
  44376=>"110100100",
  44377=>"000011000",
  44378=>"110111000",
  44379=>"100011000",
  44380=>"111001011",
  44381=>"000111000",
  44382=>"110101011",
  44383=>"001011010",
  44384=>"000110001",
  44385=>"101000101",
  44386=>"100010000",
  44387=>"000101000",
  44388=>"001101001",
  44389=>"001100110",
  44390=>"010111110",
  44391=>"110110000",
  44392=>"001000010",
  44393=>"011110011",
  44394=>"100110011",
  44395=>"100010010",
  44396=>"001010100",
  44397=>"011100101",
  44398=>"000011000",
  44399=>"000100001",
  44400=>"000101001",
  44401=>"111000101",
  44402=>"110110001",
  44403=>"011011010",
  44404=>"110101011",
  44405=>"011000000",
  44406=>"101001001",
  44407=>"010011011",
  44408=>"101010010",
  44409=>"001110001",
  44410=>"000101101",
  44411=>"000001000",
  44412=>"011101011",
  44413=>"101001011",
  44414=>"010101111",
  44415=>"101000101",
  44416=>"010010111",
  44417=>"000100110",
  44418=>"010110101",
  44419=>"011100000",
  44420=>"110000111",
  44421=>"011100011",
  44422=>"110101001",
  44423=>"111001000",
  44424=>"110001111",
  44425=>"001011001",
  44426=>"100110010",
  44427=>"001011011",
  44428=>"011001101",
  44429=>"110100101",
  44430=>"011001000",
  44431=>"110110010",
  44432=>"011100111",
  44433=>"101100101",
  44434=>"000100011",
  44435=>"101101100",
  44436=>"110111111",
  44437=>"001010010",
  44438=>"001010011",
  44439=>"001101111",
  44440=>"101011011",
  44441=>"000100110",
  44442=>"101011000",
  44443=>"111000111",
  44444=>"000010001",
  44445=>"111111000",
  44446=>"000010001",
  44447=>"110000100",
  44448=>"110000001",
  44449=>"010100010",
  44450=>"000010001",
  44451=>"001101010",
  44452=>"111010011",
  44453=>"010000100",
  44454=>"000000001",
  44455=>"000001111",
  44456=>"000111100",
  44457=>"010111001",
  44458=>"011100101",
  44459=>"000001010",
  44460=>"010001010",
  44461=>"011010010",
  44462=>"000111101",
  44463=>"111111001",
  44464=>"011100100",
  44465=>"001100110",
  44466=>"111001001",
  44467=>"110101111",
  44468=>"100110101",
  44469=>"101000011",
  44470=>"000001011",
  44471=>"001000000",
  44472=>"111011101",
  44473=>"110101101",
  44474=>"000010110",
  44475=>"101010010",
  44476=>"000111000",
  44477=>"110110001",
  44478=>"111011111",
  44479=>"110011000",
  44480=>"111000110",
  44481=>"100101000",
  44482=>"010010100",
  44483=>"010010100",
  44484=>"110101001",
  44485=>"100010111",
  44486=>"101100010",
  44487=>"000000001",
  44488=>"101100001",
  44489=>"011011010",
  44490=>"111100011",
  44491=>"011010110",
  44492=>"000001100",
  44493=>"111101101",
  44494=>"000110110",
  44495=>"110100101",
  44496=>"110111110",
  44497=>"000101001",
  44498=>"011101001",
  44499=>"111001100",
  44500=>"110111110",
  44501=>"010001100",
  44502=>"000000111",
  44503=>"101010011",
  44504=>"101110010",
  44505=>"100111011",
  44506=>"110010110",
  44507=>"100110011",
  44508=>"011010110",
  44509=>"001011100",
  44510=>"011010010",
  44511=>"111101011",
  44512=>"100101011",
  44513=>"001101000",
  44514=>"010000010",
  44515=>"110011001",
  44516=>"010110000",
  44517=>"011101011",
  44518=>"001101101",
  44519=>"001000000",
  44520=>"111001111",
  44521=>"110111011",
  44522=>"000110101",
  44523=>"111001001",
  44524=>"100010100",
  44525=>"001100000",
  44526=>"010010000",
  44527=>"100010101",
  44528=>"011010011",
  44529=>"100111001",
  44530=>"000100110",
  44531=>"000100111",
  44532=>"111101111",
  44533=>"101100110",
  44534=>"011001000",
  44535=>"101101011",
  44536=>"000101110",
  44537=>"101101001",
  44538=>"010100101",
  44539=>"000101001",
  44540=>"010010101",
  44541=>"011001010",
  44542=>"110111110",
  44543=>"100001101",
  44544=>"101101001",
  44545=>"011110001",
  44546=>"101111000",
  44547=>"010110011",
  44548=>"101101001",
  44549=>"110000001",
  44550=>"011000011",
  44551=>"101001100",
  44552=>"101110100",
  44553=>"001100010",
  44554=>"110001110",
  44555=>"100100010",
  44556=>"100011100",
  44557=>"111000101",
  44558=>"010001001",
  44559=>"010001111",
  44560=>"111101011",
  44561=>"101101010",
  44562=>"101111010",
  44563=>"101110011",
  44564=>"110010001",
  44565=>"111001110",
  44566=>"110111101",
  44567=>"011101110",
  44568=>"011110011",
  44569=>"010111101",
  44570=>"001000000",
  44571=>"010100111",
  44572=>"010110001",
  44573=>"010100111",
  44574=>"111101111",
  44575=>"100010010",
  44576=>"111011111",
  44577=>"000100000",
  44578=>"000011101",
  44579=>"000000010",
  44580=>"111111001",
  44581=>"010110010",
  44582=>"011110000",
  44583=>"001000000",
  44584=>"001000000",
  44585=>"000101010",
  44586=>"101001110",
  44587=>"110010110",
  44588=>"010011011",
  44589=>"000110111",
  44590=>"110110000",
  44591=>"000101010",
  44592=>"100000110",
  44593=>"010101001",
  44594=>"100010101",
  44595=>"000010010",
  44596=>"111111101",
  44597=>"110111110",
  44598=>"100001010",
  44599=>"110101101",
  44600=>"111011100",
  44601=>"010001111",
  44602=>"010110001",
  44603=>"100011001",
  44604=>"000110101",
  44605=>"010100001",
  44606=>"100100110",
  44607=>"100001110",
  44608=>"010100100",
  44609=>"111101100",
  44610=>"011001110",
  44611=>"001111100",
  44612=>"000001010",
  44613=>"000000010",
  44614=>"011000001",
  44615=>"000000110",
  44616=>"110001100",
  44617=>"111101110",
  44618=>"010010001",
  44619=>"100000000",
  44620=>"110100110",
  44621=>"010101101",
  44622=>"110111000",
  44623=>"000000100",
  44624=>"110011101",
  44625=>"100110101",
  44626=>"011110010",
  44627=>"001101110",
  44628=>"100010101",
  44629=>"110111100",
  44630=>"110010111",
  44631=>"000111101",
  44632=>"000000010",
  44633=>"101000000",
  44634=>"101110010",
  44635=>"100000011",
  44636=>"101000110",
  44637=>"010110101",
  44638=>"101100100",
  44639=>"111010011",
  44640=>"001111000",
  44641=>"010010110",
  44642=>"101111100",
  44643=>"000111000",
  44644=>"000000101",
  44645=>"101001101",
  44646=>"100101011",
  44647=>"100010011",
  44648=>"100000000",
  44649=>"000111001",
  44650=>"011010011",
  44651=>"001000011",
  44652=>"000001101",
  44653=>"000011010",
  44654=>"110101100",
  44655=>"110000110",
  44656=>"000111000",
  44657=>"000000010",
  44658=>"101011000",
  44659=>"011100101",
  44660=>"000011011",
  44661=>"100001001",
  44662=>"101000110",
  44663=>"010010000",
  44664=>"100110001",
  44665=>"111000111",
  44666=>"011110111",
  44667=>"011110100",
  44668=>"000110101",
  44669=>"100000100",
  44670=>"111000010",
  44671=>"110000100",
  44672=>"111011000",
  44673=>"110010100",
  44674=>"010010010",
  44675=>"111000110",
  44676=>"000001100",
  44677=>"101000000",
  44678=>"011110100",
  44679=>"110001000",
  44680=>"001100100",
  44681=>"011011100",
  44682=>"011011111",
  44683=>"100010000",
  44684=>"000000000",
  44685=>"001110011",
  44686=>"111101001",
  44687=>"100111101",
  44688=>"101100101",
  44689=>"110011001",
  44690=>"010110101",
  44691=>"001110111",
  44692=>"101101110",
  44693=>"111111110",
  44694=>"101101101",
  44695=>"110011100",
  44696=>"001110000",
  44697=>"011111011",
  44698=>"001110000",
  44699=>"011001001",
  44700=>"011001010",
  44701=>"011100011",
  44702=>"100100010",
  44703=>"011101100",
  44704=>"101001011",
  44705=>"010011001",
  44706=>"000110111",
  44707=>"111100001",
  44708=>"000110011",
  44709=>"010101011",
  44710=>"000010011",
  44711=>"001000001",
  44712=>"100100111",
  44713=>"110111000",
  44714=>"010100101",
  44715=>"111101001",
  44716=>"001010000",
  44717=>"100001011",
  44718=>"111000001",
  44719=>"110010001",
  44720=>"100001011",
  44721=>"001110110",
  44722=>"111011001",
  44723=>"010001000",
  44724=>"011011111",
  44725=>"010001101",
  44726=>"110101000",
  44727=>"011000100",
  44728=>"100101111",
  44729=>"100111000",
  44730=>"011011101",
  44731=>"010010001",
  44732=>"010010010",
  44733=>"011011110",
  44734=>"010000010",
  44735=>"000010010",
  44736=>"111100001",
  44737=>"101001111",
  44738=>"010100001",
  44739=>"101110010",
  44740=>"101101010",
  44741=>"111001110",
  44742=>"101011100",
  44743=>"011111110",
  44744=>"101101111",
  44745=>"011001001",
  44746=>"001111001",
  44747=>"111101110",
  44748=>"001011101",
  44749=>"111011000",
  44750=>"111100111",
  44751=>"000111001",
  44752=>"000011101",
  44753=>"100011110",
  44754=>"011100111",
  44755=>"100010110",
  44756=>"110011111",
  44757=>"000010011",
  44758=>"011100011",
  44759=>"001100000",
  44760=>"001110010",
  44761=>"011000110",
  44762=>"110000001",
  44763=>"110100001",
  44764=>"100111011",
  44765=>"101110001",
  44766=>"101010011",
  44767=>"011000101",
  44768=>"111100100",
  44769=>"100011011",
  44770=>"000010111",
  44771=>"011001111",
  44772=>"100100000",
  44773=>"011000001",
  44774=>"001001001",
  44775=>"100101100",
  44776=>"101111110",
  44777=>"100100011",
  44778=>"111101011",
  44779=>"011000001",
  44780=>"010010111",
  44781=>"010110011",
  44782=>"101001110",
  44783=>"110010100",
  44784=>"011011100",
  44785=>"010100001",
  44786=>"111111001",
  44787=>"101111010",
  44788=>"100000000",
  44789=>"101001000",
  44790=>"111111000",
  44791=>"010001100",
  44792=>"011111011",
  44793=>"111110101",
  44794=>"110011000",
  44795=>"000100001",
  44796=>"011101100",
  44797=>"000100000",
  44798=>"110100011",
  44799=>"101100000",
  44800=>"101101101",
  44801=>"100001000",
  44802=>"111100010",
  44803=>"001011010",
  44804=>"100101001",
  44805=>"100001010",
  44806=>"000100010",
  44807=>"100101111",
  44808=>"011010111",
  44809=>"010100011",
  44810=>"001111111",
  44811=>"001101011",
  44812=>"101010101",
  44813=>"011011011",
  44814=>"011000101",
  44815=>"110011110",
  44816=>"001010100",
  44817=>"001101110",
  44818=>"110001100",
  44819=>"001010010",
  44820=>"000000001",
  44821=>"000011001",
  44822=>"010010000",
  44823=>"101101010",
  44824=>"010001100",
  44825=>"000000010",
  44826=>"100011100",
  44827=>"111011101",
  44828=>"011110011",
  44829=>"001101100",
  44830=>"101010010",
  44831=>"110110000",
  44832=>"110000000",
  44833=>"111000111",
  44834=>"001000001",
  44835=>"100111101",
  44836=>"000100000",
  44837=>"101100011",
  44838=>"111100010",
  44839=>"111110001",
  44840=>"000110011",
  44841=>"100010001",
  44842=>"111010111",
  44843=>"100110110",
  44844=>"101111011",
  44845=>"100000001",
  44846=>"011011000",
  44847=>"110010110",
  44848=>"010010111",
  44849=>"111101011",
  44850=>"000100100",
  44851=>"001111111",
  44852=>"011111110",
  44853=>"101000101",
  44854=>"001101000",
  44855=>"000010111",
  44856=>"000110001",
  44857=>"101001000",
  44858=>"010111011",
  44859=>"001101000",
  44860=>"101000001",
  44861=>"010000100",
  44862=>"100000000",
  44863=>"100101010",
  44864=>"000010101",
  44865=>"111001110",
  44866=>"010111100",
  44867=>"100110111",
  44868=>"001001100",
  44869=>"110101111",
  44870=>"111100101",
  44871=>"010011011",
  44872=>"100110110",
  44873=>"110001000",
  44874=>"100001111",
  44875=>"010001001",
  44876=>"110011000",
  44877=>"110100001",
  44878=>"010101000",
  44879=>"110000110",
  44880=>"010110110",
  44881=>"010110010",
  44882=>"100110001",
  44883=>"000010101",
  44884=>"100010010",
  44885=>"111111111",
  44886=>"010101011",
  44887=>"011010110",
  44888=>"101001100",
  44889=>"100100101",
  44890=>"111111110",
  44891=>"100000100",
  44892=>"100001111",
  44893=>"111000000",
  44894=>"111110011",
  44895=>"000100111",
  44896=>"000111100",
  44897=>"000011010",
  44898=>"111000011",
  44899=>"110010111",
  44900=>"010000111",
  44901=>"001001011",
  44902=>"101000011",
  44903=>"101101111",
  44904=>"001000111",
  44905=>"000011001",
  44906=>"100010111",
  44907=>"111101000",
  44908=>"100001111",
  44909=>"011110000",
  44910=>"101011101",
  44911=>"110010011",
  44912=>"101001000",
  44913=>"010000010",
  44914=>"011110011",
  44915=>"001001100",
  44916=>"011100010",
  44917=>"000101000",
  44918=>"000000000",
  44919=>"001111000",
  44920=>"100110011",
  44921=>"011110111",
  44922=>"000011000",
  44923=>"111011011",
  44924=>"001001010",
  44925=>"010101000",
  44926=>"101110000",
  44927=>"000010101",
  44928=>"000000101",
  44929=>"101011111",
  44930=>"001010000",
  44931=>"110000011",
  44932=>"110000010",
  44933=>"100100110",
  44934=>"001000011",
  44935=>"100100110",
  44936=>"010111110",
  44937=>"011110001",
  44938=>"110111101",
  44939=>"101101111",
  44940=>"111001011",
  44941=>"001010001",
  44942=>"100100010",
  44943=>"001111111",
  44944=>"001001101",
  44945=>"011110000",
  44946=>"001000111",
  44947=>"111001011",
  44948=>"101001000",
  44949=>"001111011",
  44950=>"110101010",
  44951=>"111111110",
  44952=>"001001010",
  44953=>"100000111",
  44954=>"001111100",
  44955=>"110100011",
  44956=>"011010000",
  44957=>"110111010",
  44958=>"110010010",
  44959=>"101111010",
  44960=>"000000011",
  44961=>"011011011",
  44962=>"000110001",
  44963=>"101011111",
  44964=>"000000100",
  44965=>"110100111",
  44966=>"101110001",
  44967=>"011011110",
  44968=>"011111111",
  44969=>"111001001",
  44970=>"011000110",
  44971=>"111111000",
  44972=>"100011000",
  44973=>"111111011",
  44974=>"010101000",
  44975=>"011001111",
  44976=>"000111001",
  44977=>"111101110",
  44978=>"000111010",
  44979=>"010000000",
  44980=>"010110010",
  44981=>"111110011",
  44982=>"101100111",
  44983=>"011000001",
  44984=>"101101110",
  44985=>"000110011",
  44986=>"100000010",
  44987=>"101001101",
  44988=>"111001101",
  44989=>"110001111",
  44990=>"100001110",
  44991=>"101000001",
  44992=>"111000011",
  44993=>"011101010",
  44994=>"111000110",
  44995=>"111011100",
  44996=>"010111010",
  44997=>"011000011",
  44998=>"001110010",
  44999=>"010101110",
  45000=>"010001000",
  45001=>"111000010",
  45002=>"000101110",
  45003=>"001111001",
  45004=>"000001010",
  45005=>"100000010",
  45006=>"000000000",
  45007=>"010011100",
  45008=>"101100100",
  45009=>"101010000",
  45010=>"101110011",
  45011=>"001000101",
  45012=>"010111110",
  45013=>"101010011",
  45014=>"001001010",
  45015=>"111110111",
  45016=>"000111101",
  45017=>"100000111",
  45018=>"100010000",
  45019=>"111100000",
  45020=>"010100011",
  45021=>"111001101",
  45022=>"000001010",
  45023=>"100110110",
  45024=>"100101010",
  45025=>"011111101",
  45026=>"111001101",
  45027=>"110010101",
  45028=>"010010010",
  45029=>"010010011",
  45030=>"001111110",
  45031=>"101110000",
  45032=>"000010001",
  45033=>"011000111",
  45034=>"101101111",
  45035=>"001110011",
  45036=>"000010010",
  45037=>"111100000",
  45038=>"010101110",
  45039=>"110100011",
  45040=>"010111101",
  45041=>"011111000",
  45042=>"101011011",
  45043=>"010101010",
  45044=>"111110001",
  45045=>"000000000",
  45046=>"011000000",
  45047=>"000111000",
  45048=>"011010100",
  45049=>"111011111",
  45050=>"101011001",
  45051=>"111010100",
  45052=>"011010111",
  45053=>"001001011",
  45054=>"111000010",
  45055=>"100010111",
  45056=>"010000110",
  45057=>"111011000",
  45058=>"111000110",
  45059=>"010010111",
  45060=>"110010011",
  45061=>"100011000",
  45062=>"011010110",
  45063=>"111001010",
  45064=>"110010010",
  45065=>"000000000",
  45066=>"010001010",
  45067=>"101011111",
  45068=>"000000111",
  45069=>"111001000",
  45070=>"100100011",
  45071=>"011111111",
  45072=>"000001011",
  45073=>"110011001",
  45074=>"001000011",
  45075=>"011000001",
  45076=>"001000100",
  45077=>"101001110",
  45078=>"110101000",
  45079=>"010001000",
  45080=>"001010010",
  45081=>"110010000",
  45082=>"000011110",
  45083=>"000110000",
  45084=>"110010111",
  45085=>"110001000",
  45086=>"010010111",
  45087=>"000101010",
  45088=>"010001000",
  45089=>"000100000",
  45090=>"001010110",
  45091=>"010011110",
  45092=>"100101011",
  45093=>"011011101",
  45094=>"000110101",
  45095=>"111111100",
  45096=>"101101011",
  45097=>"111110101",
  45098=>"100110101",
  45099=>"111100011",
  45100=>"011011000",
  45101=>"000000000",
  45102=>"111011000",
  45103=>"111111111",
  45104=>"010101111",
  45105=>"010011111",
  45106=>"001110100",
  45107=>"111101110",
  45108=>"000010011",
  45109=>"101111011",
  45110=>"001011101",
  45111=>"111100011",
  45112=>"010011101",
  45113=>"000000010",
  45114=>"000000111",
  45115=>"111101000",
  45116=>"101101001",
  45117=>"101100000",
  45118=>"001101111",
  45119=>"000101111",
  45120=>"011000011",
  45121=>"000000011",
  45122=>"111111001",
  45123=>"101101110",
  45124=>"111111110",
  45125=>"001000110",
  45126=>"111110100",
  45127=>"011100011",
  45128=>"011001001",
  45129=>"001101110",
  45130=>"100011101",
  45131=>"000110110",
  45132=>"110101001",
  45133=>"010011101",
  45134=>"011000001",
  45135=>"011111101",
  45136=>"010011101",
  45137=>"011011111",
  45138=>"000111111",
  45139=>"001011000",
  45140=>"011100100",
  45141=>"001001001",
  45142=>"010101101",
  45143=>"000111010",
  45144=>"111011101",
  45145=>"000011111",
  45146=>"101000000",
  45147=>"000001111",
  45148=>"001010111",
  45149=>"000111100",
  45150=>"000001110",
  45151=>"000010000",
  45152=>"000001001",
  45153=>"001000001",
  45154=>"001010101",
  45155=>"001000010",
  45156=>"001101001",
  45157=>"110110000",
  45158=>"100001000",
  45159=>"110010101",
  45160=>"011010000",
  45161=>"110100010",
  45162=>"000111111",
  45163=>"110001000",
  45164=>"101110111",
  45165=>"000100100",
  45166=>"110010010",
  45167=>"000110000",
  45168=>"110001100",
  45169=>"001111100",
  45170=>"101010011",
  45171=>"001101001",
  45172=>"000000000",
  45173=>"100100100",
  45174=>"101011111",
  45175=>"111111101",
  45176=>"001001111",
  45177=>"010000111",
  45178=>"100100011",
  45179=>"010111001",
  45180=>"001000001",
  45181=>"110001100",
  45182=>"001110000",
  45183=>"000110111",
  45184=>"000101111",
  45185=>"101100100",
  45186=>"011010110",
  45187=>"010010101",
  45188=>"001101110",
  45189=>"111111011",
  45190=>"010001011",
  45191=>"110010101",
  45192=>"101010011",
  45193=>"101010111",
  45194=>"101011000",
  45195=>"001110001",
  45196=>"101101011",
  45197=>"110100110",
  45198=>"000100110",
  45199=>"101101010",
  45200=>"010110101",
  45201=>"001001110",
  45202=>"000000110",
  45203=>"010101010",
  45204=>"111101011",
  45205=>"000001010",
  45206=>"111001001",
  45207=>"011100001",
  45208=>"000011110",
  45209=>"111001110",
  45210=>"110111010",
  45211=>"011110111",
  45212=>"010010111",
  45213=>"000100111",
  45214=>"111011100",
  45215=>"100011100",
  45216=>"100111101",
  45217=>"111000011",
  45218=>"100100111",
  45219=>"001100101",
  45220=>"101011010",
  45221=>"101100110",
  45222=>"110101010",
  45223=>"110000000",
  45224=>"101100110",
  45225=>"000101111",
  45226=>"011101111",
  45227=>"110010110",
  45228=>"100000111",
  45229=>"011111000",
  45230=>"101110100",
  45231=>"011110101",
  45232=>"001100000",
  45233=>"011001110",
  45234=>"011111010",
  45235=>"000101000",
  45236=>"110101001",
  45237=>"101011000",
  45238=>"111100011",
  45239=>"001111011",
  45240=>"110101101",
  45241=>"001111111",
  45242=>"111001001",
  45243=>"111111001",
  45244=>"100010000",
  45245=>"101011100",
  45246=>"100100001",
  45247=>"001011000",
  45248=>"100001001",
  45249=>"100000111",
  45250=>"111001001",
  45251=>"110010110",
  45252=>"100001001",
  45253=>"010010010",
  45254=>"011011000",
  45255=>"000000000",
  45256=>"111100111",
  45257=>"100000111",
  45258=>"011101111",
  45259=>"000100011",
  45260=>"110111010",
  45261=>"111011000",
  45262=>"111100010",
  45263=>"000101001",
  45264=>"001100110",
  45265=>"111110110",
  45266=>"010011100",
  45267=>"111000110",
  45268=>"101001101",
  45269=>"110011001",
  45270=>"000110000",
  45271=>"111111111",
  45272=>"101001011",
  45273=>"000000100",
  45274=>"100010110",
  45275=>"000001000",
  45276=>"010100001",
  45277=>"010011100",
  45278=>"011000010",
  45279=>"000101101",
  45280=>"000010011",
  45281=>"000110000",
  45282=>"010111101",
  45283=>"100000001",
  45284=>"100011110",
  45285=>"110111001",
  45286=>"100111101",
  45287=>"010111001",
  45288=>"110111000",
  45289=>"001000110",
  45290=>"100100100",
  45291=>"110000001",
  45292=>"000000010",
  45293=>"010011110",
  45294=>"011000001",
  45295=>"111000001",
  45296=>"110000000",
  45297=>"101111011",
  45298=>"000010000",
  45299=>"011001011",
  45300=>"111110101",
  45301=>"000011010",
  45302=>"101101100",
  45303=>"011100100",
  45304=>"100000110",
  45305=>"000110111",
  45306=>"100010101",
  45307=>"011011001",
  45308=>"110000010",
  45309=>"010111010",
  45310=>"000100101",
  45311=>"101111000",
  45312=>"101101000",
  45313=>"110110101",
  45314=>"010101101",
  45315=>"101101110",
  45316=>"111100001",
  45317=>"001000111",
  45318=>"001111011",
  45319=>"000010111",
  45320=>"010100010",
  45321=>"001110110",
  45322=>"001100110",
  45323=>"000001100",
  45324=>"110111110",
  45325=>"000110100",
  45326=>"101011010",
  45327=>"000001011",
  45328=>"001100111",
  45329=>"101100001",
  45330=>"001000110",
  45331=>"100111001",
  45332=>"000100100",
  45333=>"001111100",
  45334=>"110001100",
  45335=>"000011111",
  45336=>"110011110",
  45337=>"101001000",
  45338=>"110100101",
  45339=>"100101111",
  45340=>"000100101",
  45341=>"011111000",
  45342=>"011000010",
  45343=>"001110010",
  45344=>"101011100",
  45345=>"110101101",
  45346=>"101111101",
  45347=>"100111001",
  45348=>"110011011",
  45349=>"100111010",
  45350=>"111101011",
  45351=>"011111101",
  45352=>"101001001",
  45353=>"001010101",
  45354=>"100100011",
  45355=>"010001010",
  45356=>"000100001",
  45357=>"001010100",
  45358=>"000101100",
  45359=>"001010101",
  45360=>"000010010",
  45361=>"000100100",
  45362=>"110101010",
  45363=>"111011000",
  45364=>"110101110",
  45365=>"010001000",
  45366=>"100101001",
  45367=>"011001001",
  45368=>"101100101",
  45369=>"101100011",
  45370=>"101000000",
  45371=>"010110101",
  45372=>"110111001",
  45373=>"111000111",
  45374=>"101101110",
  45375=>"110001110",
  45376=>"101010111",
  45377=>"000100010",
  45378=>"011010010",
  45379=>"010010000",
  45380=>"101001110",
  45381=>"100011011",
  45382=>"001001101",
  45383=>"110100100",
  45384=>"010011100",
  45385=>"000100010",
  45386=>"101101101",
  45387=>"110000011",
  45388=>"100010001",
  45389=>"100101000",
  45390=>"010000111",
  45391=>"111111111",
  45392=>"000011101",
  45393=>"111101101",
  45394=>"011101000",
  45395=>"010100100",
  45396=>"010100100",
  45397=>"001001110",
  45398=>"010100110",
  45399=>"011101000",
  45400=>"010110100",
  45401=>"110100110",
  45402=>"110100110",
  45403=>"010000000",
  45404=>"100010000",
  45405=>"010000110",
  45406=>"111101001",
  45407=>"001101011",
  45408=>"110110001",
  45409=>"000010010",
  45410=>"101010001",
  45411=>"010111011",
  45412=>"010010010",
  45413=>"101110101",
  45414=>"110011111",
  45415=>"011011011",
  45416=>"101101101",
  45417=>"110110110",
  45418=>"111111010",
  45419=>"000111011",
  45420=>"100000101",
  45421=>"110001111",
  45422=>"010010101",
  45423=>"000001100",
  45424=>"110010111",
  45425=>"000101111",
  45426=>"101111111",
  45427=>"101010100",
  45428=>"011100110",
  45429=>"001100111",
  45430=>"110111111",
  45431=>"001001001",
  45432=>"000011001",
  45433=>"011111000",
  45434=>"100101111",
  45435=>"010111100",
  45436=>"101100000",
  45437=>"011110101",
  45438=>"110011111",
  45439=>"001001010",
  45440=>"111110001",
  45441=>"101000011",
  45442=>"001110001",
  45443=>"011100111",
  45444=>"100000001",
  45445=>"101001011",
  45446=>"100111011",
  45447=>"111010000",
  45448=>"111001111",
  45449=>"111000011",
  45450=>"000010011",
  45451=>"000111001",
  45452=>"110100110",
  45453=>"100111110",
  45454=>"110101111",
  45455=>"000000111",
  45456=>"011111000",
  45457=>"101000011",
  45458=>"001011001",
  45459=>"001000110",
  45460=>"111110110",
  45461=>"001000110",
  45462=>"000001011",
  45463=>"111110110",
  45464=>"100100111",
  45465=>"001111000",
  45466=>"000110001",
  45467=>"100011000",
  45468=>"101101011",
  45469=>"101011000",
  45470=>"111110011",
  45471=>"011101010",
  45472=>"010110101",
  45473=>"010101111",
  45474=>"110011000",
  45475=>"011111000",
  45476=>"010101100",
  45477=>"111011000",
  45478=>"100111100",
  45479=>"011111111",
  45480=>"110101101",
  45481=>"101100011",
  45482=>"110010100",
  45483=>"101100101",
  45484=>"011000100",
  45485=>"000111000",
  45486=>"000110100",
  45487=>"100001110",
  45488=>"110000000",
  45489=>"110000100",
  45490=>"111101001",
  45491=>"000000001",
  45492=>"100001000",
  45493=>"010010010",
  45494=>"111110000",
  45495=>"010101101",
  45496=>"111101000",
  45497=>"100011001",
  45498=>"000011010",
  45499=>"011101001",
  45500=>"011000001",
  45501=>"100111111",
  45502=>"100101110",
  45503=>"001100110",
  45504=>"001010101",
  45505=>"010000100",
  45506=>"010010111",
  45507=>"100011110",
  45508=>"000000011",
  45509=>"101010101",
  45510=>"100001101",
  45511=>"001101001",
  45512=>"111010110",
  45513=>"001001110",
  45514=>"011000011",
  45515=>"001110100",
  45516=>"000001101",
  45517=>"101101101",
  45518=>"111010011",
  45519=>"110110111",
  45520=>"110110011",
  45521=>"100100010",
  45522=>"010001100",
  45523=>"000110000",
  45524=>"111110001",
  45525=>"010101010",
  45526=>"101101101",
  45527=>"011011000",
  45528=>"101000011",
  45529=>"010010100",
  45530=>"101010011",
  45531=>"101010110",
  45532=>"100100010",
  45533=>"011101000",
  45534=>"110001111",
  45535=>"000111011",
  45536=>"010100000",
  45537=>"011001100",
  45538=>"111010010",
  45539=>"011001110",
  45540=>"101000010",
  45541=>"111100100",
  45542=>"111110100",
  45543=>"110100011",
  45544=>"000100110",
  45545=>"001000000",
  45546=>"100110001",
  45547=>"011001101",
  45548=>"001100110",
  45549=>"010001111",
  45550=>"011100000",
  45551=>"101011000",
  45552=>"111111001",
  45553=>"101101100",
  45554=>"111100011",
  45555=>"110010111",
  45556=>"010001000",
  45557=>"110010100",
  45558=>"010110011",
  45559=>"010000000",
  45560=>"001001101",
  45561=>"110000111",
  45562=>"100000110",
  45563=>"101001010",
  45564=>"010110000",
  45565=>"010000101",
  45566=>"010010001",
  45567=>"101100000",
  45568=>"000000000",
  45569=>"101001110",
  45570=>"011110111",
  45571=>"010011101",
  45572=>"110000110",
  45573=>"000001100",
  45574=>"100111111",
  45575=>"111000011",
  45576=>"111000000",
  45577=>"011111001",
  45578=>"010110110",
  45579=>"001001101",
  45580=>"111101000",
  45581=>"011110001",
  45582=>"011100111",
  45583=>"001101110",
  45584=>"011100011",
  45585=>"111001011",
  45586=>"000101111",
  45587=>"011010100",
  45588=>"101011001",
  45589=>"000000001",
  45590=>"001100001",
  45591=>"100111111",
  45592=>"111101100",
  45593=>"011010111",
  45594=>"100110010",
  45595=>"101001111",
  45596=>"110000101",
  45597=>"011011010",
  45598=>"011010010",
  45599=>"111111111",
  45600=>"111111010",
  45601=>"010001000",
  45602=>"000000011",
  45603=>"111010001",
  45604=>"101000011",
  45605=>"101000101",
  45606=>"110000111",
  45607=>"110110011",
  45608=>"110110111",
  45609=>"011100011",
  45610=>"000100011",
  45611=>"000011101",
  45612=>"101100001",
  45613=>"101110111",
  45614=>"111100001",
  45615=>"010101001",
  45616=>"010010111",
  45617=>"110111001",
  45618=>"100001000",
  45619=>"011110110",
  45620=>"101100110",
  45621=>"000010011",
  45622=>"010101011",
  45623=>"111100000",
  45624=>"110100010",
  45625=>"011001011",
  45626=>"011000101",
  45627=>"101000011",
  45628=>"101001011",
  45629=>"010000001",
  45630=>"111010000",
  45631=>"100100000",
  45632=>"001101011",
  45633=>"000011101",
  45634=>"111000000",
  45635=>"111111110",
  45636=>"111100100",
  45637=>"010110001",
  45638=>"000010110",
  45639=>"111101111",
  45640=>"101011101",
  45641=>"101100010",
  45642=>"111101101",
  45643=>"001000000",
  45644=>"010110101",
  45645=>"011000011",
  45646=>"111110000",
  45647=>"010010001",
  45648=>"000011111",
  45649=>"111101111",
  45650=>"000110111",
  45651=>"110111110",
  45652=>"001000110",
  45653=>"001011000",
  45654=>"111111101",
  45655=>"111101100",
  45656=>"101001101",
  45657=>"110001000",
  45658=>"100011100",
  45659=>"010111000",
  45660=>"001110011",
  45661=>"100000010",
  45662=>"000010000",
  45663=>"000100100",
  45664=>"011111011",
  45665=>"110111000",
  45666=>"110101110",
  45667=>"011010001",
  45668=>"000100111",
  45669=>"000111001",
  45670=>"101010111",
  45671=>"110111111",
  45672=>"000111001",
  45673=>"000100000",
  45674=>"001001111",
  45675=>"010011111",
  45676=>"110111100",
  45677=>"111001010",
  45678=>"101000010",
  45679=>"010110111",
  45680=>"001110000",
  45681=>"000000010",
  45682=>"101011100",
  45683=>"101110101",
  45684=>"001010100",
  45685=>"001000001",
  45686=>"100010011",
  45687=>"000001110",
  45688=>"001001011",
  45689=>"100000000",
  45690=>"111101100",
  45691=>"001100011",
  45692=>"011000011",
  45693=>"000000010",
  45694=>"000001001",
  45695=>"011111110",
  45696=>"001000011",
  45697=>"000111001",
  45698=>"101111010",
  45699=>"010011110",
  45700=>"000011110",
  45701=>"111010011",
  45702=>"101000100",
  45703=>"101110110",
  45704=>"000010001",
  45705=>"001111101",
  45706=>"111101101",
  45707=>"110110000",
  45708=>"110110000",
  45709=>"000010000",
  45710=>"011010110",
  45711=>"110011001",
  45712=>"001010101",
  45713=>"101001111",
  45714=>"000000111",
  45715=>"111010011",
  45716=>"000100101",
  45717=>"101010010",
  45718=>"010100101",
  45719=>"111110100",
  45720=>"001111000",
  45721=>"000000000",
  45722=>"001000110",
  45723=>"111011111",
  45724=>"101010110",
  45725=>"000001000",
  45726=>"101101000",
  45727=>"011011111",
  45728=>"011001111",
  45729=>"110100100",
  45730=>"000110011",
  45731=>"010100111",
  45732=>"001000001",
  45733=>"111100000",
  45734=>"111100000",
  45735=>"001010111",
  45736=>"000110111",
  45737=>"001000011",
  45738=>"001000100",
  45739=>"000100001",
  45740=>"101101011",
  45741=>"011100101",
  45742=>"000100101",
  45743=>"001000111",
  45744=>"011011111",
  45745=>"001110110",
  45746=>"010111111",
  45747=>"100011001",
  45748=>"111101001",
  45749=>"000101000",
  45750=>"111111111",
  45751=>"101111100",
  45752=>"000000111",
  45753=>"010111001",
  45754=>"001111110",
  45755=>"000000110",
  45756=>"011101011",
  45757=>"101001001",
  45758=>"000101011",
  45759=>"001111110",
  45760=>"011110111",
  45761=>"010010101",
  45762=>"011001010",
  45763=>"111100111",
  45764=>"111111100",
  45765=>"101110011",
  45766=>"000110110",
  45767=>"000001111",
  45768=>"101000110",
  45769=>"100000101",
  45770=>"011010010",
  45771=>"110101011",
  45772=>"101101000",
  45773=>"010000111",
  45774=>"101000011",
  45775=>"110110010",
  45776=>"001000111",
  45777=>"111111001",
  45778=>"110110001",
  45779=>"010101011",
  45780=>"111101000",
  45781=>"111110011",
  45782=>"111000110",
  45783=>"101000011",
  45784=>"110011111",
  45785=>"011100010",
  45786=>"000010000",
  45787=>"100011101",
  45788=>"100110110",
  45789=>"001110111",
  45790=>"101000010",
  45791=>"000000111",
  45792=>"101011110",
  45793=>"000000001",
  45794=>"000000100",
  45795=>"101000011",
  45796=>"001010010",
  45797=>"110011000",
  45798=>"110110101",
  45799=>"000100110",
  45800=>"101011101",
  45801=>"111001011",
  45802=>"111010011",
  45803=>"001001111",
  45804=>"011110100",
  45805=>"110001001",
  45806=>"010011100",
  45807=>"001000100",
  45808=>"000010000",
  45809=>"001001101",
  45810=>"001111110",
  45811=>"111011011",
  45812=>"101110001",
  45813=>"010111100",
  45814=>"100001101",
  45815=>"111000011",
  45816=>"000101100",
  45817=>"000111001",
  45818=>"011100011",
  45819=>"010101110",
  45820=>"010101011",
  45821=>"101000011",
  45822=>"101000101",
  45823=>"100110001",
  45824=>"000110000",
  45825=>"100001011",
  45826=>"111111000",
  45827=>"000011111",
  45828=>"011101011",
  45829=>"100110011",
  45830=>"010000111",
  45831=>"100000011",
  45832=>"101001011",
  45833=>"000001010",
  45834=>"111000110",
  45835=>"111001011",
  45836=>"111001000",
  45837=>"000100000",
  45838=>"010111000",
  45839=>"101010101",
  45840=>"100010100",
  45841=>"100010011",
  45842=>"100100100",
  45843=>"000001111",
  45844=>"001110111",
  45845=>"101101111",
  45846=>"110001100",
  45847=>"101111111",
  45848=>"101011011",
  45849=>"001101001",
  45850=>"011000101",
  45851=>"110001010",
  45852=>"001000100",
  45853=>"011100111",
  45854=>"001001010",
  45855=>"100000011",
  45856=>"011010111",
  45857=>"000111110",
  45858=>"011010111",
  45859=>"101000111",
  45860=>"011110011",
  45861=>"000001010",
  45862=>"000110111",
  45863=>"111010011",
  45864=>"001001110",
  45865=>"011000110",
  45866=>"111001111",
  45867=>"111111101",
  45868=>"010010001",
  45869=>"011001110",
  45870=>"011000100",
  45871=>"111000001",
  45872=>"011111100",
  45873=>"011001001",
  45874=>"100010110",
  45875=>"101101100",
  45876=>"010011010",
  45877=>"100111101",
  45878=>"000011110",
  45879=>"000000111",
  45880=>"100111001",
  45881=>"100100011",
  45882=>"101010001",
  45883=>"101011101",
  45884=>"001010001",
  45885=>"000001000",
  45886=>"001111000",
  45887=>"011110110",
  45888=>"100011100",
  45889=>"001111111",
  45890=>"011000010",
  45891=>"100100110",
  45892=>"100011100",
  45893=>"111010011",
  45894=>"010111101",
  45895=>"000011110",
  45896=>"111110100",
  45897=>"101011110",
  45898=>"000110000",
  45899=>"010101000",
  45900=>"100101110",
  45901=>"000111001",
  45902=>"101101110",
  45903=>"100011000",
  45904=>"001000101",
  45905=>"101111111",
  45906=>"000101100",
  45907=>"011110001",
  45908=>"101110000",
  45909=>"101100000",
  45910=>"111000001",
  45911=>"000100110",
  45912=>"110011110",
  45913=>"010111010",
  45914=>"100100110",
  45915=>"100000110",
  45916=>"111010000",
  45917=>"010100000",
  45918=>"010111110",
  45919=>"001000111",
  45920=>"000001000",
  45921=>"001010000",
  45922=>"000001100",
  45923=>"100100111",
  45924=>"111011101",
  45925=>"011000000",
  45926=>"000010001",
  45927=>"101010100",
  45928=>"011100001",
  45929=>"110001011",
  45930=>"101111011",
  45931=>"011010110",
  45932=>"001111011",
  45933=>"001011000",
  45934=>"100010000",
  45935=>"011001101",
  45936=>"100111000",
  45937=>"101000010",
  45938=>"110101000",
  45939=>"110001111",
  45940=>"001100100",
  45941=>"000010011",
  45942=>"010000011",
  45943=>"110000000",
  45944=>"101000010",
  45945=>"011001000",
  45946=>"110101110",
  45947=>"001001100",
  45948=>"011011010",
  45949=>"101110101",
  45950=>"101110011",
  45951=>"011011100",
  45952=>"001010101",
  45953=>"010001000",
  45954=>"110001011",
  45955=>"111000101",
  45956=>"000110001",
  45957=>"101010011",
  45958=>"001110110",
  45959=>"011010010",
  45960=>"101101101",
  45961=>"111111010",
  45962=>"110110101",
  45963=>"101001011",
  45964=>"100001111",
  45965=>"011101111",
  45966=>"011110111",
  45967=>"010111101",
  45968=>"101100000",
  45969=>"000101000",
  45970=>"100110011",
  45971=>"110101011",
  45972=>"000001100",
  45973=>"101011011",
  45974=>"110010111",
  45975=>"010001110",
  45976=>"010100010",
  45977=>"101111101",
  45978=>"000100001",
  45979=>"101000001",
  45980=>"000110110",
  45981=>"000011110",
  45982=>"000101000",
  45983=>"100111101",
  45984=>"111111011",
  45985=>"011011001",
  45986=>"011000111",
  45987=>"110000111",
  45988=>"000001110",
  45989=>"110101110",
  45990=>"101011101",
  45991=>"111100111",
  45992=>"001011101",
  45993=>"010010000",
  45994=>"100110111",
  45995=>"000110110",
  45996=>"000111111",
  45997=>"000010000",
  45998=>"100001010",
  45999=>"100100011",
  46000=>"111101110",
  46001=>"101110110",
  46002=>"000110101",
  46003=>"100100011",
  46004=>"011101001",
  46005=>"111101010",
  46006=>"100001110",
  46007=>"000001110",
  46008=>"101011110",
  46009=>"011100010",
  46010=>"100010111",
  46011=>"000110101",
  46012=>"001110001",
  46013=>"000101100",
  46014=>"010100000",
  46015=>"001001000",
  46016=>"101000000",
  46017=>"101011011",
  46018=>"010101011",
  46019=>"011100011",
  46020=>"001011010",
  46021=>"111101111",
  46022=>"101000111",
  46023=>"001000011",
  46024=>"011011011",
  46025=>"111000111",
  46026=>"100010010",
  46027=>"000000010",
  46028=>"101111010",
  46029=>"001111110",
  46030=>"000100101",
  46031=>"101101111",
  46032=>"000110100",
  46033=>"000000111",
  46034=>"110001011",
  46035=>"011101011",
  46036=>"000100001",
  46037=>"011100101",
  46038=>"001000100",
  46039=>"101010110",
  46040=>"001111000",
  46041=>"100010111",
  46042=>"111010110",
  46043=>"101000000",
  46044=>"000010101",
  46045=>"001011101",
  46046=>"000001100",
  46047=>"001110111",
  46048=>"010000000",
  46049=>"100000100",
  46050=>"001110111",
  46051=>"111111101",
  46052=>"100110001",
  46053=>"010111000",
  46054=>"100010000",
  46055=>"101101001",
  46056=>"101111010",
  46057=>"101011001",
  46058=>"110011100",
  46059=>"110111001",
  46060=>"110101000",
  46061=>"001100010",
  46062=>"101001100",
  46063=>"110011111",
  46064=>"010111001",
  46065=>"010011100",
  46066=>"010111111",
  46067=>"110100110",
  46068=>"001001111",
  46069=>"011001110",
  46070=>"000001010",
  46071=>"100111110",
  46072=>"100011000",
  46073=>"111100000",
  46074=>"110011111",
  46075=>"100011011",
  46076=>"001001000",
  46077=>"101001100",
  46078=>"001101001",
  46079=>"001100111",
  46080=>"111101110",
  46081=>"000111001",
  46082=>"000101100",
  46083=>"011100101",
  46084=>"111100111",
  46085=>"111010001",
  46086=>"100101101",
  46087=>"011001111",
  46088=>"010101100",
  46089=>"011000000",
  46090=>"000000010",
  46091=>"110011111",
  46092=>"000111000",
  46093=>"110111000",
  46094=>"011101111",
  46095=>"000011000",
  46096=>"111000000",
  46097=>"100111100",
  46098=>"000110011",
  46099=>"111010111",
  46100=>"000011101",
  46101=>"100010011",
  46102=>"011010010",
  46103=>"101000111",
  46104=>"110001100",
  46105=>"001110100",
  46106=>"001010011",
  46107=>"011100001",
  46108=>"011010010",
  46109=>"100101111",
  46110=>"010110111",
  46111=>"101101110",
  46112=>"110010111",
  46113=>"100000101",
  46114=>"011111100",
  46115=>"111111100",
  46116=>"101011110",
  46117=>"010110110",
  46118=>"101101110",
  46119=>"010000110",
  46120=>"111111000",
  46121=>"110101101",
  46122=>"010010110",
  46123=>"011000010",
  46124=>"111001000",
  46125=>"110010101",
  46126=>"011100010",
  46127=>"010110001",
  46128=>"001011100",
  46129=>"101100111",
  46130=>"000010110",
  46131=>"111111111",
  46132=>"011011010",
  46133=>"110111000",
  46134=>"011000111",
  46135=>"101001011",
  46136=>"000000111",
  46137=>"011000010",
  46138=>"100110010",
  46139=>"001101000",
  46140=>"000110110",
  46141=>"010011000",
  46142=>"100000110",
  46143=>"000111111",
  46144=>"101100000",
  46145=>"110011011",
  46146=>"001101110",
  46147=>"011101001",
  46148=>"000000101",
  46149=>"110111010",
  46150=>"000111011",
  46151=>"000000101",
  46152=>"101000110",
  46153=>"100011001",
  46154=>"001111010",
  46155=>"000101111",
  46156=>"001111101",
  46157=>"001100111",
  46158=>"111110111",
  46159=>"111111011",
  46160=>"000101000",
  46161=>"001010010",
  46162=>"111001110",
  46163=>"101000000",
  46164=>"001110010",
  46165=>"101001100",
  46166=>"001100011",
  46167=>"101001101",
  46168=>"101011111",
  46169=>"001100110",
  46170=>"101111010",
  46171=>"010001011",
  46172=>"010100110",
  46173=>"000101010",
  46174=>"100011001",
  46175=>"100100010",
  46176=>"110111011",
  46177=>"101001001",
  46178=>"001100011",
  46179=>"000011010",
  46180=>"110101111",
  46181=>"010111010",
  46182=>"111000110",
  46183=>"011111000",
  46184=>"111111101",
  46185=>"110100000",
  46186=>"111001111",
  46187=>"100011111",
  46188=>"000001011",
  46189=>"100100100",
  46190=>"000010010",
  46191=>"111101111",
  46192=>"011011110",
  46193=>"000001111",
  46194=>"111110101",
  46195=>"010011000",
  46196=>"001011100",
  46197=>"010101000",
  46198=>"000010010",
  46199=>"000001010",
  46200=>"001110001",
  46201=>"000011000",
  46202=>"100111001",
  46203=>"101000010",
  46204=>"101100010",
  46205=>"100010101",
  46206=>"111100100",
  46207=>"110000001",
  46208=>"001011001",
  46209=>"010010000",
  46210=>"000110101",
  46211=>"101011010",
  46212=>"010101110",
  46213=>"011111011",
  46214=>"011100000",
  46215=>"111111000",
  46216=>"011001011",
  46217=>"010111101",
  46218=>"110001000",
  46219=>"100110111",
  46220=>"000101111",
  46221=>"110101110",
  46222=>"111110011",
  46223=>"111011001",
  46224=>"011110001",
  46225=>"001110011",
  46226=>"010111110",
  46227=>"000100110",
  46228=>"110111000",
  46229=>"101001100",
  46230=>"110001010",
  46231=>"111100001",
  46232=>"001100000",
  46233=>"010001100",
  46234=>"010111010",
  46235=>"110001000",
  46236=>"000100100",
  46237=>"111000011",
  46238=>"110101010",
  46239=>"010000100",
  46240=>"100000100",
  46241=>"000100001",
  46242=>"100000010",
  46243=>"111111011",
  46244=>"110010011",
  46245=>"111010011",
  46246=>"101011100",
  46247=>"110010011",
  46248=>"111011100",
  46249=>"010000100",
  46250=>"011100000",
  46251=>"011000010",
  46252=>"110111010",
  46253=>"110100010",
  46254=>"100111110",
  46255=>"111000001",
  46256=>"001110111",
  46257=>"110100001",
  46258=>"011111000",
  46259=>"110001001",
  46260=>"000100101",
  46261=>"100011001",
  46262=>"111100011",
  46263=>"010101010",
  46264=>"010101100",
  46265=>"101100101",
  46266=>"000100000",
  46267=>"111111010",
  46268=>"111001100",
  46269=>"000111010",
  46270=>"011010010",
  46271=>"011110010",
  46272=>"010000110",
  46273=>"111001001",
  46274=>"101101100",
  46275=>"000011010",
  46276=>"111111110",
  46277=>"010000000",
  46278=>"011011110",
  46279=>"000011010",
  46280=>"011101101",
  46281=>"001101010",
  46282=>"100011001",
  46283=>"010001010",
  46284=>"000111110",
  46285=>"111010110",
  46286=>"111010111",
  46287=>"111101000",
  46288=>"011011011",
  46289=>"100100010",
  46290=>"101110101",
  46291=>"011111000",
  46292=>"100100010",
  46293=>"111100001",
  46294=>"110001111",
  46295=>"011111010",
  46296=>"110100100",
  46297=>"000000010",
  46298=>"010100111",
  46299=>"000100111",
  46300=>"100011100",
  46301=>"101000001",
  46302=>"111100111",
  46303=>"010111111",
  46304=>"001001000",
  46305=>"110111011",
  46306=>"011010110",
  46307=>"001000010",
  46308=>"100000011",
  46309=>"010001111",
  46310=>"011000011",
  46311=>"010100010",
  46312=>"000101111",
  46313=>"111110000",
  46314=>"011001100",
  46315=>"101001010",
  46316=>"011110100",
  46317=>"101110111",
  46318=>"110110111",
  46319=>"010100110",
  46320=>"011100001",
  46321=>"011000100",
  46322=>"010101101",
  46323=>"101001111",
  46324=>"111011000",
  46325=>"100010000",
  46326=>"001001001",
  46327=>"001010110",
  46328=>"000001110",
  46329=>"110010001",
  46330=>"100110010",
  46331=>"001111000",
  46332=>"000100100",
  46333=>"000100101",
  46334=>"001000010",
  46335=>"101011000",
  46336=>"111010000",
  46337=>"100101001",
  46338=>"111000010",
  46339=>"001000101",
  46340=>"110100011",
  46341=>"101100111",
  46342=>"101100101",
  46343=>"111001111",
  46344=>"011111100",
  46345=>"000000100",
  46346=>"010100100",
  46347=>"010001100",
  46348=>"000001101",
  46349=>"111101011",
  46350=>"010111110",
  46351=>"001111010",
  46352=>"110000000",
  46353=>"100000000",
  46354=>"011000000",
  46355=>"001001101",
  46356=>"111011010",
  46357=>"000000001",
  46358=>"111011101",
  46359=>"011101100",
  46360=>"111111000",
  46361=>"110011001",
  46362=>"001001100",
  46363=>"111000100",
  46364=>"101001110",
  46365=>"111111011",
  46366=>"100001000",
  46367=>"000001001",
  46368=>"111110111",
  46369=>"001000001",
  46370=>"101010000",
  46371=>"001001100",
  46372=>"111110100",
  46373=>"111011011",
  46374=>"011000001",
  46375=>"111111110",
  46376=>"101010110",
  46377=>"011101101",
  46378=>"010100101",
  46379=>"000100000",
  46380=>"111101111",
  46381=>"100101100",
  46382=>"101101010",
  46383=>"100110111",
  46384=>"110010101",
  46385=>"100000110",
  46386=>"100111011",
  46387=>"000010000",
  46388=>"111000100",
  46389=>"000110100",
  46390=>"000011000",
  46391=>"111000000",
  46392=>"001100111",
  46393=>"010001101",
  46394=>"111100001",
  46395=>"010100111",
  46396=>"001100010",
  46397=>"000000011",
  46398=>"000001001",
  46399=>"001100001",
  46400=>"001110000",
  46401=>"000000001",
  46402=>"000100111",
  46403=>"111000101",
  46404=>"100000001",
  46405=>"111001000",
  46406=>"011111111",
  46407=>"110110110",
  46408=>"011000010",
  46409=>"101001100",
  46410=>"110101100",
  46411=>"100001000",
  46412=>"001000000",
  46413=>"000110101",
  46414=>"110110010",
  46415=>"111110100",
  46416=>"111001010",
  46417=>"110011000",
  46418=>"110000100",
  46419=>"011111011",
  46420=>"101111001",
  46421=>"111001111",
  46422=>"101111100",
  46423=>"000001001",
  46424=>"001101101",
  46425=>"000101000",
  46426=>"011100110",
  46427=>"000101111",
  46428=>"001001100",
  46429=>"110110001",
  46430=>"101011111",
  46431=>"000110100",
  46432=>"000010110",
  46433=>"011101001",
  46434=>"010001111",
  46435=>"101100011",
  46436=>"100101001",
  46437=>"110101001",
  46438=>"111011011",
  46439=>"010011110",
  46440=>"010001001",
  46441=>"000101101",
  46442=>"011111010",
  46443=>"100010001",
  46444=>"000011011",
  46445=>"000111111",
  46446=>"010110010",
  46447=>"100001101",
  46448=>"010111001",
  46449=>"110110001",
  46450=>"011000100",
  46451=>"101000101",
  46452=>"001101110",
  46453=>"001011111",
  46454=>"101011110",
  46455=>"001101100",
  46456=>"000110000",
  46457=>"101000111",
  46458=>"111011110",
  46459=>"100100111",
  46460=>"101000000",
  46461=>"001000010",
  46462=>"011011111",
  46463=>"000100100",
  46464=>"100010000",
  46465=>"111000001",
  46466=>"001101101",
  46467=>"110011001",
  46468=>"111100100",
  46469=>"110010111",
  46470=>"101000101",
  46471=>"010010001",
  46472=>"100010000",
  46473=>"111010110",
  46474=>"111100101",
  46475=>"100000100",
  46476=>"011000011",
  46477=>"000000110",
  46478=>"011000010",
  46479=>"111010101",
  46480=>"101101011",
  46481=>"001001000",
  46482=>"000101011",
  46483=>"101100101",
  46484=>"100110100",
  46485=>"110111000",
  46486=>"011000101",
  46487=>"101011110",
  46488=>"100011010",
  46489=>"000001000",
  46490=>"000100010",
  46491=>"011010111",
  46492=>"111011010",
  46493=>"100001000",
  46494=>"101000100",
  46495=>"000111111",
  46496=>"101101001",
  46497=>"101000111",
  46498=>"011110101",
  46499=>"001001100",
  46500=>"100101000",
  46501=>"001000000",
  46502=>"000100001",
  46503=>"100101011",
  46504=>"000011010",
  46505=>"010110111",
  46506=>"000101001",
  46507=>"100100011",
  46508=>"110000010",
  46509=>"111010010",
  46510=>"111111100",
  46511=>"010011111",
  46512=>"101110100",
  46513=>"011101010",
  46514=>"011000001",
  46515=>"000011111",
  46516=>"111011111",
  46517=>"011111011",
  46518=>"000000010",
  46519=>"100001100",
  46520=>"010001000",
  46521=>"000101110",
  46522=>"000110101",
  46523=>"101011011",
  46524=>"011110010",
  46525=>"000001111",
  46526=>"001100001",
  46527=>"100010011",
  46528=>"101001101",
  46529=>"011010000",
  46530=>"011100000",
  46531=>"111111111",
  46532=>"010000100",
  46533=>"101001110",
  46534=>"000100000",
  46535=>"010000000",
  46536=>"110011001",
  46537=>"101101101",
  46538=>"010010010",
  46539=>"110000110",
  46540=>"000100111",
  46541=>"011011000",
  46542=>"001100111",
  46543=>"100011111",
  46544=>"001100100",
  46545=>"000011101",
  46546=>"011111000",
  46547=>"110110100",
  46548=>"000001111",
  46549=>"001111011",
  46550=>"111011000",
  46551=>"101110110",
  46552=>"011100111",
  46553=>"000000011",
  46554=>"110001001",
  46555=>"011011011",
  46556=>"010001111",
  46557=>"010011010",
  46558=>"100101000",
  46559=>"010101101",
  46560=>"000010011",
  46561=>"001011110",
  46562=>"001000110",
  46563=>"011011011",
  46564=>"100000010",
  46565=>"101101110",
  46566=>"010101000",
  46567=>"011100000",
  46568=>"000100001",
  46569=>"010100110",
  46570=>"111100101",
  46571=>"101010110",
  46572=>"100010100",
  46573=>"000110110",
  46574=>"010111011",
  46575=>"101101001",
  46576=>"110011000",
  46577=>"010101010",
  46578=>"101110010",
  46579=>"101110000",
  46580=>"100010010",
  46581=>"110110100",
  46582=>"001101001",
  46583=>"100110010",
  46584=>"011011000",
  46585=>"100101111",
  46586=>"111111101",
  46587=>"001111000",
  46588=>"011010110",
  46589=>"000011100",
  46590=>"101100010",
  46591=>"001000001",
  46592=>"010101101",
  46593=>"100001011",
  46594=>"000100010",
  46595=>"111101111",
  46596=>"110000100",
  46597=>"010100011",
  46598=>"100010000",
  46599=>"100111000",
  46600=>"001000000",
  46601=>"100100001",
  46602=>"000100100",
  46603=>"000111011",
  46604=>"100101011",
  46605=>"000000001",
  46606=>"111100101",
  46607=>"001001010",
  46608=>"000110110",
  46609=>"000010001",
  46610=>"000011101",
  46611=>"010101110",
  46612=>"110001100",
  46613=>"011010010",
  46614=>"101011001",
  46615=>"101001110",
  46616=>"000110101",
  46617=>"001000010",
  46618=>"011111010",
  46619=>"111110010",
  46620=>"110111000",
  46621=>"011001000",
  46622=>"011000101",
  46623=>"011000111",
  46624=>"110101110",
  46625=>"000011110",
  46626=>"000000011",
  46627=>"110010000",
  46628=>"011010101",
  46629=>"101000111",
  46630=>"001010100",
  46631=>"100010001",
  46632=>"110100000",
  46633=>"001010100",
  46634=>"000011000",
  46635=>"000000011",
  46636=>"010000001",
  46637=>"110100100",
  46638=>"111110110",
  46639=>"001101111",
  46640=>"101110010",
  46641=>"111110110",
  46642=>"101000100",
  46643=>"010110100",
  46644=>"011101101",
  46645=>"010011011",
  46646=>"001111110",
  46647=>"011110101",
  46648=>"011110111",
  46649=>"001101111",
  46650=>"010101110",
  46651=>"100010001",
  46652=>"011101000",
  46653=>"111111011",
  46654=>"011011100",
  46655=>"001010000",
  46656=>"100000111",
  46657=>"000000111",
  46658=>"101010111",
  46659=>"011010110",
  46660=>"110100010",
  46661=>"010001010",
  46662=>"001101110",
  46663=>"110010000",
  46664=>"111000101",
  46665=>"000111001",
  46666=>"101101000",
  46667=>"011011001",
  46668=>"011110101",
  46669=>"110100101",
  46670=>"101001001",
  46671=>"001100100",
  46672=>"111001110",
  46673=>"100001000",
  46674=>"010110001",
  46675=>"001111010",
  46676=>"000010100",
  46677=>"000010011",
  46678=>"000110000",
  46679=>"111110101",
  46680=>"110001111",
  46681=>"001001010",
  46682=>"101011001",
  46683=>"001010000",
  46684=>"000000000",
  46685=>"100101010",
  46686=>"101111011",
  46687=>"101111000",
  46688=>"100011001",
  46689=>"100001010",
  46690=>"100111100",
  46691=>"011001111",
  46692=>"010011011",
  46693=>"000111100",
  46694=>"001111100",
  46695=>"110100100",
  46696=>"010000011",
  46697=>"101001000",
  46698=>"111101111",
  46699=>"110100100",
  46700=>"100100111",
  46701=>"011101001",
  46702=>"111101001",
  46703=>"101110111",
  46704=>"100111100",
  46705=>"001000000",
  46706=>"001011101",
  46707=>"101010111",
  46708=>"001110011",
  46709=>"111100110",
  46710=>"000111000",
  46711=>"100011010",
  46712=>"110001000",
  46713=>"100001101",
  46714=>"101011111",
  46715=>"000010001",
  46716=>"000000100",
  46717=>"110000111",
  46718=>"011000101",
  46719=>"111111001",
  46720=>"101011000",
  46721=>"111001001",
  46722=>"110011011",
  46723=>"100001111",
  46724=>"011100010",
  46725=>"000010010",
  46726=>"011000011",
  46727=>"100101000",
  46728=>"000110001",
  46729=>"001001001",
  46730=>"011011010",
  46731=>"000010100",
  46732=>"000000101",
  46733=>"110101001",
  46734=>"110010100",
  46735=>"101100111",
  46736=>"010100001",
  46737=>"011101110",
  46738=>"011101100",
  46739=>"101101101",
  46740=>"100011000",
  46741=>"100011111",
  46742=>"000100111",
  46743=>"010101000",
  46744=>"111010010",
  46745=>"101000010",
  46746=>"100001100",
  46747=>"011010011",
  46748=>"101110111",
  46749=>"101010001",
  46750=>"010011000",
  46751=>"110000000",
  46752=>"011011010",
  46753=>"010100010",
  46754=>"100010111",
  46755=>"110101000",
  46756=>"000011110",
  46757=>"011011101",
  46758=>"000101101",
  46759=>"110011000",
  46760=>"000000011",
  46761=>"000001000",
  46762=>"000000000",
  46763=>"100001110",
  46764=>"111100101",
  46765=>"000101010",
  46766=>"011011100",
  46767=>"110101000",
  46768=>"010000110",
  46769=>"011100010",
  46770=>"100000001",
  46771=>"011010111",
  46772=>"001111011",
  46773=>"111010110",
  46774=>"100110001",
  46775=>"111011011",
  46776=>"110010101",
  46777=>"111010101",
  46778=>"111000010",
  46779=>"011101000",
  46780=>"001100110",
  46781=>"101010000",
  46782=>"101001001",
  46783=>"110111011",
  46784=>"100000110",
  46785=>"011110011",
  46786=>"110101000",
  46787=>"100011000",
  46788=>"111111110",
  46789=>"011011010",
  46790=>"010100010",
  46791=>"010000000",
  46792=>"111100100",
  46793=>"001000111",
  46794=>"100000011",
  46795=>"111101110",
  46796=>"001001011",
  46797=>"001000101",
  46798=>"110100100",
  46799=>"011011100",
  46800=>"100010011",
  46801=>"101000010",
  46802=>"111111010",
  46803=>"011111100",
  46804=>"000101101",
  46805=>"111010111",
  46806=>"011111000",
  46807=>"100001000",
  46808=>"000011101",
  46809=>"010001100",
  46810=>"101001111",
  46811=>"001000111",
  46812=>"101001010",
  46813=>"011101000",
  46814=>"010100101",
  46815=>"100011011",
  46816=>"110011100",
  46817=>"100100110",
  46818=>"111011100",
  46819=>"101000000",
  46820=>"100101001",
  46821=>"001000110",
  46822=>"000110011",
  46823=>"101011010",
  46824=>"100100111",
  46825=>"110101001",
  46826=>"110011011",
  46827=>"010010011",
  46828=>"101101011",
  46829=>"101111000",
  46830=>"111011111",
  46831=>"000110100",
  46832=>"010110100",
  46833=>"000110011",
  46834=>"011110010",
  46835=>"101000101",
  46836=>"000010110",
  46837=>"000001110",
  46838=>"011010111",
  46839=>"111110100",
  46840=>"011001001",
  46841=>"100001100",
  46842=>"000101010",
  46843=>"110010110",
  46844=>"100001001",
  46845=>"000100110",
  46846=>"010011011",
  46847=>"111111011",
  46848=>"101011100",
  46849=>"010101100",
  46850=>"011000001",
  46851=>"111000001",
  46852=>"110111100",
  46853=>"000010011",
  46854=>"010010000",
  46855=>"110011100",
  46856=>"011111000",
  46857=>"101011000",
  46858=>"101010000",
  46859=>"101000100",
  46860=>"011001000",
  46861=>"011111011",
  46862=>"010010011",
  46863=>"000110000",
  46864=>"000110001",
  46865=>"000110000",
  46866=>"001010011",
  46867=>"101110101",
  46868=>"101110000",
  46869=>"010011000",
  46870=>"000001010",
  46871=>"101000011",
  46872=>"111001111",
  46873=>"001110000",
  46874=>"100111001",
  46875=>"000000011",
  46876=>"010010110",
  46877=>"010011110",
  46878=>"110100101",
  46879=>"110011011",
  46880=>"110010001",
  46881=>"111111000",
  46882=>"111010110",
  46883=>"100000001",
  46884=>"100101111",
  46885=>"111100101",
  46886=>"010100110",
  46887=>"101100000",
  46888=>"010001000",
  46889=>"101010001",
  46890=>"101011000",
  46891=>"000010001",
  46892=>"110111011",
  46893=>"111110111",
  46894=>"010000101",
  46895=>"110100111",
  46896=>"000001010",
  46897=>"110100100",
  46898=>"001011001",
  46899=>"000001111",
  46900=>"101000111",
  46901=>"110010100",
  46902=>"100011100",
  46903=>"010010110",
  46904=>"100111011",
  46905=>"111110110",
  46906=>"000010100",
  46907=>"111011101",
  46908=>"111101100",
  46909=>"101110111",
  46910=>"001001110",
  46911=>"100011100",
  46912=>"010011011",
  46913=>"000000000",
  46914=>"101100001",
  46915=>"100100100",
  46916=>"101011010",
  46917=>"011111111",
  46918=>"010000100",
  46919=>"000010001",
  46920=>"101010100",
  46921=>"001000100",
  46922=>"010001111",
  46923=>"011100010",
  46924=>"101011100",
  46925=>"110110001",
  46926=>"010011110",
  46927=>"001001100",
  46928=>"101110110",
  46929=>"110000100",
  46930=>"111100101",
  46931=>"101001101",
  46932=>"000000110",
  46933=>"010000001",
  46934=>"011100010",
  46935=>"010010100",
  46936=>"111100000",
  46937=>"011101010",
  46938=>"100011100",
  46939=>"111001111",
  46940=>"101001010",
  46941=>"100011011",
  46942=>"111000000",
  46943=>"000100111",
  46944=>"000101011",
  46945=>"011001100",
  46946=>"000111011",
  46947=>"101010110",
  46948=>"011101000",
  46949=>"000101110",
  46950=>"111110111",
  46951=>"011111111",
  46952=>"010110100",
  46953=>"100111011",
  46954=>"010010000",
  46955=>"110101111",
  46956=>"111011000",
  46957=>"010000100",
  46958=>"001111100",
  46959=>"110011111",
  46960=>"110010001",
  46961=>"111101011",
  46962=>"110000101",
  46963=>"000000001",
  46964=>"010000110",
  46965=>"100110001",
  46966=>"000111011",
  46967=>"110001111",
  46968=>"000101000",
  46969=>"101100101",
  46970=>"111110011",
  46971=>"000101011",
  46972=>"111001000",
  46973=>"100011100",
  46974=>"110110111",
  46975=>"010011010",
  46976=>"010001011",
  46977=>"001101111",
  46978=>"011100001",
  46979=>"100100111",
  46980=>"000100111",
  46981=>"100001101",
  46982=>"000101100",
  46983=>"011111011",
  46984=>"101010001",
  46985=>"010000001",
  46986=>"000000101",
  46987=>"111001011",
  46988=>"001110111",
  46989=>"101011110",
  46990=>"101101010",
  46991=>"111001011",
  46992=>"111101111",
  46993=>"110001101",
  46994=>"000000010",
  46995=>"110110101",
  46996=>"101000001",
  46997=>"111100010",
  46998=>"110111001",
  46999=>"000111011",
  47000=>"100000110",
  47001=>"100011010",
  47002=>"001101000",
  47003=>"110101111",
  47004=>"011101111",
  47005=>"001101110",
  47006=>"000010110",
  47007=>"011110001",
  47008=>"100110001",
  47009=>"111010000",
  47010=>"010100111",
  47011=>"100001111",
  47012=>"100000101",
  47013=>"010000110",
  47014=>"110111001",
  47015=>"110110101",
  47016=>"010110100",
  47017=>"100001011",
  47018=>"101011111",
  47019=>"111010100",
  47020=>"000001001",
  47021=>"011111111",
  47022=>"100011000",
  47023=>"001101000",
  47024=>"111010011",
  47025=>"010101011",
  47026=>"111000110",
  47027=>"001110000",
  47028=>"111110010",
  47029=>"100010010",
  47030=>"010010010",
  47031=>"010010000",
  47032=>"100100010",
  47033=>"011000110",
  47034=>"110101000",
  47035=>"111100110",
  47036=>"100100111",
  47037=>"010100100",
  47038=>"101010110",
  47039=>"000101011",
  47040=>"010110000",
  47041=>"001001101",
  47042=>"110011001",
  47043=>"111000100",
  47044=>"100011110",
  47045=>"110011110",
  47046=>"011111011",
  47047=>"101001100",
  47048=>"110011111",
  47049=>"000110110",
  47050=>"000100100",
  47051=>"111001010",
  47052=>"000011111",
  47053=>"100100111",
  47054=>"000011111",
  47055=>"001100111",
  47056=>"010111110",
  47057=>"001010011",
  47058=>"111101010",
  47059=>"110111111",
  47060=>"000010111",
  47061=>"000010111",
  47062=>"100111101",
  47063=>"001110111",
  47064=>"001000000",
  47065=>"101110011",
  47066=>"001000000",
  47067=>"110100110",
  47068=>"101111111",
  47069=>"110011011",
  47070=>"111101101",
  47071=>"111001010",
  47072=>"001111001",
  47073=>"010101100",
  47074=>"110110000",
  47075=>"000101101",
  47076=>"011110011",
  47077=>"011001100",
  47078=>"110011110",
  47079=>"000100101",
  47080=>"000000101",
  47081=>"100111101",
  47082=>"010001101",
  47083=>"110100100",
  47084=>"101101111",
  47085=>"110011100",
  47086=>"000000010",
  47087=>"001101100",
  47088=>"101111101",
  47089=>"001001111",
  47090=>"101110010",
  47091=>"001011000",
  47092=>"010000100",
  47093=>"101111000",
  47094=>"100001101",
  47095=>"001111010",
  47096=>"011011111",
  47097=>"100100101",
  47098=>"100001011",
  47099=>"111101001",
  47100=>"100011111",
  47101=>"010100011",
  47102=>"001100101",
  47103=>"011101011",
  47104=>"101101110",
  47105=>"111101110",
  47106=>"010110010",
  47107=>"001100010",
  47108=>"100101000",
  47109=>"010111011",
  47110=>"011111010",
  47111=>"111110101",
  47112=>"100100101",
  47113=>"100000100",
  47114=>"111101111",
  47115=>"010100001",
  47116=>"011010111",
  47117=>"101000001",
  47118=>"111001100",
  47119=>"100101010",
  47120=>"100000001",
  47121=>"001001001",
  47122=>"001000010",
  47123=>"000110110",
  47124=>"011011011",
  47125=>"101101111",
  47126=>"100010001",
  47127=>"101011110",
  47128=>"111011110",
  47129=>"101000011",
  47130=>"100110011",
  47131=>"011110110",
  47132=>"001011010",
  47133=>"101011000",
  47134=>"000010001",
  47135=>"100110000",
  47136=>"010010100",
  47137=>"000101111",
  47138=>"111000001",
  47139=>"101110110",
  47140=>"010000101",
  47141=>"101010101",
  47142=>"001110010",
  47143=>"110001000",
  47144=>"000011100",
  47145=>"100101111",
  47146=>"000000010",
  47147=>"001001101",
  47148=>"010010001",
  47149=>"001101011",
  47150=>"011111001",
  47151=>"010011011",
  47152=>"100000000",
  47153=>"010001111",
  47154=>"011001001",
  47155=>"100110111",
  47156=>"110011001",
  47157=>"010100101",
  47158=>"001101011",
  47159=>"001110000",
  47160=>"111100001",
  47161=>"110000101",
  47162=>"100100010",
  47163=>"101000101",
  47164=>"000011101",
  47165=>"011011001",
  47166=>"110001110",
  47167=>"100001011",
  47168=>"011101001",
  47169=>"001100101",
  47170=>"111101010",
  47171=>"011101000",
  47172=>"111110110",
  47173=>"010100101",
  47174=>"010110110",
  47175=>"001101001",
  47176=>"010010110",
  47177=>"011110100",
  47178=>"111000011",
  47179=>"101101001",
  47180=>"011110011",
  47181=>"110100110",
  47182=>"010110101",
  47183=>"001001001",
  47184=>"001110010",
  47185=>"000110101",
  47186=>"100110101",
  47187=>"101101001",
  47188=>"010111100",
  47189=>"101101010",
  47190=>"011101111",
  47191=>"100000100",
  47192=>"101001001",
  47193=>"001110011",
  47194=>"001001010",
  47195=>"111001110",
  47196=>"010010000",
  47197=>"110110011",
  47198=>"000010111",
  47199=>"110100010",
  47200=>"111100010",
  47201=>"100000111",
  47202=>"001000000",
  47203=>"001010111",
  47204=>"010001010",
  47205=>"111011001",
  47206=>"000110100",
  47207=>"000110010",
  47208=>"000010101",
  47209=>"110101101",
  47210=>"011001110",
  47211=>"101001101",
  47212=>"100111001",
  47213=>"111111001",
  47214=>"001011000",
  47215=>"100100100",
  47216=>"000001011",
  47217=>"100110010",
  47218=>"010011100",
  47219=>"010111111",
  47220=>"111111100",
  47221=>"110111001",
  47222=>"111011000",
  47223=>"111110001",
  47224=>"010101101",
  47225=>"100001011",
  47226=>"011011100",
  47227=>"001100001",
  47228=>"010001010",
  47229=>"101000001",
  47230=>"001001100",
  47231=>"100000101",
  47232=>"010000100",
  47233=>"101111000",
  47234=>"010011100",
  47235=>"111000110",
  47236=>"000101111",
  47237=>"100000100",
  47238=>"000010010",
  47239=>"011010110",
  47240=>"100110010",
  47241=>"001011101",
  47242=>"101100110",
  47243=>"111000010",
  47244=>"101010010",
  47245=>"101000000",
  47246=>"010000000",
  47247=>"101111100",
  47248=>"101000110",
  47249=>"011010001",
  47250=>"110100010",
  47251=>"111111110",
  47252=>"011110000",
  47253=>"001100001",
  47254=>"000000101",
  47255=>"000000001",
  47256=>"001110111",
  47257=>"010110001",
  47258=>"000111001",
  47259=>"000110110",
  47260=>"001000000",
  47261=>"101111101",
  47262=>"111111101",
  47263=>"001000101",
  47264=>"011110001",
  47265=>"000111000",
  47266=>"010111111",
  47267=>"111000011",
  47268=>"110100110",
  47269=>"101100000",
  47270=>"111011110",
  47271=>"001101011",
  47272=>"000110001",
  47273=>"100101000",
  47274=>"100001101",
  47275=>"101011011",
  47276=>"110101101",
  47277=>"100001100",
  47278=>"001010110",
  47279=>"101111001",
  47280=>"100110101",
  47281=>"111001100",
  47282=>"100000100",
  47283=>"001111101",
  47284=>"011100001",
  47285=>"000101100",
  47286=>"110110110",
  47287=>"111010100",
  47288=>"110010101",
  47289=>"111110110",
  47290=>"011000101",
  47291=>"110011101",
  47292=>"000101101",
  47293=>"110111110",
  47294=>"110110110",
  47295=>"100010111",
  47296=>"001001000",
  47297=>"010011101",
  47298=>"000011101",
  47299=>"100110100",
  47300=>"001110000",
  47301=>"101101100",
  47302=>"100001011",
  47303=>"001110010",
  47304=>"110010101",
  47305=>"000110100",
  47306=>"100101110",
  47307=>"100101000",
  47308=>"100010100",
  47309=>"000101111",
  47310=>"001011011",
  47311=>"010000010",
  47312=>"110000001",
  47313=>"011101100",
  47314=>"011111110",
  47315=>"011101010",
  47316=>"110100110",
  47317=>"011100010",
  47318=>"100110100",
  47319=>"101101011",
  47320=>"001110000",
  47321=>"111100001",
  47322=>"000011111",
  47323=>"111100001",
  47324=>"100001000",
  47325=>"100111111",
  47326=>"111011101",
  47327=>"111110100",
  47328=>"010000110",
  47329=>"000001100",
  47330=>"010100000",
  47331=>"000110000",
  47332=>"100011101",
  47333=>"011001110",
  47334=>"100010001",
  47335=>"110010011",
  47336=>"011111110",
  47337=>"001100110",
  47338=>"000001010",
  47339=>"100101010",
  47340=>"001010000",
  47341=>"101000000",
  47342=>"010100100",
  47343=>"010101100",
  47344=>"111001001",
  47345=>"000011001",
  47346=>"100011001",
  47347=>"010011111",
  47348=>"100111110",
  47349=>"100111101",
  47350=>"000000011",
  47351=>"010001011",
  47352=>"111101011",
  47353=>"111000011",
  47354=>"101011001",
  47355=>"100100010",
  47356=>"011100111",
  47357=>"000001100",
  47358=>"111011000",
  47359=>"101101100",
  47360=>"010101001",
  47361=>"100010101",
  47362=>"101101100",
  47363=>"011100111",
  47364=>"101111011",
  47365=>"000100010",
  47366=>"000110000",
  47367=>"000100110",
  47368=>"011111101",
  47369=>"111100011",
  47370=>"010000101",
  47371=>"111010100",
  47372=>"111111001",
  47373=>"001011000",
  47374=>"011110011",
  47375=>"010101010",
  47376=>"011100101",
  47377=>"110111001",
  47378=>"110000101",
  47379=>"111111111",
  47380=>"110101111",
  47381=>"100011111",
  47382=>"000100001",
  47383=>"110011101",
  47384=>"101010000",
  47385=>"001001000",
  47386=>"010000101",
  47387=>"010000000",
  47388=>"011111011",
  47389=>"110010111",
  47390=>"101110110",
  47391=>"000100000",
  47392=>"100101101",
  47393=>"110001000",
  47394=>"010100100",
  47395=>"110010000",
  47396=>"101010011",
  47397=>"011101101",
  47398=>"010110111",
  47399=>"011010111",
  47400=>"000000000",
  47401=>"100110100",
  47402=>"101001000",
  47403=>"000001110",
  47404=>"100010101",
  47405=>"000010100",
  47406=>"100010010",
  47407=>"010011011",
  47408=>"010010010",
  47409=>"010000000",
  47410=>"010011000",
  47411=>"011010001",
  47412=>"101111100",
  47413=>"000000101",
  47414=>"101010110",
  47415=>"110111101",
  47416=>"000001011",
  47417=>"011101110",
  47418=>"110000101",
  47419=>"011111000",
  47420=>"000000100",
  47421=>"110011011",
  47422=>"000100100",
  47423=>"111011111",
  47424=>"111111010",
  47425=>"111111110",
  47426=>"110101000",
  47427=>"010101000",
  47428=>"101100010",
  47429=>"011101101",
  47430=>"100000001",
  47431=>"100111011",
  47432=>"010001110",
  47433=>"010010111",
  47434=>"001110011",
  47435=>"010000111",
  47436=>"000000001",
  47437=>"001000000",
  47438=>"001010111",
  47439=>"001100011",
  47440=>"110100011",
  47441=>"011011001",
  47442=>"101101000",
  47443=>"000110010",
  47444=>"110000010",
  47445=>"110111111",
  47446=>"101100000",
  47447=>"000100111",
  47448=>"000100000",
  47449=>"100111010",
  47450=>"011000011",
  47451=>"000011011",
  47452=>"001100001",
  47453=>"000010000",
  47454=>"001011010",
  47455=>"000011111",
  47456=>"111100000",
  47457=>"001010101",
  47458=>"011000101",
  47459=>"000000010",
  47460=>"101110110",
  47461=>"100111000",
  47462=>"110101110",
  47463=>"010100000",
  47464=>"001011101",
  47465=>"011011100",
  47466=>"001000111",
  47467=>"100100111",
  47468=>"000000010",
  47469=>"110100011",
  47470=>"101101100",
  47471=>"010001001",
  47472=>"000000100",
  47473=>"111000001",
  47474=>"101001000",
  47475=>"110000011",
  47476=>"010001011",
  47477=>"010000011",
  47478=>"011011111",
  47479=>"001100001",
  47480=>"000000111",
  47481=>"010110101",
  47482=>"011111111",
  47483=>"110101111",
  47484=>"100001100",
  47485=>"011100001",
  47486=>"011110001",
  47487=>"010110100",
  47488=>"100000001",
  47489=>"001000111",
  47490=>"010111111",
  47491=>"011110010",
  47492=>"111100011",
  47493=>"100111001",
  47494=>"110110110",
  47495=>"110010111",
  47496=>"110111101",
  47497=>"100111111",
  47498=>"110000011",
  47499=>"000000000",
  47500=>"111001011",
  47501=>"000111100",
  47502=>"000100000",
  47503=>"000100110",
  47504=>"100000000",
  47505=>"000100000",
  47506=>"110011011",
  47507=>"010100100",
  47508=>"001011011",
  47509=>"010001100",
  47510=>"000111101",
  47511=>"110001111",
  47512=>"111110101",
  47513=>"110011110",
  47514=>"101111101",
  47515=>"000011111",
  47516=>"001111100",
  47517=>"011011001",
  47518=>"010000010",
  47519=>"011111101",
  47520=>"110000011",
  47521=>"010101000",
  47522=>"111111010",
  47523=>"010010000",
  47524=>"000000100",
  47525=>"011000010",
  47526=>"111101011",
  47527=>"111000100",
  47528=>"001110000",
  47529=>"110000100",
  47530=>"000101101",
  47531=>"100011100",
  47532=>"010110110",
  47533=>"101111100",
  47534=>"000011100",
  47535=>"101100011",
  47536=>"011100101",
  47537=>"000011111",
  47538=>"011101011",
  47539=>"011010011",
  47540=>"001001100",
  47541=>"000111000",
  47542=>"101111001",
  47543=>"100100111",
  47544=>"100110011",
  47545=>"000000010",
  47546=>"100001110",
  47547=>"101011011",
  47548=>"111100100",
  47549=>"001110000",
  47550=>"111101000",
  47551=>"011001101",
  47552=>"010001011",
  47553=>"001000000",
  47554=>"110010010",
  47555=>"111110100",
  47556=>"000011001",
  47557=>"101010100",
  47558=>"000001011",
  47559=>"011100000",
  47560=>"110110111",
  47561=>"001110110",
  47562=>"001000111",
  47563=>"001011010",
  47564=>"000010000",
  47565=>"011001000",
  47566=>"100100010",
  47567=>"111000111",
  47568=>"010101110",
  47569=>"000110000",
  47570=>"110110111",
  47571=>"110111100",
  47572=>"101111111",
  47573=>"000011110",
  47574=>"110001011",
  47575=>"011001010",
  47576=>"011110110",
  47577=>"101100101",
  47578=>"111010100",
  47579=>"100110001",
  47580=>"111111010",
  47581=>"100100000",
  47582=>"000111000",
  47583=>"001010100",
  47584=>"100100000",
  47585=>"000110010",
  47586=>"111001000",
  47587=>"001010100",
  47588=>"111001000",
  47589=>"101001101",
  47590=>"101000011",
  47591=>"000000111",
  47592=>"011111111",
  47593=>"010001101",
  47594=>"010101000",
  47595=>"001101000",
  47596=>"010101000",
  47597=>"000000101",
  47598=>"100000101",
  47599=>"101001000",
  47600=>"010001110",
  47601=>"100101101",
  47602=>"000111100",
  47603=>"111111001",
  47604=>"110011001",
  47605=>"100100101",
  47606=>"111100110",
  47607=>"010010111",
  47608=>"100000001",
  47609=>"111011001",
  47610=>"101111000",
  47611=>"000011001",
  47612=>"011101010",
  47613=>"000000111",
  47614=>"100011111",
  47615=>"011110111",
  47616=>"001000000",
  47617=>"000000101",
  47618=>"111011110",
  47619=>"000110110",
  47620=>"111100110",
  47621=>"011011000",
  47622=>"111111011",
  47623=>"100100001",
  47624=>"100001101",
  47625=>"110001101",
  47626=>"101000101",
  47627=>"011101100",
  47628=>"110101100",
  47629=>"110110001",
  47630=>"101001001",
  47631=>"010011001",
  47632=>"000010001",
  47633=>"111101110",
  47634=>"000000111",
  47635=>"100101110",
  47636=>"100101010",
  47637=>"011011001",
  47638=>"110011100",
  47639=>"101000000",
  47640=>"010011111",
  47641=>"001011000",
  47642=>"001011011",
  47643=>"000100101",
  47644=>"001110000",
  47645=>"000010000",
  47646=>"100011111",
  47647=>"110110110",
  47648=>"001011101",
  47649=>"000011000",
  47650=>"000101101",
  47651=>"011011101",
  47652=>"011001011",
  47653=>"010110101",
  47654=>"111110000",
  47655=>"010110010",
  47656=>"000101000",
  47657=>"011110000",
  47658=>"101101000",
  47659=>"001011010",
  47660=>"000110111",
  47661=>"001010011",
  47662=>"100000111",
  47663=>"100111111",
  47664=>"001101111",
  47665=>"001101100",
  47666=>"100011100",
  47667=>"100011110",
  47668=>"001000000",
  47669=>"000010000",
  47670=>"000000111",
  47671=>"010001011",
  47672=>"001001101",
  47673=>"010001110",
  47674=>"101001001",
  47675=>"011101000",
  47676=>"000001101",
  47677=>"011011000",
  47678=>"111010000",
  47679=>"011011110",
  47680=>"000000111",
  47681=>"110101010",
  47682=>"101000111",
  47683=>"001100111",
  47684=>"000011000",
  47685=>"110010101",
  47686=>"110100000",
  47687=>"111010111",
  47688=>"000110110",
  47689=>"111110100",
  47690=>"110011110",
  47691=>"100100011",
  47692=>"011111100",
  47693=>"001101100",
  47694=>"110100011",
  47695=>"011001000",
  47696=>"111001011",
  47697=>"111001001",
  47698=>"101110111",
  47699=>"010101111",
  47700=>"011000111",
  47701=>"100100100",
  47702=>"000001000",
  47703=>"011100000",
  47704=>"011101011",
  47705=>"111111101",
  47706=>"100100101",
  47707=>"010011010",
  47708=>"011000100",
  47709=>"100010110",
  47710=>"101110011",
  47711=>"011000101",
  47712=>"111000001",
  47713=>"010110000",
  47714=>"111110111",
  47715=>"001001100",
  47716=>"011111011",
  47717=>"101011100",
  47718=>"001100110",
  47719=>"111010110",
  47720=>"010110111",
  47721=>"010100011",
  47722=>"010111111",
  47723=>"110110110",
  47724=>"010001001",
  47725=>"101001100",
  47726=>"110001101",
  47727=>"101100011",
  47728=>"110100010",
  47729=>"011110101",
  47730=>"110011000",
  47731=>"110111100",
  47732=>"010100011",
  47733=>"111111000",
  47734=>"000111100",
  47735=>"110010000",
  47736=>"010010011",
  47737=>"111001010",
  47738=>"011010110",
  47739=>"000010110",
  47740=>"111111101",
  47741=>"001000111",
  47742=>"011011100",
  47743=>"100111111",
  47744=>"001010110",
  47745=>"011011101",
  47746=>"010110110",
  47747=>"101000000",
  47748=>"100111111",
  47749=>"000011001",
  47750=>"000010001",
  47751=>"001011110",
  47752=>"001010010",
  47753=>"111101111",
  47754=>"011000111",
  47755=>"101101011",
  47756=>"110110001",
  47757=>"000111010",
  47758=>"011001110",
  47759=>"101010111",
  47760=>"000000011",
  47761=>"101101011",
  47762=>"010011011",
  47763=>"010010101",
  47764=>"110101000",
  47765=>"011111000",
  47766=>"110011010",
  47767=>"100000101",
  47768=>"110111111",
  47769=>"011100111",
  47770=>"101110001",
  47771=>"101011101",
  47772=>"000101000",
  47773=>"101011101",
  47774=>"000110100",
  47775=>"111001110",
  47776=>"101101010",
  47777=>"000010001",
  47778=>"100101111",
  47779=>"001110000",
  47780=>"111101000",
  47781=>"000100110",
  47782=>"100111000",
  47783=>"001101101",
  47784=>"110111001",
  47785=>"001011101",
  47786=>"101000001",
  47787=>"111100011",
  47788=>"110110001",
  47789=>"000111111",
  47790=>"111111101",
  47791=>"100100010",
  47792=>"001001000",
  47793=>"011111000",
  47794=>"111111111",
  47795=>"111000000",
  47796=>"010110111",
  47797=>"110010111",
  47798=>"001000001",
  47799=>"010101001",
  47800=>"010000110",
  47801=>"111000010",
  47802=>"101000101",
  47803=>"101110000",
  47804=>"011100010",
  47805=>"001111111",
  47806=>"010100010",
  47807=>"110101010",
  47808=>"011111001",
  47809=>"010011101",
  47810=>"111011111",
  47811=>"010000010",
  47812=>"001000100",
  47813=>"001000001",
  47814=>"100011000",
  47815=>"111001111",
  47816=>"110000110",
  47817=>"011110100",
  47818=>"111101110",
  47819=>"001000001",
  47820=>"110010010",
  47821=>"010100000",
  47822=>"110101100",
  47823=>"000000010",
  47824=>"111101010",
  47825=>"000100100",
  47826=>"111100000",
  47827=>"001001011",
  47828=>"010001111",
  47829=>"011101111",
  47830=>"000000011",
  47831=>"000110010",
  47832=>"101111011",
  47833=>"111101010",
  47834=>"000101001",
  47835=>"001001010",
  47836=>"110001101",
  47837=>"110110110",
  47838=>"011010100",
  47839=>"101001011",
  47840=>"010000110",
  47841=>"001010100",
  47842=>"010011010",
  47843=>"001010111",
  47844=>"110010100",
  47845=>"010010001",
  47846=>"011010111",
  47847=>"011110110",
  47848=>"100100100",
  47849=>"011111111",
  47850=>"111110011",
  47851=>"010000101",
  47852=>"010001001",
  47853=>"111011001",
  47854=>"000110000",
  47855=>"011001100",
  47856=>"100100010",
  47857=>"110001001",
  47858=>"000101010",
  47859=>"101100100",
  47860=>"011011111",
  47861=>"111011011",
  47862=>"000100010",
  47863=>"011101001",
  47864=>"101100110",
  47865=>"011011000",
  47866=>"111011001",
  47867=>"100100001",
  47868=>"000001111",
  47869=>"100101111",
  47870=>"011001000",
  47871=>"001101000",
  47872=>"101110110",
  47873=>"000111110",
  47874=>"001010100",
  47875=>"101101100",
  47876=>"110111110",
  47877=>"100100010",
  47878=>"110101000",
  47879=>"000101111",
  47880=>"100011010",
  47881=>"000010011",
  47882=>"001001001",
  47883=>"000100010",
  47884=>"000000100",
  47885=>"111011110",
  47886=>"100100001",
  47887=>"101001011",
  47888=>"101110110",
  47889=>"011001100",
  47890=>"000100111",
  47891=>"000110100",
  47892=>"010001010",
  47893=>"001010001",
  47894=>"110000111",
  47895=>"010100101",
  47896=>"100100111",
  47897=>"010111100",
  47898=>"011101111",
  47899=>"110000100",
  47900=>"110011011",
  47901=>"011010011",
  47902=>"010111110",
  47903=>"011100001",
  47904=>"010101000",
  47905=>"110010111",
  47906=>"100100000",
  47907=>"001001100",
  47908=>"100010100",
  47909=>"111110000",
  47910=>"010100111",
  47911=>"011000010",
  47912=>"111101010",
  47913=>"101000001",
  47914=>"110100111",
  47915=>"100010000",
  47916=>"010001101",
  47917=>"111111100",
  47918=>"010010101",
  47919=>"110110010",
  47920=>"101000000",
  47921=>"000010010",
  47922=>"100010111",
  47923=>"001111001",
  47924=>"001000111",
  47925=>"011000110",
  47926=>"101100101",
  47927=>"111110111",
  47928=>"100110101",
  47929=>"010111100",
  47930=>"100001110",
  47931=>"000100001",
  47932=>"111011001",
  47933=>"100000110",
  47934=>"000110001",
  47935=>"011101101",
  47936=>"101000010",
  47937=>"100011010",
  47938=>"111001001",
  47939=>"000111110",
  47940=>"100011110",
  47941=>"101111100",
  47942=>"100100100",
  47943=>"111010011",
  47944=>"001111111",
  47945=>"011100111",
  47946=>"011011010",
  47947=>"011000111",
  47948=>"101010000",
  47949=>"100010011",
  47950=>"100100000",
  47951=>"101110001",
  47952=>"100001010",
  47953=>"110110101",
  47954=>"100011111",
  47955=>"101111111",
  47956=>"000110000",
  47957=>"100000100",
  47958=>"000100111",
  47959=>"010110000",
  47960=>"010101110",
  47961=>"011111110",
  47962=>"110010000",
  47963=>"110110011",
  47964=>"011111001",
  47965=>"011000001",
  47966=>"011110101",
  47967=>"011110011",
  47968=>"010001111",
  47969=>"011001110",
  47970=>"111110010",
  47971=>"011001001",
  47972=>"001100001",
  47973=>"010010101",
  47974=>"010010100",
  47975=>"011011001",
  47976=>"010011101",
  47977=>"101101000",
  47978=>"100011110",
  47979=>"111000101",
  47980=>"011110110",
  47981=>"001110001",
  47982=>"110000000",
  47983=>"110100100",
  47984=>"111101101",
  47985=>"001100001",
  47986=>"001010101",
  47987=>"101111111",
  47988=>"110111010",
  47989=>"110101101",
  47990=>"001000100",
  47991=>"011110011",
  47992=>"101110100",
  47993=>"101010010",
  47994=>"100011110",
  47995=>"110100000",
  47996=>"000011100",
  47997=>"100101000",
  47998=>"110011100",
  47999=>"111011110",
  48000=>"100001001",
  48001=>"000100101",
  48002=>"110110111",
  48003=>"011100101",
  48004=>"011010000",
  48005=>"001111011",
  48006=>"010110100",
  48007=>"101100110",
  48008=>"111011111",
  48009=>"110000111",
  48010=>"100100111",
  48011=>"100001101",
  48012=>"100000100",
  48013=>"100111111",
  48014=>"101100001",
  48015=>"000100011",
  48016=>"001001011",
  48017=>"110111100",
  48018=>"000110100",
  48019=>"010000101",
  48020=>"111010000",
  48021=>"000110011",
  48022=>"010111000",
  48023=>"011100101",
  48024=>"010000110",
  48025=>"101110100",
  48026=>"100011111",
  48027=>"011011011",
  48028=>"100100111",
  48029=>"010011000",
  48030=>"110100001",
  48031=>"011000000",
  48032=>"010010100",
  48033=>"000100110",
  48034=>"100101100",
  48035=>"010100010",
  48036=>"100101011",
  48037=>"001011100",
  48038=>"101111000",
  48039=>"100101001",
  48040=>"101110001",
  48041=>"000110110",
  48042=>"000111110",
  48043=>"110011101",
  48044=>"111111111",
  48045=>"001011100",
  48046=>"111111010",
  48047=>"000101001",
  48048=>"000101100",
  48049=>"110110101",
  48050=>"011110111",
  48051=>"110100010",
  48052=>"111001101",
  48053=>"111000111",
  48054=>"011000001",
  48055=>"110000001",
  48056=>"111000110",
  48057=>"010011110",
  48058=>"000111010",
  48059=>"111010101",
  48060=>"011100101",
  48061=>"110110010",
  48062=>"101011100",
  48063=>"011101110",
  48064=>"000010111",
  48065=>"110110110",
  48066=>"000110010",
  48067=>"101010010",
  48068=>"101000010",
  48069=>"111010111",
  48070=>"111110101",
  48071=>"011111111",
  48072=>"000000001",
  48073=>"010011110",
  48074=>"100110010",
  48075=>"101100010",
  48076=>"001011110",
  48077=>"100001110",
  48078=>"101101110",
  48079=>"111011101",
  48080=>"010100110",
  48081=>"100110111",
  48082=>"101111011",
  48083=>"011001000",
  48084=>"011101001",
  48085=>"000100110",
  48086=>"001001001",
  48087=>"001111111",
  48088=>"111000000",
  48089=>"010000011",
  48090=>"011010101",
  48091=>"111010110",
  48092=>"001011000",
  48093=>"111011000",
  48094=>"110110011",
  48095=>"001101010",
  48096=>"001001011",
  48097=>"000000101",
  48098=>"000001100",
  48099=>"010001101",
  48100=>"010101010",
  48101=>"100001000",
  48102=>"111010011",
  48103=>"000100111",
  48104=>"100100000",
  48105=>"100110011",
  48106=>"100000101",
  48107=>"010111101",
  48108=>"011011111",
  48109=>"101110010",
  48110=>"101110101",
  48111=>"000001110",
  48112=>"100100010",
  48113=>"001101111",
  48114=>"101110001",
  48115=>"001101110",
  48116=>"101110011",
  48117=>"010110111",
  48118=>"111110110",
  48119=>"101111010",
  48120=>"111000101",
  48121=>"010110101",
  48122=>"110101111",
  48123=>"000000111",
  48124=>"010100011",
  48125=>"010000110",
  48126=>"001000010",
  48127=>"011100001",
  48128=>"111110101",
  48129=>"110000001",
  48130=>"011000101",
  48131=>"111011110",
  48132=>"010111110",
  48133=>"001100111",
  48134=>"111000111",
  48135=>"001001000",
  48136=>"010110100",
  48137=>"000101001",
  48138=>"000100011",
  48139=>"100101010",
  48140=>"010111000",
  48141=>"001011011",
  48142=>"100101000",
  48143=>"000001111",
  48144=>"100111011",
  48145=>"011110000",
  48146=>"010100111",
  48147=>"101111100",
  48148=>"110101111",
  48149=>"100000100",
  48150=>"011010101",
  48151=>"000000011",
  48152=>"011111110",
  48153=>"000000001",
  48154=>"010100000",
  48155=>"010011100",
  48156=>"100011011",
  48157=>"111011010",
  48158=>"110101101",
  48159=>"100110101",
  48160=>"011001010",
  48161=>"000010110",
  48162=>"111001011",
  48163=>"111100000",
  48164=>"100000110",
  48165=>"101000100",
  48166=>"110011011",
  48167=>"101011101",
  48168=>"110011011",
  48169=>"010100101",
  48170=>"111001101",
  48171=>"111011111",
  48172=>"110101010",
  48173=>"011000110",
  48174=>"111000001",
  48175=>"100010110",
  48176=>"111111011",
  48177=>"000110000",
  48178=>"001101100",
  48179=>"101000100",
  48180=>"101110100",
  48181=>"001001001",
  48182=>"000110101",
  48183=>"000010100",
  48184=>"010001101",
  48185=>"110100110",
  48186=>"110110111",
  48187=>"101110001",
  48188=>"111100111",
  48189=>"111100101",
  48190=>"111010001",
  48191=>"101000011",
  48192=>"111000001",
  48193=>"111000001",
  48194=>"100011000",
  48195=>"100101110",
  48196=>"010000101",
  48197=>"100100010",
  48198=>"011010100",
  48199=>"010011100",
  48200=>"111111111",
  48201=>"000100011",
  48202=>"011100000",
  48203=>"011010100",
  48204=>"001001110",
  48205=>"101111011",
  48206=>"110011101",
  48207=>"011101010",
  48208=>"110110101",
  48209=>"000110000",
  48210=>"000111100",
  48211=>"011101110",
  48212=>"100101001",
  48213=>"001001010",
  48214=>"111110011",
  48215=>"110100001",
  48216=>"100011101",
  48217=>"101000110",
  48218=>"010000100",
  48219=>"111011010",
  48220=>"010010010",
  48221=>"011111100",
  48222=>"000000001",
  48223=>"011100111",
  48224=>"111100100",
  48225=>"001001000",
  48226=>"011000100",
  48227=>"001101001",
  48228=>"111000010",
  48229=>"011111011",
  48230=>"010011011",
  48231=>"101001010",
  48232=>"111111101",
  48233=>"000001011",
  48234=>"110111011",
  48235=>"000001001",
  48236=>"010100101",
  48237=>"101101100",
  48238=>"010100000",
  48239=>"010110010",
  48240=>"101111001",
  48241=>"110000000",
  48242=>"001001111",
  48243=>"000110010",
  48244=>"110100110",
  48245=>"000111011",
  48246=>"110001111",
  48247=>"111011011",
  48248=>"001101011",
  48249=>"101110110",
  48250=>"100100100",
  48251=>"011000111",
  48252=>"110111001",
  48253=>"110010100",
  48254=>"110000100",
  48255=>"110010111",
  48256=>"011101010",
  48257=>"000100000",
  48258=>"110010001",
  48259=>"000010111",
  48260=>"011111110",
  48261=>"000100101",
  48262=>"010100001",
  48263=>"100111001",
  48264=>"111101110",
  48265=>"101110111",
  48266=>"100010111",
  48267=>"101101001",
  48268=>"010011100",
  48269=>"011011001",
  48270=>"001101111",
  48271=>"011000011",
  48272=>"100010011",
  48273=>"010101111",
  48274=>"010100100",
  48275=>"101101000",
  48276=>"000001000",
  48277=>"110001001",
  48278=>"011100100",
  48279=>"000101110",
  48280=>"011010001",
  48281=>"010001110",
  48282=>"011011100",
  48283=>"111001110",
  48284=>"101100100",
  48285=>"110101111",
  48286=>"011110010",
  48287=>"010101011",
  48288=>"010001100",
  48289=>"011101110",
  48290=>"011110100",
  48291=>"011000111",
  48292=>"111111111",
  48293=>"001100011",
  48294=>"010100011",
  48295=>"100111101",
  48296=>"000000001",
  48297=>"000010000",
  48298=>"110010100",
  48299=>"101101110",
  48300=>"011101100",
  48301=>"101001011",
  48302=>"110100111",
  48303=>"111101101",
  48304=>"001101101",
  48305=>"010001010",
  48306=>"100111011",
  48307=>"100111101",
  48308=>"100111011",
  48309=>"001011001",
  48310=>"001000111",
  48311=>"001101010",
  48312=>"101000110",
  48313=>"101001011",
  48314=>"101101001",
  48315=>"101011000",
  48316=>"001011010",
  48317=>"101110000",
  48318=>"110100100",
  48319=>"111110001",
  48320=>"000011010",
  48321=>"111100001",
  48322=>"110001010",
  48323=>"000001111",
  48324=>"001111010",
  48325=>"100000110",
  48326=>"010100000",
  48327=>"110000010",
  48328=>"111110011",
  48329=>"000010100",
  48330=>"110100000",
  48331=>"100101110",
  48332=>"110010000",
  48333=>"110101101",
  48334=>"110000000",
  48335=>"010001111",
  48336=>"110100010",
  48337=>"011100101",
  48338=>"011110101",
  48339=>"110110011",
  48340=>"001100000",
  48341=>"101000100",
  48342=>"000010010",
  48343=>"111010100",
  48344=>"111001111",
  48345=>"010010110",
  48346=>"001000000",
  48347=>"001100100",
  48348=>"001000000",
  48349=>"110111010",
  48350=>"101000100",
  48351=>"010001010",
  48352=>"000001110",
  48353=>"000100100",
  48354=>"100010101",
  48355=>"100110001",
  48356=>"001000101",
  48357=>"000000111",
  48358=>"100100101",
  48359=>"000010001",
  48360=>"110000011",
  48361=>"100111100",
  48362=>"001111000",
  48363=>"110000100",
  48364=>"010011110",
  48365=>"100100001",
  48366=>"100011001",
  48367=>"110001001",
  48368=>"010001110",
  48369=>"100101101",
  48370=>"000011001",
  48371=>"000111001",
  48372=>"111111010",
  48373=>"111101100",
  48374=>"101000101",
  48375=>"100001000",
  48376=>"000001101",
  48377=>"010110001",
  48378=>"011001010",
  48379=>"001000000",
  48380=>"101001010",
  48381=>"110101001",
  48382=>"111011001",
  48383=>"010110111",
  48384=>"001101011",
  48385=>"110010101",
  48386=>"001011010",
  48387=>"000110101",
  48388=>"101110110",
  48389=>"110001000",
  48390=>"011000101",
  48391=>"101011100",
  48392=>"100101000",
  48393=>"100000011",
  48394=>"010111110",
  48395=>"111111001",
  48396=>"100000111",
  48397=>"111100001",
  48398=>"101100100",
  48399=>"001110011",
  48400=>"100100111",
  48401=>"010100100",
  48402=>"001010101",
  48403=>"010100000",
  48404=>"000011111",
  48405=>"101011011",
  48406=>"010111111",
  48407=>"010001011",
  48408=>"000110110",
  48409=>"010000001",
  48410=>"000000011",
  48411=>"110001110",
  48412=>"110000010",
  48413=>"101000001",
  48414=>"111110100",
  48415=>"010000110",
  48416=>"001000011",
  48417=>"110110001",
  48418=>"110001110",
  48419=>"110010001",
  48420=>"111100000",
  48421=>"010001001",
  48422=>"000000001",
  48423=>"111010011",
  48424=>"111110100",
  48425=>"101111011",
  48426=>"000101111",
  48427=>"010101011",
  48428=>"111000100",
  48429=>"100110110",
  48430=>"000101000",
  48431=>"110111010",
  48432=>"010110100",
  48433=>"101011111",
  48434=>"011111111",
  48435=>"010000110",
  48436=>"011001011",
  48437=>"100010000",
  48438=>"011111001",
  48439=>"111011100",
  48440=>"101000001",
  48441=>"110001111",
  48442=>"100100110",
  48443=>"110000111",
  48444=>"000000010",
  48445=>"010100111",
  48446=>"010011111",
  48447=>"011100001",
  48448=>"010011111",
  48449=>"011010110",
  48450=>"101001101",
  48451=>"001101011",
  48452=>"100111001",
  48453=>"110100100",
  48454=>"000101101",
  48455=>"111111100",
  48456=>"000011011",
  48457=>"100000101",
  48458=>"000001100",
  48459=>"000111100",
  48460=>"111100101",
  48461=>"111010111",
  48462=>"011100110",
  48463=>"010101011",
  48464=>"111000100",
  48465=>"101101111",
  48466=>"000111100",
  48467=>"110001110",
  48468=>"011011000",
  48469=>"110001101",
  48470=>"110100111",
  48471=>"101000101",
  48472=>"000111001",
  48473=>"101101100",
  48474=>"000110111",
  48475=>"111100100",
  48476=>"100000011",
  48477=>"110110000",
  48478=>"110011010",
  48479=>"010000000",
  48480=>"110101101",
  48481=>"011001110",
  48482=>"110110101",
  48483=>"010001100",
  48484=>"001000111",
  48485=>"100100010",
  48486=>"110111100",
  48487=>"100110111",
  48488=>"010101001",
  48489=>"101010100",
  48490=>"001011110",
  48491=>"010111010",
  48492=>"111101011",
  48493=>"110001100",
  48494=>"110000000",
  48495=>"000100000",
  48496=>"000100000",
  48497=>"100001000",
  48498=>"111010100",
  48499=>"111010011",
  48500=>"010110110",
  48501=>"000110110",
  48502=>"111110111",
  48503=>"100000001",
  48504=>"001111011",
  48505=>"001011111",
  48506=>"001111010",
  48507=>"100110011",
  48508=>"010101110",
  48509=>"010010010",
  48510=>"010000101",
  48511=>"110110010",
  48512=>"000100100",
  48513=>"001111111",
  48514=>"001001100",
  48515=>"100011111",
  48516=>"000111010",
  48517=>"100001011",
  48518=>"100011111",
  48519=>"001000110",
  48520=>"101110111",
  48521=>"000010100",
  48522=>"000001001",
  48523=>"001010000",
  48524=>"000111011",
  48525=>"101000001",
  48526=>"010111000",
  48527=>"100000101",
  48528=>"001000001",
  48529=>"101000100",
  48530=>"010010101",
  48531=>"010000011",
  48532=>"011100110",
  48533=>"001000110",
  48534=>"110010000",
  48535=>"111011001",
  48536=>"101010101",
  48537=>"000101011",
  48538=>"010111100",
  48539=>"011011110",
  48540=>"111101110",
  48541=>"111101100",
  48542=>"011000000",
  48543=>"010101011",
  48544=>"111001001",
  48545=>"010000000",
  48546=>"111111010",
  48547=>"000100111",
  48548=>"011011001",
  48549=>"011100000",
  48550=>"111111111",
  48551=>"011101101",
  48552=>"110101010",
  48553=>"010101010",
  48554=>"000000100",
  48555=>"011000101",
  48556=>"000110000",
  48557=>"111111000",
  48558=>"100001011",
  48559=>"111000011",
  48560=>"110111100",
  48561=>"111110111",
  48562=>"110001000",
  48563=>"001001011",
  48564=>"110010000",
  48565=>"001111000",
  48566=>"100110110",
  48567=>"100100100",
  48568=>"111011001",
  48569=>"010001100",
  48570=>"000010111",
  48571=>"011110101",
  48572=>"110110111",
  48573=>"111011001",
  48574=>"101001011",
  48575=>"011000011",
  48576=>"111001100",
  48577=>"110000111",
  48578=>"011000100",
  48579=>"010001101",
  48580=>"000011101",
  48581=>"111000100",
  48582=>"100001000",
  48583=>"101000000",
  48584=>"010001111",
  48585=>"100000110",
  48586=>"011000101",
  48587=>"010001100",
  48588=>"000001000",
  48589=>"111001110",
  48590=>"110000110",
  48591=>"101110010",
  48592=>"101011011",
  48593=>"011001101",
  48594=>"001111110",
  48595=>"110011111",
  48596=>"000000100",
  48597=>"001111000",
  48598=>"110001000",
  48599=>"000100000",
  48600=>"001110001",
  48601=>"111111011",
  48602=>"100001011",
  48603=>"111000011",
  48604=>"000111110",
  48605=>"011011111",
  48606=>"001110100",
  48607=>"100101101",
  48608=>"000100011",
  48609=>"100111011",
  48610=>"111010101",
  48611=>"001010111",
  48612=>"110110111",
  48613=>"010000101",
  48614=>"111000010",
  48615=>"001101010",
  48616=>"100011110",
  48617=>"100000011",
  48618=>"110101001",
  48619=>"111110111",
  48620=>"101100100",
  48621=>"010100010",
  48622=>"111011101",
  48623=>"100101001",
  48624=>"010100100",
  48625=>"001111011",
  48626=>"110110111",
  48627=>"101001001",
  48628=>"101100111",
  48629=>"111110100",
  48630=>"101110000",
  48631=>"010011011",
  48632=>"111001100",
  48633=>"011111001",
  48634=>"010000111",
  48635=>"000000101",
  48636=>"001101000",
  48637=>"001111010",
  48638=>"001101101",
  48639=>"110011001",
  48640=>"010101101",
  48641=>"000001001",
  48642=>"110111000",
  48643=>"111011001",
  48644=>"011111110",
  48645=>"111000000",
  48646=>"110111101",
  48647=>"101000000",
  48648=>"011001110",
  48649=>"011000100",
  48650=>"000001011",
  48651=>"011001100",
  48652=>"001110001",
  48653=>"101111000",
  48654=>"100010010",
  48655=>"111100010",
  48656=>"100010100",
  48657=>"110100000",
  48658=>"110000110",
  48659=>"000010101",
  48660=>"010001001",
  48661=>"110001101",
  48662=>"101111110",
  48663=>"010010001",
  48664=>"101101110",
  48665=>"000011110",
  48666=>"110010011",
  48667=>"011010110",
  48668=>"100110001",
  48669=>"101010001",
  48670=>"000010010",
  48671=>"010111001",
  48672=>"001001101",
  48673=>"111100010",
  48674=>"110000001",
  48675=>"001000100",
  48676=>"101111101",
  48677=>"100110110",
  48678=>"101011010",
  48679=>"111011000",
  48680=>"111000100",
  48681=>"110000011",
  48682=>"001011011",
  48683=>"110101010",
  48684=>"110000100",
  48685=>"110100111",
  48686=>"011001100",
  48687=>"101000011",
  48688=>"001101011",
  48689=>"010110101",
  48690=>"001111111",
  48691=>"001110110",
  48692=>"110000100",
  48693=>"010000010",
  48694=>"101101000",
  48695=>"010000110",
  48696=>"000010110",
  48697=>"100010011",
  48698=>"000111010",
  48699=>"001001110",
  48700=>"100000000",
  48701=>"000010010",
  48702=>"011000011",
  48703=>"111001000",
  48704=>"101100000",
  48705=>"110000010",
  48706=>"011000011",
  48707=>"101111111",
  48708=>"000101010",
  48709=>"011000001",
  48710=>"111001001",
  48711=>"110001001",
  48712=>"000000010",
  48713=>"101110010",
  48714=>"001111111",
  48715=>"000110001",
  48716=>"101110011",
  48717=>"011101101",
  48718=>"011011000",
  48719=>"111101011",
  48720=>"100010000",
  48721=>"000001000",
  48722=>"010111101",
  48723=>"011000000",
  48724=>"000010010",
  48725=>"111000010",
  48726=>"001010011",
  48727=>"001010000",
  48728=>"010111111",
  48729=>"101100011",
  48730=>"101000101",
  48731=>"001011001",
  48732=>"111110011",
  48733=>"010000010",
  48734=>"000000011",
  48735=>"110001110",
  48736=>"011101000",
  48737=>"101100000",
  48738=>"011011110",
  48739=>"010110110",
  48740=>"111111111",
  48741=>"000010011",
  48742=>"100010011",
  48743=>"100000111",
  48744=>"111011001",
  48745=>"000001001",
  48746=>"010000100",
  48747=>"100110001",
  48748=>"000100110",
  48749=>"101111010",
  48750=>"001100000",
  48751=>"000010001",
  48752=>"101001110",
  48753=>"000001011",
  48754=>"011000011",
  48755=>"010000110",
  48756=>"010110111",
  48757=>"010010000",
  48758=>"110100101",
  48759=>"011110110",
  48760=>"010010010",
  48761=>"110011100",
  48762=>"111110000",
  48763=>"100110010",
  48764=>"000011000",
  48765=>"011000100",
  48766=>"011110001",
  48767=>"100110100",
  48768=>"110000011",
  48769=>"000110001",
  48770=>"000110010",
  48771=>"000010100",
  48772=>"101100001",
  48773=>"110000000",
  48774=>"100011001",
  48775=>"001101111",
  48776=>"001010001",
  48777=>"101000010",
  48778=>"001111010",
  48779=>"101100001",
  48780=>"011000000",
  48781=>"100000110",
  48782=>"111111100",
  48783=>"101110001",
  48784=>"010111001",
  48785=>"111100001",
  48786=>"111010101",
  48787=>"100110111",
  48788=>"000001100",
  48789=>"000101110",
  48790=>"100111100",
  48791=>"101110111",
  48792=>"111010100",
  48793=>"011001101",
  48794=>"011011110",
  48795=>"000001000",
  48796=>"011011000",
  48797=>"110110111",
  48798=>"010001000",
  48799=>"010001011",
  48800=>"101110111",
  48801=>"101111100",
  48802=>"110111000",
  48803=>"101111010",
  48804=>"100110100",
  48805=>"000000000",
  48806=>"000101011",
  48807=>"001111101",
  48808=>"000001101",
  48809=>"000000110",
  48810=>"010100100",
  48811=>"101101100",
  48812=>"001010011",
  48813=>"100010010",
  48814=>"101111000",
  48815=>"000001110",
  48816=>"100000101",
  48817=>"100000101",
  48818=>"111111001",
  48819=>"010011101",
  48820=>"110111111",
  48821=>"010101110",
  48822=>"000110011",
  48823=>"011111101",
  48824=>"111100110",
  48825=>"010111010",
  48826=>"001101100",
  48827=>"110100011",
  48828=>"011010000",
  48829=>"100110111",
  48830=>"011101000",
  48831=>"000001111",
  48832=>"110000000",
  48833=>"101010001",
  48834=>"001010111",
  48835=>"101001001",
  48836=>"110100111",
  48837=>"111110101",
  48838=>"101011011",
  48839=>"000010100",
  48840=>"101101011",
  48841=>"010110001",
  48842=>"100111000",
  48843=>"001010010",
  48844=>"010111111",
  48845=>"101111011",
  48846=>"111000111",
  48847=>"110001001",
  48848=>"011111111",
  48849=>"110000000",
  48850=>"001101110",
  48851=>"110010011",
  48852=>"000010101",
  48853=>"100000001",
  48854=>"110111101",
  48855=>"110101001",
  48856=>"001011010",
  48857=>"110110111",
  48858=>"010110010",
  48859=>"111000001",
  48860=>"011001101",
  48861=>"010110011",
  48862=>"100000001",
  48863=>"010100111",
  48864=>"000001001",
  48865=>"111001100",
  48866=>"010110010",
  48867=>"001110001",
  48868=>"000100011",
  48869=>"010101000",
  48870=>"010010010",
  48871=>"101100001",
  48872=>"110110111",
  48873=>"011100000",
  48874=>"010010110",
  48875=>"010100010",
  48876=>"011111111",
  48877=>"010000001",
  48878=>"101100110",
  48879=>"100011000",
  48880=>"100100111",
  48881=>"000010111",
  48882=>"011001011",
  48883=>"110010101",
  48884=>"011010011",
  48885=>"101100011",
  48886=>"001111110",
  48887=>"001010011",
  48888=>"000001111",
  48889=>"000000000",
  48890=>"101010111",
  48891=>"010111011",
  48892=>"011001101",
  48893=>"110010111",
  48894=>"011110110",
  48895=>"010011101",
  48896=>"010011000",
  48897=>"101101011",
  48898=>"000110111",
  48899=>"100010001",
  48900=>"011010000",
  48901=>"000111101",
  48902=>"111111101",
  48903=>"010000011",
  48904=>"000000011",
  48905=>"110110001",
  48906=>"000100000",
  48907=>"001001000",
  48908=>"110111111",
  48909=>"101100101",
  48910=>"101110111",
  48911=>"111110111",
  48912=>"101001101",
  48913=>"111000000",
  48914=>"100110111",
  48915=>"011100111",
  48916=>"001001010",
  48917=>"010101101",
  48918=>"000000101",
  48919=>"010000001",
  48920=>"110000011",
  48921=>"110110011",
  48922=>"011011000",
  48923=>"001110100",
  48924=>"000000000",
  48925=>"011100100",
  48926=>"010110010",
  48927=>"111100000",
  48928=>"110010010",
  48929=>"111100000",
  48930=>"110011100",
  48931=>"111001101",
  48932=>"100110111",
  48933=>"101000001",
  48934=>"000001111",
  48935=>"110101001",
  48936=>"010011110",
  48937=>"111010100",
  48938=>"010011011",
  48939=>"110101001",
  48940=>"001010101",
  48941=>"000000000",
  48942=>"000100010",
  48943=>"010111000",
  48944=>"001000111",
  48945=>"101100000",
  48946=>"110111010",
  48947=>"100111011",
  48948=>"111001001",
  48949=>"010010101",
  48950=>"111111000",
  48951=>"100001000",
  48952=>"101100011",
  48953=>"100000011",
  48954=>"101010001",
  48955=>"001000111",
  48956=>"101100110",
  48957=>"010010010",
  48958=>"000101000",
  48959=>"101110000",
  48960=>"111111010",
  48961=>"010100111",
  48962=>"100110101",
  48963=>"110101110",
  48964=>"010101110",
  48965=>"011101101",
  48966=>"010001001",
  48967=>"101010100",
  48968=>"011011010",
  48969=>"000110010",
  48970=>"111111111",
  48971=>"000011000",
  48972=>"110111010",
  48973=>"010111000",
  48974=>"010110100",
  48975=>"001100100",
  48976=>"101111011",
  48977=>"010001111",
  48978=>"010100110",
  48979=>"011000000",
  48980=>"011110100",
  48981=>"010001001",
  48982=>"111011000",
  48983=>"011010001",
  48984=>"001111001",
  48985=>"110110100",
  48986=>"010101010",
  48987=>"011001001",
  48988=>"101101100",
  48989=>"111101011",
  48990=>"000111110",
  48991=>"000011000",
  48992=>"100010010",
  48993=>"110001000",
  48994=>"000010110",
  48995=>"111111011",
  48996=>"010100000",
  48997=>"110010001",
  48998=>"101011010",
  48999=>"010110011",
  49000=>"111100100",
  49001=>"101110010",
  49002=>"011010010",
  49003=>"101001010",
  49004=>"101001110",
  49005=>"000000111",
  49006=>"000011000",
  49007=>"001010010",
  49008=>"110100001",
  49009=>"110001110",
  49010=>"101001111",
  49011=>"010010001",
  49012=>"100010000",
  49013=>"100000101",
  49014=>"100100011",
  49015=>"110001111",
  49016=>"001100100",
  49017=>"000100000",
  49018=>"010011011",
  49019=>"010110111",
  49020=>"001110011",
  49021=>"110000011",
  49022=>"010100111",
  49023=>"100011010",
  49024=>"011111110",
  49025=>"111111001",
  49026=>"000111011",
  49027=>"110110111",
  49028=>"010111000",
  49029=>"101111000",
  49030=>"100001010",
  49031=>"110011100",
  49032=>"110111000",
  49033=>"011110000",
  49034=>"011010010",
  49035=>"101010011",
  49036=>"000010110",
  49037=>"111100101",
  49038=>"000101001",
  49039=>"010011101",
  49040=>"101001001",
  49041=>"011000110",
  49042=>"111000100",
  49043=>"011011000",
  49044=>"100110011",
  49045=>"000111100",
  49046=>"000111101",
  49047=>"111111110",
  49048=>"000010110",
  49049=>"100101000",
  49050=>"100000111",
  49051=>"110011000",
  49052=>"010000001",
  49053=>"110001110",
  49054=>"011110010",
  49055=>"110000011",
  49056=>"010011010",
  49057=>"111110111",
  49058=>"111001101",
  49059=>"000010001",
  49060=>"011000110",
  49061=>"011011101",
  49062=>"000001111",
  49063=>"110111000",
  49064=>"001111011",
  49065=>"011111010",
  49066=>"111011001",
  49067=>"010011000",
  49068=>"111111010",
  49069=>"010001010",
  49070=>"010100011",
  49071=>"110101110",
  49072=>"000101110",
  49073=>"011101001",
  49074=>"000101000",
  49075=>"110000110",
  49076=>"001111000",
  49077=>"010010011",
  49078=>"011101111",
  49079=>"110011101",
  49080=>"110111011",
  49081=>"100011000",
  49082=>"110111011",
  49083=>"110101101",
  49084=>"101000001",
  49085=>"100111010",
  49086=>"110011010",
  49087=>"101010110",
  49088=>"110111111",
  49089=>"110001111",
  49090=>"011100001",
  49091=>"011111100",
  49092=>"101010001",
  49093=>"000110110",
  49094=>"100110000",
  49095=>"101011001",
  49096=>"001010110",
  49097=>"100010101",
  49098=>"110110010",
  49099=>"010100110",
  49100=>"011110110",
  49101=>"100110111",
  49102=>"010000001",
  49103=>"111000011",
  49104=>"001001101",
  49105=>"100000000",
  49106=>"100000000",
  49107=>"101110011",
  49108=>"000110000",
  49109=>"011110001",
  49110=>"011101110",
  49111=>"001100011",
  49112=>"010101110",
  49113=>"110001110",
  49114=>"111111001",
  49115=>"001001001",
  49116=>"000000110",
  49117=>"101101100",
  49118=>"110110001",
  49119=>"100000011",
  49120=>"001111111",
  49121=>"000111100",
  49122=>"011110001",
  49123=>"000110100",
  49124=>"011101010",
  49125=>"111010001",
  49126=>"000011110",
  49127=>"101000100",
  49128=>"111000001",
  49129=>"111011001",
  49130=>"111010111",
  49131=>"000100001",
  49132=>"011000111",
  49133=>"111110111",
  49134=>"111110100",
  49135=>"011001101",
  49136=>"000000100",
  49137=>"110111000",
  49138=>"001101101",
  49139=>"001011000",
  49140=>"111100100",
  49141=>"111110100",
  49142=>"000000000",
  49143=>"110001110",
  49144=>"010001001",
  49145=>"011101110",
  49146=>"011011100",
  49147=>"101110010",
  49148=>"010000110",
  49149=>"111101010",
  49150=>"000010011",
  49151=>"001001111",
  49152=>"000001010",
  49153=>"111001011",
  49154=>"101111111",
  49155=>"001010100",
  49156=>"101111001",
  49157=>"001001000",
  49158=>"110111011",
  49159=>"111001101",
  49160=>"101000001",
  49161=>"101000110",
  49162=>"001110001",
  49163=>"101011111",
  49164=>"101111101",
  49165=>"110011110",
  49166=>"111110010",
  49167=>"110000001",
  49168=>"111010010",
  49169=>"110001100",
  49170=>"000010100",
  49171=>"000010001",
  49172=>"000000101",
  49173=>"000100001",
  49174=>"011000110",
  49175=>"010000010",
  49176=>"001011110",
  49177=>"101101111",
  49178=>"011001111",
  49179=>"010101011",
  49180=>"000101000",
  49181=>"000001001",
  49182=>"110100011",
  49183=>"100011001",
  49184=>"001110000",
  49185=>"101111111",
  49186=>"000100101",
  49187=>"001100101",
  49188=>"101010110",
  49189=>"000010100",
  49190=>"111111111",
  49191=>"011011001",
  49192=>"010101100",
  49193=>"110000010",
  49194=>"000001001",
  49195=>"011001011",
  49196=>"011110111",
  49197=>"100100111",
  49198=>"110101001",
  49199=>"001100110",
  49200=>"011110100",
  49201=>"000111100",
  49202=>"100101000",
  49203=>"010001010",
  49204=>"001011011",
  49205=>"010001111",
  49206=>"000110110",
  49207=>"111010001",
  49208=>"101110000",
  49209=>"100101110",
  49210=>"111110001",
  49211=>"101000010",
  49212=>"000110111",
  49213=>"101101100",
  49214=>"010100001",
  49215=>"001000100",
  49216=>"001100010",
  49217=>"000010100",
  49218=>"000101010",
  49219=>"100001001",
  49220=>"001100001",
  49221=>"000111011",
  49222=>"011011100",
  49223=>"101011010",
  49224=>"001001000",
  49225=>"010100011",
  49226=>"011000100",
  49227=>"111111000",
  49228=>"000010010",
  49229=>"001001001",
  49230=>"000111110",
  49231=>"001110110",
  49232=>"110101001",
  49233=>"001010010",
  49234=>"011100001",
  49235=>"010101110",
  49236=>"110011100",
  49237=>"010010110",
  49238=>"111000101",
  49239=>"111100010",
  49240=>"100001101",
  49241=>"110010111",
  49242=>"011001011",
  49243=>"000110001",
  49244=>"000000000",
  49245=>"101000110",
  49246=>"101011110",
  49247=>"011011101",
  49248=>"111110000",
  49249=>"100011100",
  49250=>"000000001",
  49251=>"000011111",
  49252=>"101101000",
  49253=>"101101101",
  49254=>"000010000",
  49255=>"011110000",
  49256=>"011010000",
  49257=>"101111111",
  49258=>"011011011",
  49259=>"100010101",
  49260=>"100010000",
  49261=>"010101111",
  49262=>"101011110",
  49263=>"111000010",
  49264=>"110011000",
  49265=>"001101111",
  49266=>"010100011",
  49267=>"101010001",
  49268=>"101110111",
  49269=>"100111101",
  49270=>"010101011",
  49271=>"001010111",
  49272=>"001011100",
  49273=>"000100001",
  49274=>"000101110",
  49275=>"001101011",
  49276=>"100010010",
  49277=>"101101111",
  49278=>"000001000",
  49279=>"001000000",
  49280=>"000000111",
  49281=>"111110000",
  49282=>"110011110",
  49283=>"001001101",
  49284=>"001000001",
  49285=>"011011100",
  49286=>"001000011",
  49287=>"011000000",
  49288=>"000101010",
  49289=>"000010000",
  49290=>"001011000",
  49291=>"101111000",
  49292=>"110111100",
  49293=>"001010001",
  49294=>"110010001",
  49295=>"111111000",
  49296=>"110111001",
  49297=>"101101100",
  49298=>"111110100",
  49299=>"110101000",
  49300=>"011101111",
  49301=>"000100001",
  49302=>"110100110",
  49303=>"111110000",
  49304=>"100111000",
  49305=>"111000110",
  49306=>"100011110",
  49307=>"111011011",
  49308=>"110010110",
  49309=>"000001111",
  49310=>"001111000",
  49311=>"100000001",
  49312=>"100010101",
  49313=>"000011001",
  49314=>"101011000",
  49315=>"100011000",
  49316=>"101001100",
  49317=>"010101111",
  49318=>"011001111",
  49319=>"111000110",
  49320=>"111110000",
  49321=>"011111100",
  49322=>"011111111",
  49323=>"111000111",
  49324=>"000010110",
  49325=>"100001000",
  49326=>"100101110",
  49327=>"000000101",
  49328=>"010010111",
  49329=>"010100111",
  49330=>"111100011",
  49331=>"010011001",
  49332=>"110100111",
  49333=>"000000001",
  49334=>"101111111",
  49335=>"011110100",
  49336=>"000000101",
  49337=>"001101000",
  49338=>"110100110",
  49339=>"110101111",
  49340=>"100001000",
  49341=>"001001101",
  49342=>"010010000",
  49343=>"010011001",
  49344=>"101100110",
  49345=>"111011111",
  49346=>"110110010",
  49347=>"110111010",
  49348=>"110001001",
  49349=>"110001101",
  49350=>"100001101",
  49351=>"111100111",
  49352=>"011101000",
  49353=>"001010100",
  49354=>"010000100",
  49355=>"001110000",
  49356=>"001101001",
  49357=>"111110110",
  49358=>"010110001",
  49359=>"000101111",
  49360=>"111010010",
  49361=>"100010001",
  49362=>"100111001",
  49363=>"001111001",
  49364=>"001100011",
  49365=>"001001110",
  49366=>"101000101",
  49367=>"110101100",
  49368=>"100000010",
  49369=>"110000100",
  49370=>"000001001",
  49371=>"011101100",
  49372=>"111000010",
  49373=>"010111110",
  49374=>"101110010",
  49375=>"011110001",
  49376=>"010000101",
  49377=>"011100111",
  49378=>"010011110",
  49379=>"111000100",
  49380=>"100100001",
  49381=>"110000001",
  49382=>"000110001",
  49383=>"110110001",
  49384=>"101001101",
  49385=>"100110100",
  49386=>"010100000",
  49387=>"111100000",
  49388=>"000110000",
  49389=>"001101010",
  49390=>"010100000",
  49391=>"011001101",
  49392=>"010100000",
  49393=>"100011110",
  49394=>"110001111",
  49395=>"101111101",
  49396=>"110010010",
  49397=>"001001001",
  49398=>"100011100",
  49399=>"000010001",
  49400=>"111011110",
  49401=>"010010100",
  49402=>"011100000",
  49403=>"010010010",
  49404=>"011011001",
  49405=>"011110101",
  49406=>"111001110",
  49407=>"111111101",
  49408=>"101111110",
  49409=>"000000101",
  49410=>"011011001",
  49411=>"110011111",
  49412=>"000011111",
  49413=>"010111111",
  49414=>"110000011",
  49415=>"000000101",
  49416=>"001000000",
  49417=>"011110101",
  49418=>"001100100",
  49419=>"000011100",
  49420=>"010000001",
  49421=>"010011101",
  49422=>"100000000",
  49423=>"000110110",
  49424=>"101101100",
  49425=>"001111100",
  49426=>"011111010",
  49427=>"011100010",
  49428=>"101011111",
  49429=>"111110000",
  49430=>"000111101",
  49431=>"110010110",
  49432=>"001100000",
  49433=>"001000011",
  49434=>"000100001",
  49435=>"111101000",
  49436=>"101000101",
  49437=>"101110011",
  49438=>"010100000",
  49439=>"111001001",
  49440=>"100001100",
  49441=>"101101000",
  49442=>"010000000",
  49443=>"110001010",
  49444=>"000101100",
  49445=>"001111001",
  49446=>"011000001",
  49447=>"010001110",
  49448=>"000111000",
  49449=>"101001010",
  49450=>"111111101",
  49451=>"100100100",
  49452=>"100010100",
  49453=>"100001111",
  49454=>"111110111",
  49455=>"101110111",
  49456=>"010110101",
  49457=>"011110111",
  49458=>"011001111",
  49459=>"110110101",
  49460=>"000000111",
  49461=>"001100000",
  49462=>"111010110",
  49463=>"010001111",
  49464=>"000001000",
  49465=>"100010000",
  49466=>"000111011",
  49467=>"110000101",
  49468=>"110011111",
  49469=>"011010111",
  49470=>"010010000",
  49471=>"000010001",
  49472=>"110011001",
  49473=>"100000100",
  49474=>"110110001",
  49475=>"000000010",
  49476=>"001001110",
  49477=>"101100000",
  49478=>"000001100",
  49479=>"110111111",
  49480=>"000011110",
  49481=>"010100001",
  49482=>"011110110",
  49483=>"100001001",
  49484=>"110010111",
  49485=>"111111100",
  49486=>"010100111",
  49487=>"011110000",
  49488=>"111000000",
  49489=>"111111100",
  49490=>"010100100",
  49491=>"010000000",
  49492=>"011111000",
  49493=>"011111111",
  49494=>"000000101",
  49495=>"110111011",
  49496=>"001100101",
  49497=>"111001010",
  49498=>"111100010",
  49499=>"110110010",
  49500=>"001000011",
  49501=>"001101010",
  49502=>"100011011",
  49503=>"100101100",
  49504=>"010100000",
  49505=>"110010010",
  49506=>"100101111",
  49507=>"000100000",
  49508=>"111110011",
  49509=>"110011000",
  49510=>"001010010",
  49511=>"100000000",
  49512=>"111001100",
  49513=>"101100100",
  49514=>"000000101",
  49515=>"100101110",
  49516=>"011001001",
  49517=>"000101110",
  49518=>"101010010",
  49519=>"000001010",
  49520=>"000000011",
  49521=>"000011101",
  49522=>"000110011",
  49523=>"000111101",
  49524=>"001101011",
  49525=>"101000001",
  49526=>"110001001",
  49527=>"000000100",
  49528=>"100100000",
  49529=>"110100010",
  49530=>"011101010",
  49531=>"111101011",
  49532=>"000110110",
  49533=>"110000110",
  49534=>"100111111",
  49535=>"000000000",
  49536=>"001001001",
  49537=>"110001010",
  49538=>"111001001",
  49539=>"100110100",
  49540=>"110001110",
  49541=>"011000100",
  49542=>"111001001",
  49543=>"000000010",
  49544=>"000000000",
  49545=>"100101110",
  49546=>"101110111",
  49547=>"001010110",
  49548=>"111000000",
  49549=>"011110101",
  49550=>"111010000",
  49551=>"010111101",
  49552=>"110111111",
  49553=>"111100110",
  49554=>"110001000",
  49555=>"000001001",
  49556=>"000011011",
  49557=>"011001001",
  49558=>"011111101",
  49559=>"101011111",
  49560=>"111000110",
  49561=>"101001111",
  49562=>"101010011",
  49563=>"000000000",
  49564=>"110111101",
  49565=>"000001011",
  49566=>"010100101",
  49567=>"000011000",
  49568=>"011100001",
  49569=>"010000110",
  49570=>"001100110",
  49571=>"110111110",
  49572=>"001110101",
  49573=>"100001101",
  49574=>"011100101",
  49575=>"101101110",
  49576=>"111101000",
  49577=>"000000001",
  49578=>"011110000",
  49579=>"000011110",
  49580=>"000000101",
  49581=>"001001001",
  49582=>"111110000",
  49583=>"001010001",
  49584=>"000010100",
  49585=>"010000001",
  49586=>"000100000",
  49587=>"101011111",
  49588=>"010001111",
  49589=>"100100000",
  49590=>"110101110",
  49591=>"010000110",
  49592=>"100001100",
  49593=>"000001000",
  49594=>"001111001",
  49595=>"001000111",
  49596=>"101101110",
  49597=>"101110100",
  49598=>"111001000",
  49599=>"011000100",
  49600=>"000000111",
  49601=>"000001110",
  49602=>"110110101",
  49603=>"110101101",
  49604=>"101000000",
  49605=>"100111000",
  49606=>"001001011",
  49607=>"000000000",
  49608=>"000001010",
  49609=>"110100001",
  49610=>"101000110",
  49611=>"110101111",
  49612=>"111000010",
  49613=>"100101110",
  49614=>"010000010",
  49615=>"000000011",
  49616=>"001101011",
  49617=>"001111001",
  49618=>"010100001",
  49619=>"010101011",
  49620=>"011100010",
  49621=>"011010000",
  49622=>"001101001",
  49623=>"010010110",
  49624=>"011001111",
  49625=>"011100111",
  49626=>"101111000",
  49627=>"010010001",
  49628=>"001111101",
  49629=>"101001100",
  49630=>"101100110",
  49631=>"001001000",
  49632=>"110101100",
  49633=>"000010111",
  49634=>"000001011",
  49635=>"000011001",
  49636=>"001010111",
  49637=>"111011010",
  49638=>"001001001",
  49639=>"101001001",
  49640=>"010011100",
  49641=>"110110111",
  49642=>"110100010",
  49643=>"000110001",
  49644=>"011010110",
  49645=>"001001110",
  49646=>"000000100",
  49647=>"000000010",
  49648=>"111111100",
  49649=>"100100011",
  49650=>"111000100",
  49651=>"100100101",
  49652=>"010110111",
  49653=>"100000001",
  49654=>"011110110",
  49655=>"101000011",
  49656=>"010101000",
  49657=>"101110101",
  49658=>"111010101",
  49659=>"011001100",
  49660=>"110111010",
  49661=>"001011101",
  49662=>"111110101",
  49663=>"011000010",
  49664=>"100110110",
  49665=>"001100000",
  49666=>"000011111",
  49667=>"010000000",
  49668=>"101000111",
  49669=>"011110101",
  49670=>"001010111",
  49671=>"000010010",
  49672=>"101001011",
  49673=>"101110001",
  49674=>"111001011",
  49675=>"001000010",
  49676=>"001100010",
  49677=>"010011010",
  49678=>"000010000",
  49679=>"111100110",
  49680=>"100111000",
  49681=>"111011011",
  49682=>"010010000",
  49683=>"110111111",
  49684=>"000000110",
  49685=>"011001001",
  49686=>"110110101",
  49687=>"010010101",
  49688=>"010011001",
  49689=>"110010101",
  49690=>"111001000",
  49691=>"101000100",
  49692=>"100100001",
  49693=>"110000001",
  49694=>"110010100",
  49695=>"111011101",
  49696=>"010001111",
  49697=>"110001110",
  49698=>"000000110",
  49699=>"000100010",
  49700=>"101101111",
  49701=>"001100000",
  49702=>"111101111",
  49703=>"001000011",
  49704=>"000110001",
  49705=>"000101000",
  49706=>"100110000",
  49707=>"101011000",
  49708=>"111010000",
  49709=>"010001001",
  49710=>"010111110",
  49711=>"010100100",
  49712=>"110100011",
  49713=>"010100001",
  49714=>"110100101",
  49715=>"110011110",
  49716=>"110110011",
  49717=>"011111001",
  49718=>"010110111",
  49719=>"100000111",
  49720=>"001101100",
  49721=>"000000001",
  49722=>"101000100",
  49723=>"001100101",
  49724=>"001000101",
  49725=>"010001101",
  49726=>"100001001",
  49727=>"010001101",
  49728=>"000101000",
  49729=>"101011101",
  49730=>"101010010",
  49731=>"011001010",
  49732=>"100011111",
  49733=>"011111011",
  49734=>"000001010",
  49735=>"011001111",
  49736=>"001100010",
  49737=>"001111110",
  49738=>"010010001",
  49739=>"010001111",
  49740=>"000011100",
  49741=>"010110010",
  49742=>"100000101",
  49743=>"101101100",
  49744=>"010110101",
  49745=>"100100000",
  49746=>"010011001",
  49747=>"001001110",
  49748=>"010101101",
  49749=>"001111010",
  49750=>"010010101",
  49751=>"101100100",
  49752=>"101001100",
  49753=>"100001101",
  49754=>"101100000",
  49755=>"010000101",
  49756=>"010100011",
  49757=>"000001011",
  49758=>"001101010",
  49759=>"111100001",
  49760=>"101001101",
  49761=>"010000110",
  49762=>"100001000",
  49763=>"100000100",
  49764=>"101101001",
  49765=>"101001100",
  49766=>"101111111",
  49767=>"001101010",
  49768=>"001010100",
  49769=>"100010111",
  49770=>"001011111",
  49771=>"001110110",
  49772=>"111100110",
  49773=>"101000010",
  49774=>"101000011",
  49775=>"111100011",
  49776=>"010000110",
  49777=>"100101100",
  49778=>"110101001",
  49779=>"010010101",
  49780=>"110111011",
  49781=>"000001010",
  49782=>"011001111",
  49783=>"111001000",
  49784=>"011011000",
  49785=>"011101100",
  49786=>"011110110",
  49787=>"001001100",
  49788=>"100110110",
  49789=>"101100101",
  49790=>"110000011",
  49791=>"111010100",
  49792=>"001011010",
  49793=>"000110001",
  49794=>"000000110",
  49795=>"000001101",
  49796=>"100110000",
  49797=>"101000001",
  49798=>"100001000",
  49799=>"101110111",
  49800=>"010001001",
  49801=>"000100000",
  49802=>"100001011",
  49803=>"000101010",
  49804=>"111001110",
  49805=>"010010000",
  49806=>"000100101",
  49807=>"111101011",
  49808=>"000010000",
  49809=>"100011010",
  49810=>"111000000",
  49811=>"110010100",
  49812=>"000000101",
  49813=>"011100010",
  49814=>"101100110",
  49815=>"010011000",
  49816=>"111111000",
  49817=>"010101111",
  49818=>"111001000",
  49819=>"110100000",
  49820=>"000010000",
  49821=>"000001111",
  49822=>"101101000",
  49823=>"100101011",
  49824=>"101101110",
  49825=>"111111010",
  49826=>"000101110",
  49827=>"101111000",
  49828=>"100101111",
  49829=>"111111110",
  49830=>"000000010",
  49831=>"010011111",
  49832=>"101101011",
  49833=>"100011011",
  49834=>"111111011",
  49835=>"000011011",
  49836=>"000110000",
  49837=>"100101000",
  49838=>"100111111",
  49839=>"010000010",
  49840=>"000010011",
  49841=>"010100011",
  49842=>"110000000",
  49843=>"010000110",
  49844=>"110000111",
  49845=>"111001110",
  49846=>"100010011",
  49847=>"110010000",
  49848=>"101111000",
  49849=>"011010110",
  49850=>"001011111",
  49851=>"111011001",
  49852=>"110100011",
  49853=>"011000000",
  49854=>"000110111",
  49855=>"100110110",
  49856=>"000010000",
  49857=>"011111001",
  49858=>"011001100",
  49859=>"111111100",
  49860=>"100011100",
  49861=>"000000100",
  49862=>"011110101",
  49863=>"100110000",
  49864=>"100010110",
  49865=>"000110100",
  49866=>"110010110",
  49867=>"111001010",
  49868=>"111110100",
  49869=>"010000101",
  49870=>"000110000",
  49871=>"110011101",
  49872=>"100100100",
  49873=>"101100011",
  49874=>"111101100",
  49875=>"100010001",
  49876=>"010000000",
  49877=>"001000001",
  49878=>"000011110",
  49879=>"100010001",
  49880=>"000011010",
  49881=>"110101100",
  49882=>"110001101",
  49883=>"000000010",
  49884=>"101101111",
  49885=>"011001011",
  49886=>"101000101",
  49887=>"101011001",
  49888=>"111100101",
  49889=>"000010001",
  49890=>"011010100",
  49891=>"101100011",
  49892=>"101001011",
  49893=>"111001000",
  49894=>"000101111",
  49895=>"000010111",
  49896=>"000000001",
  49897=>"000111011",
  49898=>"010010110",
  49899=>"111001010",
  49900=>"000001010",
  49901=>"100000111",
  49902=>"100100110",
  49903=>"110001110",
  49904=>"000110111",
  49905=>"000100110",
  49906=>"111000000",
  49907=>"011011011",
  49908=>"100010000",
  49909=>"000100001",
  49910=>"010100010",
  49911=>"010101100",
  49912=>"111001111",
  49913=>"000100001",
  49914=>"010010111",
  49915=>"100001111",
  49916=>"000011110",
  49917=>"110011100",
  49918=>"000101101",
  49919=>"000000001",
  49920=>"000011110",
  49921=>"110001011",
  49922=>"110000101",
  49923=>"011111100",
  49924=>"010100000",
  49925=>"000000110",
  49926=>"011011100",
  49927=>"001011011",
  49928=>"000011000",
  49929=>"010100100",
  49930=>"111011111",
  49931=>"000010000",
  49932=>"110110010",
  49933=>"111101001",
  49934=>"010111010",
  49935=>"101110010",
  49936=>"111100001",
  49937=>"000000101",
  49938=>"111100101",
  49939=>"001011010",
  49940=>"111110000",
  49941=>"000011000",
  49942=>"011011000",
  49943=>"111000000",
  49944=>"100010000",
  49945=>"000001110",
  49946=>"000000101",
  49947=>"000101001",
  49948=>"011110100",
  49949=>"010101000",
  49950=>"000110001",
  49951=>"000101001",
  49952=>"110001000",
  49953=>"111101001",
  49954=>"101100000",
  49955=>"111101111",
  49956=>"110111001",
  49957=>"000100101",
  49958=>"101000000",
  49959=>"100101000",
  49960=>"110011010",
  49961=>"100111101",
  49962=>"101000100",
  49963=>"100001101",
  49964=>"010110100",
  49965=>"100101101",
  49966=>"110001110",
  49967=>"000100011",
  49968=>"111111010",
  49969=>"111111111",
  49970=>"100111001",
  49971=>"111101010",
  49972=>"100001111",
  49973=>"010100011",
  49974=>"110101111",
  49975=>"111001110",
  49976=>"110000001",
  49977=>"100111111",
  49978=>"000001100",
  49979=>"101111010",
  49980=>"101110000",
  49981=>"101110110",
  49982=>"111101110",
  49983=>"000000010",
  49984=>"101011101",
  49985=>"000010111",
  49986=>"111011000",
  49987=>"010110001",
  49988=>"110110110",
  49989=>"011011111",
  49990=>"001011000",
  49991=>"111110101",
  49992=>"001001100",
  49993=>"010001010",
  49994=>"011011011",
  49995=>"000000101",
  49996=>"101111000",
  49997=>"011010001",
  49998=>"100111100",
  49999=>"001110101",
  50000=>"011110010",
  50001=>"000011111",
  50002=>"001010001",
  50003=>"001110010",
  50004=>"000010011",
  50005=>"010001001",
  50006=>"001000101",
  50007=>"000001110",
  50008=>"011010011",
  50009=>"000001100",
  50010=>"001111000",
  50011=>"000101001",
  50012=>"111111110",
  50013=>"000001100",
  50014=>"001111011",
  50015=>"001101100",
  50016=>"011000100",
  50017=>"010111000",
  50018=>"111000000",
  50019=>"001011011",
  50020=>"110101000",
  50021=>"111110010",
  50022=>"111111011",
  50023=>"110110100",
  50024=>"111010110",
  50025=>"000010101",
  50026=>"111000010",
  50027=>"111101100",
  50028=>"000000010",
  50029=>"110011110",
  50030=>"000111001",
  50031=>"100100111",
  50032=>"010011100",
  50033=>"001001110",
  50034=>"011001100",
  50035=>"000101010",
  50036=>"100010000",
  50037=>"000011000",
  50038=>"010110011",
  50039=>"110111111",
  50040=>"010000111",
  50041=>"001011110",
  50042=>"101100011",
  50043=>"011110110",
  50044=>"000100110",
  50045=>"011001000",
  50046=>"101001101",
  50047=>"011101100",
  50048=>"110001010",
  50049=>"110111111",
  50050=>"100100011",
  50051=>"101001010",
  50052=>"111011010",
  50053=>"101011111",
  50054=>"011110101",
  50055=>"000100100",
  50056=>"101010111",
  50057=>"000000011",
  50058=>"000110111",
  50059=>"111010111",
  50060=>"001010110",
  50061=>"001001001",
  50062=>"010111110",
  50063=>"111111000",
  50064=>"100010011",
  50065=>"010100001",
  50066=>"010110000",
  50067=>"110011110",
  50068=>"001011010",
  50069=>"011011110",
  50070=>"000110110",
  50071=>"001110110",
  50072=>"101101111",
  50073=>"100101010",
  50074=>"011100100",
  50075=>"110001110",
  50076=>"110011111",
  50077=>"011010010",
  50078=>"101100001",
  50079=>"100010000",
  50080=>"011111100",
  50081=>"100001111",
  50082=>"100110100",
  50083=>"001000000",
  50084=>"100011000",
  50085=>"110110100",
  50086=>"011111011",
  50087=>"001110001",
  50088=>"101100000",
  50089=>"000110001",
  50090=>"011101110",
  50091=>"011010011",
  50092=>"110000100",
  50093=>"101100000",
  50094=>"110011001",
  50095=>"000000001",
  50096=>"001000001",
  50097=>"011011010",
  50098=>"000101000",
  50099=>"101101011",
  50100=>"111110000",
  50101=>"010011111",
  50102=>"100101011",
  50103=>"001111001",
  50104=>"101001000",
  50105=>"000111111",
  50106=>"101101011",
  50107=>"101110111",
  50108=>"010000010",
  50109=>"001001110",
  50110=>"100101010",
  50111=>"000000111",
  50112=>"101010110",
  50113=>"111010000",
  50114=>"000101111",
  50115=>"000111011",
  50116=>"000000001",
  50117=>"111000101",
  50118=>"011110011",
  50119=>"000111000",
  50120=>"011000100",
  50121=>"010111011",
  50122=>"100100011",
  50123=>"011101011",
  50124=>"011010101",
  50125=>"010100101",
  50126=>"001111111",
  50127=>"101000111",
  50128=>"100111100",
  50129=>"000101001",
  50130=>"010100111",
  50131=>"001101000",
  50132=>"101011110",
  50133=>"100100011",
  50134=>"101101100",
  50135=>"001101010",
  50136=>"111101011",
  50137=>"101001100",
  50138=>"101100110",
  50139=>"000000111",
  50140=>"111101010",
  50141=>"010111101",
  50142=>"000100001",
  50143=>"111101110",
  50144=>"111110100",
  50145=>"000101011",
  50146=>"110010001",
  50147=>"110100100",
  50148=>"010000011",
  50149=>"111010000",
  50150=>"001101101",
  50151=>"101111001",
  50152=>"111001111",
  50153=>"101100110",
  50154=>"010000000",
  50155=>"111100010",
  50156=>"111001100",
  50157=>"001001110",
  50158=>"010010010",
  50159=>"000010110",
  50160=>"111111010",
  50161=>"000010100",
  50162=>"111001110",
  50163=>"111111101",
  50164=>"011011010",
  50165=>"011000011",
  50166=>"000100001",
  50167=>"000100000",
  50168=>"100011010",
  50169=>"000011101",
  50170=>"111011011",
  50171=>"000001001",
  50172=>"000000000",
  50173=>"011110100",
  50174=>"000000010",
  50175=>"100001101",
  50176=>"011011011",
  50177=>"101110001",
  50178=>"000100010",
  50179=>"101101010",
  50180=>"011000110",
  50181=>"000001110",
  50182=>"011111001",
  50183=>"111100011",
  50184=>"100101010",
  50185=>"010010101",
  50186=>"010001100",
  50187=>"011001000",
  50188=>"110011011",
  50189=>"010001000",
  50190=>"000011010",
  50191=>"010010111",
  50192=>"001011011",
  50193=>"010000010",
  50194=>"011011101",
  50195=>"000010001",
  50196=>"101000101",
  50197=>"111111110",
  50198=>"100001111",
  50199=>"011000110",
  50200=>"001010110",
  50201=>"111110011",
  50202=>"010110010",
  50203=>"110110010",
  50204=>"000101100",
  50205=>"000101001",
  50206=>"111100100",
  50207=>"111011011",
  50208=>"000000100",
  50209=>"011000010",
  50210=>"010110010",
  50211=>"111100111",
  50212=>"000111001",
  50213=>"001111000",
  50214=>"010001001",
  50215=>"010001011",
  50216=>"111100011",
  50217=>"010001001",
  50218=>"111011111",
  50219=>"001001110",
  50220=>"001111000",
  50221=>"111110101",
  50222=>"001011111",
  50223=>"111110111",
  50224=>"110100000",
  50225=>"011011001",
  50226=>"100110110",
  50227=>"000110111",
  50228=>"001101111",
  50229=>"011011111",
  50230=>"110011001",
  50231=>"010100111",
  50232=>"101101000",
  50233=>"101111111",
  50234=>"101100000",
  50235=>"110000000",
  50236=>"111001011",
  50237=>"000110001",
  50238=>"111001110",
  50239=>"000011100",
  50240=>"100001000",
  50241=>"001000001",
  50242=>"000000110",
  50243=>"111101011",
  50244=>"010001110",
  50245=>"011111000",
  50246=>"010100000",
  50247=>"010111010",
  50248=>"110101111",
  50249=>"101111010",
  50250=>"110101110",
  50251=>"101001011",
  50252=>"111001000",
  50253=>"111111011",
  50254=>"010000001",
  50255=>"011111100",
  50256=>"000111111",
  50257=>"000101010",
  50258=>"100100000",
  50259=>"110000010",
  50260=>"000000001",
  50261=>"011001011",
  50262=>"100111001",
  50263=>"111011011",
  50264=>"011111101",
  50265=>"000100110",
  50266=>"100111011",
  50267=>"001110111",
  50268=>"010111011",
  50269=>"011111011",
  50270=>"011100100",
  50271=>"111100000",
  50272=>"100111100",
  50273=>"110010110",
  50274=>"001101001",
  50275=>"100001010",
  50276=>"010001011",
  50277=>"010011001",
  50278=>"011110110",
  50279=>"010010100",
  50280=>"101011010",
  50281=>"100101100",
  50282=>"000101111",
  50283=>"010010010",
  50284=>"100100010",
  50285=>"011111100",
  50286=>"100100111",
  50287=>"000011111",
  50288=>"101100001",
  50289=>"011000100",
  50290=>"010100001",
  50291=>"111101000",
  50292=>"010010101",
  50293=>"001001001",
  50294=>"110010000",
  50295=>"001000101",
  50296=>"101100010",
  50297=>"001110001",
  50298=>"011111000",
  50299=>"000000111",
  50300=>"001101001",
  50301=>"000011101",
  50302=>"101111011",
  50303=>"010111000",
  50304=>"110011110",
  50305=>"111000011",
  50306=>"101010110",
  50307=>"101111001",
  50308=>"010110010",
  50309=>"000011111",
  50310=>"010110010",
  50311=>"100001110",
  50312=>"110001100",
  50313=>"000110100",
  50314=>"001000110",
  50315=>"100001011",
  50316=>"000100010",
  50317=>"110111101",
  50318=>"111000001",
  50319=>"110110001",
  50320=>"110100101",
  50321=>"110111111",
  50322=>"110011111",
  50323=>"100111010",
  50324=>"010011010",
  50325=>"100100110",
  50326=>"011111101",
  50327=>"100101100",
  50328=>"110111100",
  50329=>"111110111",
  50330=>"110000101",
  50331=>"000011000",
  50332=>"011011011",
  50333=>"111110111",
  50334=>"111011101",
  50335=>"000000111",
  50336=>"111000111",
  50337=>"000110100",
  50338=>"010010001",
  50339=>"010000010",
  50340=>"110010110",
  50341=>"000010011",
  50342=>"100111100",
  50343=>"010100110",
  50344=>"011111011",
  50345=>"110110110",
  50346=>"011100011",
  50347=>"010011000",
  50348=>"110010111",
  50349=>"011101001",
  50350=>"000100010",
  50351=>"110110100",
  50352=>"010100010",
  50353=>"101000001",
  50354=>"001011100",
  50355=>"110110011",
  50356=>"000110101",
  50357=>"111011100",
  50358=>"010100000",
  50359=>"001001001",
  50360=>"110110101",
  50361=>"111110001",
  50362=>"110110001",
  50363=>"001000011",
  50364=>"010101100",
  50365=>"000011011",
  50366=>"001110110",
  50367=>"001110000",
  50368=>"111110011",
  50369=>"111111010",
  50370=>"100101100",
  50371=>"000101010",
  50372=>"000011101",
  50373=>"010100100",
  50374=>"011111111",
  50375=>"010100001",
  50376=>"100011110",
  50377=>"110001111",
  50378=>"001110110",
  50379=>"011101111",
  50380=>"101110011",
  50381=>"000010001",
  50382=>"011001010",
  50383=>"000000100",
  50384=>"100011010",
  50385=>"011001111",
  50386=>"111111011",
  50387=>"001100001",
  50388=>"100010001",
  50389=>"110101101",
  50390=>"111100000",
  50391=>"011011111",
  50392=>"111111110",
  50393=>"010011100",
  50394=>"110011110",
  50395=>"111100111",
  50396=>"011001100",
  50397=>"111111101",
  50398=>"110100110",
  50399=>"001001011",
  50400=>"111000100",
  50401=>"000010011",
  50402=>"000011111",
  50403=>"010110111",
  50404=>"110000110",
  50405=>"100000100",
  50406=>"010001111",
  50407=>"101100101",
  50408=>"010001111",
  50409=>"011110101",
  50410=>"110111111",
  50411=>"010111100",
  50412=>"110000010",
  50413=>"010101010",
  50414=>"101110111",
  50415=>"110100100",
  50416=>"010001110",
  50417=>"111110110",
  50418=>"111110110",
  50419=>"111011101",
  50420=>"010100101",
  50421=>"010010011",
  50422=>"100000011",
  50423=>"100111010",
  50424=>"000010100",
  50425=>"101010001",
  50426=>"000011010",
  50427=>"010001110",
  50428=>"000011001",
  50429=>"101011111",
  50430=>"010000101",
  50431=>"000100101",
  50432=>"010101110",
  50433=>"001101001",
  50434=>"110000110",
  50435=>"011010011",
  50436=>"100011010",
  50437=>"101110101",
  50438=>"001100000",
  50439=>"111010111",
  50440=>"011111000",
  50441=>"111010110",
  50442=>"101110111",
  50443=>"000010011",
  50444=>"010101110",
  50445=>"110010111",
  50446=>"111110110",
  50447=>"101110111",
  50448=>"100110101",
  50449=>"010001000",
  50450=>"010111000",
  50451=>"001110100",
  50452=>"100110010",
  50453=>"001111100",
  50454=>"001110101",
  50455=>"100000110",
  50456=>"000000111",
  50457=>"111111110",
  50458=>"111011011",
  50459=>"001010010",
  50460=>"101010000",
  50461=>"101110001",
  50462=>"111111100",
  50463=>"001100101",
  50464=>"011000011",
  50465=>"111110000",
  50466=>"010011011",
  50467=>"000011101",
  50468=>"011101011",
  50469=>"100000101",
  50470=>"010011101",
  50471=>"011010100",
  50472=>"010000000",
  50473=>"011100011",
  50474=>"010101100",
  50475=>"101000000",
  50476=>"001111001",
  50477=>"010110110",
  50478=>"011011000",
  50479=>"001010011",
  50480=>"100101110",
  50481=>"101001110",
  50482=>"111101111",
  50483=>"101011110",
  50484=>"011000011",
  50485=>"100110010",
  50486=>"001001111",
  50487=>"111100010",
  50488=>"111111111",
  50489=>"100111111",
  50490=>"000010000",
  50491=>"010100011",
  50492=>"000010011",
  50493=>"010001000",
  50494=>"101010001",
  50495=>"000000100",
  50496=>"111000100",
  50497=>"100010111",
  50498=>"000100110",
  50499=>"011101110",
  50500=>"011001010",
  50501=>"010011110",
  50502=>"000111101",
  50503=>"111110011",
  50504=>"010000101",
  50505=>"010101110",
  50506=>"011000100",
  50507=>"011011101",
  50508=>"100010100",
  50509=>"010100101",
  50510=>"000011111",
  50511=>"000010000",
  50512=>"111100000",
  50513=>"011110111",
  50514=>"110110110",
  50515=>"100000000",
  50516=>"111010000",
  50517=>"011100110",
  50518=>"010010110",
  50519=>"100011110",
  50520=>"111010111",
  50521=>"001111110",
  50522=>"001101110",
  50523=>"000001001",
  50524=>"000011100",
  50525=>"000011100",
  50526=>"010101000",
  50527=>"000111000",
  50528=>"001100011",
  50529=>"011001111",
  50530=>"101100010",
  50531=>"110000011",
  50532=>"000101101",
  50533=>"001111101",
  50534=>"111110010",
  50535=>"001111010",
  50536=>"000110110",
  50537=>"111010000",
  50538=>"111010110",
  50539=>"100001100",
  50540=>"001010101",
  50541=>"010110011",
  50542=>"101101000",
  50543=>"111111100",
  50544=>"000000010",
  50545=>"010000001",
  50546=>"000011111",
  50547=>"011010111",
  50548=>"000111100",
  50549=>"000100100",
  50550=>"101111110",
  50551=>"110001010",
  50552=>"010100101",
  50553=>"010010001",
  50554=>"111101101",
  50555=>"011001111",
  50556=>"101111101",
  50557=>"011011101",
  50558=>"110110100",
  50559=>"111011001",
  50560=>"111001000",
  50561=>"100111101",
  50562=>"011101101",
  50563=>"101000010",
  50564=>"001011111",
  50565=>"011111101",
  50566=>"100011101",
  50567=>"101011101",
  50568=>"111110110",
  50569=>"010000010",
  50570=>"110101100",
  50571=>"110101001",
  50572=>"100110011",
  50573=>"110111111",
  50574=>"110101010",
  50575=>"101011100",
  50576=>"001101011",
  50577=>"010001010",
  50578=>"111010101",
  50579=>"101100101",
  50580=>"000101010",
  50581=>"011111011",
  50582=>"011000100",
  50583=>"001110001",
  50584=>"010001101",
  50585=>"110000000",
  50586=>"101011110",
  50587=>"011110111",
  50588=>"111001100",
  50589=>"010011110",
  50590=>"111011111",
  50591=>"000100101",
  50592=>"100111010",
  50593=>"110011010",
  50594=>"111011111",
  50595=>"000001000",
  50596=>"100000001",
  50597=>"111001101",
  50598=>"110111110",
  50599=>"010111011",
  50600=>"000011000",
  50601=>"110111001",
  50602=>"010000100",
  50603=>"111110100",
  50604=>"110100001",
  50605=>"001100110",
  50606=>"100100101",
  50607=>"100101001",
  50608=>"111010111",
  50609=>"100101001",
  50610=>"010011011",
  50611=>"111100101",
  50612=>"101001001",
  50613=>"000101011",
  50614=>"111111101",
  50615=>"110110011",
  50616=>"100000001",
  50617=>"110011101",
  50618=>"110100111",
  50619=>"010010001",
  50620=>"011010001",
  50621=>"001110101",
  50622=>"101100110",
  50623=>"010110111",
  50624=>"110100111",
  50625=>"111010011",
  50626=>"110110111",
  50627=>"111111101",
  50628=>"111001001",
  50629=>"010101001",
  50630=>"011000011",
  50631=>"000101111",
  50632=>"111000101",
  50633=>"101101011",
  50634=>"111101100",
  50635=>"010010101",
  50636=>"011101001",
  50637=>"001101111",
  50638=>"001100000",
  50639=>"100001111",
  50640=>"111110000",
  50641=>"100010100",
  50642=>"001011000",
  50643=>"010111000",
  50644=>"000010100",
  50645=>"110111010",
  50646=>"011011000",
  50647=>"111110001",
  50648=>"001011100",
  50649=>"011011101",
  50650=>"101001111",
  50651=>"101110111",
  50652=>"000000111",
  50653=>"001110100",
  50654=>"010111111",
  50655=>"101001100",
  50656=>"111111101",
  50657=>"111001000",
  50658=>"110111000",
  50659=>"100111111",
  50660=>"001001001",
  50661=>"000101110",
  50662=>"000010110",
  50663=>"001110100",
  50664=>"000001001",
  50665=>"011001111",
  50666=>"101010010",
  50667=>"100110011",
  50668=>"001001110",
  50669=>"101110000",
  50670=>"110110111",
  50671=>"011111000",
  50672=>"011011001",
  50673=>"001100111",
  50674=>"000010001",
  50675=>"010010111",
  50676=>"011100100",
  50677=>"100011111",
  50678=>"110111100",
  50679=>"111001001",
  50680=>"110110001",
  50681=>"110110111",
  50682=>"000001010",
  50683=>"000100100",
  50684=>"010110110",
  50685=>"100111100",
  50686=>"111111010",
  50687=>"110110000",
  50688=>"001100000",
  50689=>"100010110",
  50690=>"100110011",
  50691=>"100101001",
  50692=>"001101001",
  50693=>"111011111",
  50694=>"111100011",
  50695=>"100110110",
  50696=>"110010111",
  50697=>"000011011",
  50698=>"110100100",
  50699=>"000010000",
  50700=>"000000000",
  50701=>"110011100",
  50702=>"010001111",
  50703=>"101010010",
  50704=>"110010000",
  50705=>"011010011",
  50706=>"001101110",
  50707=>"111010100",
  50708=>"111010011",
  50709=>"000011101",
  50710=>"010011011",
  50711=>"111001010",
  50712=>"010001110",
  50713=>"011111001",
  50714=>"001111110",
  50715=>"001011111",
  50716=>"101000000",
  50717=>"110011111",
  50718=>"001110001",
  50719=>"001001110",
  50720=>"011010111",
  50721=>"110101000",
  50722=>"001011010",
  50723=>"011111010",
  50724=>"111000011",
  50725=>"001000010",
  50726=>"001011010",
  50727=>"110100100",
  50728=>"111101111",
  50729=>"010011010",
  50730=>"111111111",
  50731=>"000000110",
  50732=>"010010111",
  50733=>"011111101",
  50734=>"001010010",
  50735=>"010000000",
  50736=>"001001000",
  50737=>"101000011",
  50738=>"010100010",
  50739=>"101000100",
  50740=>"110000111",
  50741=>"010100111",
  50742=>"100001001",
  50743=>"001111110",
  50744=>"011101001",
  50745=>"000100111",
  50746=>"100100000",
  50747=>"000000010",
  50748=>"101111000",
  50749=>"101000111",
  50750=>"100101011",
  50751=>"011111000",
  50752=>"011010010",
  50753=>"010000101",
  50754=>"000110001",
  50755=>"110010001",
  50756=>"011111001",
  50757=>"011011100",
  50758=>"111110010",
  50759=>"110001010",
  50760=>"100010100",
  50761=>"100010011",
  50762=>"010100010",
  50763=>"110100000",
  50764=>"110101010",
  50765=>"011101011",
  50766=>"111100111",
  50767=>"110101110",
  50768=>"100001000",
  50769=>"110100101",
  50770=>"110101000",
  50771=>"000110100",
  50772=>"001010000",
  50773=>"100011011",
  50774=>"110000010",
  50775=>"000111011",
  50776=>"101110010",
  50777=>"001111001",
  50778=>"000000101",
  50779=>"001100100",
  50780=>"000010110",
  50781=>"010111000",
  50782=>"111111100",
  50783=>"101000001",
  50784=>"100110011",
  50785=>"100110111",
  50786=>"100011111",
  50787=>"100111011",
  50788=>"011011000",
  50789=>"101101011",
  50790=>"111001101",
  50791=>"100001000",
  50792=>"010101111",
  50793=>"101010101",
  50794=>"101111100",
  50795=>"110000000",
  50796=>"010100011",
  50797=>"010010100",
  50798=>"111000000",
  50799=>"110101011",
  50800=>"100010111",
  50801=>"111111111",
  50802=>"100100011",
  50803=>"000011101",
  50804=>"101000000",
  50805=>"110001101",
  50806=>"011101000",
  50807=>"111100110",
  50808=>"111111011",
  50809=>"100101011",
  50810=>"111111101",
  50811=>"110001100",
  50812=>"001001010",
  50813=>"111010000",
  50814=>"100011000",
  50815=>"000100100",
  50816=>"111101100",
  50817=>"101101001",
  50818=>"101001100",
  50819=>"111111111",
  50820=>"111111111",
  50821=>"111010011",
  50822=>"001001110",
  50823=>"011100001",
  50824=>"100000110",
  50825=>"111010000",
  50826=>"010010110",
  50827=>"100101000",
  50828=>"101100000",
  50829=>"111011101",
  50830=>"111011101",
  50831=>"000100011",
  50832=>"000001011",
  50833=>"101100001",
  50834=>"101100001",
  50835=>"010001111",
  50836=>"011001001",
  50837=>"000101100",
  50838=>"101000001",
  50839=>"100101110",
  50840=>"010011110",
  50841=>"010001100",
  50842=>"001101101",
  50843=>"010100000",
  50844=>"001001110",
  50845=>"111110001",
  50846=>"100010000",
  50847=>"001000011",
  50848=>"111000111",
  50849=>"011110001",
  50850=>"000110011",
  50851=>"111111010",
  50852=>"011010000",
  50853=>"110101110",
  50854=>"011000011",
  50855=>"101100100",
  50856=>"011010000",
  50857=>"010000101",
  50858=>"101100111",
  50859=>"000111110",
  50860=>"001101011",
  50861=>"010111011",
  50862=>"111010100",
  50863=>"000100001",
  50864=>"101111111",
  50865=>"000110010",
  50866=>"100011001",
  50867=>"110000000",
  50868=>"000101101",
  50869=>"110000000",
  50870=>"100101010",
  50871=>"010111110",
  50872=>"000100000",
  50873=>"110111100",
  50874=>"100110010",
  50875=>"101101001",
  50876=>"010010000",
  50877=>"100001000",
  50878=>"100110110",
  50879=>"101011001",
  50880=>"000001101",
  50881=>"111011111",
  50882=>"000110001",
  50883=>"010010011",
  50884=>"001110100",
  50885=>"111001100",
  50886=>"001000010",
  50887=>"111110010",
  50888=>"100110101",
  50889=>"011100101",
  50890=>"010010100",
  50891=>"011000011",
  50892=>"010011110",
  50893=>"011110010",
  50894=>"110111111",
  50895=>"110100101",
  50896=>"101101000",
  50897=>"111111001",
  50898=>"111011111",
  50899=>"111100001",
  50900=>"100101100",
  50901=>"000010111",
  50902=>"001111101",
  50903=>"101100101",
  50904=>"000101000",
  50905=>"110000111",
  50906=>"110111101",
  50907=>"100010000",
  50908=>"111011011",
  50909=>"000000111",
  50910=>"110100010",
  50911=>"101110000",
  50912=>"100111000",
  50913=>"011010111",
  50914=>"011001111",
  50915=>"001110111",
  50916=>"101110101",
  50917=>"010111101",
  50918=>"111011111",
  50919=>"110101011",
  50920=>"111111111",
  50921=>"101010011",
  50922=>"110111101",
  50923=>"111001010",
  50924=>"111000110",
  50925=>"000111010",
  50926=>"101100001",
  50927=>"101010101",
  50928=>"000011111",
  50929=>"000100111",
  50930=>"001110110",
  50931=>"110010101",
  50932=>"010011011",
  50933=>"000100100",
  50934=>"100100011",
  50935=>"010001001",
  50936=>"011011110",
  50937=>"001100000",
  50938=>"000010001",
  50939=>"010100011",
  50940=>"000111010",
  50941=>"110000000",
  50942=>"110110110",
  50943=>"101101001",
  50944=>"010000010",
  50945=>"111110000",
  50946=>"001001110",
  50947=>"100010110",
  50948=>"101001110",
  50949=>"110111101",
  50950=>"010011110",
  50951=>"100001001",
  50952=>"101111010",
  50953=>"000110001",
  50954=>"010011110",
  50955=>"010000100",
  50956=>"000111011",
  50957=>"000100001",
  50958=>"001010101",
  50959=>"001110101",
  50960=>"000011011",
  50961=>"110111111",
  50962=>"001101011",
  50963=>"100000110",
  50964=>"001111001",
  50965=>"110110101",
  50966=>"110111111",
  50967=>"111011110",
  50968=>"110100111",
  50969=>"000110011",
  50970=>"000110101",
  50971=>"011011100",
  50972=>"101101000",
  50973=>"110011111",
  50974=>"011010001",
  50975=>"100110011",
  50976=>"111010111",
  50977=>"100010100",
  50978=>"011011000",
  50979=>"110110110",
  50980=>"000000000",
  50981=>"001100000",
  50982=>"101011010",
  50983=>"110010010",
  50984=>"100001011",
  50985=>"000110010",
  50986=>"100011000",
  50987=>"011111011",
  50988=>"101001011",
  50989=>"101010000",
  50990=>"000101010",
  50991=>"000010001",
  50992=>"011111110",
  50993=>"101111110",
  50994=>"000100111",
  50995=>"000001110",
  50996=>"110101010",
  50997=>"001011010",
  50998=>"011011110",
  50999=>"010110111",
  51000=>"011111001",
  51001=>"011000010",
  51002=>"000001010",
  51003=>"010101011",
  51004=>"110011111",
  51005=>"111100010",
  51006=>"100001000",
  51007=>"011100100",
  51008=>"101101100",
  51009=>"101011010",
  51010=>"100100101",
  51011=>"111101101",
  51012=>"101101011",
  51013=>"100000000",
  51014=>"000000101",
  51015=>"110000111",
  51016=>"100110011",
  51017=>"101010101",
  51018=>"001111011",
  51019=>"101111111",
  51020=>"001001001",
  51021=>"111101101",
  51022=>"000101111",
  51023=>"000010100",
  51024=>"100010110",
  51025=>"110010010",
  51026=>"010011110",
  51027=>"111100001",
  51028=>"000101101",
  51029=>"001100100",
  51030=>"100010110",
  51031=>"011100011",
  51032=>"111101110",
  51033=>"011001111",
  51034=>"101011010",
  51035=>"111111101",
  51036=>"100000111",
  51037=>"111111011",
  51038=>"010000101",
  51039=>"010011010",
  51040=>"111000000",
  51041=>"011111010",
  51042=>"010100011",
  51043=>"111100111",
  51044=>"000000010",
  51045=>"011001111",
  51046=>"001010111",
  51047=>"011111011",
  51048=>"110000111",
  51049=>"101001101",
  51050=>"011110100",
  51051=>"001000101",
  51052=>"100011101",
  51053=>"110100000",
  51054=>"010101000",
  51055=>"010101111",
  51056=>"011001101",
  51057=>"011101111",
  51058=>"111111010",
  51059=>"011111000",
  51060=>"110101001",
  51061=>"011110111",
  51062=>"111110100",
  51063=>"010011010",
  51064=>"001101001",
  51065=>"010001011",
  51066=>"000001001",
  51067=>"110010111",
  51068=>"011111101",
  51069=>"101100110",
  51070=>"101011101",
  51071=>"111000001",
  51072=>"000010111",
  51073=>"110000000",
  51074=>"110110000",
  51075=>"011011011",
  51076=>"110011011",
  51077=>"010010101",
  51078=>"110000100",
  51079=>"010101100",
  51080=>"001111000",
  51081=>"001111000",
  51082=>"010100011",
  51083=>"110011111",
  51084=>"010010111",
  51085=>"100100000",
  51086=>"000111111",
  51087=>"111001010",
  51088=>"000100111",
  51089=>"100011001",
  51090=>"111000011",
  51091=>"000010110",
  51092=>"110100100",
  51093=>"101000000",
  51094=>"110000100",
  51095=>"111010110",
  51096=>"100001011",
  51097=>"110000011",
  51098=>"101101110",
  51099=>"101111001",
  51100=>"110000000",
  51101=>"001110010",
  51102=>"101111011",
  51103=>"110001110",
  51104=>"010000000",
  51105=>"110101101",
  51106=>"100101110",
  51107=>"111111000",
  51108=>"101010101",
  51109=>"011000010",
  51110=>"011011110",
  51111=>"110011111",
  51112=>"000101110",
  51113=>"110100111",
  51114=>"000100000",
  51115=>"100100010",
  51116=>"101001000",
  51117=>"011000001",
  51118=>"110010010",
  51119=>"111101110",
  51120=>"110101100",
  51121=>"001110000",
  51122=>"001110011",
  51123=>"010010011",
  51124=>"000110110",
  51125=>"100010100",
  51126=>"000100011",
  51127=>"100011010",
  51128=>"111110010",
  51129=>"110010101",
  51130=>"111101011",
  51131=>"100011010",
  51132=>"100011110",
  51133=>"101101000",
  51134=>"001001101",
  51135=>"111011101",
  51136=>"101010000",
  51137=>"110011101",
  51138=>"110101100",
  51139=>"111001101",
  51140=>"110111101",
  51141=>"010010000",
  51142=>"010101101",
  51143=>"110011000",
  51144=>"011100001",
  51145=>"011011001",
  51146=>"010100011",
  51147=>"100101100",
  51148=>"110000010",
  51149=>"101101101",
  51150=>"100110111",
  51151=>"100111001",
  51152=>"010010001",
  51153=>"101111011",
  51154=>"010011101",
  51155=>"001101000",
  51156=>"100011100",
  51157=>"100011100",
  51158=>"010111110",
  51159=>"000010111",
  51160=>"010011100",
  51161=>"110100010",
  51162=>"110010001",
  51163=>"111101110",
  51164=>"000110110",
  51165=>"010011001",
  51166=>"011001001",
  51167=>"101011111",
  51168=>"111100100",
  51169=>"100011000",
  51170=>"000011101",
  51171=>"001101011",
  51172=>"010100110",
  51173=>"110111011",
  51174=>"101010010",
  51175=>"011101010",
  51176=>"111001000",
  51177=>"001111001",
  51178=>"010010011",
  51179=>"010000000",
  51180=>"010101110",
  51181=>"111001111",
  51182=>"010100000",
  51183=>"011110001",
  51184=>"101111101",
  51185=>"010011010",
  51186=>"001100101",
  51187=>"000110010",
  51188=>"110001001",
  51189=>"010100111",
  51190=>"101100101",
  51191=>"010100111",
  51192=>"000101011",
  51193=>"111100100",
  51194=>"101101111",
  51195=>"011110111",
  51196=>"101100001",
  51197=>"010010011",
  51198=>"101110110",
  51199=>"000000100",
  51200=>"001111101",
  51201=>"000111000",
  51202=>"100111110",
  51203=>"110111011",
  51204=>"111011011",
  51205=>"101011000",
  51206=>"001001111",
  51207=>"010100111",
  51208=>"011111101",
  51209=>"101010000",
  51210=>"111100001",
  51211=>"110110010",
  51212=>"010110101",
  51213=>"100100000",
  51214=>"100110011",
  51215=>"010110110",
  51216=>"100110000",
  51217=>"001111011",
  51218=>"010000011",
  51219=>"110111011",
  51220=>"010100000",
  51221=>"011111000",
  51222=>"011011111",
  51223=>"101010101",
  51224=>"110011010",
  51225=>"010101100",
  51226=>"111010111",
  51227=>"010001011",
  51228=>"111011011",
  51229=>"001101011",
  51230=>"000011000",
  51231=>"000011101",
  51232=>"110111111",
  51233=>"010101011",
  51234=>"011110100",
  51235=>"100011000",
  51236=>"011110010",
  51237=>"000001110",
  51238=>"010001000",
  51239=>"111100000",
  51240=>"100000010",
  51241=>"011010111",
  51242=>"010110100",
  51243=>"110011011",
  51244=>"001100011",
  51245=>"111011010",
  51246=>"000100011",
  51247=>"111011000",
  51248=>"010011101",
  51249=>"010101100",
  51250=>"101101010",
  51251=>"111011101",
  51252=>"010101000",
  51253=>"001011011",
  51254=>"101010000",
  51255=>"010000010",
  51256=>"000000101",
  51257=>"110101110",
  51258=>"100000110",
  51259=>"010011111",
  51260=>"110111000",
  51261=>"111010111",
  51262=>"110011000",
  51263=>"110000001",
  51264=>"011001000",
  51265=>"110010000",
  51266=>"001011011",
  51267=>"101010010",
  51268=>"101011001",
  51269=>"111010000",
  51270=>"111100001",
  51271=>"101000000",
  51272=>"000101101",
  51273=>"000000010",
  51274=>"001010000",
  51275=>"010000100",
  51276=>"000001101",
  51277=>"011001001",
  51278=>"001110001",
  51279=>"000110001",
  51280=>"010000100",
  51281=>"111010100",
  51282=>"001011001",
  51283=>"101111011",
  51284=>"000011010",
  51285=>"111100001",
  51286=>"010111100",
  51287=>"011110000",
  51288=>"101011000",
  51289=>"011110111",
  51290=>"101100101",
  51291=>"111100101",
  51292=>"111111010",
  51293=>"011101110",
  51294=>"000111101",
  51295=>"110100101",
  51296=>"001000000",
  51297=>"100100000",
  51298=>"101110011",
  51299=>"001010101",
  51300=>"100000101",
  51301=>"001101001",
  51302=>"110001101",
  51303=>"101001010",
  51304=>"100000111",
  51305=>"000011100",
  51306=>"111011111",
  51307=>"100101100",
  51308=>"000010011",
  51309=>"010001101",
  51310=>"001111000",
  51311=>"111101110",
  51312=>"010101001",
  51313=>"010100000",
  51314=>"111000100",
  51315=>"101100101",
  51316=>"001101111",
  51317=>"010100001",
  51318=>"000001101",
  51319=>"101110110",
  51320=>"110110110",
  51321=>"110100010",
  51322=>"101111100",
  51323=>"001010000",
  51324=>"111100011",
  51325=>"001100110",
  51326=>"011110101",
  51327=>"110001100",
  51328=>"101000010",
  51329=>"000111101",
  51330=>"011111111",
  51331=>"110101011",
  51332=>"111101110",
  51333=>"110110111",
  51334=>"011000010",
  51335=>"001101111",
  51336=>"100000110",
  51337=>"100111010",
  51338=>"011100001",
  51339=>"110001000",
  51340=>"000111110",
  51341=>"010100111",
  51342=>"111011101",
  51343=>"001011000",
  51344=>"101110100",
  51345=>"011111001",
  51346=>"111100101",
  51347=>"010010111",
  51348=>"000000010",
  51349=>"000100110",
  51350=>"111111000",
  51351=>"101101111",
  51352=>"101000011",
  51353=>"100100100",
  51354=>"110100011",
  51355=>"000000001",
  51356=>"110000100",
  51357=>"110010110",
  51358=>"001010000",
  51359=>"101001100",
  51360=>"011011100",
  51361=>"110101100",
  51362=>"011110110",
  51363=>"110110100",
  51364=>"011100000",
  51365=>"111000101",
  51366=>"111101001",
  51367=>"000100001",
  51368=>"001101000",
  51369=>"110100001",
  51370=>"000100000",
  51371=>"000010110",
  51372=>"100100011",
  51373=>"000001010",
  51374=>"110101001",
  51375=>"100111011",
  51376=>"000011011",
  51377=>"000000111",
  51378=>"000110010",
  51379=>"110000100",
  51380=>"001110000",
  51381=>"110010110",
  51382=>"111010001",
  51383=>"111101111",
  51384=>"100101101",
  51385=>"000000000",
  51386=>"110001001",
  51387=>"101110000",
  51388=>"001001101",
  51389=>"010001010",
  51390=>"001011001",
  51391=>"010001000",
  51392=>"010111000",
  51393=>"011111101",
  51394=>"101010110",
  51395=>"011111011",
  51396=>"001001011",
  51397=>"111011000",
  51398=>"110000011",
  51399=>"111001110",
  51400=>"010100000",
  51401=>"011110000",
  51402=>"110000000",
  51403=>"000001000",
  51404=>"110010100",
  51405=>"011100110",
  51406=>"010100111",
  51407=>"001000100",
  51408=>"001100011",
  51409=>"110110111",
  51410=>"001111101",
  51411=>"010101111",
  51412=>"001110101",
  51413=>"000111011",
  51414=>"111100001",
  51415=>"100111001",
  51416=>"000000100",
  51417=>"111001001",
  51418=>"011000100",
  51419=>"111100001",
  51420=>"101111101",
  51421=>"000011010",
  51422=>"111100101",
  51423=>"101011001",
  51424=>"110110110",
  51425=>"011111010",
  51426=>"000110000",
  51427=>"100011001",
  51428=>"111111000",
  51429=>"011011111",
  51430=>"101111001",
  51431=>"011101111",
  51432=>"000111011",
  51433=>"001001111",
  51434=>"101000001",
  51435=>"110101000",
  51436=>"000101010",
  51437=>"000101111",
  51438=>"001100001",
  51439=>"010000001",
  51440=>"000111111",
  51441=>"000100100",
  51442=>"001101010",
  51443=>"100101111",
  51444=>"010000001",
  51445=>"111100101",
  51446=>"000001110",
  51447=>"010010010",
  51448=>"101000011",
  51449=>"001000110",
  51450=>"101110010",
  51451=>"000110011",
  51452=>"101011101",
  51453=>"110111111",
  51454=>"110110100",
  51455=>"010000100",
  51456=>"010010111",
  51457=>"001110010",
  51458=>"111110100",
  51459=>"010000101",
  51460=>"010101100",
  51461=>"010011001",
  51462=>"001011101",
  51463=>"000000101",
  51464=>"001101010",
  51465=>"110101110",
  51466=>"010010111",
  51467=>"010110111",
  51468=>"011011001",
  51469=>"000100001",
  51470=>"111010110",
  51471=>"100001011",
  51472=>"101011011",
  51473=>"011010100",
  51474=>"011110001",
  51475=>"101110010",
  51476=>"011111010",
  51477=>"110101111",
  51478=>"101111111",
  51479=>"000111101",
  51480=>"010100110",
  51481=>"110010100",
  51482=>"110101101",
  51483=>"110011101",
  51484=>"001100110",
  51485=>"011000011",
  51486=>"100000000",
  51487=>"011110100",
  51488=>"001000100",
  51489=>"011100010",
  51490=>"111101100",
  51491=>"010100101",
  51492=>"101011000",
  51493=>"111001001",
  51494=>"101101101",
  51495=>"101100001",
  51496=>"000001110",
  51497=>"110001001",
  51498=>"110010000",
  51499=>"011010101",
  51500=>"110110101",
  51501=>"101110110",
  51502=>"001110010",
  51503=>"011111111",
  51504=>"000101101",
  51505=>"001001110",
  51506=>"111110011",
  51507=>"101110100",
  51508=>"011111010",
  51509=>"100100110",
  51510=>"010101100",
  51511=>"111010010",
  51512=>"110110011",
  51513=>"000110101",
  51514=>"110100010",
  51515=>"111111100",
  51516=>"011010100",
  51517=>"011011010",
  51518=>"000011010",
  51519=>"101011011",
  51520=>"010111010",
  51521=>"110000010",
  51522=>"111110101",
  51523=>"101010100",
  51524=>"001111110",
  51525=>"001010111",
  51526=>"100101000",
  51527=>"101100111",
  51528=>"000110011",
  51529=>"111011001",
  51530=>"100000011",
  51531=>"000111100",
  51532=>"001011000",
  51533=>"000100011",
  51534=>"010001010",
  51535=>"011001001",
  51536=>"110111001",
  51537=>"101110011",
  51538=>"100000111",
  51539=>"111010011",
  51540=>"000110000",
  51541=>"100010010",
  51542=>"010001111",
  51543=>"000010111",
  51544=>"110010000",
  51545=>"100001000",
  51546=>"000101000",
  51547=>"011011010",
  51548=>"100001001",
  51549=>"000110101",
  51550=>"100010001",
  51551=>"111110110",
  51552=>"100011100",
  51553=>"010011110",
  51554=>"010000001",
  51555=>"101100000",
  51556=>"001000101",
  51557=>"111110111",
  51558=>"000011010",
  51559=>"101101011",
  51560=>"010000000",
  51561=>"110001101",
  51562=>"010100001",
  51563=>"011000001",
  51564=>"010101011",
  51565=>"111010111",
  51566=>"100000000",
  51567=>"110100101",
  51568=>"100111101",
  51569=>"011101000",
  51570=>"001011111",
  51571=>"100110000",
  51572=>"110111001",
  51573=>"100011010",
  51574=>"100101111",
  51575=>"011010000",
  51576=>"100101111",
  51577=>"110111101",
  51578=>"001101111",
  51579=>"110000101",
  51580=>"000110011",
  51581=>"101101000",
  51582=>"111000000",
  51583=>"101001001",
  51584=>"101011000",
  51585=>"010001100",
  51586=>"111001111",
  51587=>"101110001",
  51588=>"100100011",
  51589=>"110001000",
  51590=>"101101110",
  51591=>"010001100",
  51592=>"001100110",
  51593=>"101100010",
  51594=>"101001110",
  51595=>"011111100",
  51596=>"011100100",
  51597=>"001000000",
  51598=>"110111000",
  51599=>"110000011",
  51600=>"011011001",
  51601=>"010000110",
  51602=>"001111101",
  51603=>"001100000",
  51604=>"000110000",
  51605=>"000011001",
  51606=>"111101111",
  51607=>"000101010",
  51608=>"000111001",
  51609=>"101001011",
  51610=>"110111001",
  51611=>"001101111",
  51612=>"101111101",
  51613=>"001100011",
  51614=>"001000100",
  51615=>"101010100",
  51616=>"100011101",
  51617=>"111101111",
  51618=>"011100001",
  51619=>"010100111",
  51620=>"111011111",
  51621=>"001110100",
  51622=>"101011100",
  51623=>"001110110",
  51624=>"100011000",
  51625=>"010010000",
  51626=>"001001101",
  51627=>"010011101",
  51628=>"011000010",
  51629=>"011001101",
  51630=>"111000100",
  51631=>"101010000",
  51632=>"100110010",
  51633=>"110000010",
  51634=>"111010111",
  51635=>"111010001",
  51636=>"101110001",
  51637=>"100000000",
  51638=>"010110110",
  51639=>"101111011",
  51640=>"100010010",
  51641=>"101101000",
  51642=>"001110110",
  51643=>"011001011",
  51644=>"101011110",
  51645=>"111101101",
  51646=>"111111100",
  51647=>"001101001",
  51648=>"100010001",
  51649=>"001010010",
  51650=>"100101010",
  51651=>"000100110",
  51652=>"001111001",
  51653=>"001110000",
  51654=>"001001101",
  51655=>"011000000",
  51656=>"111011111",
  51657=>"011100000",
  51658=>"100101011",
  51659=>"101101001",
  51660=>"001010000",
  51661=>"001110010",
  51662=>"100100101",
  51663=>"010011101",
  51664=>"110000010",
  51665=>"001100111",
  51666=>"000111011",
  51667=>"000101101",
  51668=>"111110110",
  51669=>"101010110",
  51670=>"010001011",
  51671=>"000010010",
  51672=>"011001111",
  51673=>"110001000",
  51674=>"111111001",
  51675=>"001000001",
  51676=>"111110110",
  51677=>"111110110",
  51678=>"000000000",
  51679=>"000001110",
  51680=>"111000111",
  51681=>"110011000",
  51682=>"010010010",
  51683=>"110111101",
  51684=>"001110000",
  51685=>"111111011",
  51686=>"111110011",
  51687=>"101001101",
  51688=>"000001110",
  51689=>"101011011",
  51690=>"010100111",
  51691=>"100101111",
  51692=>"001101111",
  51693=>"000001000",
  51694=>"001101010",
  51695=>"100011000",
  51696=>"000110111",
  51697=>"110110000",
  51698=>"010101010",
  51699=>"101001010",
  51700=>"011011011",
  51701=>"111001001",
  51702=>"101101100",
  51703=>"101111110",
  51704=>"001100101",
  51705=>"001011111",
  51706=>"111000011",
  51707=>"111010110",
  51708=>"011111010",
  51709=>"010111111",
  51710=>"001010111",
  51711=>"010011100",
  51712=>"000010010",
  51713=>"010010010",
  51714=>"010101010",
  51715=>"111100100",
  51716=>"010000001",
  51717=>"101111111",
  51718=>"010111000",
  51719=>"100000010",
  51720=>"101111011",
  51721=>"000111001",
  51722=>"000000101",
  51723=>"110101010",
  51724=>"111010001",
  51725=>"001110011",
  51726=>"110111010",
  51727=>"110110111",
  51728=>"101111010",
  51729=>"110011010",
  51730=>"011000000",
  51731=>"110000001",
  51732=>"100011000",
  51733=>"010111001",
  51734=>"000101110",
  51735=>"000001101",
  51736=>"110111111",
  51737=>"111100101",
  51738=>"111000000",
  51739=>"000010001",
  51740=>"101000001",
  51741=>"101111111",
  51742=>"000111011",
  51743=>"011111001",
  51744=>"000000111",
  51745=>"001010100",
  51746=>"111101000",
  51747=>"011001001",
  51748=>"001011010",
  51749=>"000110001",
  51750=>"010110010",
  51751=>"011001100",
  51752=>"000000101",
  51753=>"000001001",
  51754=>"000110100",
  51755=>"110111001",
  51756=>"010000101",
  51757=>"001010100",
  51758=>"000110111",
  51759=>"111001111",
  51760=>"001010000",
  51761=>"011111110",
  51762=>"001110101",
  51763=>"110100100",
  51764=>"010010110",
  51765=>"111010111",
  51766=>"011011000",
  51767=>"000101101",
  51768=>"000010011",
  51769=>"011001000",
  51770=>"011010001",
  51771=>"011010101",
  51772=>"101111111",
  51773=>"000101101",
  51774=>"110000000",
  51775=>"000001000",
  51776=>"110100111",
  51777=>"100101010",
  51778=>"111001110",
  51779=>"010111101",
  51780=>"000111110",
  51781=>"111100010",
  51782=>"101001110",
  51783=>"000000000",
  51784=>"010111000",
  51785=>"010100111",
  51786=>"000001000",
  51787=>"101011000",
  51788=>"100000000",
  51789=>"010110111",
  51790=>"000100101",
  51791=>"001011101",
  51792=>"101000010",
  51793=>"010001000",
  51794=>"000111111",
  51795=>"101001100",
  51796=>"001110101",
  51797=>"011110110",
  51798=>"001010100",
  51799=>"100101001",
  51800=>"110101000",
  51801=>"111100100",
  51802=>"110000001",
  51803=>"001001000",
  51804=>"110010100",
  51805=>"011010011",
  51806=>"010100111",
  51807=>"000011110",
  51808=>"110010000",
  51809=>"100010111",
  51810=>"000000011",
  51811=>"011011111",
  51812=>"101000011",
  51813=>"000010101",
  51814=>"101111110",
  51815=>"100001001",
  51816=>"101011101",
  51817=>"111100101",
  51818=>"110001011",
  51819=>"101000111",
  51820=>"101001011",
  51821=>"010111110",
  51822=>"111111000",
  51823=>"100011001",
  51824=>"100000001",
  51825=>"001011001",
  51826=>"001001101",
  51827=>"010100111",
  51828=>"011111101",
  51829=>"001100010",
  51830=>"011010011",
  51831=>"011010110",
  51832=>"100011100",
  51833=>"000001011",
  51834=>"001011100",
  51835=>"100111001",
  51836=>"110010100",
  51837=>"001000000",
  51838=>"111011010",
  51839=>"010110100",
  51840=>"101010100",
  51841=>"011101000",
  51842=>"011111001",
  51843=>"011100000",
  51844=>"100011010",
  51845=>"100001011",
  51846=>"110101000",
  51847=>"010101000",
  51848=>"000011100",
  51849=>"100000000",
  51850=>"010100101",
  51851=>"010010000",
  51852=>"100010000",
  51853=>"010101010",
  51854=>"011100100",
  51855=>"011101101",
  51856=>"011111111",
  51857=>"010110110",
  51858=>"110011101",
  51859=>"010001111",
  51860=>"000011001",
  51861=>"101000100",
  51862=>"000010010",
  51863=>"010100101",
  51864=>"110010011",
  51865=>"000000111",
  51866=>"010101111",
  51867=>"000000111",
  51868=>"001011001",
  51869=>"001111101",
  51870=>"111110100",
  51871=>"110100100",
  51872=>"001101110",
  51873=>"000001000",
  51874=>"000000011",
  51875=>"001111000",
  51876=>"111101101",
  51877=>"101011100",
  51878=>"001110110",
  51879=>"100100111",
  51880=>"111001101",
  51881=>"111100110",
  51882=>"011000110",
  51883=>"010111001",
  51884=>"010110110",
  51885=>"000001111",
  51886=>"111110111",
  51887=>"001001100",
  51888=>"101101100",
  51889=>"000011111",
  51890=>"001001000",
  51891=>"001110111",
  51892=>"000110110",
  51893=>"111011011",
  51894=>"110110000",
  51895=>"110011011",
  51896=>"001000001",
  51897=>"000100011",
  51898=>"011111010",
  51899=>"011110000",
  51900=>"101101001",
  51901=>"000110101",
  51902=>"010001101",
  51903=>"111011100",
  51904=>"001000000",
  51905=>"011001011",
  51906=>"101010000",
  51907=>"110001001",
  51908=>"000110010",
  51909=>"101111001",
  51910=>"101110100",
  51911=>"001011001",
  51912=>"101111011",
  51913=>"101001011",
  51914=>"010100000",
  51915=>"110001010",
  51916=>"110110100",
  51917=>"000000100",
  51918=>"011000101",
  51919=>"011010001",
  51920=>"110110111",
  51921=>"000001010",
  51922=>"111011100",
  51923=>"011010010",
  51924=>"010111111",
  51925=>"011100010",
  51926=>"010110011",
  51927=>"010110010",
  51928=>"100000111",
  51929=>"011000111",
  51930=>"100010000",
  51931=>"111111001",
  51932=>"000100011",
  51933=>"101111110",
  51934=>"000010000",
  51935=>"100001101",
  51936=>"111000000",
  51937=>"100001100",
  51938=>"110011001",
  51939=>"001010100",
  51940=>"001101000",
  51941=>"110110000",
  51942=>"010111110",
  51943=>"010100100",
  51944=>"100100001",
  51945=>"111011010",
  51946=>"010100101",
  51947=>"101010000",
  51948=>"110111011",
  51949=>"011111111",
  51950=>"001101011",
  51951=>"010110111",
  51952=>"111101101",
  51953=>"010011000",
  51954=>"011111000",
  51955=>"000100010",
  51956=>"110000000",
  51957=>"011010001",
  51958=>"100011010",
  51959=>"101010010",
  51960=>"010101000",
  51961=>"000000111",
  51962=>"010110000",
  51963=>"001111001",
  51964=>"010111000",
  51965=>"011111111",
  51966=>"110001011",
  51967=>"111100010",
  51968=>"110111100",
  51969=>"011100011",
  51970=>"010010000",
  51971=>"110100101",
  51972=>"100001001",
  51973=>"000100000",
  51974=>"000000001",
  51975=>"000010000",
  51976=>"000111010",
  51977=>"010101011",
  51978=>"011011001",
  51979=>"001100010",
  51980=>"000000111",
  51981=>"010101011",
  51982=>"011111110",
  51983=>"010110000",
  51984=>"111100101",
  51985=>"000000000",
  51986=>"001001001",
  51987=>"001111010",
  51988=>"100010001",
  51989=>"000000010",
  51990=>"011101100",
  51991=>"110100010",
  51992=>"011110101",
  51993=>"000010010",
  51994=>"111000101",
  51995=>"111100011",
  51996=>"001100100",
  51997=>"101001110",
  51998=>"111001111",
  51999=>"000111100",
  52000=>"000001001",
  52001=>"001001011",
  52002=>"010010111",
  52003=>"110110001",
  52004=>"101100011",
  52005=>"111110111",
  52006=>"110010011",
  52007=>"101000010",
  52008=>"001001100",
  52009=>"000101001",
  52010=>"011110111",
  52011=>"000001001",
  52012=>"100111011",
  52013=>"001010110",
  52014=>"011001100",
  52015=>"011001000",
  52016=>"101110010",
  52017=>"111010001",
  52018=>"000010001",
  52019=>"100100011",
  52020=>"101000101",
  52021=>"100101110",
  52022=>"110111011",
  52023=>"001110010",
  52024=>"010001110",
  52025=>"011011100",
  52026=>"001011101",
  52027=>"011001110",
  52028=>"000011000",
  52029=>"111000101",
  52030=>"100101000",
  52031=>"000011001",
  52032=>"001101101",
  52033=>"110111101",
  52034=>"111111001",
  52035=>"111010100",
  52036=>"101010000",
  52037=>"001110010",
  52038=>"010100011",
  52039=>"111011101",
  52040=>"110010111",
  52041=>"010110110",
  52042=>"011010110",
  52043=>"110000110",
  52044=>"011001101",
  52045=>"000000001",
  52046=>"010101011",
  52047=>"000000111",
  52048=>"111001001",
  52049=>"010001010",
  52050=>"111100101",
  52051=>"100000000",
  52052=>"111101100",
  52053=>"010110100",
  52054=>"011010100",
  52055=>"111000011",
  52056=>"100111100",
  52057=>"100010110",
  52058=>"010011011",
  52059=>"110011001",
  52060=>"000000001",
  52061=>"000000011",
  52062=>"011001010",
  52063=>"111111101",
  52064=>"010010101",
  52065=>"111100001",
  52066=>"110110001",
  52067=>"101111100",
  52068=>"001011111",
  52069=>"000011111",
  52070=>"101100111",
  52071=>"010100100",
  52072=>"101111011",
  52073=>"001101110",
  52074=>"100111110",
  52075=>"100011110",
  52076=>"101110000",
  52077=>"000000111",
  52078=>"110111010",
  52079=>"111111100",
  52080=>"100011000",
  52081=>"101010000",
  52082=>"111110101",
  52083=>"101100001",
  52084=>"100100100",
  52085=>"000000010",
  52086=>"010110100",
  52087=>"110101001",
  52088=>"110100011",
  52089=>"011101100",
  52090=>"011010110",
  52091=>"111010001",
  52092=>"100100100",
  52093=>"010110011",
  52094=>"010110011",
  52095=>"001110011",
  52096=>"010111111",
  52097=>"100000111",
  52098=>"010001001",
  52099=>"000111100",
  52100=>"011001111",
  52101=>"110100101",
  52102=>"000101000",
  52103=>"001111111",
  52104=>"011111111",
  52105=>"101111110",
  52106=>"111111100",
  52107=>"000011100",
  52108=>"011010000",
  52109=>"101011111",
  52110=>"011010011",
  52111=>"011001011",
  52112=>"111000000",
  52113=>"001111101",
  52114=>"111001001",
  52115=>"000100101",
  52116=>"101011000",
  52117=>"001101101",
  52118=>"010011111",
  52119=>"101000001",
  52120=>"110111101",
  52121=>"011011000",
  52122=>"010100101",
  52123=>"000100010",
  52124=>"100000010",
  52125=>"110001000",
  52126=>"010111010",
  52127=>"011000011",
  52128=>"000011101",
  52129=>"011111001",
  52130=>"000011000",
  52131=>"001111001",
  52132=>"111100110",
  52133=>"101110011",
  52134=>"101101101",
  52135=>"111011001",
  52136=>"101001110",
  52137=>"010010000",
  52138=>"000111111",
  52139=>"010011011",
  52140=>"010010010",
  52141=>"101011010",
  52142=>"101111000",
  52143=>"100100011",
  52144=>"001110001",
  52145=>"010101100",
  52146=>"011110100",
  52147=>"000100100",
  52148=>"101110101",
  52149=>"110001110",
  52150=>"110011010",
  52151=>"110100001",
  52152=>"100010010",
  52153=>"010000100",
  52154=>"010100000",
  52155=>"000011010",
  52156=>"100001010",
  52157=>"111101110",
  52158=>"111101000",
  52159=>"110110011",
  52160=>"100011111",
  52161=>"011101011",
  52162=>"010110110",
  52163=>"001100011",
  52164=>"101110110",
  52165=>"001000100",
  52166=>"000110000",
  52167=>"001000000",
  52168=>"011001111",
  52169=>"011001110",
  52170=>"100011001",
  52171=>"001101001",
  52172=>"101111111",
  52173=>"010111011",
  52174=>"011111110",
  52175=>"111110011",
  52176=>"000010110",
  52177=>"100001011",
  52178=>"111001110",
  52179=>"110010110",
  52180=>"110100111",
  52181=>"000011100",
  52182=>"111100111",
  52183=>"111111110",
  52184=>"100010000",
  52185=>"000010101",
  52186=>"011110011",
  52187=>"000000011",
  52188=>"000000100",
  52189=>"101100000",
  52190=>"011010111",
  52191=>"010001001",
  52192=>"010110001",
  52193=>"001010011",
  52194=>"111110110",
  52195=>"011001110",
  52196=>"111100000",
  52197=>"011100111",
  52198=>"110001000",
  52199=>"110010100",
  52200=>"001010011",
  52201=>"000001001",
  52202=>"010100111",
  52203=>"100110100",
  52204=>"010110010",
  52205=>"101100000",
  52206=>"001010011",
  52207=>"110001010",
  52208=>"000010010",
  52209=>"101101111",
  52210=>"100101001",
  52211=>"101111011",
  52212=>"001001100",
  52213=>"000000010",
  52214=>"101110110",
  52215=>"011011100",
  52216=>"001001000",
  52217=>"101000111",
  52218=>"101110100",
  52219=>"111101101",
  52220=>"110010110",
  52221=>"110111001",
  52222=>"111100011",
  52223=>"011101100",
  52224=>"111110111",
  52225=>"111000110",
  52226=>"000100110",
  52227=>"111110010",
  52228=>"010100000",
  52229=>"000101001",
  52230=>"000110000",
  52231=>"001000100",
  52232=>"101000000",
  52233=>"001111100",
  52234=>"100101110",
  52235=>"111000010",
  52236=>"000101000",
  52237=>"001000100",
  52238=>"010010100",
  52239=>"001101011",
  52240=>"101000101",
  52241=>"101011111",
  52242=>"111011000",
  52243=>"100110111",
  52244=>"010010001",
  52245=>"101010101",
  52246=>"101000001",
  52247=>"111101100",
  52248=>"000101111",
  52249=>"001000100",
  52250=>"110110000",
  52251=>"101010110",
  52252=>"011101000",
  52253=>"010010101",
  52254=>"110010100",
  52255=>"100101010",
  52256=>"100110001",
  52257=>"000101000",
  52258=>"011011000",
  52259=>"101110101",
  52260=>"000100000",
  52261=>"000110110",
  52262=>"101111001",
  52263=>"101100101",
  52264=>"011010100",
  52265=>"001110001",
  52266=>"000111101",
  52267=>"110011001",
  52268=>"100000001",
  52269=>"000010000",
  52270=>"000000010",
  52271=>"001111010",
  52272=>"011001100",
  52273=>"111010100",
  52274=>"101111011",
  52275=>"011110101",
  52276=>"001001101",
  52277=>"001010011",
  52278=>"000101001",
  52279=>"101010011",
  52280=>"000111000",
  52281=>"100100001",
  52282=>"100101111",
  52283=>"110101011",
  52284=>"011101110",
  52285=>"110011111",
  52286=>"000110010",
  52287=>"100001010",
  52288=>"010010111",
  52289=>"110100101",
  52290=>"100000010",
  52291=>"001001000",
  52292=>"010010101",
  52293=>"101000001",
  52294=>"011111101",
  52295=>"111010000",
  52296=>"101001100",
  52297=>"010100000",
  52298=>"000011111",
  52299=>"010010100",
  52300=>"110101000",
  52301=>"111110000",
  52302=>"011110000",
  52303=>"010010100",
  52304=>"110100100",
  52305=>"100101100",
  52306=>"011111100",
  52307=>"111000101",
  52308=>"110110010",
  52309=>"111100111",
  52310=>"100000100",
  52311=>"001101100",
  52312=>"101100000",
  52313=>"000000101",
  52314=>"100111011",
  52315=>"100001100",
  52316=>"010101101",
  52317=>"110111001",
  52318=>"001101000",
  52319=>"100001011",
  52320=>"000011101",
  52321=>"111110010",
  52322=>"011011110",
  52323=>"001011011",
  52324=>"010111101",
  52325=>"110010000",
  52326=>"101010111",
  52327=>"100000000",
  52328=>"001100000",
  52329=>"010011110",
  52330=>"000000111",
  52331=>"000000000",
  52332=>"011110100",
  52333=>"011100111",
  52334=>"110100110",
  52335=>"111100111",
  52336=>"100010011",
  52337=>"101000110",
  52338=>"011000111",
  52339=>"100100111",
  52340=>"011001101",
  52341=>"100001010",
  52342=>"101000111",
  52343=>"111111011",
  52344=>"110101101",
  52345=>"100011001",
  52346=>"011010000",
  52347=>"011000010",
  52348=>"111100100",
  52349=>"100010000",
  52350=>"001100111",
  52351=>"100001011",
  52352=>"000000100",
  52353=>"011001111",
  52354=>"101011001",
  52355=>"000111100",
  52356=>"000101010",
  52357=>"001101011",
  52358=>"101000100",
  52359=>"101111000",
  52360=>"001010111",
  52361=>"000100111",
  52362=>"001000111",
  52363=>"111100101",
  52364=>"100011011",
  52365=>"100111011",
  52366=>"111011111",
  52367=>"111111010",
  52368=>"110110101",
  52369=>"101011110",
  52370=>"011111101",
  52371=>"101001000",
  52372=>"100001011",
  52373=>"010110011",
  52374=>"000101001",
  52375=>"001110000",
  52376=>"011110000",
  52377=>"011110001",
  52378=>"011000010",
  52379=>"001101111",
  52380=>"101000100",
  52381=>"101110101",
  52382=>"001011010",
  52383=>"101011110",
  52384=>"010001001",
  52385=>"111000010",
  52386=>"110110111",
  52387=>"111001001",
  52388=>"100011000",
  52389=>"101001000",
  52390=>"010010010",
  52391=>"111111101",
  52392=>"100111101",
  52393=>"001011111",
  52394=>"000111011",
  52395=>"000000010",
  52396=>"000111100",
  52397=>"010111011",
  52398=>"000001011",
  52399=>"000100010",
  52400=>"100000010",
  52401=>"101111010",
  52402=>"011001110",
  52403=>"100111101",
  52404=>"011010101",
  52405=>"010110000",
  52406=>"100110110",
  52407=>"110011011",
  52408=>"011100010",
  52409=>"000011001",
  52410=>"100011001",
  52411=>"000101001",
  52412=>"101001110",
  52413=>"101000101",
  52414=>"111000110",
  52415=>"101111000",
  52416=>"101010000",
  52417=>"001111101",
  52418=>"001111000",
  52419=>"011111110",
  52420=>"111001110",
  52421=>"110011010",
  52422=>"100111110",
  52423=>"001101001",
  52424=>"101011011",
  52425=>"111001010",
  52426=>"001011100",
  52427=>"111101111",
  52428=>"111100110",
  52429=>"000101010",
  52430=>"011001110",
  52431=>"101000011",
  52432=>"111101011",
  52433=>"101000101",
  52434=>"101110000",
  52435=>"100110100",
  52436=>"000000101",
  52437=>"010100110",
  52438=>"100000111",
  52439=>"101110010",
  52440=>"011111011",
  52441=>"011001011",
  52442=>"101010011",
  52443=>"010100101",
  52444=>"001000110",
  52445=>"100111101",
  52446=>"010100100",
  52447=>"011001100",
  52448=>"101010100",
  52449=>"101011001",
  52450=>"111001101",
  52451=>"111100101",
  52452=>"101011110",
  52453=>"000000000",
  52454=>"000110111",
  52455=>"100101001",
  52456=>"011101110",
  52457=>"010011110",
  52458=>"001000000",
  52459=>"010110001",
  52460=>"000000111",
  52461=>"011110111",
  52462=>"100001101",
  52463=>"010100101",
  52464=>"100110101",
  52465=>"001110001",
  52466=>"101110000",
  52467=>"101001000",
  52468=>"010010010",
  52469=>"111111100",
  52470=>"011001100",
  52471=>"000000111",
  52472=>"011110101",
  52473=>"001000100",
  52474=>"100111110",
  52475=>"111101010",
  52476=>"100101011",
  52477=>"010010001",
  52478=>"001001001",
  52479=>"110001011",
  52480=>"011111000",
  52481=>"101111100",
  52482=>"101100001",
  52483=>"000010010",
  52484=>"100010100",
  52485=>"111010101",
  52486=>"100010111",
  52487=>"111111111",
  52488=>"111011010",
  52489=>"001101011",
  52490=>"100100011",
  52491=>"011100110",
  52492=>"011111001",
  52493=>"011101010",
  52494=>"001101110",
  52495=>"001010001",
  52496=>"001011101",
  52497=>"110111111",
  52498=>"111111100",
  52499=>"000011010",
  52500=>"111001001",
  52501=>"111100001",
  52502=>"001110011",
  52503=>"011110001",
  52504=>"100011001",
  52505=>"010010000",
  52506=>"011111101",
  52507=>"001001011",
  52508=>"011111000",
  52509=>"101100000",
  52510=>"010101001",
  52511=>"101011111",
  52512=>"011101011",
  52513=>"000001001",
  52514=>"010000001",
  52515=>"110010110",
  52516=>"000000011",
  52517=>"100110100",
  52518=>"001010110",
  52519=>"111011010",
  52520=>"101100110",
  52521=>"110101011",
  52522=>"111000101",
  52523=>"111101111",
  52524=>"011110001",
  52525=>"000111001",
  52526=>"000010010",
  52527=>"111101010",
  52528=>"100001110",
  52529=>"101011111",
  52530=>"111011111",
  52531=>"110000111",
  52532=>"011101111",
  52533=>"010010111",
  52534=>"100011100",
  52535=>"010101010",
  52536=>"001111110",
  52537=>"100100110",
  52538=>"110111001",
  52539=>"011000010",
  52540=>"110011101",
  52541=>"101110010",
  52542=>"001001101",
  52543=>"111111010",
  52544=>"100111111",
  52545=>"000001001",
  52546=>"100011100",
  52547=>"110111010",
  52548=>"000110011",
  52549=>"111010001",
  52550=>"001011110",
  52551=>"000101110",
  52552=>"000110101",
  52553=>"110100101",
  52554=>"001111001",
  52555=>"001101101",
  52556=>"000011010",
  52557=>"010001000",
  52558=>"111111100",
  52559=>"100100100",
  52560=>"110101010",
  52561=>"011110010",
  52562=>"001000110",
  52563=>"010111001",
  52564=>"001000100",
  52565=>"001110011",
  52566=>"011010010",
  52567=>"111111100",
  52568=>"100001010",
  52569=>"001011110",
  52570=>"000010010",
  52571=>"000100111",
  52572=>"111111101",
  52573=>"011101011",
  52574=>"000111000",
  52575=>"001010100",
  52576=>"100000000",
  52577=>"100011111",
  52578=>"101010111",
  52579=>"000100111",
  52580=>"111010101",
  52581=>"010011110",
  52582=>"010010000",
  52583=>"100001111",
  52584=>"101111110",
  52585=>"010111011",
  52586=>"000110100",
  52587=>"101001011",
  52588=>"110000001",
  52589=>"001110100",
  52590=>"010100001",
  52591=>"010110010",
  52592=>"011011010",
  52593=>"011000101",
  52594=>"011011110",
  52595=>"110010100",
  52596=>"101011001",
  52597=>"110110110",
  52598=>"001101101",
  52599=>"001010001",
  52600=>"101100000",
  52601=>"001011001",
  52602=>"110111001",
  52603=>"001100111",
  52604=>"001110010",
  52605=>"001010001",
  52606=>"000110001",
  52607=>"100001000",
  52608=>"111111011",
  52609=>"101110000",
  52610=>"111001110",
  52611=>"000100001",
  52612=>"000111100",
  52613=>"010000100",
  52614=>"111011101",
  52615=>"010100001",
  52616=>"000100001",
  52617=>"111101011",
  52618=>"111110100",
  52619=>"000100101",
  52620=>"111110100",
  52621=>"110110001",
  52622=>"000101000",
  52623=>"100111000",
  52624=>"001101000",
  52625=>"001010000",
  52626=>"011010101",
  52627=>"000110001",
  52628=>"011110101",
  52629=>"111100011",
  52630=>"000011101",
  52631=>"011101110",
  52632=>"101001011",
  52633=>"101001110",
  52634=>"101000110",
  52635=>"110001100",
  52636=>"110100101",
  52637=>"111111011",
  52638=>"111100100",
  52639=>"001010101",
  52640=>"111001100",
  52641=>"010101011",
  52642=>"001111010",
  52643=>"001101111",
  52644=>"100011001",
  52645=>"111000010",
  52646=>"011000100",
  52647=>"000000010",
  52648=>"000000011",
  52649=>"011011001",
  52650=>"100110101",
  52651=>"011001001",
  52652=>"010010000",
  52653=>"111110011",
  52654=>"000011101",
  52655=>"100111010",
  52656=>"001100001",
  52657=>"000011010",
  52658=>"010100101",
  52659=>"101111001",
  52660=>"011010001",
  52661=>"110110111",
  52662=>"001110111",
  52663=>"100001001",
  52664=>"001101001",
  52665=>"000001101",
  52666=>"010100101",
  52667=>"011100101",
  52668=>"101010010",
  52669=>"010010010",
  52670=>"111110110",
  52671=>"110101111",
  52672=>"010100001",
  52673=>"011010110",
  52674=>"001111011",
  52675=>"100010100",
  52676=>"111101001",
  52677=>"000010000",
  52678=>"101101111",
  52679=>"000110110",
  52680=>"111111101",
  52681=>"101110110",
  52682=>"111110110",
  52683=>"111000110",
  52684=>"100011000",
  52685=>"000111110",
  52686=>"110111011",
  52687=>"110000010",
  52688=>"100011000",
  52689=>"100001110",
  52690=>"100101000",
  52691=>"111011010",
  52692=>"101100010",
  52693=>"100000010",
  52694=>"101111110",
  52695=>"101010011",
  52696=>"011111111",
  52697=>"011111010",
  52698=>"100100110",
  52699=>"001000100",
  52700=>"011111101",
  52701=>"010110110",
  52702=>"010010110",
  52703=>"000101101",
  52704=>"010101010",
  52705=>"110111010",
  52706=>"100110101",
  52707=>"111011100",
  52708=>"111101101",
  52709=>"111111101",
  52710=>"001100110",
  52711=>"111101100",
  52712=>"010000101",
  52713=>"111001011",
  52714=>"111100001",
  52715=>"001011111",
  52716=>"111001011",
  52717=>"001010111",
  52718=>"101100000",
  52719=>"000001110",
  52720=>"101101001",
  52721=>"110010100",
  52722=>"101110110",
  52723=>"110110100",
  52724=>"101011010",
  52725=>"111100101",
  52726=>"100010001",
  52727=>"101010111",
  52728=>"001110010",
  52729=>"000100110",
  52730=>"000010110",
  52731=>"111100001",
  52732=>"001100100",
  52733=>"010000100",
  52734=>"010001010",
  52735=>"000000101",
  52736=>"000101110",
  52737=>"010011000",
  52738=>"010111100",
  52739=>"000000111",
  52740=>"111110100",
  52741=>"110000010",
  52742=>"011001111",
  52743=>"101111000",
  52744=>"001111011",
  52745=>"001111111",
  52746=>"111101011",
  52747=>"000110110",
  52748=>"010001110",
  52749=>"110111001",
  52750=>"011110101",
  52751=>"011010011",
  52752=>"011011000",
  52753=>"111010011",
  52754=>"010111001",
  52755=>"111010100",
  52756=>"011100001",
  52757=>"011100101",
  52758=>"110001100",
  52759=>"000011111",
  52760=>"010111011",
  52761=>"111101011",
  52762=>"000010100",
  52763=>"100001101",
  52764=>"011101000",
  52765=>"011010000",
  52766=>"101011101",
  52767=>"100111010",
  52768=>"111010010",
  52769=>"000101010",
  52770=>"111111101",
  52771=>"110011100",
  52772=>"100010100",
  52773=>"001100000",
  52774=>"101001011",
  52775=>"000101100",
  52776=>"000111011",
  52777=>"001111010",
  52778=>"101011011",
  52779=>"100111000",
  52780=>"010010100",
  52781=>"110111000",
  52782=>"001000110",
  52783=>"000101111",
  52784=>"000001101",
  52785=>"010110100",
  52786=>"100100011",
  52787=>"100011100",
  52788=>"110000011",
  52789=>"110000101",
  52790=>"011000110",
  52791=>"100010100",
  52792=>"110101111",
  52793=>"010001010",
  52794=>"101100000",
  52795=>"001110001",
  52796=>"110001001",
  52797=>"000011010",
  52798=>"111101010",
  52799=>"010010000",
  52800=>"011111001",
  52801=>"100111011",
  52802=>"001110100",
  52803=>"010111111",
  52804=>"001100000",
  52805=>"101100111",
  52806=>"110101011",
  52807=>"000111110",
  52808=>"010010100",
  52809=>"111111110",
  52810=>"110010010",
  52811=>"011010011",
  52812=>"110010001",
  52813=>"000010010",
  52814=>"100001111",
  52815=>"000010011",
  52816=>"110010110",
  52817=>"100100000",
  52818=>"000100000",
  52819=>"100111010",
  52820=>"111100000",
  52821=>"110010001",
  52822=>"110000011",
  52823=>"100110111",
  52824=>"110111110",
  52825=>"010000100",
  52826=>"111111011",
  52827=>"001011000",
  52828=>"101100011",
  52829=>"000100111",
  52830=>"111101000",
  52831=>"111101000",
  52832=>"110101001",
  52833=>"100100010",
  52834=>"101101001",
  52835=>"010011110",
  52836=>"001011001",
  52837=>"011101100",
  52838=>"010001010",
  52839=>"000010110",
  52840=>"100110100",
  52841=>"100111110",
  52842=>"111010011",
  52843=>"011010001",
  52844=>"000110101",
  52845=>"000111100",
  52846=>"100110001",
  52847=>"100110111",
  52848=>"000110010",
  52849=>"100101001",
  52850=>"010001001",
  52851=>"100100100",
  52852=>"101110010",
  52853=>"101010111",
  52854=>"001011100",
  52855=>"111001001",
  52856=>"001111000",
  52857=>"110010101",
  52858=>"111011110",
  52859=>"000001100",
  52860=>"101000000",
  52861=>"000011011",
  52862=>"101111001",
  52863=>"110011111",
  52864=>"000010110",
  52865=>"010001101",
  52866=>"111101000",
  52867=>"001101000",
  52868=>"001001000",
  52869=>"000101011",
  52870=>"100100100",
  52871=>"100001011",
  52872=>"100100011",
  52873=>"000110010",
  52874=>"111101100",
  52875=>"101100110",
  52876=>"100001000",
  52877=>"100111010",
  52878=>"111101110",
  52879=>"110000111",
  52880=>"011101010",
  52881=>"110111000",
  52882=>"000011000",
  52883=>"111111011",
  52884=>"001001100",
  52885=>"101100010",
  52886=>"000011011",
  52887=>"001100111",
  52888=>"010100101",
  52889=>"111011000",
  52890=>"010010111",
  52891=>"100110000",
  52892=>"100001101",
  52893=>"111001000",
  52894=>"101101011",
  52895=>"101110101",
  52896=>"101010011",
  52897=>"110100000",
  52898=>"000110111",
  52899=>"010000011",
  52900=>"111111101",
  52901=>"110000010",
  52902=>"110011100",
  52903=>"101101011",
  52904=>"110001111",
  52905=>"011011100",
  52906=>"000101110",
  52907=>"001001001",
  52908=>"000001111",
  52909=>"001000110",
  52910=>"100111101",
  52911=>"000001101",
  52912=>"100100110",
  52913=>"010110101",
  52914=>"001010110",
  52915=>"001101000",
  52916=>"110001111",
  52917=>"110100110",
  52918=>"111010111",
  52919=>"000110110",
  52920=>"110000001",
  52921=>"110100111",
  52922=>"111000111",
  52923=>"011100111",
  52924=>"001111010",
  52925=>"000000000",
  52926=>"010011101",
  52927=>"001111101",
  52928=>"110110000",
  52929=>"001000110",
  52930=>"010011100",
  52931=>"001100100",
  52932=>"000100011",
  52933=>"101110001",
  52934=>"111000100",
  52935=>"000111101",
  52936=>"101110010",
  52937=>"010010110",
  52938=>"010101100",
  52939=>"000111100",
  52940=>"111111010",
  52941=>"010100010",
  52942=>"111111011",
  52943=>"110111101",
  52944=>"001010100",
  52945=>"100000101",
  52946=>"101010101",
  52947=>"100001010",
  52948=>"000101000",
  52949=>"010011100",
  52950=>"010110011",
  52951=>"110001001",
  52952=>"001111011",
  52953=>"011111110",
  52954=>"010110111",
  52955=>"001010001",
  52956=>"101110000",
  52957=>"000100111",
  52958=>"111001000",
  52959=>"111101010",
  52960=>"101111111",
  52961=>"110011101",
  52962=>"100111000",
  52963=>"000100011",
  52964=>"101110000",
  52965=>"110101000",
  52966=>"101010011",
  52967=>"000000110",
  52968=>"010110101",
  52969=>"011000010",
  52970=>"010000100",
  52971=>"100011111",
  52972=>"110011110",
  52973=>"001100100",
  52974=>"011011000",
  52975=>"110011010",
  52976=>"110000111",
  52977=>"010011101",
  52978=>"011101101",
  52979=>"001001101",
  52980=>"101000010",
  52981=>"000000010",
  52982=>"110111100",
  52983=>"010011110",
  52984=>"001010110",
  52985=>"100001111",
  52986=>"000000101",
  52987=>"001001011",
  52988=>"101000011",
  52989=>"001101010",
  52990=>"011100111",
  52991=>"000111111",
  52992=>"000000101",
  52993=>"100000100",
  52994=>"010100100",
  52995=>"000100000",
  52996=>"001110111",
  52997=>"011000111",
  52998=>"001011000",
  52999=>"111111001",
  53000=>"101011111",
  53001=>"001001010",
  53002=>"101010010",
  53003=>"111100011",
  53004=>"010101000",
  53005=>"101000001",
  53006=>"111110101",
  53007=>"111110100",
  53008=>"111111111",
  53009=>"010111000",
  53010=>"011001111",
  53011=>"110001000",
  53012=>"000100001",
  53013=>"110111011",
  53014=>"000101100",
  53015=>"110111111",
  53016=>"011101110",
  53017=>"000110011",
  53018=>"100001011",
  53019=>"111111111",
  53020=>"000110111",
  53021=>"011010010",
  53022=>"011011111",
  53023=>"001110000",
  53024=>"010001101",
  53025=>"111110010",
  53026=>"000100100",
  53027=>"010000001",
  53028=>"001010111",
  53029=>"001110101",
  53030=>"010011101",
  53031=>"100010010",
  53032=>"110111011",
  53033=>"000101001",
  53034=>"111111001",
  53035=>"110000011",
  53036=>"010000000",
  53037=>"011101000",
  53038=>"001100000",
  53039=>"000010100",
  53040=>"001110000",
  53041=>"001110110",
  53042=>"010101100",
  53043=>"000001000",
  53044=>"111010000",
  53045=>"101001111",
  53046=>"010110001",
  53047=>"010000000",
  53048=>"101011100",
  53049=>"110001001",
  53050=>"000001100",
  53051=>"000001100",
  53052=>"101010100",
  53053=>"000001000",
  53054=>"010011100",
  53055=>"010000100",
  53056=>"010101010",
  53057=>"001000000",
  53058=>"110010011",
  53059=>"001011110",
  53060=>"111101110",
  53061=>"010010110",
  53062=>"101100011",
  53063=>"000010010",
  53064=>"011011000",
  53065=>"100100111",
  53066=>"011001001",
  53067=>"111110010",
  53068=>"000111111",
  53069=>"000000110",
  53070=>"111100011",
  53071=>"001111001",
  53072=>"110000001",
  53073=>"100010101",
  53074=>"111101010",
  53075=>"011000111",
  53076=>"000001000",
  53077=>"101010110",
  53078=>"101001110",
  53079=>"001010110",
  53080=>"000110000",
  53081=>"100100101",
  53082=>"010001001",
  53083=>"001001111",
  53084=>"100010010",
  53085=>"001000011",
  53086=>"110110010",
  53087=>"100111111",
  53088=>"111001100",
  53089=>"111011100",
  53090=>"001000100",
  53091=>"000001010",
  53092=>"011100101",
  53093=>"010011000",
  53094=>"000101111",
  53095=>"100110001",
  53096=>"111110100",
  53097=>"101101101",
  53098=>"101010110",
  53099=>"100110100",
  53100=>"000001100",
  53101=>"010011111",
  53102=>"000000110",
  53103=>"011111110",
  53104=>"010011110",
  53105=>"010101000",
  53106=>"000001010",
  53107=>"010001010",
  53108=>"000110000",
  53109=>"001011010",
  53110=>"100000000",
  53111=>"111000000",
  53112=>"101100001",
  53113=>"010110001",
  53114=>"100000100",
  53115=>"011101101",
  53116=>"110100001",
  53117=>"111000110",
  53118=>"101100010",
  53119=>"101110111",
  53120=>"101100111",
  53121=>"100000101",
  53122=>"000000010",
  53123=>"011110101",
  53124=>"110111111",
  53125=>"010001110",
  53126=>"110101111",
  53127=>"001101010",
  53128=>"100111111",
  53129=>"011110110",
  53130=>"110110111",
  53131=>"010101100",
  53132=>"001010010",
  53133=>"010101000",
  53134=>"010101000",
  53135=>"001110001",
  53136=>"001010110",
  53137=>"100010011",
  53138=>"001111001",
  53139=>"011010100",
  53140=>"011000110",
  53141=>"111010001",
  53142=>"101111100",
  53143=>"110001100",
  53144=>"101100010",
  53145=>"110011000",
  53146=>"100000000",
  53147=>"001000010",
  53148=>"100100111",
  53149=>"010110010",
  53150=>"000100101",
  53151=>"000111110",
  53152=>"101111100",
  53153=>"000111000",
  53154=>"111011101",
  53155=>"100111110",
  53156=>"001110010",
  53157=>"001101010",
  53158=>"110110100",
  53159=>"001101000",
  53160=>"100101110",
  53161=>"000001110",
  53162=>"010000011",
  53163=>"100000100",
  53164=>"010101111",
  53165=>"101000011",
  53166=>"101010000",
  53167=>"100010101",
  53168=>"010000111",
  53169=>"010000110",
  53170=>"001111010",
  53171=>"101010011",
  53172=>"110000101",
  53173=>"001001110",
  53174=>"010101010",
  53175=>"100100111",
  53176=>"000010111",
  53177=>"011111010",
  53178=>"100000111",
  53179=>"111001100",
  53180=>"110101111",
  53181=>"000101100",
  53182=>"110101010",
  53183=>"000101100",
  53184=>"110101011",
  53185=>"111000010",
  53186=>"001010000",
  53187=>"000110110",
  53188=>"110011001",
  53189=>"001000011",
  53190=>"010100010",
  53191=>"011101110",
  53192=>"110101000",
  53193=>"111001010",
  53194=>"011000110",
  53195=>"100111011",
  53196=>"000110100",
  53197=>"000100000",
  53198=>"101010010",
  53199=>"001011101",
  53200=>"010000110",
  53201=>"111001011",
  53202=>"011101011",
  53203=>"010011000",
  53204=>"000111101",
  53205=>"001010101",
  53206=>"111000000",
  53207=>"001111011",
  53208=>"101110011",
  53209=>"110000000",
  53210=>"010001111",
  53211=>"010011001",
  53212=>"110000110",
  53213=>"101011111",
  53214=>"111010101",
  53215=>"110101110",
  53216=>"101001101",
  53217=>"110001111",
  53218=>"111111101",
  53219=>"110110110",
  53220=>"100001100",
  53221=>"100101111",
  53222=>"111010000",
  53223=>"110001000",
  53224=>"100010000",
  53225=>"010110101",
  53226=>"010110101",
  53227=>"001101001",
  53228=>"110010110",
  53229=>"110110001",
  53230=>"001110101",
  53231=>"000011101",
  53232=>"111010001",
  53233=>"100000001",
  53234=>"100111101",
  53235=>"001000101",
  53236=>"111110101",
  53237=>"000111101",
  53238=>"010110010",
  53239=>"110011000",
  53240=>"001101001",
  53241=>"001010011",
  53242=>"111101010",
  53243=>"111010101",
  53244=>"110000001",
  53245=>"010000010",
  53246=>"111101110",
  53247=>"011101111",
  53248=>"111100000",
  53249=>"000101001",
  53250=>"111110111",
  53251=>"000100100",
  53252=>"001111001",
  53253=>"011111111",
  53254=>"110010010",
  53255=>"001001101",
  53256=>"110110011",
  53257=>"010101111",
  53258=>"010001001",
  53259=>"101010101",
  53260=>"110110111",
  53261=>"100000010",
  53262=>"111010001",
  53263=>"000010100",
  53264=>"101110011",
  53265=>"010000110",
  53266=>"111101000",
  53267=>"100110110",
  53268=>"010111001",
  53269=>"110010111",
  53270=>"001111011",
  53271=>"111000000",
  53272=>"110010111",
  53273=>"101000000",
  53274=>"100101100",
  53275=>"101101110",
  53276=>"101111101",
  53277=>"101001001",
  53278=>"111000011",
  53279=>"110110100",
  53280=>"001001001",
  53281=>"101001001",
  53282=>"111001110",
  53283=>"111011111",
  53284=>"110111111",
  53285=>"010001101",
  53286=>"111110100",
  53287=>"101011111",
  53288=>"000001010",
  53289=>"000001100",
  53290=>"010001010",
  53291=>"000110111",
  53292=>"100100000",
  53293=>"011111001",
  53294=>"101010001",
  53295=>"101110111",
  53296=>"111011100",
  53297=>"100110000",
  53298=>"010000010",
  53299=>"011110110",
  53300=>"010000010",
  53301=>"001010010",
  53302=>"110111111",
  53303=>"110001000",
  53304=>"010110111",
  53305=>"100110000",
  53306=>"101000101",
  53307=>"001111111",
  53308=>"000010010",
  53309=>"101111001",
  53310=>"011000100",
  53311=>"001000000",
  53312=>"011011001",
  53313=>"010000100",
  53314=>"001011110",
  53315=>"001001010",
  53316=>"000111100",
  53317=>"000110110",
  53318=>"010011010",
  53319=>"110110011",
  53320=>"010011000",
  53321=>"011010000",
  53322=>"000001011",
  53323=>"001010000",
  53324=>"111110000",
  53325=>"111010010",
  53326=>"010001100",
  53327=>"010100100",
  53328=>"010010011",
  53329=>"001101101",
  53330=>"000001100",
  53331=>"111111100",
  53332=>"000110100",
  53333=>"001011110",
  53334=>"000001110",
  53335=>"010010000",
  53336=>"000011001",
  53337=>"010000000",
  53338=>"000001111",
  53339=>"101100011",
  53340=>"001101010",
  53341=>"000000111",
  53342=>"000010111",
  53343=>"111110101",
  53344=>"000111101",
  53345=>"111001111",
  53346=>"100101100",
  53347=>"001110000",
  53348=>"000110000",
  53349=>"011110110",
  53350=>"111011100",
  53351=>"011111010",
  53352=>"000110101",
  53353=>"011100001",
  53354=>"010000011",
  53355=>"011101101",
  53356=>"100100001",
  53357=>"101101010",
  53358=>"001001110",
  53359=>"100001011",
  53360=>"000100101",
  53361=>"001001001",
  53362=>"001011001",
  53363=>"111110111",
  53364=>"001011101",
  53365=>"110110010",
  53366=>"000100100",
  53367=>"011000010",
  53368=>"101100010",
  53369=>"100100001",
  53370=>"010110011",
  53371=>"110110001",
  53372=>"011101101",
  53373=>"010101111",
  53374=>"000110101",
  53375=>"010101110",
  53376=>"010011000",
  53377=>"001001001",
  53378=>"011000100",
  53379=>"011100000",
  53380=>"110010111",
  53381=>"101011010",
  53382=>"100010110",
  53383=>"101010111",
  53384=>"101001110",
  53385=>"010111011",
  53386=>"010111110",
  53387=>"001010000",
  53388=>"010110001",
  53389=>"101000011",
  53390=>"111111100",
  53391=>"110000011",
  53392=>"010001000",
  53393=>"110110111",
  53394=>"101000101",
  53395=>"111110011",
  53396=>"111011000",
  53397=>"011000011",
  53398=>"100101101",
  53399=>"000000101",
  53400=>"100000010",
  53401=>"110011001",
  53402=>"101110010",
  53403=>"001001000",
  53404=>"110100101",
  53405=>"010111111",
  53406=>"101111000",
  53407=>"011110111",
  53408=>"001000010",
  53409=>"111100100",
  53410=>"110110001",
  53411=>"101001101",
  53412=>"010011010",
  53413=>"000000011",
  53414=>"101101001",
  53415=>"111001111",
  53416=>"110111000",
  53417=>"000000000",
  53418=>"111101111",
  53419=>"101000110",
  53420=>"000111101",
  53421=>"010100001",
  53422=>"001110010",
  53423=>"101110101",
  53424=>"001101100",
  53425=>"110111000",
  53426=>"010001011",
  53427=>"100000001",
  53428=>"101100010",
  53429=>"101000110",
  53430=>"000110001",
  53431=>"001101000",
  53432=>"000000101",
  53433=>"110001010",
  53434=>"010001001",
  53435=>"010111011",
  53436=>"100011101",
  53437=>"001011101",
  53438=>"101010000",
  53439=>"101110110",
  53440=>"000000010",
  53441=>"100101100",
  53442=>"100001010",
  53443=>"000011000",
  53444=>"101110000",
  53445=>"110111011",
  53446=>"011100001",
  53447=>"111111111",
  53448=>"111101100",
  53449=>"111111011",
  53450=>"110110111",
  53451=>"101010001",
  53452=>"100011001",
  53453=>"000100001",
  53454=>"000010101",
  53455=>"111010111",
  53456=>"001000111",
  53457=>"101010010",
  53458=>"000000011",
  53459=>"011001101",
  53460=>"111001000",
  53461=>"100111100",
  53462=>"000100011",
  53463=>"010110011",
  53464=>"000000100",
  53465=>"000001100",
  53466=>"000001100",
  53467=>"110000001",
  53468=>"110000101",
  53469=>"001110101",
  53470=>"111101101",
  53471=>"110111010",
  53472=>"100011100",
  53473=>"000110101",
  53474=>"001101010",
  53475=>"101110000",
  53476=>"000101010",
  53477=>"001001101",
  53478=>"001001001",
  53479=>"101101001",
  53480=>"001011010",
  53481=>"011101111",
  53482=>"101110010",
  53483=>"000001111",
  53484=>"100000000",
  53485=>"001111011",
  53486=>"111101000",
  53487=>"000100001",
  53488=>"010010000",
  53489=>"011101010",
  53490=>"110110000",
  53491=>"101100101",
  53492=>"000100110",
  53493=>"100011110",
  53494=>"010110100",
  53495=>"100100000",
  53496=>"000111101",
  53497=>"100111110",
  53498=>"001001010",
  53499=>"001101001",
  53500=>"110000010",
  53501=>"001110010",
  53502=>"111011001",
  53503=>"100100111",
  53504=>"101000111",
  53505=>"001001001",
  53506=>"000000010",
  53507=>"000100001",
  53508=>"000101111",
  53509=>"000101101",
  53510=>"000101100",
  53511=>"100011111",
  53512=>"000100100",
  53513=>"001001010",
  53514=>"010001111",
  53515=>"111010011",
  53516=>"110000001",
  53517=>"000000101",
  53518=>"101110000",
  53519=>"110000101",
  53520=>"010100010",
  53521=>"000000000",
  53522=>"000011010",
  53523=>"101011101",
  53524=>"001010001",
  53525=>"001011110",
  53526=>"100110100",
  53527=>"000101001",
  53528=>"011111001",
  53529=>"010110100",
  53530=>"000001011",
  53531=>"000100100",
  53532=>"010010101",
  53533=>"110110000",
  53534=>"110100010",
  53535=>"000111110",
  53536=>"101010010",
  53537=>"110010010",
  53538=>"000100001",
  53539=>"011001111",
  53540=>"000000000",
  53541=>"100011000",
  53542=>"100000010",
  53543=>"110111011",
  53544=>"100000100",
  53545=>"000001110",
  53546=>"111000000",
  53547=>"011000010",
  53548=>"011011110",
  53549=>"001100111",
  53550=>"101010101",
  53551=>"010111001",
  53552=>"010001101",
  53553=>"011001000",
  53554=>"000100011",
  53555=>"010100001",
  53556=>"111100101",
  53557=>"110100101",
  53558=>"001011011",
  53559=>"111001101",
  53560=>"000001001",
  53561=>"010110110",
  53562=>"001010110",
  53563=>"110110110",
  53564=>"101100101",
  53565=>"111110011",
  53566=>"010110100",
  53567=>"001001111",
  53568=>"111101111",
  53569=>"101111010",
  53570=>"111111111",
  53571=>"011011001",
  53572=>"101010101",
  53573=>"100011110",
  53574=>"000000001",
  53575=>"010100100",
  53576=>"110011110",
  53577=>"100010001",
  53578=>"010011010",
  53579=>"000000110",
  53580=>"010101101",
  53581=>"011101000",
  53582=>"000010100",
  53583=>"110001011",
  53584=>"110011010",
  53585=>"100001010",
  53586=>"101101101",
  53587=>"100100111",
  53588=>"111111011",
  53589=>"101011110",
  53590=>"110011100",
  53591=>"101100101",
  53592=>"001001101",
  53593=>"001011000",
  53594=>"101100111",
  53595=>"101110011",
  53596=>"011000110",
  53597=>"110010111",
  53598=>"000001010",
  53599=>"000011001",
  53600=>"001011100",
  53601=>"000100010",
  53602=>"001010100",
  53603=>"000000100",
  53604=>"000100100",
  53605=>"110010100",
  53606=>"111001000",
  53607=>"111111000",
  53608=>"011110000",
  53609=>"100000101",
  53610=>"000101010",
  53611=>"001010100",
  53612=>"011111010",
  53613=>"110101011",
  53614=>"001101000",
  53615=>"001111100",
  53616=>"001000100",
  53617=>"010010101",
  53618=>"100011110",
  53619=>"001110001",
  53620=>"100010111",
  53621=>"000100011",
  53622=>"100001111",
  53623=>"000000101",
  53624=>"010110111",
  53625=>"000111001",
  53626=>"000101100",
  53627=>"001101010",
  53628=>"000111010",
  53629=>"111111110",
  53630=>"011111110",
  53631=>"011100100",
  53632=>"000110000",
  53633=>"001010110",
  53634=>"100111111",
  53635=>"001100111",
  53636=>"100101000",
  53637=>"001010001",
  53638=>"101101110",
  53639=>"111000110",
  53640=>"000000010",
  53641=>"010000011",
  53642=>"111100100",
  53643=>"101000111",
  53644=>"000110100",
  53645=>"101111011",
  53646=>"100101001",
  53647=>"110001010",
  53648=>"000000000",
  53649=>"000000011",
  53650=>"000000110",
  53651=>"111110111",
  53652=>"011010000",
  53653=>"110010111",
  53654=>"110101101",
  53655=>"010100100",
  53656=>"000111000",
  53657=>"110000100",
  53658=>"110011110",
  53659=>"010001101",
  53660=>"000111000",
  53661=>"010101001",
  53662=>"011000011",
  53663=>"111011111",
  53664=>"110100100",
  53665=>"001011100",
  53666=>"000100010",
  53667=>"011101010",
  53668=>"110111100",
  53669=>"110100110",
  53670=>"110111101",
  53671=>"111100000",
  53672=>"110110010",
  53673=>"100111010",
  53674=>"100110100",
  53675=>"011000001",
  53676=>"100111110",
  53677=>"110010110",
  53678=>"000101010",
  53679=>"100010100",
  53680=>"100101101",
  53681=>"110101110",
  53682=>"101111100",
  53683=>"011110110",
  53684=>"100010100",
  53685=>"000110100",
  53686=>"000111101",
  53687=>"101010001",
  53688=>"100010000",
  53689=>"010010110",
  53690=>"101100000",
  53691=>"000001000",
  53692=>"111110010",
  53693=>"101001111",
  53694=>"000000100",
  53695=>"011000111",
  53696=>"110101001",
  53697=>"011011100",
  53698=>"011010001",
  53699=>"010010110",
  53700=>"101011000",
  53701=>"111110001",
  53702=>"110111101",
  53703=>"010000011",
  53704=>"110001101",
  53705=>"111101111",
  53706=>"110100110",
  53707=>"010011000",
  53708=>"110011010",
  53709=>"010111001",
  53710=>"000000000",
  53711=>"000000110",
  53712=>"000001110",
  53713=>"011001001",
  53714=>"001100010",
  53715=>"000100101",
  53716=>"101011000",
  53717=>"101110111",
  53718=>"000111100",
  53719=>"001001100",
  53720=>"000101001",
  53721=>"001101010",
  53722=>"001110110",
  53723=>"010100101",
  53724=>"010010100",
  53725=>"110101010",
  53726=>"110111110",
  53727=>"101101110",
  53728=>"001101101",
  53729=>"001110110",
  53730=>"101001110",
  53731=>"111001000",
  53732=>"100101001",
  53733=>"100101001",
  53734=>"000110011",
  53735=>"111011100",
  53736=>"011101001",
  53737=>"110010111",
  53738=>"111110000",
  53739=>"011010011",
  53740=>"111100101",
  53741=>"011011100",
  53742=>"110010100",
  53743=>"001000000",
  53744=>"000000100",
  53745=>"101010010",
  53746=>"010010000",
  53747=>"001100010",
  53748=>"011101111",
  53749=>"011001111",
  53750=>"100011010",
  53751=>"011100011",
  53752=>"011101101",
  53753=>"001110000",
  53754=>"000100011",
  53755=>"111001111",
  53756=>"011100111",
  53757=>"000010111",
  53758=>"001011101",
  53759=>"101000000",
  53760=>"010011000",
  53761=>"100000111",
  53762=>"110000111",
  53763=>"110000000",
  53764=>"110100111",
  53765=>"010001000",
  53766=>"111011101",
  53767=>"110111000",
  53768=>"101000000",
  53769=>"011111000",
  53770=>"111010111",
  53771=>"000100100",
  53772=>"011010010",
  53773=>"110001110",
  53774=>"111000000",
  53775=>"001000110",
  53776=>"011011011",
  53777=>"011110011",
  53778=>"010110111",
  53779=>"010110001",
  53780=>"111010001",
  53781=>"011011000",
  53782=>"100101011",
  53783=>"001011000",
  53784=>"101001010",
  53785=>"100010000",
  53786=>"101000001",
  53787=>"110011100",
  53788=>"100000010",
  53789=>"001100010",
  53790=>"100111110",
  53791=>"010011111",
  53792=>"101000001",
  53793=>"010000000",
  53794=>"100010001",
  53795=>"111001010",
  53796=>"110000101",
  53797=>"001100011",
  53798=>"101001100",
  53799=>"110101000",
  53800=>"000111010",
  53801=>"111000011",
  53802=>"010100101",
  53803=>"100001111",
  53804=>"000100000",
  53805=>"110001110",
  53806=>"110010010",
  53807=>"100011101",
  53808=>"010100010",
  53809=>"110111111",
  53810=>"100001100",
  53811=>"010101000",
  53812=>"000101011",
  53813=>"011011111",
  53814=>"000101100",
  53815=>"111001111",
  53816=>"101001110",
  53817=>"110101110",
  53818=>"010101011",
  53819=>"011001001",
  53820=>"001100100",
  53821=>"000010111",
  53822=>"101110000",
  53823=>"001010110",
  53824=>"111101011",
  53825=>"000111001",
  53826=>"111100101",
  53827=>"101100001",
  53828=>"010110110",
  53829=>"001010110",
  53830=>"100110110",
  53831=>"101100101",
  53832=>"110001100",
  53833=>"001010010",
  53834=>"101001110",
  53835=>"101100001",
  53836=>"101001011",
  53837=>"111110000",
  53838=>"100011101",
  53839=>"100000001",
  53840=>"100110011",
  53841=>"000100100",
  53842=>"111100110",
  53843=>"011010000",
  53844=>"010010010",
  53845=>"010101010",
  53846=>"010101100",
  53847=>"011000000",
  53848=>"001100011",
  53849=>"011000010",
  53850=>"000010010",
  53851=>"000011000",
  53852=>"111001011",
  53853=>"001100111",
  53854=>"011001111",
  53855=>"111101100",
  53856=>"000010101",
  53857=>"001110101",
  53858=>"010011000",
  53859=>"100011010",
  53860=>"111010111",
  53861=>"001001011",
  53862=>"010110001",
  53863=>"011100000",
  53864=>"001010011",
  53865=>"001101101",
  53866=>"111111001",
  53867=>"111100110",
  53868=>"100100001",
  53869=>"000100010",
  53870=>"101010000",
  53871=>"010010001",
  53872=>"010110110",
  53873=>"000000000",
  53874=>"010100110",
  53875=>"101101101",
  53876=>"000001101",
  53877=>"101101010",
  53878=>"110111110",
  53879=>"000100111",
  53880=>"001001000",
  53881=>"110001100",
  53882=>"011011111",
  53883=>"100001001",
  53884=>"100010001",
  53885=>"111000100",
  53886=>"110101111",
  53887=>"110110110",
  53888=>"000100100",
  53889=>"011100111",
  53890=>"101111110",
  53891=>"100000000",
  53892=>"010000111",
  53893=>"000110000",
  53894=>"111011010",
  53895=>"001110001",
  53896=>"100111101",
  53897=>"100000001",
  53898=>"011001110",
  53899=>"011100010",
  53900=>"000101100",
  53901=>"110111001",
  53902=>"001100000",
  53903=>"110111111",
  53904=>"000011101",
  53905=>"011111000",
  53906=>"111000000",
  53907=>"001110011",
  53908=>"001101100",
  53909=>"111101001",
  53910=>"110110010",
  53911=>"010000000",
  53912=>"110100100",
  53913=>"011001010",
  53914=>"101111111",
  53915=>"011000101",
  53916=>"101000000",
  53917=>"010011100",
  53918=>"000010100",
  53919=>"010110010",
  53920=>"101001111",
  53921=>"011100001",
  53922=>"011001010",
  53923=>"001100101",
  53924=>"000101001",
  53925=>"110100100",
  53926=>"001000000",
  53927=>"010100011",
  53928=>"100110100",
  53929=>"111010101",
  53930=>"100111111",
  53931=>"001001101",
  53932=>"000001001",
  53933=>"010010010",
  53934=>"011000111",
  53935=>"010010001",
  53936=>"001011001",
  53937=>"110111100",
  53938=>"110101111",
  53939=>"001000000",
  53940=>"101000010",
  53941=>"001100011",
  53942=>"110110001",
  53943=>"111010100",
  53944=>"010101010",
  53945=>"110010011",
  53946=>"000001111",
  53947=>"001110010",
  53948=>"010110111",
  53949=>"100100100",
  53950=>"101010100",
  53951=>"111100111",
  53952=>"010111110",
  53953=>"100001001",
  53954=>"110110010",
  53955=>"010010011",
  53956=>"010011101",
  53957=>"111101000",
  53958=>"000101110",
  53959=>"111001100",
  53960=>"001111110",
  53961=>"000101011",
  53962=>"110110100",
  53963=>"010101101",
  53964=>"111101000",
  53965=>"100111010",
  53966=>"000110011",
  53967=>"011101111",
  53968=>"110110010",
  53969=>"110001011",
  53970=>"110011111",
  53971=>"011000000",
  53972=>"001101101",
  53973=>"010000010",
  53974=>"010100111",
  53975=>"001100011",
  53976=>"010001100",
  53977=>"110011011",
  53978=>"000001110",
  53979=>"000001000",
  53980=>"011000010",
  53981=>"000010111",
  53982=>"000101101",
  53983=>"111011100",
  53984=>"011100101",
  53985=>"010101011",
  53986=>"110000010",
  53987=>"111011011",
  53988=>"011111010",
  53989=>"100111110",
  53990=>"001100000",
  53991=>"011100000",
  53992=>"000000001",
  53993=>"011101000",
  53994=>"011010000",
  53995=>"111111101",
  53996=>"000011000",
  53997=>"001000011",
  53998=>"110111001",
  53999=>"000001010",
  54000=>"000000111",
  54001=>"101101110",
  54002=>"100000111",
  54003=>"110110001",
  54004=>"110010000",
  54005=>"001011001",
  54006=>"000000001",
  54007=>"100011111",
  54008=>"010010100",
  54009=>"101101110",
  54010=>"111101101",
  54011=>"100100110",
  54012=>"100101111",
  54013=>"010110001",
  54014=>"000110001",
  54015=>"010101000",
  54016=>"011100001",
  54017=>"000100100",
  54018=>"110101100",
  54019=>"111100101",
  54020=>"111110101",
  54021=>"001000011",
  54022=>"010111010",
  54023=>"101101011",
  54024=>"110011011",
  54025=>"101101100",
  54026=>"111000010",
  54027=>"110000101",
  54028=>"111011000",
  54029=>"001111111",
  54030=>"110010101",
  54031=>"001011110",
  54032=>"111001101",
  54033=>"100000100",
  54034=>"000100101",
  54035=>"001011100",
  54036=>"011111011",
  54037=>"001000100",
  54038=>"011011101",
  54039=>"010100010",
  54040=>"110000100",
  54041=>"001011001",
  54042=>"010000001",
  54043=>"000110011",
  54044=>"111010000",
  54045=>"110010011",
  54046=>"111011110",
  54047=>"011010101",
  54048=>"100011000",
  54049=>"001110100",
  54050=>"110001101",
  54051=>"100110100",
  54052=>"100000100",
  54053=>"010100110",
  54054=>"001011001",
  54055=>"110111010",
  54056=>"101101001",
  54057=>"010000010",
  54058=>"100110011",
  54059=>"011110001",
  54060=>"101111100",
  54061=>"001000010",
  54062=>"101101110",
  54063=>"101100111",
  54064=>"010000001",
  54065=>"101101010",
  54066=>"000100100",
  54067=>"010001011",
  54068=>"100100110",
  54069=>"000101110",
  54070=>"100011000",
  54071=>"011101000",
  54072=>"110001011",
  54073=>"101110110",
  54074=>"011000011",
  54075=>"100100000",
  54076=>"111100011",
  54077=>"101011001",
  54078=>"111001100",
  54079=>"110000011",
  54080=>"000010111",
  54081=>"111011111",
  54082=>"110111010",
  54083=>"101010010",
  54084=>"100110101",
  54085=>"100010111",
  54086=>"000011000",
  54087=>"100110110",
  54088=>"000010000",
  54089=>"110011101",
  54090=>"101110011",
  54091=>"100101101",
  54092=>"011010100",
  54093=>"100111010",
  54094=>"110010100",
  54095=>"011101110",
  54096=>"100110100",
  54097=>"001110001",
  54098=>"001001100",
  54099=>"111011100",
  54100=>"000111011",
  54101=>"111000001",
  54102=>"001000100",
  54103=>"001111000",
  54104=>"100011000",
  54105=>"101000011",
  54106=>"100110101",
  54107=>"010011000",
  54108=>"001101110",
  54109=>"110001011",
  54110=>"100111111",
  54111=>"000000110",
  54112=>"101101000",
  54113=>"011101101",
  54114=>"000100001",
  54115=>"101111001",
  54116=>"110110000",
  54117=>"100010110",
  54118=>"001010100",
  54119=>"101100000",
  54120=>"011111011",
  54121=>"111111001",
  54122=>"111110001",
  54123=>"110110001",
  54124=>"110110111",
  54125=>"100111111",
  54126=>"111100110",
  54127=>"110011100",
  54128=>"100100101",
  54129=>"110000010",
  54130=>"110100110",
  54131=>"001101110",
  54132=>"110100010",
  54133=>"010111001",
  54134=>"110110000",
  54135=>"000011110",
  54136=>"110011110",
  54137=>"111001100",
  54138=>"101111001",
  54139=>"001110100",
  54140=>"001110100",
  54141=>"010101010",
  54142=>"111111111",
  54143=>"011011010",
  54144=>"000010001",
  54145=>"111010110",
  54146=>"000101010",
  54147=>"100101010",
  54148=>"011110101",
  54149=>"010001010",
  54150=>"100100110",
  54151=>"110101011",
  54152=>"111001111",
  54153=>"011100001",
  54154=>"010101111",
  54155=>"101011001",
  54156=>"011110111",
  54157=>"111111011",
  54158=>"101100001",
  54159=>"000001111",
  54160=>"100011111",
  54161=>"010000111",
  54162=>"110110110",
  54163=>"101001101",
  54164=>"001010110",
  54165=>"111111100",
  54166=>"110010101",
  54167=>"111110010",
  54168=>"110101010",
  54169=>"100010011",
  54170=>"110011000",
  54171=>"110101100",
  54172=>"100100010",
  54173=>"000010001",
  54174=>"110000100",
  54175=>"111010011",
  54176=>"110000000",
  54177=>"110010101",
  54178=>"001011010",
  54179=>"001110011",
  54180=>"000011101",
  54181=>"001101111",
  54182=>"100000100",
  54183=>"000001011",
  54184=>"001100000",
  54185=>"100110011",
  54186=>"111000011",
  54187=>"010101110",
  54188=>"100011010",
  54189=>"101011000",
  54190=>"001111001",
  54191=>"111110010",
  54192=>"000110101",
  54193=>"001100100",
  54194=>"000000000",
  54195=>"101010011",
  54196=>"011000001",
  54197=>"111000110",
  54198=>"010011111",
  54199=>"011111110",
  54200=>"110100010",
  54201=>"011111010",
  54202=>"110011110",
  54203=>"110110001",
  54204=>"111000010",
  54205=>"101011101",
  54206=>"011010101",
  54207=>"111100100",
  54208=>"110100110",
  54209=>"000000111",
  54210=>"101011000",
  54211=>"101110110",
  54212=>"000010100",
  54213=>"100010001",
  54214=>"110101100",
  54215=>"101000011",
  54216=>"100000110",
  54217=>"100110011",
  54218=>"111000111",
  54219=>"110111100",
  54220=>"101011111",
  54221=>"000010010",
  54222=>"011110000",
  54223=>"100100100",
  54224=>"000000101",
  54225=>"001011100",
  54226=>"000000100",
  54227=>"011000000",
  54228=>"001000000",
  54229=>"101110000",
  54230=>"001100100",
  54231=>"000000110",
  54232=>"011000101",
  54233=>"110110010",
  54234=>"001011111",
  54235=>"010011010",
  54236=>"001000011",
  54237=>"101111111",
  54238=>"011010000",
  54239=>"110011011",
  54240=>"000010111",
  54241=>"101011110",
  54242=>"011010110",
  54243=>"000110000",
  54244=>"100111000",
  54245=>"000110000",
  54246=>"110110110",
  54247=>"011001111",
  54248=>"100100010",
  54249=>"000110000",
  54250=>"000111000",
  54251=>"001010110",
  54252=>"011101000",
  54253=>"000110111",
  54254=>"001001011",
  54255=>"100010100",
  54256=>"000011100",
  54257=>"101111100",
  54258=>"010000100",
  54259=>"010110000",
  54260=>"110110110",
  54261=>"010101110",
  54262=>"011110100",
  54263=>"111111100",
  54264=>"011001011",
  54265=>"011111000",
  54266=>"101010110",
  54267=>"011110111",
  54268=>"100110010",
  54269=>"001110001",
  54270=>"111010100",
  54271=>"000111000",
  54272=>"101011011",
  54273=>"001101101",
  54274=>"001000001",
  54275=>"111110101",
  54276=>"001010110",
  54277=>"111100011",
  54278=>"011011111",
  54279=>"100111010",
  54280=>"110011111",
  54281=>"100010000",
  54282=>"110011100",
  54283=>"010100101",
  54284=>"001000111",
  54285=>"001100111",
  54286=>"000001100",
  54287=>"011000011",
  54288=>"000010101",
  54289=>"110011001",
  54290=>"100101110",
  54291=>"011110111",
  54292=>"111101011",
  54293=>"100111111",
  54294=>"111110100",
  54295=>"101000010",
  54296=>"100110111",
  54297=>"011001110",
  54298=>"011011101",
  54299=>"001101111",
  54300=>"011011011",
  54301=>"011111001",
  54302=>"111101011",
  54303=>"111010111",
  54304=>"001000100",
  54305=>"011000101",
  54306=>"010000001",
  54307=>"111001100",
  54308=>"011100101",
  54309=>"001101010",
  54310=>"101000001",
  54311=>"100011010",
  54312=>"000001001",
  54313=>"011001110",
  54314=>"101000001",
  54315=>"011000011",
  54316=>"111111111",
  54317=>"011100010",
  54318=>"100101010",
  54319=>"010011110",
  54320=>"101110000",
  54321=>"110100111",
  54322=>"110000111",
  54323=>"000001111",
  54324=>"001000101",
  54325=>"100000110",
  54326=>"100111111",
  54327=>"000111010",
  54328=>"000011001",
  54329=>"110011000",
  54330=>"110110000",
  54331=>"111110110",
  54332=>"000000110",
  54333=>"010110100",
  54334=>"001011000",
  54335=>"001011010",
  54336=>"011000011",
  54337=>"010100010",
  54338=>"111101000",
  54339=>"000011010",
  54340=>"001001011",
  54341=>"100110010",
  54342=>"001001110",
  54343=>"110110101",
  54344=>"000001111",
  54345=>"100000011",
  54346=>"100111011",
  54347=>"000111111",
  54348=>"011001100",
  54349=>"001010010",
  54350=>"011101001",
  54351=>"110010001",
  54352=>"011000001",
  54353=>"011011010",
  54354=>"110100010",
  54355=>"011000000",
  54356=>"000011000",
  54357=>"101101011",
  54358=>"101111001",
  54359=>"100110000",
  54360=>"111010001",
  54361=>"100001010",
  54362=>"110001010",
  54363=>"111010011",
  54364=>"010101111",
  54365=>"001000000",
  54366=>"111010001",
  54367=>"000010010",
  54368=>"110101110",
  54369=>"110010000",
  54370=>"010001101",
  54371=>"100001011",
  54372=>"001010110",
  54373=>"001010010",
  54374=>"100001101",
  54375=>"001010101",
  54376=>"011111110",
  54377=>"000111001",
  54378=>"110101111",
  54379=>"011010100",
  54380=>"110000011",
  54381=>"110110101",
  54382=>"010101001",
  54383=>"100011000",
  54384=>"001001110",
  54385=>"100011000",
  54386=>"000011001",
  54387=>"001000011",
  54388=>"110111011",
  54389=>"010000100",
  54390=>"111011001",
  54391=>"010100101",
  54392=>"010010100",
  54393=>"011000110",
  54394=>"010011110",
  54395=>"000100100",
  54396=>"000100010",
  54397=>"000111101",
  54398=>"001000111",
  54399=>"010110100",
  54400=>"010101100",
  54401=>"001101111",
  54402=>"001110000",
  54403=>"001000000",
  54404=>"111001000",
  54405=>"110101010",
  54406=>"111010111",
  54407=>"011001011",
  54408=>"110010010",
  54409=>"101001100",
  54410=>"011110111",
  54411=>"011000010",
  54412=>"011010010",
  54413=>"110000111",
  54414=>"100001110",
  54415=>"001111110",
  54416=>"110110110",
  54417=>"111100011",
  54418=>"110100111",
  54419=>"001010110",
  54420=>"110111100",
  54421=>"100011110",
  54422=>"000011101",
  54423=>"010000111",
  54424=>"000100110",
  54425=>"110001000",
  54426=>"110111100",
  54427=>"111000000",
  54428=>"000101101",
  54429=>"001111111",
  54430=>"111100101",
  54431=>"111010000",
  54432=>"100101110",
  54433=>"010001001",
  54434=>"010110111",
  54435=>"110010101",
  54436=>"001100111",
  54437=>"000000100",
  54438=>"110110110",
  54439=>"000100111",
  54440=>"111111001",
  54441=>"110011100",
  54442=>"000001101",
  54443=>"001010010",
  54444=>"101100100",
  54445=>"100001001",
  54446=>"001101110",
  54447=>"110110110",
  54448=>"101101001",
  54449=>"111110111",
  54450=>"000010011",
  54451=>"000001001",
  54452=>"100100011",
  54453=>"010011001",
  54454=>"101010100",
  54455=>"111111100",
  54456=>"100111010",
  54457=>"101101011",
  54458=>"110001110",
  54459=>"000101011",
  54460=>"101100010",
  54461=>"000111000",
  54462=>"110011111",
  54463=>"011001100",
  54464=>"111011011",
  54465=>"010011011",
  54466=>"100000100",
  54467=>"000101011",
  54468=>"101001000",
  54469=>"000001100",
  54470=>"111110101",
  54471=>"111000100",
  54472=>"000111010",
  54473=>"000001011",
  54474=>"001110011",
  54475=>"011111010",
  54476=>"011001001",
  54477=>"000110010",
  54478=>"011000010",
  54479=>"010010100",
  54480=>"011001111",
  54481=>"100011111",
  54482=>"001100100",
  54483=>"001010100",
  54484=>"110011110",
  54485=>"110111010",
  54486=>"111010111",
  54487=>"001010000",
  54488=>"111010100",
  54489=>"111000001",
  54490=>"001000010",
  54491=>"110110101",
  54492=>"100001111",
  54493=>"000001111",
  54494=>"000100000",
  54495=>"110110111",
  54496=>"010011111",
  54497=>"000010110",
  54498=>"100110001",
  54499=>"111000110",
  54500=>"000010100",
  54501=>"110110111",
  54502=>"110000100",
  54503=>"110101101",
  54504=>"000010011",
  54505=>"100001010",
  54506=>"100010001",
  54507=>"011111101",
  54508=>"000110101",
  54509=>"110100001",
  54510=>"111011001",
  54511=>"011100010",
  54512=>"000000101",
  54513=>"101101100",
  54514=>"101000000",
  54515=>"001110000",
  54516=>"110011011",
  54517=>"101010101",
  54518=>"101011110",
  54519=>"110000001",
  54520=>"010001101",
  54521=>"011111010",
  54522=>"110001110",
  54523=>"111000101",
  54524=>"001101111",
  54525=>"011001010",
  54526=>"101111000",
  54527=>"101111001",
  54528=>"011110111",
  54529=>"000101001",
  54530=>"010110101",
  54531=>"011011010",
  54532=>"011001111",
  54533=>"001101111",
  54534=>"010101111",
  54535=>"110010000",
  54536=>"011110110",
  54537=>"000011001",
  54538=>"110101101",
  54539=>"110011101",
  54540=>"010000001",
  54541=>"011010101",
  54542=>"110111111",
  54543=>"001101010",
  54544=>"001000011",
  54545=>"101011000",
  54546=>"111011010",
  54547=>"100100101",
  54548=>"000110001",
  54549=>"000001101",
  54550=>"101001000",
  54551=>"110011101",
  54552=>"001000010",
  54553=>"101101001",
  54554=>"111100010",
  54555=>"001000001",
  54556=>"011001111",
  54557=>"000011111",
  54558=>"011111010",
  54559=>"111100000",
  54560=>"000011010",
  54561=>"111111101",
  54562=>"111111101",
  54563=>"110010111",
  54564=>"001001011",
  54565=>"101010111",
  54566=>"011100110",
  54567=>"000000110",
  54568=>"110111101",
  54569=>"100010011",
  54570=>"010110100",
  54571=>"010010100",
  54572=>"000101111",
  54573=>"110001101",
  54574=>"111101110",
  54575=>"010001110",
  54576=>"101001011",
  54577=>"000100010",
  54578=>"000010111",
  54579=>"110001101",
  54580=>"110111111",
  54581=>"111100000",
  54582=>"111011101",
  54583=>"111100010",
  54584=>"101111101",
  54585=>"110101101",
  54586=>"001000001",
  54587=>"000101111",
  54588=>"000100111",
  54589=>"100111010",
  54590=>"111101000",
  54591=>"011110111",
  54592=>"010101110",
  54593=>"010100010",
  54594=>"001001010",
  54595=>"110111111",
  54596=>"001101000",
  54597=>"010110000",
  54598=>"110000010",
  54599=>"111101100",
  54600=>"101100110",
  54601=>"101011100",
  54602=>"011001011",
  54603=>"011101001",
  54604=>"101001111",
  54605=>"001100001",
  54606=>"011010111",
  54607=>"100110110",
  54608=>"000111100",
  54609=>"100001001",
  54610=>"111101101",
  54611=>"111111011",
  54612=>"000100100",
  54613=>"100111000",
  54614=>"001110010",
  54615=>"111110100",
  54616=>"000101001",
  54617=>"010110101",
  54618=>"000000100",
  54619=>"111101010",
  54620=>"100010101",
  54621=>"110101001",
  54622=>"001101011",
  54623=>"011000111",
  54624=>"101101101",
  54625=>"001011001",
  54626=>"101000101",
  54627=>"100111011",
  54628=>"100100100",
  54629=>"111100101",
  54630=>"110010010",
  54631=>"111110100",
  54632=>"011111011",
  54633=>"111000110",
  54634=>"000101001",
  54635=>"110000111",
  54636=>"100011101",
  54637=>"010100101",
  54638=>"111000001",
  54639=>"111100001",
  54640=>"011101000",
  54641=>"010001010",
  54642=>"001110110",
  54643=>"110100110",
  54644=>"010000001",
  54645=>"110101010",
  54646=>"111111011",
  54647=>"111111011",
  54648=>"000000110",
  54649=>"000101111",
  54650=>"010101010",
  54651=>"100111011",
  54652=>"111100010",
  54653=>"001101101",
  54654=>"000000110",
  54655=>"000111010",
  54656=>"111010001",
  54657=>"111010110",
  54658=>"000000001",
  54659=>"001011111",
  54660=>"001111100",
  54661=>"110010001",
  54662=>"101000101",
  54663=>"101000000",
  54664=>"111000110",
  54665=>"110001010",
  54666=>"000110001",
  54667=>"000100001",
  54668=>"110010101",
  54669=>"101101111",
  54670=>"101000100",
  54671=>"101000111",
  54672=>"011010101",
  54673=>"000000011",
  54674=>"101110001",
  54675=>"101001011",
  54676=>"101110111",
  54677=>"010010100",
  54678=>"011011000",
  54679=>"111101110",
  54680=>"110101101",
  54681=>"000001010",
  54682=>"111111011",
  54683=>"110010000",
  54684=>"000110001",
  54685=>"111011100",
  54686=>"000101011",
  54687=>"000100101",
  54688=>"000011110",
  54689=>"111010001",
  54690=>"010110111",
  54691=>"001101100",
  54692=>"001011101",
  54693=>"100001111",
  54694=>"110010111",
  54695=>"000111110",
  54696=>"100101010",
  54697=>"000111001",
  54698=>"110011111",
  54699=>"100100001",
  54700=>"111101101",
  54701=>"101010000",
  54702=>"101011111",
  54703=>"111110000",
  54704=>"111111111",
  54705=>"000100010",
  54706=>"001000011",
  54707=>"110100111",
  54708=>"010001011",
  54709=>"100100011",
  54710=>"010001100",
  54711=>"110010000",
  54712=>"000110010",
  54713=>"111001111",
  54714=>"000100100",
  54715=>"110011110",
  54716=>"100111110",
  54717=>"001010100",
  54718=>"001000110",
  54719=>"001001011",
  54720=>"110010001",
  54721=>"000001110",
  54722=>"011011101",
  54723=>"111101100",
  54724=>"001001011",
  54725=>"011011110",
  54726=>"111110110",
  54727=>"000101111",
  54728=>"110100001",
  54729=>"001111011",
  54730=>"111110001",
  54731=>"010110100",
  54732=>"011101011",
  54733=>"001111101",
  54734=>"001100011",
  54735=>"100010100",
  54736=>"100101000",
  54737=>"100100100",
  54738=>"111101000",
  54739=>"101001110",
  54740=>"100110011",
  54741=>"001110110",
  54742=>"001111000",
  54743=>"011000001",
  54744=>"100010100",
  54745=>"000100000",
  54746=>"000000001",
  54747=>"111001011",
  54748=>"101011010",
  54749=>"101000101",
  54750=>"001011100",
  54751=>"101000011",
  54752=>"001101010",
  54753=>"010111010",
  54754=>"011010011",
  54755=>"100101011",
  54756=>"000011101",
  54757=>"111011000",
  54758=>"100010101",
  54759=>"011101010",
  54760=>"100100001",
  54761=>"010001110",
  54762=>"011110001",
  54763=>"101100000",
  54764=>"010011001",
  54765=>"110100000",
  54766=>"111100001",
  54767=>"011101111",
  54768=>"101001111",
  54769=>"011011101",
  54770=>"000110100",
  54771=>"100011101",
  54772=>"010010001",
  54773=>"110111011",
  54774=>"011001100",
  54775=>"000100010",
  54776=>"101010010",
  54777=>"011011001",
  54778=>"100000101",
  54779=>"000101011",
  54780=>"000000000",
  54781=>"011011010",
  54782=>"000111000",
  54783=>"111001110",
  54784=>"011011010",
  54785=>"101100000",
  54786=>"111110110",
  54787=>"000111100",
  54788=>"000010010",
  54789=>"111110010",
  54790=>"010001000",
  54791=>"011010101",
  54792=>"101011010",
  54793=>"011011100",
  54794=>"100101011",
  54795=>"000000010",
  54796=>"111111110",
  54797=>"001001110",
  54798=>"111010000",
  54799=>"101001001",
  54800=>"110111100",
  54801=>"101110100",
  54802=>"010111100",
  54803=>"000011011",
  54804=>"010001001",
  54805=>"110100000",
  54806=>"010001001",
  54807=>"001100011",
  54808=>"111001111",
  54809=>"101100011",
  54810=>"100001110",
  54811=>"001001001",
  54812=>"101000000",
  54813=>"100110100",
  54814=>"101101101",
  54815=>"111001011",
  54816=>"000100100",
  54817=>"010100101",
  54818=>"000001100",
  54819=>"110110111",
  54820=>"101000011",
  54821=>"110100101",
  54822=>"101110001",
  54823=>"111011110",
  54824=>"000001010",
  54825=>"010111111",
  54826=>"111111001",
  54827=>"011110111",
  54828=>"110100001",
  54829=>"011111111",
  54830=>"101111101",
  54831=>"110000101",
  54832=>"001011110",
  54833=>"111100111",
  54834=>"001110101",
  54835=>"011100100",
  54836=>"010001010",
  54837=>"001100010",
  54838=>"110000010",
  54839=>"001000111",
  54840=>"101011011",
  54841=>"101110101",
  54842=>"000001100",
  54843=>"000101000",
  54844=>"001001101",
  54845=>"011110111",
  54846=>"001001101",
  54847=>"000110100",
  54848=>"100110000",
  54849=>"110011100",
  54850=>"101100000",
  54851=>"000100100",
  54852=>"010101100",
  54853=>"101001100",
  54854=>"001010110",
  54855=>"111111001",
  54856=>"000011011",
  54857=>"010110110",
  54858=>"111110001",
  54859=>"010110011",
  54860=>"101111111",
  54861=>"001100101",
  54862=>"111111111",
  54863=>"110101001",
  54864=>"010100010",
  54865=>"001110000",
  54866=>"101010000",
  54867=>"011101110",
  54868=>"100110010",
  54869=>"111011000",
  54870=>"001001011",
  54871=>"011000011",
  54872=>"000000000",
  54873=>"100011000",
  54874=>"010011110",
  54875=>"010000011",
  54876=>"111011111",
  54877=>"010010111",
  54878=>"010001101",
  54879=>"101000010",
  54880=>"111110101",
  54881=>"011011101",
  54882=>"001101011",
  54883=>"110000101",
  54884=>"101111110",
  54885=>"000001100",
  54886=>"001000101",
  54887=>"100110011",
  54888=>"110010011",
  54889=>"010001110",
  54890=>"001101110",
  54891=>"001000100",
  54892=>"000010101",
  54893=>"000000100",
  54894=>"001100110",
  54895=>"100011111",
  54896=>"001011110",
  54897=>"110100110",
  54898=>"111000011",
  54899=>"001110011",
  54900=>"101111011",
  54901=>"011000000",
  54902=>"110111101",
  54903=>"111111111",
  54904=>"010011000",
  54905=>"011101111",
  54906=>"011000111",
  54907=>"000101101",
  54908=>"100001000",
  54909=>"100011011",
  54910=>"100110000",
  54911=>"101101100",
  54912=>"000001100",
  54913=>"001100101",
  54914=>"101100111",
  54915=>"001100001",
  54916=>"001000001",
  54917=>"000001011",
  54918=>"001111011",
  54919=>"010010101",
  54920=>"000110011",
  54921=>"000001111",
  54922=>"100110111",
  54923=>"011010011",
  54924=>"101101010",
  54925=>"010100001",
  54926=>"011100100",
  54927=>"110111000",
  54928=>"011011010",
  54929=>"111111011",
  54930=>"010101000",
  54931=>"111100101",
  54932=>"010111001",
  54933=>"010100011",
  54934=>"111001101",
  54935=>"110101111",
  54936=>"100010110",
  54937=>"111001010",
  54938=>"100000010",
  54939=>"010101110",
  54940=>"110011010",
  54941=>"101010000",
  54942=>"101110011",
  54943=>"100000011",
  54944=>"011001011",
  54945=>"101011110",
  54946=>"111111000",
  54947=>"101000011",
  54948=>"000011000",
  54949=>"011111111",
  54950=>"011000100",
  54951=>"000110010",
  54952=>"101010000",
  54953=>"000100100",
  54954=>"010011110",
  54955=>"100010001",
  54956=>"000000010",
  54957=>"110110100",
  54958=>"010110100",
  54959=>"000000010",
  54960=>"100110010",
  54961=>"111011000",
  54962=>"111101110",
  54963=>"001000000",
  54964=>"011000100",
  54965=>"011100010",
  54966=>"001010101",
  54967=>"101100011",
  54968=>"110001001",
  54969=>"010001010",
  54970=>"100001010",
  54971=>"001000001",
  54972=>"101000111",
  54973=>"000011001",
  54974=>"111011000",
  54975=>"101001110",
  54976=>"110110110",
  54977=>"010001101",
  54978=>"111000111",
  54979=>"111110111",
  54980=>"000010110",
  54981=>"111000001",
  54982=>"001110001",
  54983=>"011001000",
  54984=>"000011000",
  54985=>"001011110",
  54986=>"111100100",
  54987=>"001111111",
  54988=>"111100101",
  54989=>"000000000",
  54990=>"111001100",
  54991=>"111011111",
  54992=>"100101000",
  54993=>"010100100",
  54994=>"000110101",
  54995=>"001000110",
  54996=>"010101100",
  54997=>"101011101",
  54998=>"110100010",
  54999=>"000010100",
  55000=>"001101101",
  55001=>"011001001",
  55002=>"111001011",
  55003=>"000111111",
  55004=>"111001001",
  55005=>"111110011",
  55006=>"111100101",
  55007=>"110011011",
  55008=>"110010101",
  55009=>"101001001",
  55010=>"001111010",
  55011=>"110000010",
  55012=>"101101100",
  55013=>"100010111",
  55014=>"010100011",
  55015=>"010000101",
  55016=>"100111010",
  55017=>"101100110",
  55018=>"011001010",
  55019=>"000000011",
  55020=>"011001011",
  55021=>"001100010",
  55022=>"001000000",
  55023=>"110110000",
  55024=>"001010101",
  55025=>"110010101",
  55026=>"101100110",
  55027=>"111011101",
  55028=>"111010100",
  55029=>"000101010",
  55030=>"011000000",
  55031=>"100100010",
  55032=>"000000011",
  55033=>"001111100",
  55034=>"101001011",
  55035=>"111111110",
  55036=>"111101110",
  55037=>"001011110",
  55038=>"101110000",
  55039=>"001000100",
  55040=>"100110010",
  55041=>"100111110",
  55042=>"011010001",
  55043=>"100010000",
  55044=>"100100101",
  55045=>"110011101",
  55046=>"100001100",
  55047=>"011101110",
  55048=>"100101001",
  55049=>"001100010",
  55050=>"001000000",
  55051=>"001000111",
  55052=>"101001010",
  55053=>"001101010",
  55054=>"100000011",
  55055=>"011111011",
  55056=>"111111111",
  55057=>"110100001",
  55058=>"101010100",
  55059=>"001011010",
  55060=>"110010000",
  55061=>"001010011",
  55062=>"110011001",
  55063=>"101001101",
  55064=>"100001101",
  55065=>"000010000",
  55066=>"000111011",
  55067=>"111001101",
  55068=>"000100110",
  55069=>"100010100",
  55070=>"110001111",
  55071=>"101010001",
  55072=>"100110001",
  55073=>"110101001",
  55074=>"000001010",
  55075=>"100111110",
  55076=>"010100011",
  55077=>"111000111",
  55078=>"011111011",
  55079=>"110010010",
  55080=>"110011000",
  55081=>"000000100",
  55082=>"101001001",
  55083=>"100010101",
  55084=>"000101010",
  55085=>"000101000",
  55086=>"110000110",
  55087=>"100111010",
  55088=>"111110000",
  55089=>"000001010",
  55090=>"011010111",
  55091=>"000101001",
  55092=>"111110111",
  55093=>"100000111",
  55094=>"010101001",
  55095=>"010100001",
  55096=>"111101000",
  55097=>"001100100",
  55098=>"001000100",
  55099=>"111110000",
  55100=>"000001101",
  55101=>"001010100",
  55102=>"101001100",
  55103=>"110110101",
  55104=>"100001110",
  55105=>"100001100",
  55106=>"001110110",
  55107=>"011001001",
  55108=>"000011101",
  55109=>"100111100",
  55110=>"010100001",
  55111=>"111110100",
  55112=>"110111110",
  55113=>"101101011",
  55114=>"011111101",
  55115=>"101111010",
  55116=>"101000100",
  55117=>"100000011",
  55118=>"100000110",
  55119=>"101110110",
  55120=>"101000011",
  55121=>"010001011",
  55122=>"111001101",
  55123=>"110000010",
  55124=>"110111000",
  55125=>"110111111",
  55126=>"100101010",
  55127=>"011111100",
  55128=>"111100000",
  55129=>"101111100",
  55130=>"111111101",
  55131=>"111001101",
  55132=>"000001011",
  55133=>"111000010",
  55134=>"000110001",
  55135=>"000000000",
  55136=>"100001001",
  55137=>"111110010",
  55138=>"100001110",
  55139=>"111011010",
  55140=>"101110010",
  55141=>"100110010",
  55142=>"000110001",
  55143=>"101001001",
  55144=>"111101101",
  55145=>"010000010",
  55146=>"110100010",
  55147=>"011100001",
  55148=>"100000110",
  55149=>"101100111",
  55150=>"001101010",
  55151=>"101010001",
  55152=>"101110010",
  55153=>"100100111",
  55154=>"000110111",
  55155=>"101011101",
  55156=>"110011111",
  55157=>"100001001",
  55158=>"110000000",
  55159=>"001101010",
  55160=>"101011111",
  55161=>"101100011",
  55162=>"000101000",
  55163=>"001010011",
  55164=>"111100101",
  55165=>"110110111",
  55166=>"111111100",
  55167=>"110110111",
  55168=>"100000110",
  55169=>"011101100",
  55170=>"101010110",
  55171=>"100111111",
  55172=>"010000101",
  55173=>"111000111",
  55174=>"001100010",
  55175=>"000010111",
  55176=>"111000001",
  55177=>"010011111",
  55178=>"111000101",
  55179=>"101111001",
  55180=>"110111011",
  55181=>"110111100",
  55182=>"101111101",
  55183=>"101010001",
  55184=>"101001011",
  55185=>"111110001",
  55186=>"011100011",
  55187=>"010011011",
  55188=>"100010101",
  55189=>"011111100",
  55190=>"001011000",
  55191=>"100001110",
  55192=>"000111011",
  55193=>"010000010",
  55194=>"111011010",
  55195=>"110011010",
  55196=>"000100011",
  55197=>"010010111",
  55198=>"101100000",
  55199=>"011000101",
  55200=>"000110101",
  55201=>"010110000",
  55202=>"011010101",
  55203=>"101000110",
  55204=>"110100110",
  55205=>"111101111",
  55206=>"101001000",
  55207=>"110010000",
  55208=>"111101100",
  55209=>"111110110",
  55210=>"000010101",
  55211=>"000100101",
  55212=>"001001011",
  55213=>"100100010",
  55214=>"111100101",
  55215=>"110000001",
  55216=>"000110001",
  55217=>"111000110",
  55218=>"011101010",
  55219=>"010101100",
  55220=>"100100001",
  55221=>"101001101",
  55222=>"000100100",
  55223=>"000101111",
  55224=>"111001010",
  55225=>"000100011",
  55226=>"101111000",
  55227=>"110011010",
  55228=>"010011111",
  55229=>"000001010",
  55230=>"000010000",
  55231=>"010101011",
  55232=>"110111001",
  55233=>"100000110",
  55234=>"001011011",
  55235=>"110111101",
  55236=>"001101110",
  55237=>"101000001",
  55238=>"010100011",
  55239=>"000011110",
  55240=>"111111100",
  55241=>"011000001",
  55242=>"101100111",
  55243=>"110100000",
  55244=>"001011011",
  55245=>"101011110",
  55246=>"111101110",
  55247=>"001010101",
  55248=>"100000100",
  55249=>"100011001",
  55250=>"101000100",
  55251=>"110101110",
  55252=>"111111111",
  55253=>"011000000",
  55254=>"101101111",
  55255=>"111100110",
  55256=>"001010001",
  55257=>"010100011",
  55258=>"010110000",
  55259=>"111010000",
  55260=>"011100110",
  55261=>"001100011",
  55262=>"010110110",
  55263=>"011000011",
  55264=>"010011011",
  55265=>"111000111",
  55266=>"000000010",
  55267=>"110011111",
  55268=>"001010011",
  55269=>"000000010",
  55270=>"110011010",
  55271=>"010000101",
  55272=>"111111000",
  55273=>"010000001",
  55274=>"110000100",
  55275=>"111110011",
  55276=>"010101100",
  55277=>"111101001",
  55278=>"010110100",
  55279=>"101100101",
  55280=>"100100011",
  55281=>"110110100",
  55282=>"001011010",
  55283=>"010000010",
  55284=>"100100110",
  55285=>"011011001",
  55286=>"111000111",
  55287=>"001010110",
  55288=>"001001111",
  55289=>"111110010",
  55290=>"101101110",
  55291=>"000111111",
  55292=>"010101000",
  55293=>"110000111",
  55294=>"010001100",
  55295=>"010011110",
  55296=>"101110100",
  55297=>"010110111",
  55298=>"000110110",
  55299=>"001100000",
  55300=>"100001100",
  55301=>"100011000",
  55302=>"000010011",
  55303=>"000100101",
  55304=>"100010001",
  55305=>"010110000",
  55306=>"010100010",
  55307=>"011001001",
  55308=>"111111100",
  55309=>"001111111",
  55310=>"000111001",
  55311=>"000101110",
  55312=>"011110011",
  55313=>"000001011",
  55314=>"001000000",
  55315=>"010001010",
  55316=>"010111101",
  55317=>"011110111",
  55318=>"101001101",
  55319=>"011111000",
  55320=>"000000000",
  55321=>"100010000",
  55322=>"101101100",
  55323=>"101011110",
  55324=>"101011011",
  55325=>"100010010",
  55326=>"001101101",
  55327=>"110110011",
  55328=>"001111111",
  55329=>"000111011",
  55330=>"000111010",
  55331=>"000000001",
  55332=>"101101011",
  55333=>"100101101",
  55334=>"100101111",
  55335=>"011010101",
  55336=>"101001111",
  55337=>"010000011",
  55338=>"110100101",
  55339=>"110010100",
  55340=>"110001001",
  55341=>"111111101",
  55342=>"010100011",
  55343=>"011100001",
  55344=>"011000011",
  55345=>"011010011",
  55346=>"011000101",
  55347=>"111011010",
  55348=>"101001000",
  55349=>"100111110",
  55350=>"111011001",
  55351=>"001011001",
  55352=>"111000101",
  55353=>"010111101",
  55354=>"111110011",
  55355=>"100011000",
  55356=>"110101111",
  55357=>"011100111",
  55358=>"101111111",
  55359=>"111101111",
  55360=>"001101110",
  55361=>"000000110",
  55362=>"110001000",
  55363=>"110100001",
  55364=>"010101101",
  55365=>"000010011",
  55366=>"101000011",
  55367=>"010101011",
  55368=>"110000001",
  55369=>"000100000",
  55370=>"000000010",
  55371=>"001110110",
  55372=>"101011111",
  55373=>"000010010",
  55374=>"110111110",
  55375=>"000100010",
  55376=>"011100100",
  55377=>"010101101",
  55378=>"000101100",
  55379=>"010111100",
  55380=>"001000001",
  55381=>"100101101",
  55382=>"100111000",
  55383=>"011101000",
  55384=>"001001110",
  55385=>"000000000",
  55386=>"000000011",
  55387=>"010100011",
  55388=>"101010011",
  55389=>"101100111",
  55390=>"111010011",
  55391=>"100101000",
  55392=>"111011000",
  55393=>"011101011",
  55394=>"101010111",
  55395=>"000011110",
  55396=>"101100101",
  55397=>"010100100",
  55398=>"000100100",
  55399=>"100000111",
  55400=>"011000001",
  55401=>"010100111",
  55402=>"010011011",
  55403=>"000100000",
  55404=>"101001001",
  55405=>"001100011",
  55406=>"100001100",
  55407=>"101111011",
  55408=>"000111000",
  55409=>"111001110",
  55410=>"100001111",
  55411=>"011111010",
  55412=>"111111011",
  55413=>"001111011",
  55414=>"111111110",
  55415=>"101001000",
  55416=>"101110011",
  55417=>"011011111",
  55418=>"010011000",
  55419=>"000001101",
  55420=>"111110101",
  55421=>"011111100",
  55422=>"111110001",
  55423=>"010001111",
  55424=>"000011001",
  55425=>"111000000",
  55426=>"110010101",
  55427=>"001111111",
  55428=>"011010011",
  55429=>"010101001",
  55430=>"000100011",
  55431=>"110100000",
  55432=>"101111000",
  55433=>"100111110",
  55434=>"101001101",
  55435=>"000001110",
  55436=>"011010001",
  55437=>"001001000",
  55438=>"001111111",
  55439=>"011101010",
  55440=>"111110000",
  55441=>"111010111",
  55442=>"111100101",
  55443=>"011110100",
  55444=>"111010110",
  55445=>"011111011",
  55446=>"100011011",
  55447=>"000101010",
  55448=>"111101100",
  55449=>"011000111",
  55450=>"101010001",
  55451=>"100011011",
  55452=>"101010001",
  55453=>"001001101",
  55454=>"011111011",
  55455=>"100011100",
  55456=>"000111101",
  55457=>"100100111",
  55458=>"111110110",
  55459=>"011000011",
  55460=>"010000100",
  55461=>"110000011",
  55462=>"001010110",
  55463=>"100110110",
  55464=>"000000110",
  55465=>"110111111",
  55466=>"001100001",
  55467=>"101101010",
  55468=>"001101000",
  55469=>"101010010",
  55470=>"001111010",
  55471=>"010011001",
  55472=>"000001111",
  55473=>"000001001",
  55474=>"010001111",
  55475=>"101101111",
  55476=>"111011101",
  55477=>"101001011",
  55478=>"010101110",
  55479=>"000001100",
  55480=>"100011000",
  55481=>"101010011",
  55482=>"101010010",
  55483=>"111011111",
  55484=>"011010001",
  55485=>"001100100",
  55486=>"110011111",
  55487=>"111000011",
  55488=>"010000110",
  55489=>"011000111",
  55490=>"010100010",
  55491=>"011110110",
  55492=>"110000111",
  55493=>"000111001",
  55494=>"010000101",
  55495=>"011110101",
  55496=>"110010011",
  55497=>"110101000",
  55498=>"000100111",
  55499=>"111001001",
  55500=>"110000000",
  55501=>"001101010",
  55502=>"000000010",
  55503=>"001111001",
  55504=>"011011011",
  55505=>"011000100",
  55506=>"110010010",
  55507=>"100101111",
  55508=>"000000000",
  55509=>"011110100",
  55510=>"101101010",
  55511=>"011110000",
  55512=>"111001110",
  55513=>"000001000",
  55514=>"011010000",
  55515=>"111100110",
  55516=>"011111101",
  55517=>"111111100",
  55518=>"111010101",
  55519=>"100100111",
  55520=>"010100101",
  55521=>"001000100",
  55522=>"010100001",
  55523=>"001011110",
  55524=>"001111101",
  55525=>"001000001",
  55526=>"100101000",
  55527=>"011010011",
  55528=>"110110111",
  55529=>"000110010",
  55530=>"101101011",
  55531=>"111010101",
  55532=>"000100100",
  55533=>"001101000",
  55534=>"111000100",
  55535=>"111101110",
  55536=>"010101001",
  55537=>"010011100",
  55538=>"010110000",
  55539=>"000000111",
  55540=>"001000101",
  55541=>"001111000",
  55542=>"011111000",
  55543=>"011101010",
  55544=>"000011010",
  55545=>"010000001",
  55546=>"100100000",
  55547=>"101101011",
  55548=>"110100011",
  55549=>"011001010",
  55550=>"010011111",
  55551=>"110101101",
  55552=>"011111000",
  55553=>"000011000",
  55554=>"110001010",
  55555=>"010111111",
  55556=>"101101101",
  55557=>"000111111",
  55558=>"101000100",
  55559=>"000110110",
  55560=>"001000000",
  55561=>"010000110",
  55562=>"010111111",
  55563=>"100111100",
  55564=>"100110010",
  55565=>"000011011",
  55566=>"001111001",
  55567=>"001010111",
  55568=>"010111101",
  55569=>"110101110",
  55570=>"001010100",
  55571=>"001101111",
  55572=>"010011001",
  55573=>"011101101",
  55574=>"111110110",
  55575=>"000011011",
  55576=>"100101110",
  55577=>"100010000",
  55578=>"010100101",
  55579=>"101011110",
  55580=>"111101101",
  55581=>"101011000",
  55582=>"111111011",
  55583=>"100001111",
  55584=>"101000101",
  55585=>"001111001",
  55586=>"000000101",
  55587=>"110111111",
  55588=>"111100001",
  55589=>"111011101",
  55590=>"001001010",
  55591=>"101100110",
  55592=>"110000011",
  55593=>"011010010",
  55594=>"101000110",
  55595=>"101110001",
  55596=>"010011011",
  55597=>"010110100",
  55598=>"111100100",
  55599=>"010101001",
  55600=>"010110111",
  55601=>"101010011",
  55602=>"001000000",
  55603=>"111010101",
  55604=>"100100000",
  55605=>"101110011",
  55606=>"001100100",
  55607=>"110010101",
  55608=>"011101111",
  55609=>"011100101",
  55610=>"010011101",
  55611=>"000101111",
  55612=>"001000001",
  55613=>"111101100",
  55614=>"101111100",
  55615=>"001001111",
  55616=>"101001011",
  55617=>"111010100",
  55618=>"011001001",
  55619=>"011011001",
  55620=>"101001000",
  55621=>"001101111",
  55622=>"011001010",
  55623=>"111111000",
  55624=>"101011110",
  55625=>"111001010",
  55626=>"011101010",
  55627=>"010011001",
  55628=>"101010010",
  55629=>"001000101",
  55630=>"000010100",
  55631=>"000000101",
  55632=>"001100101",
  55633=>"001110001",
  55634=>"100011011",
  55635=>"101100110",
  55636=>"101000001",
  55637=>"110110110",
  55638=>"001101111",
  55639=>"000101110",
  55640=>"100110001",
  55641=>"111111111",
  55642=>"010111010",
  55643=>"000000101",
  55644=>"101111011",
  55645=>"011000100",
  55646=>"111111101",
  55647=>"011110111",
  55648=>"101001101",
  55649=>"100111011",
  55650=>"000011001",
  55651=>"000101111",
  55652=>"100000000",
  55653=>"011101100",
  55654=>"110101000",
  55655=>"111110010",
  55656=>"111111011",
  55657=>"000100000",
  55658=>"000100001",
  55659=>"000101110",
  55660=>"000111000",
  55661=>"010101110",
  55662=>"100110111",
  55663=>"000111011",
  55664=>"011010000",
  55665=>"001001000",
  55666=>"101000101",
  55667=>"110010111",
  55668=>"010110000",
  55669=>"111111101",
  55670=>"100111010",
  55671=>"011010010",
  55672=>"010010000",
  55673=>"000101110",
  55674=>"010010110",
  55675=>"101001000",
  55676=>"101110000",
  55677=>"111011011",
  55678=>"001001000",
  55679=>"111001000",
  55680=>"000010011",
  55681=>"100110011",
  55682=>"000101000",
  55683=>"100010101",
  55684=>"101001100",
  55685=>"000010011",
  55686=>"111101011",
  55687=>"001011010",
  55688=>"100001011",
  55689=>"011110111",
  55690=>"010010100",
  55691=>"101001000",
  55692=>"010110001",
  55693=>"110100110",
  55694=>"100100100",
  55695=>"011111001",
  55696=>"110000110",
  55697=>"011000001",
  55698=>"111001000",
  55699=>"010000010",
  55700=>"110011110",
  55701=>"000100000",
  55702=>"001000100",
  55703=>"011000001",
  55704=>"001001100",
  55705=>"011111000",
  55706=>"110010010",
  55707=>"101000011",
  55708=>"011010101",
  55709=>"101100111",
  55710=>"010001011",
  55711=>"001100111",
  55712=>"000111001",
  55713=>"000100001",
  55714=>"100110111",
  55715=>"110100100",
  55716=>"001010111",
  55717=>"111010001",
  55718=>"011110111",
  55719=>"001000110",
  55720=>"001100001",
  55721=>"110010001",
  55722=>"000000011",
  55723=>"011011111",
  55724=>"000010000",
  55725=>"111100001",
  55726=>"110010111",
  55727=>"110011000",
  55728=>"111110101",
  55729=>"100001110",
  55730=>"110100010",
  55731=>"100011111",
  55732=>"101010100",
  55733=>"010101111",
  55734=>"100111010",
  55735=>"000100010",
  55736=>"100001000",
  55737=>"000100001",
  55738=>"101010000",
  55739=>"110111010",
  55740=>"101001001",
  55741=>"101110000",
  55742=>"100000011",
  55743=>"011111000",
  55744=>"000001011",
  55745=>"011100010",
  55746=>"100010101",
  55747=>"010101000",
  55748=>"000110101",
  55749=>"110001000",
  55750=>"010000000",
  55751=>"111011000",
  55752=>"011110010",
  55753=>"100100011",
  55754=>"001100000",
  55755=>"011111110",
  55756=>"101011111",
  55757=>"110100000",
  55758=>"011000010",
  55759=>"100000010",
  55760=>"001101111",
  55761=>"001111001",
  55762=>"101000001",
  55763=>"010111000",
  55764=>"100111110",
  55765=>"000100001",
  55766=>"111111110",
  55767=>"100000011",
  55768=>"111010000",
  55769=>"110001011",
  55770=>"100101001",
  55771=>"111010111",
  55772=>"100001000",
  55773=>"011010010",
  55774=>"111100110",
  55775=>"100100100",
  55776=>"010100000",
  55777=>"111101111",
  55778=>"101000000",
  55779=>"001011001",
  55780=>"110100011",
  55781=>"001001100",
  55782=>"101001011",
  55783=>"101111111",
  55784=>"000001101",
  55785=>"101110001",
  55786=>"000100000",
  55787=>"101111010",
  55788=>"111101111",
  55789=>"101000111",
  55790=>"101000111",
  55791=>"111010111",
  55792=>"010110010",
  55793=>"100000000",
  55794=>"101001000",
  55795=>"011111100",
  55796=>"010010100",
  55797=>"111101101",
  55798=>"010110101",
  55799=>"101010000",
  55800=>"000101000",
  55801=>"000000001",
  55802=>"100011101",
  55803=>"110101000",
  55804=>"000010101",
  55805=>"100011000",
  55806=>"001010000",
  55807=>"101001001",
  55808=>"111110011",
  55809=>"100010111",
  55810=>"011011110",
  55811=>"100000001",
  55812=>"001000000",
  55813=>"101001110",
  55814=>"111111000",
  55815=>"000011001",
  55816=>"001100000",
  55817=>"000100010",
  55818=>"001010101",
  55819=>"001110100",
  55820=>"111000010",
  55821=>"000110010",
  55822=>"010010100",
  55823=>"001000000",
  55824=>"110110000",
  55825=>"111111011",
  55826=>"010111001",
  55827=>"100010010",
  55828=>"110101101",
  55829=>"001010000",
  55830=>"111101100",
  55831=>"101101000",
  55832=>"000000110",
  55833=>"101110010",
  55834=>"100011010",
  55835=>"100000001",
  55836=>"111011100",
  55837=>"111111011",
  55838=>"010000111",
  55839=>"011011101",
  55840=>"011011011",
  55841=>"110110101",
  55842=>"000111111",
  55843=>"101011000",
  55844=>"111111001",
  55845=>"001100100",
  55846=>"100111001",
  55847=>"100011001",
  55848=>"101000100",
  55849=>"111111101",
  55850=>"011011010",
  55851=>"110111011",
  55852=>"011101111",
  55853=>"011100001",
  55854=>"000000110",
  55855=>"000010000",
  55856=>"110001111",
  55857=>"100000111",
  55858=>"111111101",
  55859=>"101001001",
  55860=>"100101111",
  55861=>"111010100",
  55862=>"110011000",
  55863=>"101101001",
  55864=>"100111110",
  55865=>"110000010",
  55866=>"010011100",
  55867=>"100110111",
  55868=>"000010010",
  55869=>"110011100",
  55870=>"000011001",
  55871=>"100111010",
  55872=>"000101101",
  55873=>"111110111",
  55874=>"000000111",
  55875=>"011100010",
  55876=>"110100001",
  55877=>"110001000",
  55878=>"111111001",
  55879=>"111011100",
  55880=>"110100010",
  55881=>"001010100",
  55882=>"111000010",
  55883=>"100110000",
  55884=>"000110011",
  55885=>"110100100",
  55886=>"000000000",
  55887=>"101111111",
  55888=>"101101011",
  55889=>"011111111",
  55890=>"101110001",
  55891=>"110111111",
  55892=>"011110110",
  55893=>"000011000",
  55894=>"010000000",
  55895=>"100111101",
  55896=>"000000000",
  55897=>"111010011",
  55898=>"100001000",
  55899=>"010110011",
  55900=>"011111111",
  55901=>"101101001",
  55902=>"101101000",
  55903=>"111111010",
  55904=>"001001100",
  55905=>"100001010",
  55906=>"001000000",
  55907=>"110100100",
  55908=>"100111011",
  55909=>"111111110",
  55910=>"110010000",
  55911=>"000100001",
  55912=>"101000011",
  55913=>"101001010",
  55914=>"011101100",
  55915=>"001000011",
  55916=>"000101011",
  55917=>"001010101",
  55918=>"101000100",
  55919=>"101010110",
  55920=>"101101011",
  55921=>"001011101",
  55922=>"010011000",
  55923=>"111110100",
  55924=>"111010010",
  55925=>"110111100",
  55926=>"000101100",
  55927=>"110010101",
  55928=>"001011111",
  55929=>"001101110",
  55930=>"010110011",
  55931=>"010010001",
  55932=>"111011110",
  55933=>"111101010",
  55934=>"000011101",
  55935=>"001100000",
  55936=>"001000000",
  55937=>"101011001",
  55938=>"011111110",
  55939=>"100001100",
  55940=>"000010010",
  55941=>"010010110",
  55942=>"100100001",
  55943=>"011000011",
  55944=>"001111001",
  55945=>"010001100",
  55946=>"001000011",
  55947=>"011000100",
  55948=>"110011100",
  55949=>"110010101",
  55950=>"111001100",
  55951=>"100111100",
  55952=>"111110110",
  55953=>"010000101",
  55954=>"000000100",
  55955=>"111010101",
  55956=>"001011100",
  55957=>"001101010",
  55958=>"010110011",
  55959=>"110110000",
  55960=>"010100011",
  55961=>"001001000",
  55962=>"110011101",
  55963=>"011011001",
  55964=>"111100000",
  55965=>"110010000",
  55966=>"001110010",
  55967=>"011101011",
  55968=>"101101001",
  55969=>"001100001",
  55970=>"111110111",
  55971=>"001001011",
  55972=>"011100001",
  55973=>"100100100",
  55974=>"011110000",
  55975=>"110100111",
  55976=>"100101010",
  55977=>"111110000",
  55978=>"011110000",
  55979=>"010111111",
  55980=>"011101000",
  55981=>"111011110",
  55982=>"001111100",
  55983=>"100110101",
  55984=>"011000000",
  55985=>"101000011",
  55986=>"110110101",
  55987=>"110011001",
  55988=>"010010011",
  55989=>"101000111",
  55990=>"100101111",
  55991=>"111001110",
  55992=>"001110000",
  55993=>"001000000",
  55994=>"100010000",
  55995=>"000101011",
  55996=>"111100111",
  55997=>"100011011",
  55998=>"011101001",
  55999=>"110000101",
  56000=>"111111100",
  56001=>"001111110",
  56002=>"000000101",
  56003=>"000100010",
  56004=>"010101001",
  56005=>"000001001",
  56006=>"000000000",
  56007=>"100100111",
  56008=>"001010000",
  56009=>"011111110",
  56010=>"101010100",
  56011=>"001010011",
  56012=>"001101010",
  56013=>"000100010",
  56014=>"111111111",
  56015=>"010001011",
  56016=>"000101100",
  56017=>"000101001",
  56018=>"010100000",
  56019=>"101011110",
  56020=>"110100100",
  56021=>"110010111",
  56022=>"011000010",
  56023=>"011001111",
  56024=>"110000110",
  56025=>"001111101",
  56026=>"000011001",
  56027=>"011110001",
  56028=>"010110101",
  56029=>"011000110",
  56030=>"100000001",
  56031=>"111011000",
  56032=>"111011000",
  56033=>"001010101",
  56034=>"100101010",
  56035=>"001110110",
  56036=>"111101110",
  56037=>"101011000",
  56038=>"011001010",
  56039=>"000110010",
  56040=>"110000100",
  56041=>"111111000",
  56042=>"101111100",
  56043=>"111011011",
  56044=>"111011000",
  56045=>"000001010",
  56046=>"011110101",
  56047=>"101101010",
  56048=>"110011101",
  56049=>"001011110",
  56050=>"010000010",
  56051=>"100000001",
  56052=>"000100111",
  56053=>"010111000",
  56054=>"001100101",
  56055=>"110100100",
  56056=>"110111110",
  56057=>"111111100",
  56058=>"110010100",
  56059=>"110010001",
  56060=>"100000111",
  56061=>"101101010",
  56062=>"101011000",
  56063=>"000000111",
  56064=>"100100100",
  56065=>"000000100",
  56066=>"000001011",
  56067=>"000001111",
  56068=>"100011010",
  56069=>"110101101",
  56070=>"101010101",
  56071=>"111111111",
  56072=>"100111011",
  56073=>"101110001",
  56074=>"011011101",
  56075=>"101011111",
  56076=>"110011000",
  56077=>"011001001",
  56078=>"100001101",
  56079=>"100010000",
  56080=>"101010111",
  56081=>"111010010",
  56082=>"010101000",
  56083=>"010001110",
  56084=>"010100101",
  56085=>"111111111",
  56086=>"011000111",
  56087=>"110101010",
  56088=>"011010000",
  56089=>"001101000",
  56090=>"001011111",
  56091=>"111100001",
  56092=>"000100010",
  56093=>"010000010",
  56094=>"101010100",
  56095=>"111110110",
  56096=>"001101111",
  56097=>"100101110",
  56098=>"100011101",
  56099=>"000000101",
  56100=>"110010110",
  56101=>"101101001",
  56102=>"000111010",
  56103=>"100000101",
  56104=>"001011010",
  56105=>"111111110",
  56106=>"001110001",
  56107=>"000001110",
  56108=>"111111001",
  56109=>"000000000",
  56110=>"111001000",
  56111=>"101000000",
  56112=>"100000110",
  56113=>"011110010",
  56114=>"111000110",
  56115=>"011011100",
  56116=>"000010101",
  56117=>"101000100",
  56118=>"000001111",
  56119=>"110011010",
  56120=>"010011111",
  56121=>"110010001",
  56122=>"001010001",
  56123=>"101100110",
  56124=>"001001001",
  56125=>"110001001",
  56126=>"011000101",
  56127=>"000011001",
  56128=>"100000110",
  56129=>"111000001",
  56130=>"010100000",
  56131=>"110100101",
  56132=>"100011101",
  56133=>"000110110",
  56134=>"010001110",
  56135=>"010011111",
  56136=>"001010011",
  56137=>"010111000",
  56138=>"111100000",
  56139=>"011100010",
  56140=>"100101101",
  56141=>"000110010",
  56142=>"101100101",
  56143=>"010100111",
  56144=>"011011011",
  56145=>"010001000",
  56146=>"100111000",
  56147=>"111000000",
  56148=>"101100010",
  56149=>"001101100",
  56150=>"101000111",
  56151=>"011110001",
  56152=>"110110001",
  56153=>"011111000",
  56154=>"100011001",
  56155=>"001100000",
  56156=>"101110101",
  56157=>"110111010",
  56158=>"010001001",
  56159=>"101100110",
  56160=>"001110111",
  56161=>"010010111",
  56162=>"010001010",
  56163=>"101100011",
  56164=>"011110000",
  56165=>"011100001",
  56166=>"010010111",
  56167=>"110110111",
  56168=>"110001011",
  56169=>"110111110",
  56170=>"111000001",
  56171=>"111010110",
  56172=>"100101111",
  56173=>"000001010",
  56174=>"001011110",
  56175=>"000100111",
  56176=>"010111000",
  56177=>"001110010",
  56178=>"111011011",
  56179=>"101010010",
  56180=>"111000101",
  56181=>"111110010",
  56182=>"001010111",
  56183=>"100000100",
  56184=>"110011011",
  56185=>"100101101",
  56186=>"100111001",
  56187=>"101001000",
  56188=>"001001100",
  56189=>"010110000",
  56190=>"111010001",
  56191=>"101111110",
  56192=>"110111011",
  56193=>"101011111",
  56194=>"111001000",
  56195=>"110001001",
  56196=>"101011001",
  56197=>"110011110",
  56198=>"100110011",
  56199=>"001110000",
  56200=>"000100101",
  56201=>"101101111",
  56202=>"110111011",
  56203=>"001101111",
  56204=>"110100010",
  56205=>"110111001",
  56206=>"110000010",
  56207=>"100001101",
  56208=>"001100111",
  56209=>"100001011",
  56210=>"111110101",
  56211=>"101100011",
  56212=>"101111001",
  56213=>"100110010",
  56214=>"011101110",
  56215=>"101000100",
  56216=>"100111011",
  56217=>"010101000",
  56218=>"010011111",
  56219=>"000010110",
  56220=>"011111101",
  56221=>"110011001",
  56222=>"110100100",
  56223=>"010011000",
  56224=>"100100111",
  56225=>"101101101",
  56226=>"010100100",
  56227=>"111100000",
  56228=>"011010000",
  56229=>"001011101",
  56230=>"110101011",
  56231=>"010101001",
  56232=>"010010100",
  56233=>"000000011",
  56234=>"110100111",
  56235=>"100111111",
  56236=>"011000101",
  56237=>"010110011",
  56238=>"100000101",
  56239=>"010000010",
  56240=>"011010010",
  56241=>"011110101",
  56242=>"011101110",
  56243=>"111101001",
  56244=>"110000110",
  56245=>"110110011",
  56246=>"101011010",
  56247=>"101010100",
  56248=>"011010000",
  56249=>"011101100",
  56250=>"010111011",
  56251=>"011010001",
  56252=>"010101001",
  56253=>"000111000",
  56254=>"111010101",
  56255=>"100101011",
  56256=>"001101111",
  56257=>"110011111",
  56258=>"000101100",
  56259=>"101100000",
  56260=>"011111010",
  56261=>"100000101",
  56262=>"101111110",
  56263=>"100100110",
  56264=>"100000010",
  56265=>"010100101",
  56266=>"111111000",
  56267=>"111110011",
  56268=>"101000001",
  56269=>"111001000",
  56270=>"100010001",
  56271=>"111011110",
  56272=>"000010000",
  56273=>"101001110",
  56274=>"110001010",
  56275=>"010101101",
  56276=>"001100001",
  56277=>"110000010",
  56278=>"000100100",
  56279=>"010111110",
  56280=>"110110111",
  56281=>"101001111",
  56282=>"110000101",
  56283=>"110110000",
  56284=>"111000010",
  56285=>"111110110",
  56286=>"001111000",
  56287=>"111000010",
  56288=>"110111000",
  56289=>"101011100",
  56290=>"011111001",
  56291=>"011101001",
  56292=>"110001101",
  56293=>"100011011",
  56294=>"101100011",
  56295=>"011110011",
  56296=>"011101110",
  56297=>"011101101",
  56298=>"110010010",
  56299=>"111011011",
  56300=>"100010010",
  56301=>"111100110",
  56302=>"011011001",
  56303=>"100101000",
  56304=>"000101101",
  56305=>"100101111",
  56306=>"000001101",
  56307=>"000100101",
  56308=>"011110100",
  56309=>"111010001",
  56310=>"101111100",
  56311=>"011110000",
  56312=>"101111100",
  56313=>"111000011",
  56314=>"110010101",
  56315=>"111110100",
  56316=>"010111100",
  56317=>"100111000",
  56318=>"011010100",
  56319=>"010010011",
  56320=>"111101101",
  56321=>"001111010",
  56322=>"100100010",
  56323=>"001001100",
  56324=>"010000011",
  56325=>"101010001",
  56326=>"110100101",
  56327=>"011101111",
  56328=>"111011111",
  56329=>"001001111",
  56330=>"100100100",
  56331=>"100001001",
  56332=>"111000111",
  56333=>"110111110",
  56334=>"101011001",
  56335=>"011101111",
  56336=>"000000111",
  56337=>"000001111",
  56338=>"011111111",
  56339=>"011011000",
  56340=>"001110001",
  56341=>"100010010",
  56342=>"110100001",
  56343=>"011000000",
  56344=>"111101010",
  56345=>"110011111",
  56346=>"100110001",
  56347=>"000100111",
  56348=>"000100101",
  56349=>"110101110",
  56350=>"010101011",
  56351=>"111011100",
  56352=>"000011100",
  56353=>"001101101",
  56354=>"111000011",
  56355=>"110100010",
  56356=>"000111000",
  56357=>"000010000",
  56358=>"001000000",
  56359=>"011010101",
  56360=>"100011101",
  56361=>"001110000",
  56362=>"111101110",
  56363=>"111110011",
  56364=>"111010000",
  56365=>"110010000",
  56366=>"100001010",
  56367=>"000000110",
  56368=>"001001011",
  56369=>"000100100",
  56370=>"110001011",
  56371=>"101111110",
  56372=>"111000010",
  56373=>"010101011",
  56374=>"110001100",
  56375=>"110000000",
  56376=>"000010001",
  56377=>"000000111",
  56378=>"001101100",
  56379=>"101000010",
  56380=>"101010000",
  56381=>"001010000",
  56382=>"101001010",
  56383=>"000010110",
  56384=>"011011100",
  56385=>"001000101",
  56386=>"000100110",
  56387=>"011111000",
  56388=>"001100001",
  56389=>"100011010",
  56390=>"101111101",
  56391=>"110010001",
  56392=>"110100110",
  56393=>"001101100",
  56394=>"001110000",
  56395=>"111010001",
  56396=>"101010001",
  56397=>"011101011",
  56398=>"101111110",
  56399=>"011110110",
  56400=>"000110100",
  56401=>"000000010",
  56402=>"110010100",
  56403=>"000010111",
  56404=>"101010101",
  56405=>"000000000",
  56406=>"001000001",
  56407=>"100010100",
  56408=>"110101111",
  56409=>"110010100",
  56410=>"010000111",
  56411=>"100101001",
  56412=>"000001001",
  56413=>"000000000",
  56414=>"010111110",
  56415=>"111001001",
  56416=>"010000100",
  56417=>"101101101",
  56418=>"000000101",
  56419=>"100110110",
  56420=>"110011001",
  56421=>"010100011",
  56422=>"001001100",
  56423=>"000101100",
  56424=>"100110101",
  56425=>"100100011",
  56426=>"011011100",
  56427=>"000110001",
  56428=>"010011100",
  56429=>"101011001",
  56430=>"001011111",
  56431=>"100111111",
  56432=>"010001010",
  56433=>"110011001",
  56434=>"010101110",
  56435=>"111111111",
  56436=>"001011101",
  56437=>"001000111",
  56438=>"111000011",
  56439=>"011111011",
  56440=>"001111100",
  56441=>"001001100",
  56442=>"111011100",
  56443=>"001010110",
  56444=>"101101101",
  56445=>"000000010",
  56446=>"111110111",
  56447=>"111100001",
  56448=>"000001010",
  56449=>"100000100",
  56450=>"110010010",
  56451=>"001000011",
  56452=>"100000001",
  56453=>"100011001",
  56454=>"110101101",
  56455=>"100000111",
  56456=>"100110110",
  56457=>"100110010",
  56458=>"110100011",
  56459=>"011101111",
  56460=>"011011101",
  56461=>"110110011",
  56462=>"111100011",
  56463=>"011101000",
  56464=>"001111000",
  56465=>"100001111",
  56466=>"001101001",
  56467=>"000110001",
  56468=>"111001011",
  56469=>"001000101",
  56470=>"011011110",
  56471=>"101110001",
  56472=>"001011110",
  56473=>"101000011",
  56474=>"000110000",
  56475=>"110101000",
  56476=>"010010111",
  56477=>"000010001",
  56478=>"000101111",
  56479=>"011111101",
  56480=>"001100101",
  56481=>"111110110",
  56482=>"000001001",
  56483=>"010111101",
  56484=>"010011110",
  56485=>"001010000",
  56486=>"000001001",
  56487=>"000000001",
  56488=>"001001011",
  56489=>"011000101",
  56490=>"010100001",
  56491=>"000111000",
  56492=>"001111011",
  56493=>"100000000",
  56494=>"101010100",
  56495=>"111101010",
  56496=>"100010101",
  56497=>"000111000",
  56498=>"001111011",
  56499=>"010111101",
  56500=>"000000110",
  56501=>"000101010",
  56502=>"110010101",
  56503=>"100100111",
  56504=>"011001001",
  56505=>"111000000",
  56506=>"000110001",
  56507=>"010010000",
  56508=>"100101111",
  56509=>"000010010",
  56510=>"110000110",
  56511=>"010111001",
  56512=>"100001101",
  56513=>"010000110",
  56514=>"111111000",
  56515=>"011001010",
  56516=>"111101111",
  56517=>"010101000",
  56518=>"110011100",
  56519=>"100010110",
  56520=>"010011110",
  56521=>"101100100",
  56522=>"100101000",
  56523=>"000111110",
  56524=>"111101110",
  56525=>"010101101",
  56526=>"000110111",
  56527=>"001000110",
  56528=>"110110101",
  56529=>"111000010",
  56530=>"110101000",
  56531=>"101111111",
  56532=>"100111000",
  56533=>"110001000",
  56534=>"111000110",
  56535=>"101101111",
  56536=>"100101000",
  56537=>"100101110",
  56538=>"010100000",
  56539=>"010011111",
  56540=>"010011110",
  56541=>"101101010",
  56542=>"000110111",
  56543=>"001000011",
  56544=>"001010010",
  56545=>"011100011",
  56546=>"010011101",
  56547=>"111111011",
  56548=>"000010001",
  56549=>"010100000",
  56550=>"001100001",
  56551=>"011111001",
  56552=>"000000000",
  56553=>"111110010",
  56554=>"100111101",
  56555=>"111011000",
  56556=>"110110111",
  56557=>"000111100",
  56558=>"110001111",
  56559=>"011100010",
  56560=>"110010111",
  56561=>"010000100",
  56562=>"000110111",
  56563=>"010101111",
  56564=>"000010000",
  56565=>"111100110",
  56566=>"011101000",
  56567=>"000011110",
  56568=>"110010100",
  56569=>"010011010",
  56570=>"000001101",
  56571=>"000110001",
  56572=>"001001001",
  56573=>"110110010",
  56574=>"110100101",
  56575=>"000010011",
  56576=>"100111011",
  56577=>"110100110",
  56578=>"011000100",
  56579=>"000101101",
  56580=>"100111110",
  56581=>"000000010",
  56582=>"011000011",
  56583=>"010001011",
  56584=>"110111100",
  56585=>"001111111",
  56586=>"111000001",
  56587=>"011000011",
  56588=>"101010000",
  56589=>"111101001",
  56590=>"101101011",
  56591=>"000101101",
  56592=>"001011001",
  56593=>"110000101",
  56594=>"001101000",
  56595=>"001101100",
  56596=>"010010001",
  56597=>"111110000",
  56598=>"001011011",
  56599=>"000111010",
  56600=>"000100101",
  56601=>"100011110",
  56602=>"100110111",
  56603=>"111010110",
  56604=>"111101000",
  56605=>"010001100",
  56606=>"100111111",
  56607=>"100000111",
  56608=>"000101000",
  56609=>"010110110",
  56610=>"100011010",
  56611=>"100011110",
  56612=>"110110001",
  56613=>"000100110",
  56614=>"100011000",
  56615=>"011001101",
  56616=>"100110100",
  56617=>"010100100",
  56618=>"010110100",
  56619=>"011011000",
  56620=>"010101000",
  56621=>"111111101",
  56622=>"010000000",
  56623=>"001011001",
  56624=>"010001111",
  56625=>"001001100",
  56626=>"010011010",
  56627=>"100101001",
  56628=>"001000010",
  56629=>"011000010",
  56630=>"001110100",
  56631=>"101011000",
  56632=>"010011010",
  56633=>"100101110",
  56634=>"111010000",
  56635=>"001110101",
  56636=>"101110011",
  56637=>"101000110",
  56638=>"000001011",
  56639=>"110100010",
  56640=>"111010000",
  56641=>"100000100",
  56642=>"000000010",
  56643=>"100110101",
  56644=>"000110110",
  56645=>"011111010",
  56646=>"001011111",
  56647=>"111010101",
  56648=>"000110001",
  56649=>"000011001",
  56650=>"010100111",
  56651=>"000111010",
  56652=>"011000110",
  56653=>"110100000",
  56654=>"010000010",
  56655=>"000100010",
  56656=>"111110000",
  56657=>"011101101",
  56658=>"000000001",
  56659=>"111110000",
  56660=>"111110000",
  56661=>"101001100",
  56662=>"010000011",
  56663=>"000001110",
  56664=>"001111001",
  56665=>"000101100",
  56666=>"110111010",
  56667=>"011100010",
  56668=>"100001001",
  56669=>"010100101",
  56670=>"001101101",
  56671=>"100110001",
  56672=>"111011110",
  56673=>"110000011",
  56674=>"111110101",
  56675=>"000001011",
  56676=>"100100010",
  56677=>"010001001",
  56678=>"001010010",
  56679=>"011010000",
  56680=>"111101000",
  56681=>"111111000",
  56682=>"010010011",
  56683=>"000011011",
  56684=>"000101010",
  56685=>"111110111",
  56686=>"101111111",
  56687=>"001000000",
  56688=>"000111000",
  56689=>"011101110",
  56690=>"000110001",
  56691=>"110111111",
  56692=>"010111011",
  56693=>"100010000",
  56694=>"110100110",
  56695=>"101110110",
  56696=>"010010100",
  56697=>"001100011",
  56698=>"111001000",
  56699=>"100010001",
  56700=>"011000110",
  56701=>"010101000",
  56702=>"011111100",
  56703=>"110100111",
  56704=>"011010110",
  56705=>"100100010",
  56706=>"011111010",
  56707=>"101010000",
  56708=>"010000001",
  56709=>"011111100",
  56710=>"111101100",
  56711=>"000110011",
  56712=>"000100100",
  56713=>"001110001",
  56714=>"100010111",
  56715=>"000101000",
  56716=>"111111011",
  56717=>"110111100",
  56718=>"011110010",
  56719=>"001000100",
  56720=>"010010010",
  56721=>"110111111",
  56722=>"000000110",
  56723=>"100110001",
  56724=>"101110010",
  56725=>"000100010",
  56726=>"110111011",
  56727=>"001011111",
  56728=>"010111110",
  56729=>"110000101",
  56730=>"011011101",
  56731=>"010000110",
  56732=>"001111001",
  56733=>"000001111",
  56734=>"111101101",
  56735=>"000010100",
  56736=>"110000010",
  56737=>"010100010",
  56738=>"011010101",
  56739=>"111011111",
  56740=>"001000111",
  56741=>"001001000",
  56742=>"010010110",
  56743=>"001001110",
  56744=>"011010101",
  56745=>"011110010",
  56746=>"110100000",
  56747=>"101101110",
  56748=>"100010001",
  56749=>"111010000",
  56750=>"010001000",
  56751=>"111100101",
  56752=>"100001110",
  56753=>"100110000",
  56754=>"011110001",
  56755=>"100011111",
  56756=>"001010110",
  56757=>"100000101",
  56758=>"010000000",
  56759=>"111001011",
  56760=>"101100011",
  56761=>"001010110",
  56762=>"111101010",
  56763=>"111000011",
  56764=>"000101000",
  56765=>"010010000",
  56766=>"000011100",
  56767=>"010001101",
  56768=>"111010101",
  56769=>"101001001",
  56770=>"010110101",
  56771=>"000100100",
  56772=>"110000000",
  56773=>"011001100",
  56774=>"000000000",
  56775=>"010000000",
  56776=>"111101011",
  56777=>"011101110",
  56778=>"100010100",
  56779=>"011011111",
  56780=>"110110100",
  56781=>"101001110",
  56782=>"000110001",
  56783=>"000100010",
  56784=>"011111110",
  56785=>"101011100",
  56786=>"101110110",
  56787=>"010101010",
  56788=>"101000101",
  56789=>"000110001",
  56790=>"000010000",
  56791=>"101101101",
  56792=>"010010100",
  56793=>"100101000",
  56794=>"100001111",
  56795=>"011011000",
  56796=>"101110010",
  56797=>"000111000",
  56798=>"110001001",
  56799=>"001001111",
  56800=>"111010111",
  56801=>"010111111",
  56802=>"000001001",
  56803=>"000100111",
  56804=>"100100100",
  56805=>"100110100",
  56806=>"001100001",
  56807=>"100011111",
  56808=>"000000010",
  56809=>"101111000",
  56810=>"000010000",
  56811=>"100101011",
  56812=>"101000101",
  56813=>"011100000",
  56814=>"110000000",
  56815=>"000010100",
  56816=>"111110101",
  56817=>"101001110",
  56818=>"100011111",
  56819=>"101000111",
  56820=>"000100111",
  56821=>"010011111",
  56822=>"001100101",
  56823=>"101100001",
  56824=>"010100011",
  56825=>"000111111",
  56826=>"111011110",
  56827=>"011111101",
  56828=>"110011100",
  56829=>"011011000",
  56830=>"100001110",
  56831=>"000111001",
  56832=>"010100000",
  56833=>"110010011",
  56834=>"000000100",
  56835=>"000010000",
  56836=>"100111000",
  56837=>"001110101",
  56838=>"001000000",
  56839=>"001011011",
  56840=>"010001000",
  56841=>"101001010",
  56842=>"000010110",
  56843=>"101100000",
  56844=>"001100010",
  56845=>"010001011",
  56846=>"000101011",
  56847=>"011101110",
  56848=>"100000000",
  56849=>"111101010",
  56850=>"000001100",
  56851=>"100101001",
  56852=>"000000011",
  56853=>"010011011",
  56854=>"010000010",
  56855=>"111100000",
  56856=>"000011010",
  56857=>"001001011",
  56858=>"101001011",
  56859=>"000011111",
  56860=>"001001000",
  56861=>"011111010",
  56862=>"110010000",
  56863=>"101101011",
  56864=>"000100111",
  56865=>"101110100",
  56866=>"111110111",
  56867=>"001000111",
  56868=>"010010101",
  56869=>"010010010",
  56870=>"111111100",
  56871=>"111111100",
  56872=>"010010001",
  56873=>"101010110",
  56874=>"101100100",
  56875=>"000000001",
  56876=>"110000100",
  56877=>"001101010",
  56878=>"001100100",
  56879=>"111100110",
  56880=>"000011000",
  56881=>"010000011",
  56882=>"011000001",
  56883=>"111111101",
  56884=>"000100010",
  56885=>"110101110",
  56886=>"110111000",
  56887=>"111101000",
  56888=>"001101110",
  56889=>"000010000",
  56890=>"110010100",
  56891=>"100111100",
  56892=>"011100101",
  56893=>"000000111",
  56894=>"110001100",
  56895=>"110101110",
  56896=>"101110011",
  56897=>"111010001",
  56898=>"100111111",
  56899=>"001101010",
  56900=>"101011110",
  56901=>"111001010",
  56902=>"000010111",
  56903=>"010001000",
  56904=>"101011111",
  56905=>"100100100",
  56906=>"011110011",
  56907=>"000000011",
  56908=>"100110001",
  56909=>"101110110",
  56910=>"010000000",
  56911=>"011000001",
  56912=>"101111110",
  56913=>"110010000",
  56914=>"100001010",
  56915=>"011001101",
  56916=>"111100000",
  56917=>"010011010",
  56918=>"101000010",
  56919=>"111101110",
  56920=>"011100111",
  56921=>"000101011",
  56922=>"111110010",
  56923=>"011010111",
  56924=>"101010000",
  56925=>"101110010",
  56926=>"100111110",
  56927=>"011110101",
  56928=>"100100100",
  56929=>"010000101",
  56930=>"100100111",
  56931=>"001110000",
  56932=>"000100111",
  56933=>"101101001",
  56934=>"001101100",
  56935=>"101011001",
  56936=>"100011011",
  56937=>"000001100",
  56938=>"101101001",
  56939=>"111111110",
  56940=>"110010111",
  56941=>"111100010",
  56942=>"010110000",
  56943=>"001111101",
  56944=>"111000100",
  56945=>"000101000",
  56946=>"100111000",
  56947=>"010010101",
  56948=>"011101111",
  56949=>"010111000",
  56950=>"000010111",
  56951=>"111011111",
  56952=>"111010001",
  56953=>"001000111",
  56954=>"101110100",
  56955=>"010100010",
  56956=>"001001110",
  56957=>"101101111",
  56958=>"011010011",
  56959=>"001000000",
  56960=>"000000101",
  56961=>"111010100",
  56962=>"001001000",
  56963=>"001000010",
  56964=>"111000100",
  56965=>"010001001",
  56966=>"001110001",
  56967=>"101100110",
  56968=>"110100000",
  56969=>"011010101",
  56970=>"111000101",
  56971=>"011000000",
  56972=>"111010110",
  56973=>"100001000",
  56974=>"000100110",
  56975=>"001100001",
  56976=>"000001001",
  56977=>"110101000",
  56978=>"011111011",
  56979=>"000000111",
  56980=>"000110010",
  56981=>"110101101",
  56982=>"100011111",
  56983=>"100011111",
  56984=>"111111101",
  56985=>"001010011",
  56986=>"101010100",
  56987=>"101010110",
  56988=>"000000110",
  56989=>"000010100",
  56990=>"011011001",
  56991=>"000010010",
  56992=>"111011101",
  56993=>"110001100",
  56994=>"100001111",
  56995=>"110110000",
  56996=>"010110110",
  56997=>"110001011",
  56998=>"101000000",
  56999=>"010000110",
  57000=>"010101011",
  57001=>"010100000",
  57002=>"100110010",
  57003=>"101001000",
  57004=>"111111110",
  57005=>"001101110",
  57006=>"111110111",
  57007=>"101110000",
  57008=>"001001010",
  57009=>"101101000",
  57010=>"010000100",
  57011=>"111101110",
  57012=>"110111101",
  57013=>"001011010",
  57014=>"001001001",
  57015=>"000011000",
  57016=>"001011011",
  57017=>"100001110",
  57018=>"010011101",
  57019=>"110000101",
  57020=>"001010101",
  57021=>"100110000",
  57022=>"111011011",
  57023=>"011001001",
  57024=>"000010111",
  57025=>"000111000",
  57026=>"100111100",
  57027=>"001010000",
  57028=>"101100111",
  57029=>"011010001",
  57030=>"011000011",
  57031=>"101110000",
  57032=>"111001000",
  57033=>"110001010",
  57034=>"110000100",
  57035=>"111000011",
  57036=>"100110001",
  57037=>"000110101",
  57038=>"010001110",
  57039=>"010010001",
  57040=>"111000000",
  57041=>"000000011",
  57042=>"000000100",
  57043=>"111110101",
  57044=>"100010011",
  57045=>"100000011",
  57046=>"001111100",
  57047=>"110001000",
  57048=>"101101100",
  57049=>"001111101",
  57050=>"101101110",
  57051=>"100001111",
  57052=>"111110111",
  57053=>"110000111",
  57054=>"110010101",
  57055=>"000110111",
  57056=>"101111011",
  57057=>"111010010",
  57058=>"111101010",
  57059=>"001010111",
  57060=>"001010000",
  57061=>"111111101",
  57062=>"000000010",
  57063=>"011000101",
  57064=>"110001000",
  57065=>"010111101",
  57066=>"000000000",
  57067=>"001011001",
  57068=>"000001110",
  57069=>"000011111",
  57070=>"111101111",
  57071=>"001001111",
  57072=>"110010001",
  57073=>"010101100",
  57074=>"110010011",
  57075=>"111101001",
  57076=>"111010000",
  57077=>"011011111",
  57078=>"011010110",
  57079=>"111000000",
  57080=>"111100010",
  57081=>"110111011",
  57082=>"010000111",
  57083=>"011001001",
  57084=>"111110100",
  57085=>"100101011",
  57086=>"010011010",
  57087=>"111111111",
  57088=>"100001000",
  57089=>"101110110",
  57090=>"101001000",
  57091=>"011110011",
  57092=>"100110011",
  57093=>"111101011",
  57094=>"001101010",
  57095=>"000010110",
  57096=>"001011000",
  57097=>"100100110",
  57098=>"100110010",
  57099=>"011011110",
  57100=>"000000100",
  57101=>"110100101",
  57102=>"001000110",
  57103=>"100001110",
  57104=>"100010000",
  57105=>"000000001",
  57106=>"001001110",
  57107=>"111111110",
  57108=>"111001111",
  57109=>"010000110",
  57110=>"111101111",
  57111=>"110010101",
  57112=>"010010111",
  57113=>"000101001",
  57114=>"001011010",
  57115=>"101010101",
  57116=>"010011001",
  57117=>"011000001",
  57118=>"110001111",
  57119=>"111001000",
  57120=>"011111011",
  57121=>"110010111",
  57122=>"110000010",
  57123=>"111000100",
  57124=>"000010001",
  57125=>"010100000",
  57126=>"111000110",
  57127=>"000000010",
  57128=>"111000101",
  57129=>"000101100",
  57130=>"001010111",
  57131=>"100011101",
  57132=>"111111001",
  57133=>"111110111",
  57134=>"101001001",
  57135=>"111100000",
  57136=>"110001000",
  57137=>"000000111",
  57138=>"101111000",
  57139=>"001011001",
  57140=>"000010000",
  57141=>"011110000",
  57142=>"111111111",
  57143=>"011110010",
  57144=>"100000001",
  57145=>"010000110",
  57146=>"000111011",
  57147=>"001100101",
  57148=>"011101011",
  57149=>"111010010",
  57150=>"001100000",
  57151=>"011001101",
  57152=>"000101000",
  57153=>"001111100",
  57154=>"100010010",
  57155=>"000110010",
  57156=>"011000111",
  57157=>"101100000",
  57158=>"100011010",
  57159=>"110110010",
  57160=>"111011001",
  57161=>"010101100",
  57162=>"111011101",
  57163=>"000100010",
  57164=>"000011111",
  57165=>"000001000",
  57166=>"000111001",
  57167=>"110001110",
  57168=>"001001001",
  57169=>"010011010",
  57170=>"111001110",
  57171=>"001101010",
  57172=>"000110000",
  57173=>"100010001",
  57174=>"110000111",
  57175=>"111010101",
  57176=>"111000010",
  57177=>"010110011",
  57178=>"010001000",
  57179=>"001111111",
  57180=>"001010111",
  57181=>"110011100",
  57182=>"110010000",
  57183=>"000100001",
  57184=>"100010011",
  57185=>"000011000",
  57186=>"101010101",
  57187=>"011001110",
  57188=>"010011111",
  57189=>"001100011",
  57190=>"100101111",
  57191=>"000010101",
  57192=>"111101110",
  57193=>"101100111",
  57194=>"101001111",
  57195=>"011101001",
  57196=>"110111001",
  57197=>"100011100",
  57198=>"101000001",
  57199=>"110110001",
  57200=>"110101000",
  57201=>"000001001",
  57202=>"011001000",
  57203=>"011010101",
  57204=>"010111010",
  57205=>"000010011",
  57206=>"111110111",
  57207=>"101000100",
  57208=>"110010010",
  57209=>"111110010",
  57210=>"101010011",
  57211=>"110101001",
  57212=>"110000000",
  57213=>"001000000",
  57214=>"111100101",
  57215=>"000111000",
  57216=>"111111100",
  57217=>"011000111",
  57218=>"001100101",
  57219=>"111101000",
  57220=>"000001100",
  57221=>"000011100",
  57222=>"100100000",
  57223=>"001100110",
  57224=>"111000000",
  57225=>"111001110",
  57226=>"110000000",
  57227=>"001000000",
  57228=>"111111010",
  57229=>"111000110",
  57230=>"011111111",
  57231=>"111110000",
  57232=>"001111001",
  57233=>"001100010",
  57234=>"000001010",
  57235=>"101101111",
  57236=>"011010110",
  57237=>"111111111",
  57238=>"000001111",
  57239=>"111111110",
  57240=>"001101001",
  57241=>"000011001",
  57242=>"101010101",
  57243=>"011110110",
  57244=>"111000110",
  57245=>"100110010",
  57246=>"110000101",
  57247=>"001111101",
  57248=>"001110010",
  57249=>"110000010",
  57250=>"011110100",
  57251=>"101001001",
  57252=>"000100111",
  57253=>"110101101",
  57254=>"111110101",
  57255=>"110111101",
  57256=>"111011100",
  57257=>"110110011",
  57258=>"011100110",
  57259=>"111111110",
  57260=>"100100100",
  57261=>"101001001",
  57262=>"001010011",
  57263=>"111101011",
  57264=>"111111100",
  57265=>"001011101",
  57266=>"100111110",
  57267=>"111001100",
  57268=>"001101010",
  57269=>"100000101",
  57270=>"110100110",
  57271=>"001111010",
  57272=>"010011000",
  57273=>"100111000",
  57274=>"100011000",
  57275=>"010010100",
  57276=>"000001101",
  57277=>"111010101",
  57278=>"000101011",
  57279=>"001100011",
  57280=>"011100100",
  57281=>"000100010",
  57282=>"111000010",
  57283=>"100000011",
  57284=>"111010010",
  57285=>"011110101",
  57286=>"111011001",
  57287=>"111110010",
  57288=>"100010111",
  57289=>"010101000",
  57290=>"010010010",
  57291=>"011000011",
  57292=>"011001000",
  57293=>"111000000",
  57294=>"000011011",
  57295=>"000000010",
  57296=>"110000001",
  57297=>"010100111",
  57298=>"111001100",
  57299=>"001101001",
  57300=>"010000010",
  57301=>"011011101",
  57302=>"101100100",
  57303=>"000110010",
  57304=>"010111000",
  57305=>"100110111",
  57306=>"101110000",
  57307=>"000001001",
  57308=>"000110001",
  57309=>"101101100",
  57310=>"101111101",
  57311=>"100011011",
  57312=>"101111111",
  57313=>"000100010",
  57314=>"010101001",
  57315=>"100100000",
  57316=>"000100101",
  57317=>"011101110",
  57318=>"100001110",
  57319=>"111011000",
  57320=>"110100010",
  57321=>"000100100",
  57322=>"111011011",
  57323=>"100101110",
  57324=>"101110101",
  57325=>"001011000",
  57326=>"001101001",
  57327=>"011010101",
  57328=>"110110110",
  57329=>"101000111",
  57330=>"101101000",
  57331=>"000011011",
  57332=>"100000111",
  57333=>"011101010",
  57334=>"001100001",
  57335=>"111000111",
  57336=>"000101101",
  57337=>"011100111",
  57338=>"001111000",
  57339=>"011100111",
  57340=>"101111001",
  57341=>"101001101",
  57342=>"111101011",
  57343=>"111100111",
  57344=>"000100101",
  57345=>"101010000",
  57346=>"110110100",
  57347=>"101110010",
  57348=>"110000001",
  57349=>"111100101",
  57350=>"010111010",
  57351=>"001001111",
  57352=>"101100000",
  57353=>"000000011",
  57354=>"000001111",
  57355=>"101011111",
  57356=>"010000111",
  57357=>"101001011",
  57358=>"010000110",
  57359=>"011001000",
  57360=>"101100011",
  57361=>"100110011",
  57362=>"101111101",
  57363=>"110101111",
  57364=>"000111110",
  57365=>"010000000",
  57366=>"111100000",
  57367=>"111111011",
  57368=>"000111110",
  57369=>"010110011",
  57370=>"001001111",
  57371=>"000101111",
  57372=>"101101010",
  57373=>"101011011",
  57374=>"101110100",
  57375=>"101010100",
  57376=>"110101000",
  57377=>"010111100",
  57378=>"100100101",
  57379=>"000110011",
  57380=>"100101100",
  57381=>"010011111",
  57382=>"111110001",
  57383=>"111011011",
  57384=>"100100011",
  57385=>"100010001",
  57386=>"010001100",
  57387=>"111111111",
  57388=>"011001001",
  57389=>"101110001",
  57390=>"110011010",
  57391=>"001010101",
  57392=>"110111000",
  57393=>"110100101",
  57394=>"111111001",
  57395=>"101101001",
  57396=>"100001100",
  57397=>"111110000",
  57398=>"000101101",
  57399=>"101000101",
  57400=>"111011100",
  57401=>"000110001",
  57402=>"000010001",
  57403=>"000110010",
  57404=>"010101010",
  57405=>"000011011",
  57406=>"110100011",
  57407=>"101101001",
  57408=>"101111110",
  57409=>"011101100",
  57410=>"111111010",
  57411=>"110011110",
  57412=>"100100111",
  57413=>"001101101",
  57414=>"011000000",
  57415=>"111111011",
  57416=>"101000011",
  57417=>"001110000",
  57418=>"100110000",
  57419=>"010101111",
  57420=>"101101000",
  57421=>"100101110",
  57422=>"011011010",
  57423=>"100100001",
  57424=>"011010100",
  57425=>"010111101",
  57426=>"001000001",
  57427=>"101000011",
  57428=>"100011001",
  57429=>"010001110",
  57430=>"100011101",
  57431=>"100101111",
  57432=>"111001000",
  57433=>"011001000",
  57434=>"111110110",
  57435=>"101001011",
  57436=>"101001001",
  57437=>"100010010",
  57438=>"011010110",
  57439=>"001001111",
  57440=>"010001100",
  57441=>"101001010",
  57442=>"000000011",
  57443=>"110110011",
  57444=>"100011001",
  57445=>"101011000",
  57446=>"001100001",
  57447=>"000100000",
  57448=>"000111111",
  57449=>"011100000",
  57450=>"101001111",
  57451=>"101001101",
  57452=>"111000011",
  57453=>"011001010",
  57454=>"101100000",
  57455=>"010010100",
  57456=>"001011111",
  57457=>"010000111",
  57458=>"101000101",
  57459=>"100111110",
  57460=>"011110001",
  57461=>"011111101",
  57462=>"010101010",
  57463=>"110100010",
  57464=>"110000000",
  57465=>"000101010",
  57466=>"101001001",
  57467=>"110110001",
  57468=>"000000100",
  57469=>"100110010",
  57470=>"001111010",
  57471=>"111011000",
  57472=>"111001101",
  57473=>"111011001",
  57474=>"101000100",
  57475=>"101011101",
  57476=>"111110110",
  57477=>"011011100",
  57478=>"110011100",
  57479=>"000110111",
  57480=>"001111010",
  57481=>"010010010",
  57482=>"100000100",
  57483=>"001110101",
  57484=>"001000001",
  57485=>"011111110",
  57486=>"011011010",
  57487=>"001111101",
  57488=>"100101010",
  57489=>"010111000",
  57490=>"000110111",
  57491=>"001010111",
  57492=>"010110100",
  57493=>"010111110",
  57494=>"001111111",
  57495=>"000001111",
  57496=>"001000110",
  57497=>"010110111",
  57498=>"011000001",
  57499=>"001101110",
  57500=>"000111000",
  57501=>"100111000",
  57502=>"100111011",
  57503=>"101011000",
  57504=>"001110110",
  57505=>"100101011",
  57506=>"000000110",
  57507=>"100001100",
  57508=>"100010011",
  57509=>"000111000",
  57510=>"101100001",
  57511=>"110110000",
  57512=>"110010110",
  57513=>"011011111",
  57514=>"110000000",
  57515=>"110001101",
  57516=>"111001110",
  57517=>"101111101",
  57518=>"110111001",
  57519=>"010110011",
  57520=>"100011000",
  57521=>"011011110",
  57522=>"111110010",
  57523=>"101100101",
  57524=>"100010110",
  57525=>"000100010",
  57526=>"001011111",
  57527=>"110100010",
  57528=>"000100100",
  57529=>"010110011",
  57530=>"110110011",
  57531=>"110001111",
  57532=>"101101010",
  57533=>"000011100",
  57534=>"111011001",
  57535=>"001111111",
  57536=>"101001010",
  57537=>"001000000",
  57538=>"111111001",
  57539=>"111101110",
  57540=>"111110100",
  57541=>"010010001",
  57542=>"010100100",
  57543=>"011000000",
  57544=>"011000010",
  57545=>"010000110",
  57546=>"101001011",
  57547=>"111000111",
  57548=>"011101101",
  57549=>"101010001",
  57550=>"001001100",
  57551=>"101001010",
  57552=>"010010101",
  57553=>"001110101",
  57554=>"001001010",
  57555=>"000001101",
  57556=>"001000100",
  57557=>"000100111",
  57558=>"101111000",
  57559=>"010101100",
  57560=>"001011000",
  57561=>"100011110",
  57562=>"110100111",
  57563=>"111110001",
  57564=>"010000100",
  57565=>"001011111",
  57566=>"101001011",
  57567=>"001111011",
  57568=>"101100111",
  57569=>"001000010",
  57570=>"000010101",
  57571=>"110111100",
  57572=>"111111100",
  57573=>"000110010",
  57574=>"110101110",
  57575=>"000101110",
  57576=>"000001001",
  57577=>"001010100",
  57578=>"000010101",
  57579=>"110000011",
  57580=>"011111001",
  57581=>"101111010",
  57582=>"110000111",
  57583=>"011111111",
  57584=>"110110100",
  57585=>"010001010",
  57586=>"000110001",
  57587=>"001011110",
  57588=>"001010101",
  57589=>"001110110",
  57590=>"001001111",
  57591=>"000000100",
  57592=>"011010111",
  57593=>"010010101",
  57594=>"111010101",
  57595=>"010010110",
  57596=>"011110110",
  57597=>"010101001",
  57598=>"111101000",
  57599=>"000100001",
  57600=>"001000101",
  57601=>"010011101",
  57602=>"011110110",
  57603=>"010000101",
  57604=>"010010011",
  57605=>"001111111",
  57606=>"110100100",
  57607=>"000100011",
  57608=>"010110111",
  57609=>"101111111",
  57610=>"000000001",
  57611=>"110100010",
  57612=>"011010000",
  57613=>"001000001",
  57614=>"011011001",
  57615=>"111110001",
  57616=>"010110001",
  57617=>"001011010",
  57618=>"111000010",
  57619=>"001110100",
  57620=>"000101101",
  57621=>"100000110",
  57622=>"010011010",
  57623=>"110101011",
  57624=>"111100101",
  57625=>"100100110",
  57626=>"010001111",
  57627=>"001010000",
  57628=>"110011101",
  57629=>"100000011",
  57630=>"101110000",
  57631=>"101110100",
  57632=>"010010010",
  57633=>"110010111",
  57634=>"001000011",
  57635=>"110001000",
  57636=>"011111011",
  57637=>"000000011",
  57638=>"001011001",
  57639=>"110010011",
  57640=>"011101100",
  57641=>"010010100",
  57642=>"000000100",
  57643=>"110010000",
  57644=>"101011010",
  57645=>"110101101",
  57646=>"000111101",
  57647=>"110000110",
  57648=>"000011101",
  57649=>"110010100",
  57650=>"110000000",
  57651=>"111111111",
  57652=>"100111101",
  57653=>"001011100",
  57654=>"011000100",
  57655=>"011001011",
  57656=>"010000000",
  57657=>"001000000",
  57658=>"011010111",
  57659=>"101001111",
  57660=>"000101110",
  57661=>"010000111",
  57662=>"001111010",
  57663=>"101010010",
  57664=>"100011010",
  57665=>"010001010",
  57666=>"000011001",
  57667=>"001100111",
  57668=>"101111001",
  57669=>"011111001",
  57670=>"101101011",
  57671=>"111101011",
  57672=>"101100010",
  57673=>"110010101",
  57674=>"101110111",
  57675=>"111111001",
  57676=>"101101100",
  57677=>"000010110",
  57678=>"000100111",
  57679=>"101010000",
  57680=>"101011011",
  57681=>"010011101",
  57682=>"101011001",
  57683=>"100011110",
  57684=>"100011010",
  57685=>"100101010",
  57686=>"001100101",
  57687=>"001010000",
  57688=>"000110001",
  57689=>"110001000",
  57690=>"010001001",
  57691=>"011111101",
  57692=>"000100011",
  57693=>"000000111",
  57694=>"110011100",
  57695=>"110111110",
  57696=>"000110011",
  57697=>"100111100",
  57698=>"101110000",
  57699=>"010100111",
  57700=>"010001001",
  57701=>"010100111",
  57702=>"101001010",
  57703=>"011000101",
  57704=>"110101111",
  57705=>"111001000",
  57706=>"011001011",
  57707=>"100100010",
  57708=>"011101111",
  57709=>"010000010",
  57710=>"001000110",
  57711=>"100010000",
  57712=>"001011110",
  57713=>"101010111",
  57714=>"000101100",
  57715=>"011110101",
  57716=>"110101000",
  57717=>"101000100",
  57718=>"110110101",
  57719=>"111100111",
  57720=>"100110101",
  57721=>"011010110",
  57722=>"101101110",
  57723=>"011100101",
  57724=>"000000111",
  57725=>"000000011",
  57726=>"000010111",
  57727=>"000010011",
  57728=>"010001011",
  57729=>"101100010",
  57730=>"001000000",
  57731=>"111001000",
  57732=>"001000111",
  57733=>"010001000",
  57734=>"011000000",
  57735=>"111111110",
  57736=>"001111100",
  57737=>"001010110",
  57738=>"010111010",
  57739=>"111010010",
  57740=>"110001100",
  57741=>"001011101",
  57742=>"100001001",
  57743=>"110100010",
  57744=>"001110010",
  57745=>"000111010",
  57746=>"011000111",
  57747=>"100101100",
  57748=>"010101000",
  57749=>"000111011",
  57750=>"101001000",
  57751=>"111000010",
  57752=>"011001110",
  57753=>"010100000",
  57754=>"010110010",
  57755=>"010010000",
  57756=>"110001010",
  57757=>"001101000",
  57758=>"100110000",
  57759=>"001101001",
  57760=>"101111100",
  57761=>"010000011",
  57762=>"010000110",
  57763=>"000011010",
  57764=>"010001101",
  57765=>"011011001",
  57766=>"111111010",
  57767=>"000111110",
  57768=>"111010010",
  57769=>"111101001",
  57770=>"000010101",
  57771=>"000110110",
  57772=>"101011110",
  57773=>"111000000",
  57774=>"110101010",
  57775=>"101111001",
  57776=>"000000001",
  57777=>"010001110",
  57778=>"001110100",
  57779=>"010011010",
  57780=>"110000111",
  57781=>"011111000",
  57782=>"111000000",
  57783=>"001011111",
  57784=>"111110010",
  57785=>"111101000",
  57786=>"000111111",
  57787=>"110101010",
  57788=>"110111111",
  57789=>"111000101",
  57790=>"111001011",
  57791=>"001000101",
  57792=>"010100011",
  57793=>"101101100",
  57794=>"000110101",
  57795=>"011111010",
  57796=>"101101011",
  57797=>"000000101",
  57798=>"001000001",
  57799=>"100100111",
  57800=>"001000011",
  57801=>"100000011",
  57802=>"110111011",
  57803=>"101101100",
  57804=>"010111101",
  57805=>"000010010",
  57806=>"011110111",
  57807=>"111011011",
  57808=>"111110001",
  57809=>"100100100",
  57810=>"101011111",
  57811=>"100101011",
  57812=>"100010010",
  57813=>"111001011",
  57814=>"100000010",
  57815=>"100010010",
  57816=>"010111000",
  57817=>"011101101",
  57818=>"011011000",
  57819=>"100001011",
  57820=>"100101011",
  57821=>"010010011",
  57822=>"100101100",
  57823=>"001100100",
  57824=>"111100111",
  57825=>"011000000",
  57826=>"100101101",
  57827=>"010101010",
  57828=>"011000100",
  57829=>"011011010",
  57830=>"011010001",
  57831=>"001011111",
  57832=>"010110000",
  57833=>"000011010",
  57834=>"011000000",
  57835=>"011101110",
  57836=>"010010001",
  57837=>"101111101",
  57838=>"111111111",
  57839=>"101010000",
  57840=>"101000010",
  57841=>"101000011",
  57842=>"110101000",
  57843=>"111101010",
  57844=>"001010100",
  57845=>"100100101",
  57846=>"001100001",
  57847=>"011011000",
  57848=>"011111110",
  57849=>"010111111",
  57850=>"001101110",
  57851=>"000110100",
  57852=>"000110110",
  57853=>"101001000",
  57854=>"110100011",
  57855=>"011011110",
  57856=>"001000011",
  57857=>"010100100",
  57858=>"100001111",
  57859=>"010011000",
  57860=>"101100011",
  57861=>"000001100",
  57862=>"000010000",
  57863=>"010010001",
  57864=>"000010100",
  57865=>"011100011",
  57866=>"001001010",
  57867=>"100100011",
  57868=>"111111000",
  57869=>"000110101",
  57870=>"111110000",
  57871=>"101011000",
  57872=>"000001001",
  57873=>"000000111",
  57874=>"000111100",
  57875=>"000001110",
  57876=>"101010100",
  57877=>"010000000",
  57878=>"111110101",
  57879=>"010001100",
  57880=>"011011011",
  57881=>"011101101",
  57882=>"011010101",
  57883=>"000100000",
  57884=>"111100001",
  57885=>"011100010",
  57886=>"100111101",
  57887=>"010010011",
  57888=>"000000101",
  57889=>"110000000",
  57890=>"000100011",
  57891=>"111000110",
  57892=>"001100100",
  57893=>"000000001",
  57894=>"001011101",
  57895=>"111111010",
  57896=>"101111001",
  57897=>"001010010",
  57898=>"100000001",
  57899=>"001101011",
  57900=>"001000011",
  57901=>"111110101",
  57902=>"101111000",
  57903=>"011011000",
  57904=>"010000101",
  57905=>"101100010",
  57906=>"000000011",
  57907=>"010110001",
  57908=>"011111101",
  57909=>"011001000",
  57910=>"110101001",
  57911=>"101001111",
  57912=>"001000111",
  57913=>"100000000",
  57914=>"100111100",
  57915=>"010001001",
  57916=>"011111010",
  57917=>"010111001",
  57918=>"111100011",
  57919=>"101101110",
  57920=>"111101111",
  57921=>"010000100",
  57922=>"001100110",
  57923=>"110000000",
  57924=>"100111111",
  57925=>"101100101",
  57926=>"111000111",
  57927=>"000111000",
  57928=>"000011000",
  57929=>"101001100",
  57930=>"111010110",
  57931=>"101011100",
  57932=>"111000101",
  57933=>"010010011",
  57934=>"110011101",
  57935=>"101110110",
  57936=>"001111100",
  57937=>"100000101",
  57938=>"011001101",
  57939=>"000101100",
  57940=>"111011100",
  57941=>"100111110",
  57942=>"000010111",
  57943=>"100010100",
  57944=>"110111100",
  57945=>"101101000",
  57946=>"101010110",
  57947=>"010110001",
  57948=>"101010011",
  57949=>"101111010",
  57950=>"100001110",
  57951=>"111111011",
  57952=>"111001010",
  57953=>"100000111",
  57954=>"001101010",
  57955=>"001001101",
  57956=>"001100110",
  57957=>"001000101",
  57958=>"101110110",
  57959=>"011101010",
  57960=>"111001010",
  57961=>"110001110",
  57962=>"100011111",
  57963=>"011010010",
  57964=>"110101101",
  57965=>"101101100",
  57966=>"111001110",
  57967=>"010100000",
  57968=>"110100001",
  57969=>"001011011",
  57970=>"111000111",
  57971=>"001010001",
  57972=>"110010001",
  57973=>"101101001",
  57974=>"111111010",
  57975=>"110101100",
  57976=>"011111110",
  57977=>"010110001",
  57978=>"011100101",
  57979=>"001000011",
  57980=>"101100000",
  57981=>"111100111",
  57982=>"000011100",
  57983=>"000100000",
  57984=>"110110010",
  57985=>"000000000",
  57986=>"101101010",
  57987=>"101110011",
  57988=>"110100111",
  57989=>"111111101",
  57990=>"111110010",
  57991=>"011111111",
  57992=>"111111101",
  57993=>"000111010",
  57994=>"000010001",
  57995=>"100111100",
  57996=>"111111011",
  57997=>"010000001",
  57998=>"110001010",
  57999=>"110000011",
  58000=>"110100101",
  58001=>"110101000",
  58002=>"110111001",
  58003=>"101101011",
  58004=>"110011010",
  58005=>"000010011",
  58006=>"100100010",
  58007=>"111101111",
  58008=>"111111000",
  58009=>"000101111",
  58010=>"110010001",
  58011=>"010100101",
  58012=>"010000111",
  58013=>"110001111",
  58014=>"110011110",
  58015=>"100100110",
  58016=>"000001001",
  58017=>"011001001",
  58018=>"010000101",
  58019=>"111000010",
  58020=>"111111111",
  58021=>"000100011",
  58022=>"011111011",
  58023=>"100000010",
  58024=>"000110011",
  58025=>"000100101",
  58026=>"011001101",
  58027=>"001100101",
  58028=>"001101000",
  58029=>"000010100",
  58030=>"011000010",
  58031=>"010001110",
  58032=>"000111111",
  58033=>"001001011",
  58034=>"000100010",
  58035=>"110100010",
  58036=>"010111000",
  58037=>"011011100",
  58038=>"110001000",
  58039=>"111001011",
  58040=>"000011101",
  58041=>"110001110",
  58042=>"011011011",
  58043=>"010110001",
  58044=>"111010000",
  58045=>"011111010",
  58046=>"101111011",
  58047=>"011011000",
  58048=>"111100010",
  58049=>"011010000",
  58050=>"101111011",
  58051=>"111001101",
  58052=>"010010101",
  58053=>"001000011",
  58054=>"010110101",
  58055=>"011101000",
  58056=>"001101111",
  58057=>"110010100",
  58058=>"001111001",
  58059=>"110011110",
  58060=>"000110000",
  58061=>"000100000",
  58062=>"011000010",
  58063=>"001001101",
  58064=>"001001111",
  58065=>"100010111",
  58066=>"100010110",
  58067=>"010000011",
  58068=>"000001001",
  58069=>"111111111",
  58070=>"111001101",
  58071=>"000010011",
  58072=>"101001011",
  58073=>"101100001",
  58074=>"110011000",
  58075=>"100000010",
  58076=>"010110100",
  58077=>"010100010",
  58078=>"011100111",
  58079=>"011111100",
  58080=>"000000111",
  58081=>"001001010",
  58082=>"000011010",
  58083=>"101101111",
  58084=>"111010010",
  58085=>"000111100",
  58086=>"001101011",
  58087=>"010001010",
  58088=>"000100110",
  58089=>"010111110",
  58090=>"100001111",
  58091=>"011111100",
  58092=>"000011101",
  58093=>"110100101",
  58094=>"110100011",
  58095=>"000001111",
  58096=>"101010100",
  58097=>"000100010",
  58098=>"001000111",
  58099=>"001100111",
  58100=>"001111100",
  58101=>"110010101",
  58102=>"111011011",
  58103=>"000000110",
  58104=>"110010110",
  58105=>"010010111",
  58106=>"101000111",
  58107=>"000101001",
  58108=>"010110001",
  58109=>"011000110",
  58110=>"010101111",
  58111=>"111001011",
  58112=>"001000001",
  58113=>"001000110",
  58114=>"011111101",
  58115=>"001001010",
  58116=>"000000100",
  58117=>"010000000",
  58118=>"100111100",
  58119=>"100111010",
  58120=>"110010100",
  58121=>"110100001",
  58122=>"000100010",
  58123=>"100111001",
  58124=>"000101000",
  58125=>"110011111",
  58126=>"111011010",
  58127=>"011001110",
  58128=>"110000100",
  58129=>"001111100",
  58130=>"001111011",
  58131=>"100101001",
  58132=>"011000100",
  58133=>"111110111",
  58134=>"011001110",
  58135=>"010000100",
  58136=>"000110000",
  58137=>"001001111",
  58138=>"111001101",
  58139=>"101001000",
  58140=>"111101000",
  58141=>"101101001",
  58142=>"010000111",
  58143=>"001110111",
  58144=>"001000010",
  58145=>"101110011",
  58146=>"001011011",
  58147=>"100011001",
  58148=>"000100101",
  58149=>"001001111",
  58150=>"011011110",
  58151=>"000111011",
  58152=>"000011110",
  58153=>"001000110",
  58154=>"100100110",
  58155=>"010101000",
  58156=>"110101110",
  58157=>"011101111",
  58158=>"000011111",
  58159=>"110010001",
  58160=>"110101001",
  58161=>"101000010",
  58162=>"111111100",
  58163=>"101010110",
  58164=>"011000101",
  58165=>"100100110",
  58166=>"110111000",
  58167=>"110010001",
  58168=>"101000000",
  58169=>"110000101",
  58170=>"000000100",
  58171=>"001110000",
  58172=>"000100111",
  58173=>"110101111",
  58174=>"010111001",
  58175=>"011100010",
  58176=>"011110000",
  58177=>"100111000",
  58178=>"111100011",
  58179=>"000000000",
  58180=>"000000000",
  58181=>"100010100",
  58182=>"100110101",
  58183=>"001110110",
  58184=>"000100100",
  58185=>"110011111",
  58186=>"100010000",
  58187=>"011100010",
  58188=>"000001111",
  58189=>"010001010",
  58190=>"011000000",
  58191=>"001011101",
  58192=>"100111001",
  58193=>"111000001",
  58194=>"011100111",
  58195=>"010000001",
  58196=>"000001011",
  58197=>"110110110",
  58198=>"101110111",
  58199=>"111011000",
  58200=>"011100000",
  58201=>"011010110",
  58202=>"011110011",
  58203=>"100101011",
  58204=>"011100000",
  58205=>"101100100",
  58206=>"011001011",
  58207=>"001101101",
  58208=>"010110111",
  58209=>"101000111",
  58210=>"100110110",
  58211=>"101010100",
  58212=>"100111010",
  58213=>"111001111",
  58214=>"100100110",
  58215=>"001000110",
  58216=>"101010100",
  58217=>"100010011",
  58218=>"001001101",
  58219=>"000000000",
  58220=>"101101001",
  58221=>"101001101",
  58222=>"100000100",
  58223=>"111001111",
  58224=>"010000000",
  58225=>"001010101",
  58226=>"111000111",
  58227=>"000011001",
  58228=>"110001101",
  58229=>"101111111",
  58230=>"110001011",
  58231=>"111100000",
  58232=>"001001011",
  58233=>"100111010",
  58234=>"011110111",
  58235=>"100001011",
  58236=>"000100010",
  58237=>"110010101",
  58238=>"001000110",
  58239=>"110111011",
  58240=>"000110100",
  58241=>"110100100",
  58242=>"101101001",
  58243=>"100001011",
  58244=>"111101101",
  58245=>"010000000",
  58246=>"001000110",
  58247=>"010001000",
  58248=>"100101010",
  58249=>"000111011",
  58250=>"000000110",
  58251=>"010001100",
  58252=>"100001010",
  58253=>"010101100",
  58254=>"001001110",
  58255=>"111110010",
  58256=>"000100100",
  58257=>"110110100",
  58258=>"110001100",
  58259=>"010011001",
  58260=>"101011001",
  58261=>"111011100",
  58262=>"001101000",
  58263=>"111001000",
  58264=>"001011101",
  58265=>"110010110",
  58266=>"010111010",
  58267=>"100111011",
  58268=>"111000011",
  58269=>"111000011",
  58270=>"001100101",
  58271=>"011100001",
  58272=>"111110000",
  58273=>"101010000",
  58274=>"111100001",
  58275=>"010100011",
  58276=>"010001010",
  58277=>"000100001",
  58278=>"101000100",
  58279=>"101001110",
  58280=>"000111011",
  58281=>"000110100",
  58282=>"110000000",
  58283=>"000110010",
  58284=>"111011001",
  58285=>"101110001",
  58286=>"100111110",
  58287=>"011000001",
  58288=>"100010011",
  58289=>"110001001",
  58290=>"000001010",
  58291=>"011010110",
  58292=>"101111111",
  58293=>"101011110",
  58294=>"111101100",
  58295=>"110110111",
  58296=>"000101000",
  58297=>"101000101",
  58298=>"101101100",
  58299=>"111000000",
  58300=>"101010111",
  58301=>"110011101",
  58302=>"100010111",
  58303=>"000100100",
  58304=>"111110111",
  58305=>"010000101",
  58306=>"100101101",
  58307=>"010000100",
  58308=>"100111110",
  58309=>"111111000",
  58310=>"111111100",
  58311=>"110110110",
  58312=>"100100010",
  58313=>"001110001",
  58314=>"110010110",
  58315=>"111100010",
  58316=>"000100110",
  58317=>"110111111",
  58318=>"000001001",
  58319=>"001011111",
  58320=>"101111010",
  58321=>"010010011",
  58322=>"011100000",
  58323=>"001101101",
  58324=>"011111110",
  58325=>"000010010",
  58326=>"101101101",
  58327=>"101000100",
  58328=>"000000110",
  58329=>"010101001",
  58330=>"011011001",
  58331=>"101010101",
  58332=>"100100010",
  58333=>"000100111",
  58334=>"110010110",
  58335=>"011111110",
  58336=>"111010111",
  58337=>"111110011",
  58338=>"011011000",
  58339=>"101101101",
  58340=>"110011001",
  58341=>"010010101",
  58342=>"001000000",
  58343=>"111011010",
  58344=>"010101111",
  58345=>"010101110",
  58346=>"110000000",
  58347=>"010011010",
  58348=>"101100110",
  58349=>"101010001",
  58350=>"100011011",
  58351=>"000010100",
  58352=>"011001000",
  58353=>"111111100",
  58354=>"111011010",
  58355=>"001100011",
  58356=>"000101011",
  58357=>"001100101",
  58358=>"001111110",
  58359=>"110101111",
  58360=>"101101010",
  58361=>"111101010",
  58362=>"001100011",
  58363=>"111101111",
  58364=>"101011111",
  58365=>"011100010",
  58366=>"100011110",
  58367=>"001000010",
  58368=>"111101111",
  58369=>"101101001",
  58370=>"111010000",
  58371=>"000010011",
  58372=>"011111101",
  58373=>"101001111",
  58374=>"000110100",
  58375=>"111111010",
  58376=>"110111001",
  58377=>"000001011",
  58378=>"100101111",
  58379=>"000111011",
  58380=>"111110010",
  58381=>"101110111",
  58382=>"111011101",
  58383=>"000001111",
  58384=>"011011001",
  58385=>"100010110",
  58386=>"011111011",
  58387=>"111010001",
  58388=>"000110001",
  58389=>"111001100",
  58390=>"100100010",
  58391=>"001001101",
  58392=>"111101111",
  58393=>"010000100",
  58394=>"101011000",
  58395=>"011010100",
  58396=>"101101110",
  58397=>"110011010",
  58398=>"010001100",
  58399=>"001001010",
  58400=>"001100011",
  58401=>"010110101",
  58402=>"110111111",
  58403=>"111101110",
  58404=>"011010100",
  58405=>"100110110",
  58406=>"101010111",
  58407=>"101110011",
  58408=>"100000001",
  58409=>"000001011",
  58410=>"110101011",
  58411=>"000001000",
  58412=>"110000110",
  58413=>"101010000",
  58414=>"010101011",
  58415=>"010010100",
  58416=>"010010000",
  58417=>"001100110",
  58418=>"111011101",
  58419=>"101000000",
  58420=>"100110000",
  58421=>"010100000",
  58422=>"100000101",
  58423=>"010001111",
  58424=>"100011101",
  58425=>"010011111",
  58426=>"000011101",
  58427=>"111010100",
  58428=>"101101011",
  58429=>"101110111",
  58430=>"111001100",
  58431=>"001011101",
  58432=>"001010110",
  58433=>"111011000",
  58434=>"011001100",
  58435=>"100001000",
  58436=>"000001010",
  58437=>"001000110",
  58438=>"011101000",
  58439=>"001111101",
  58440=>"111011100",
  58441=>"001111111",
  58442=>"100101110",
  58443=>"110000000",
  58444=>"110100100",
  58445=>"011010000",
  58446=>"001110000",
  58447=>"001000011",
  58448=>"111101100",
  58449=>"111110110",
  58450=>"000110000",
  58451=>"100100100",
  58452=>"011101000",
  58453=>"001010100",
  58454=>"110011011",
  58455=>"100111111",
  58456=>"011010010",
  58457=>"101001100",
  58458=>"011000011",
  58459=>"000001010",
  58460=>"000101101",
  58461=>"011001001",
  58462=>"010010000",
  58463=>"110011110",
  58464=>"011000100",
  58465=>"001110010",
  58466=>"011111111",
  58467=>"010011010",
  58468=>"110001010",
  58469=>"000101000",
  58470=>"110111011",
  58471=>"000000100",
  58472=>"110111011",
  58473=>"110001101",
  58474=>"000001011",
  58475=>"100011011",
  58476=>"110101110",
  58477=>"100001010",
  58478=>"011100001",
  58479=>"011101001",
  58480=>"110001100",
  58481=>"111010111",
  58482=>"000001100",
  58483=>"010100011",
  58484=>"010000100",
  58485=>"001000100",
  58486=>"111000000",
  58487=>"111010101",
  58488=>"111111000",
  58489=>"111011010",
  58490=>"111110100",
  58491=>"000000011",
  58492=>"000000001",
  58493=>"110000100",
  58494=>"101100011",
  58495=>"010101000",
  58496=>"111010010",
  58497=>"101001101",
  58498=>"010000100",
  58499=>"100101011",
  58500=>"110001110",
  58501=>"001100001",
  58502=>"011110010",
  58503=>"111010111",
  58504=>"101100101",
  58505=>"101011110",
  58506=>"111000100",
  58507=>"010011111",
  58508=>"100110111",
  58509=>"011110011",
  58510=>"101001110",
  58511=>"001101010",
  58512=>"100111001",
  58513=>"001000111",
  58514=>"100100000",
  58515=>"001110111",
  58516=>"011100100",
  58517=>"001101101",
  58518=>"110010011",
  58519=>"001111111",
  58520=>"100000011",
  58521=>"111101101",
  58522=>"010110010",
  58523=>"101111100",
  58524=>"100111110",
  58525=>"011111000",
  58526=>"010010110",
  58527=>"110100010",
  58528=>"100100101",
  58529=>"000110100",
  58530=>"001110110",
  58531=>"010111110",
  58532=>"100111011",
  58533=>"111110100",
  58534=>"101001100",
  58535=>"000100010",
  58536=>"001100101",
  58537=>"100010001",
  58538=>"101011000",
  58539=>"101011101",
  58540=>"001001001",
  58541=>"100000010",
  58542=>"001010011",
  58543=>"010111011",
  58544=>"000011100",
  58545=>"010011101",
  58546=>"100001010",
  58547=>"000111001",
  58548=>"101101011",
  58549=>"111001110",
  58550=>"101010111",
  58551=>"011011010",
  58552=>"011100010",
  58553=>"000011000",
  58554=>"111001100",
  58555=>"111101111",
  58556=>"100111011",
  58557=>"101111110",
  58558=>"111110110",
  58559=>"101011110",
  58560=>"110111110",
  58561=>"000101111",
  58562=>"010100010",
  58563=>"111101110",
  58564=>"001010010",
  58565=>"000010011",
  58566=>"010100101",
  58567=>"011110111",
  58568=>"101011001",
  58569=>"000111000",
  58570=>"010001100",
  58571=>"110101111",
  58572=>"011001001",
  58573=>"111101000",
  58574=>"100001011",
  58575=>"000110110",
  58576=>"111011011",
  58577=>"011010100",
  58578=>"110110110",
  58579=>"010000000",
  58580=>"111001010",
  58581=>"011000001",
  58582=>"101000010",
  58583=>"010011010",
  58584=>"010101000",
  58585=>"110110000",
  58586=>"010100011",
  58587=>"110011011",
  58588=>"000011010",
  58589=>"101000100",
  58590=>"111001100",
  58591=>"110110000",
  58592=>"110010101",
  58593=>"010110101",
  58594=>"100001001",
  58595=>"010001100",
  58596=>"100100101",
  58597=>"011101010",
  58598=>"011000010",
  58599=>"100001011",
  58600=>"001101100",
  58601=>"000110011",
  58602=>"110110010",
  58603=>"100110111",
  58604=>"000011100",
  58605=>"010100011",
  58606=>"101001010",
  58607=>"001000011",
  58608=>"111001001",
  58609=>"001011000",
  58610=>"111000101",
  58611=>"101000000",
  58612=>"000110010",
  58613=>"000001000",
  58614=>"000001110",
  58615=>"000001110",
  58616=>"000011001",
  58617=>"001100010",
  58618=>"001011000",
  58619=>"011100111",
  58620=>"001000100",
  58621=>"001000001",
  58622=>"011011011",
  58623=>"000011010",
  58624=>"110011101",
  58625=>"000101101",
  58626=>"111111001",
  58627=>"001000100",
  58628=>"010001001",
  58629=>"010111111",
  58630=>"000000100",
  58631=>"101111110",
  58632=>"010001111",
  58633=>"001111100",
  58634=>"011011101",
  58635=>"010110010",
  58636=>"000111110",
  58637=>"100110010",
  58638=>"011111100",
  58639=>"100101100",
  58640=>"001110000",
  58641=>"011110101",
  58642=>"010110111",
  58643=>"010000111",
  58644=>"010001001",
  58645=>"011001011",
  58646=>"100001001",
  58647=>"100000100",
  58648=>"111111101",
  58649=>"010100100",
  58650=>"010001110",
  58651=>"111110110",
  58652=>"001000000",
  58653=>"101100010",
  58654=>"110111110",
  58655=>"010000000",
  58656=>"000100100",
  58657=>"110001110",
  58658=>"101011000",
  58659=>"101110000",
  58660=>"100100100",
  58661=>"000011001",
  58662=>"101000101",
  58663=>"000010110",
  58664=>"001110100",
  58665=>"100010011",
  58666=>"011111001",
  58667=>"100001010",
  58668=>"001000100",
  58669=>"011111010",
  58670=>"000001101",
  58671=>"101010011",
  58672=>"000001101",
  58673=>"001111101",
  58674=>"000011101",
  58675=>"000110101",
  58676=>"010000101",
  58677=>"111100101",
  58678=>"100001110",
  58679=>"000010000",
  58680=>"111000000",
  58681=>"101001111",
  58682=>"000001111",
  58683=>"011011010",
  58684=>"111011101",
  58685=>"011001110",
  58686=>"011110001",
  58687=>"101110010",
  58688=>"011111001",
  58689=>"011010000",
  58690=>"111101100",
  58691=>"100011101",
  58692=>"011101111",
  58693=>"101110011",
  58694=>"101000100",
  58695=>"111111110",
  58696=>"001100011",
  58697=>"101001000",
  58698=>"110000000",
  58699=>"101100100",
  58700=>"110100010",
  58701=>"000111110",
  58702=>"110110111",
  58703=>"111110100",
  58704=>"010100100",
  58705=>"000010110",
  58706=>"111001000",
  58707=>"001100101",
  58708=>"010100100",
  58709=>"010001010",
  58710=>"101000111",
  58711=>"011001011",
  58712=>"001111110",
  58713=>"100010100",
  58714=>"100000010",
  58715=>"111000000",
  58716=>"101011011",
  58717=>"011110101",
  58718=>"100000110",
  58719=>"011011010",
  58720=>"001101110",
  58721=>"110111110",
  58722=>"111001101",
  58723=>"100000101",
  58724=>"001100110",
  58725=>"001001001",
  58726=>"101011101",
  58727=>"000100011",
  58728=>"100111101",
  58729=>"100010000",
  58730=>"100000101",
  58731=>"000101000",
  58732=>"110100100",
  58733=>"001101011",
  58734=>"010010111",
  58735=>"001101111",
  58736=>"000111100",
  58737=>"100011111",
  58738=>"010110100",
  58739=>"000111000",
  58740=>"000011100",
  58741=>"010111011",
  58742=>"100010111",
  58743=>"000111000",
  58744=>"010000000",
  58745=>"001100111",
  58746=>"000011001",
  58747=>"001111111",
  58748=>"001101000",
  58749=>"101100011",
  58750=>"001110100",
  58751=>"010100001",
  58752=>"010000000",
  58753=>"011010011",
  58754=>"000010000",
  58755=>"000000111",
  58756=>"001010010",
  58757=>"011010111",
  58758=>"101010110",
  58759=>"000100011",
  58760=>"110100001",
  58761=>"101110101",
  58762=>"011000011",
  58763=>"101010000",
  58764=>"110110100",
  58765=>"100110110",
  58766=>"111101010",
  58767=>"101001000",
  58768=>"011111100",
  58769=>"101000111",
  58770=>"100011000",
  58771=>"100010001",
  58772=>"000110010",
  58773=>"010011101",
  58774=>"101100010",
  58775=>"011111000",
  58776=>"110000001",
  58777=>"000001011",
  58778=>"101100101",
  58779=>"000111111",
  58780=>"000001011",
  58781=>"101111011",
  58782=>"001100001",
  58783=>"011001000",
  58784=>"111000000",
  58785=>"101000001",
  58786=>"111111111",
  58787=>"000001000",
  58788=>"110101101",
  58789=>"010011101",
  58790=>"110101101",
  58791=>"010101000",
  58792=>"000100101",
  58793=>"100011110",
  58794=>"100010111",
  58795=>"011110010",
  58796=>"111000110",
  58797=>"011111011",
  58798=>"001110100",
  58799=>"110001110",
  58800=>"001000100",
  58801=>"000100111",
  58802=>"000100000",
  58803=>"100000100",
  58804=>"001011000",
  58805=>"101110000",
  58806=>"011111111",
  58807=>"110110111",
  58808=>"100101100",
  58809=>"000011000",
  58810=>"101011001",
  58811=>"100011110",
  58812=>"111011011",
  58813=>"110100010",
  58814=>"001111001",
  58815=>"100011110",
  58816=>"110011000",
  58817=>"100010101",
  58818=>"101110001",
  58819=>"011000011",
  58820=>"001100111",
  58821=>"011101001",
  58822=>"101101001",
  58823=>"111011000",
  58824=>"100001000",
  58825=>"010111101",
  58826=>"110110001",
  58827=>"010000111",
  58828=>"000111011",
  58829=>"111110100",
  58830=>"110111011",
  58831=>"101110111",
  58832=>"000100110",
  58833=>"111100001",
  58834=>"100101000",
  58835=>"001111001",
  58836=>"011110011",
  58837=>"001000100",
  58838=>"011101110",
  58839=>"101001100",
  58840=>"101010011",
  58841=>"001110011",
  58842=>"000111010",
  58843=>"110000110",
  58844=>"011100110",
  58845=>"000101011",
  58846=>"101010001",
  58847=>"011100111",
  58848=>"100001000",
  58849=>"010010110",
  58850=>"100100000",
  58851=>"110000010",
  58852=>"011000000",
  58853=>"010100001",
  58854=>"011000001",
  58855=>"101100010",
  58856=>"110111101",
  58857=>"111010011",
  58858=>"101001010",
  58859=>"001111010",
  58860=>"010110000",
  58861=>"101000110",
  58862=>"110000000",
  58863=>"001100101",
  58864=>"010000011",
  58865=>"000101111",
  58866=>"111110011",
  58867=>"110110110",
  58868=>"000101111",
  58869=>"000000110",
  58870=>"001000011",
  58871=>"001101000",
  58872=>"110101001",
  58873=>"101100000",
  58874=>"011100101",
  58875=>"000010110",
  58876=>"011001110",
  58877=>"010001000",
  58878=>"010100010",
  58879=>"101001101",
  58880=>"101111111",
  58881=>"111110100",
  58882=>"011001000",
  58883=>"101110001",
  58884=>"110011111",
  58885=>"010011000",
  58886=>"111001110",
  58887=>"000110001",
  58888=>"001100100",
  58889=>"100101001",
  58890=>"101101001",
  58891=>"000000100",
  58892=>"001001100",
  58893=>"100101000",
  58894=>"001001111",
  58895=>"011110000",
  58896=>"000011111",
  58897=>"100111010",
  58898=>"000111101",
  58899=>"110010100",
  58900=>"111000001",
  58901=>"010011011",
  58902=>"010100111",
  58903=>"010001000",
  58904=>"011100000",
  58905=>"011010001",
  58906=>"101001011",
  58907=>"011101001",
  58908=>"110101000",
  58909=>"101111101",
  58910=>"000010010",
  58911=>"100110100",
  58912=>"100111110",
  58913=>"010111011",
  58914=>"000100010",
  58915=>"111101001",
  58916=>"101010111",
  58917=>"001011101",
  58918=>"011111001",
  58919=>"101100000",
  58920=>"111001101",
  58921=>"010001100",
  58922=>"011100100",
  58923=>"000010001",
  58924=>"011101101",
  58925=>"100011100",
  58926=>"101001001",
  58927=>"001011100",
  58928=>"111000101",
  58929=>"100101001",
  58930=>"010101100",
  58931=>"001110100",
  58932=>"111100000",
  58933=>"001000000",
  58934=>"011010011",
  58935=>"100000101",
  58936=>"101011110",
  58937=>"000000111",
  58938=>"100111110",
  58939=>"010110010",
  58940=>"000011001",
  58941=>"111011001",
  58942=>"100000010",
  58943=>"101100100",
  58944=>"110001011",
  58945=>"100000101",
  58946=>"000001101",
  58947=>"011000010",
  58948=>"110110111",
  58949=>"011010001",
  58950=>"011111010",
  58951=>"001001110",
  58952=>"100000101",
  58953=>"011111101",
  58954=>"001111001",
  58955=>"010001110",
  58956=>"100101100",
  58957=>"011000011",
  58958=>"011011110",
  58959=>"111001010",
  58960=>"011101001",
  58961=>"111010111",
  58962=>"100101100",
  58963=>"010001011",
  58964=>"100100001",
  58965=>"000010110",
  58966=>"010100110",
  58967=>"110100011",
  58968=>"001010111",
  58969=>"100110000",
  58970=>"011001100",
  58971=>"000000001",
  58972=>"111000101",
  58973=>"000011000",
  58974=>"010010000",
  58975=>"111100010",
  58976=>"110011100",
  58977=>"111111111",
  58978=>"001001011",
  58979=>"001011101",
  58980=>"111000010",
  58981=>"111000010",
  58982=>"110010000",
  58983=>"000111100",
  58984=>"000010000",
  58985=>"001110100",
  58986=>"011000101",
  58987=>"011000101",
  58988=>"000100110",
  58989=>"010110101",
  58990=>"101101101",
  58991=>"100111101",
  58992=>"001000111",
  58993=>"001100100",
  58994=>"011011101",
  58995=>"000000001",
  58996=>"110011111",
  58997=>"000110111",
  58998=>"110011000",
  58999=>"000111100",
  59000=>"010000000",
  59001=>"010011111",
  59002=>"100111100",
  59003=>"000110010",
  59004=>"101000111",
  59005=>"111010001",
  59006=>"001100001",
  59007=>"101010111",
  59008=>"011010000",
  59009=>"001111111",
  59010=>"101110100",
  59011=>"011000000",
  59012=>"100000100",
  59013=>"111000001",
  59014=>"111011100",
  59015=>"000001000",
  59016=>"001001010",
  59017=>"011000001",
  59018=>"010011101",
  59019=>"110101001",
  59020=>"010010001",
  59021=>"000001111",
  59022=>"011001011",
  59023=>"110101111",
  59024=>"111100111",
  59025=>"101100110",
  59026=>"011011011",
  59027=>"011110100",
  59028=>"010101100",
  59029=>"101110111",
  59030=>"111110001",
  59031=>"001101000",
  59032=>"010111011",
  59033=>"101001110",
  59034=>"011001110",
  59035=>"000110001",
  59036=>"110001101",
  59037=>"000111011",
  59038=>"100011010",
  59039=>"111000111",
  59040=>"101001100",
  59041=>"001101001",
  59042=>"100001111",
  59043=>"010001010",
  59044=>"010011111",
  59045=>"111010011",
  59046=>"100101010",
  59047=>"101101100",
  59048=>"011100001",
  59049=>"000101101",
  59050=>"101101111",
  59051=>"110001111",
  59052=>"001110101",
  59053=>"101111001",
  59054=>"101111111",
  59055=>"111011010",
  59056=>"101011111",
  59057=>"110100110",
  59058=>"010001100",
  59059=>"110001000",
  59060=>"001111100",
  59061=>"010011000",
  59062=>"110010100",
  59063=>"000001001",
  59064=>"110110100",
  59065=>"100101011",
  59066=>"000101000",
  59067=>"010100001",
  59068=>"010010010",
  59069=>"011100000",
  59070=>"001000011",
  59071=>"001001000",
  59072=>"100001000",
  59073=>"000011011",
  59074=>"001011001",
  59075=>"010111110",
  59076=>"100101000",
  59077=>"000001111",
  59078=>"101101110",
  59079=>"011101100",
  59080=>"111011111",
  59081=>"011101101",
  59082=>"100010101",
  59083=>"100001011",
  59084=>"100101001",
  59085=>"110011111",
  59086=>"010011111",
  59087=>"010110111",
  59088=>"011001110",
  59089=>"010010011",
  59090=>"100100010",
  59091=>"111011000",
  59092=>"110000100",
  59093=>"100000100",
  59094=>"000011001",
  59095=>"001100101",
  59096=>"001111001",
  59097=>"110111100",
  59098=>"010000111",
  59099=>"111010010",
  59100=>"100101101",
  59101=>"000111100",
  59102=>"010111111",
  59103=>"110100011",
  59104=>"000100100",
  59105=>"110110000",
  59106=>"110001101",
  59107=>"000101101",
  59108=>"101000000",
  59109=>"000110101",
  59110=>"000000101",
  59111=>"111010110",
  59112=>"011001111",
  59113=>"100011011",
  59114=>"011101100",
  59115=>"100000110",
  59116=>"001010011",
  59117=>"011100110",
  59118=>"001001000",
  59119=>"001110001",
  59120=>"101111111",
  59121=>"100011101",
  59122=>"100010000",
  59123=>"010101100",
  59124=>"011100000",
  59125=>"100100100",
  59126=>"001111110",
  59127=>"000001000",
  59128=>"010011101",
  59129=>"010010000",
  59130=>"100111010",
  59131=>"100101010",
  59132=>"000100110",
  59133=>"010011000",
  59134=>"110100001",
  59135=>"110001111",
  59136=>"111101010",
  59137=>"111110001",
  59138=>"000100110",
  59139=>"100011010",
  59140=>"010111010",
  59141=>"110001100",
  59142=>"101001010",
  59143=>"010110001",
  59144=>"000100111",
  59145=>"110101001",
  59146=>"011111001",
  59147=>"011010001",
  59148=>"100011110",
  59149=>"001000100",
  59150=>"001010011",
  59151=>"100010001",
  59152=>"011111110",
  59153=>"011011000",
  59154=>"001011011",
  59155=>"101011000",
  59156=>"111000010",
  59157=>"110010100",
  59158=>"100010000",
  59159=>"010000000",
  59160=>"111011110",
  59161=>"111111101",
  59162=>"000001110",
  59163=>"100000110",
  59164=>"110001001",
  59165=>"001111011",
  59166=>"100001110",
  59167=>"011111100",
  59168=>"101001000",
  59169=>"101000100",
  59170=>"000110101",
  59171=>"010010111",
  59172=>"010001010",
  59173=>"000000011",
  59174=>"101001110",
  59175=>"100000111",
  59176=>"110110111",
  59177=>"001011001",
  59178=>"111101001",
  59179=>"010101101",
  59180=>"100111011",
  59181=>"000000000",
  59182=>"100000111",
  59183=>"011001100",
  59184=>"001100011",
  59185=>"000001111",
  59186=>"100010010",
  59187=>"100101101",
  59188=>"011010000",
  59189=>"001000011",
  59190=>"100111010",
  59191=>"011000000",
  59192=>"011110010",
  59193=>"000010110",
  59194=>"000101111",
  59195=>"010110011",
  59196=>"011101111",
  59197=>"011001011",
  59198=>"110101100",
  59199=>"100110101",
  59200=>"110011101",
  59201=>"011110101",
  59202=>"111110110",
  59203=>"101110011",
  59204=>"010110100",
  59205=>"001001010",
  59206=>"101101011",
  59207=>"011010011",
  59208=>"011100100",
  59209=>"000110011",
  59210=>"010100000",
  59211=>"110000000",
  59212=>"010111101",
  59213=>"110000100",
  59214=>"011100001",
  59215=>"000010010",
  59216=>"111110001",
  59217=>"011110110",
  59218=>"011101011",
  59219=>"010111011",
  59220=>"101010001",
  59221=>"000000111",
  59222=>"110000010",
  59223=>"100110001",
  59224=>"010100100",
  59225=>"010111010",
  59226=>"111111011",
  59227=>"000101011",
  59228=>"010110111",
  59229=>"110100101",
  59230=>"101111101",
  59231=>"000000100",
  59232=>"001100011",
  59233=>"111011110",
  59234=>"000011110",
  59235=>"101101100",
  59236=>"111011001",
  59237=>"001010110",
  59238=>"111101100",
  59239=>"111110000",
  59240=>"101000001",
  59241=>"001010110",
  59242=>"100000010",
  59243=>"110000000",
  59244=>"000101110",
  59245=>"110111101",
  59246=>"101100101",
  59247=>"011110110",
  59248=>"000110101",
  59249=>"010011001",
  59250=>"101110001",
  59251=>"101011000",
  59252=>"000000011",
  59253=>"000000010",
  59254=>"100111010",
  59255=>"101101010",
  59256=>"110110100",
  59257=>"000010100",
  59258=>"111000001",
  59259=>"011111110",
  59260=>"011100001",
  59261=>"110001111",
  59262=>"010111000",
  59263=>"010101101",
  59264=>"111001100",
  59265=>"001001010",
  59266=>"000000011",
  59267=>"111100011",
  59268=>"001010010",
  59269=>"111001101",
  59270=>"001000000",
  59271=>"101000111",
  59272=>"100000000",
  59273=>"100101010",
  59274=>"000110101",
  59275=>"111010100",
  59276=>"011110001",
  59277=>"001011001",
  59278=>"111111101",
  59279=>"111000011",
  59280=>"010110011",
  59281=>"110101001",
  59282=>"111000010",
  59283=>"111101110",
  59284=>"000101010",
  59285=>"010111000",
  59286=>"111111111",
  59287=>"111001111",
  59288=>"000000111",
  59289=>"010101100",
  59290=>"010110000",
  59291=>"010100011",
  59292=>"000010001",
  59293=>"011001110",
  59294=>"000000101",
  59295=>"000100000",
  59296=>"111010100",
  59297=>"110111101",
  59298=>"000100001",
  59299=>"000010101",
  59300=>"011101100",
  59301=>"111111110",
  59302=>"110101011",
  59303=>"101111110",
  59304=>"000111111",
  59305=>"011011010",
  59306=>"001110101",
  59307=>"111101111",
  59308=>"000110100",
  59309=>"101110010",
  59310=>"110111001",
  59311=>"010101011",
  59312=>"111100100",
  59313=>"110101001",
  59314=>"000000101",
  59315=>"100011110",
  59316=>"000100111",
  59317=>"001111010",
  59318=>"110001001",
  59319=>"000010000",
  59320=>"011001111",
  59321=>"101011111",
  59322=>"100011000",
  59323=>"100010110",
  59324=>"110000110",
  59325=>"011001110",
  59326=>"011000110",
  59327=>"001011000",
  59328=>"110001110",
  59329=>"001100111",
  59330=>"100111111",
  59331=>"101111111",
  59332=>"001111110",
  59333=>"101100111",
  59334=>"111000011",
  59335=>"101111111",
  59336=>"001000010",
  59337=>"100101001",
  59338=>"111010110",
  59339=>"001010000",
  59340=>"010101001",
  59341=>"010001001",
  59342=>"000010000",
  59343=>"010111100",
  59344=>"010000100",
  59345=>"001011110",
  59346=>"001000000",
  59347=>"110100000",
  59348=>"101011100",
  59349=>"110010001",
  59350=>"011101001",
  59351=>"010000100",
  59352=>"100010110",
  59353=>"000101101",
  59354=>"000101010",
  59355=>"111011101",
  59356=>"111101100",
  59357=>"110100101",
  59358=>"111000101",
  59359=>"111001000",
  59360=>"100000010",
  59361=>"110101001",
  59362=>"001010001",
  59363=>"010001111",
  59364=>"010010000",
  59365=>"111110001",
  59366=>"000001000",
  59367=>"111110110",
  59368=>"101000000",
  59369=>"000000000",
  59370=>"001001111",
  59371=>"000000111",
  59372=>"000010010",
  59373=>"100101100",
  59374=>"101000100",
  59375=>"111001001",
  59376=>"010101001",
  59377=>"010010110",
  59378=>"101100011",
  59379=>"000011000",
  59380=>"010100010",
  59381=>"011101000",
  59382=>"110000101",
  59383=>"010010110",
  59384=>"111000110",
  59385=>"101000010",
  59386=>"101010100",
  59387=>"011111011",
  59388=>"111000110",
  59389=>"011110001",
  59390=>"011101110",
  59391=>"000111110",
  59392=>"111111100",
  59393=>"100000000",
  59394=>"011011001",
  59395=>"001011011",
  59396=>"101001110",
  59397=>"100101111",
  59398=>"111011101",
  59399=>"100001100",
  59400=>"110011100",
  59401=>"100110100",
  59402=>"110010111",
  59403=>"111101000",
  59404=>"110100100",
  59405=>"000010101",
  59406=>"001110000",
  59407=>"011001100",
  59408=>"011111001",
  59409=>"001001011",
  59410=>"000111010",
  59411=>"000010100",
  59412=>"001010100",
  59413=>"100011100",
  59414=>"111011000",
  59415=>"111000000",
  59416=>"000111100",
  59417=>"010100101",
  59418=>"011101001",
  59419=>"000000110",
  59420=>"110100011",
  59421=>"001000011",
  59422=>"111100110",
  59423=>"110101011",
  59424=>"001001010",
  59425=>"011011000",
  59426=>"001100101",
  59427=>"111111101",
  59428=>"001010110",
  59429=>"010111111",
  59430=>"110001101",
  59431=>"011011110",
  59432=>"110101101",
  59433=>"000010010",
  59434=>"011110001",
  59435=>"110010001",
  59436=>"011000100",
  59437=>"111011101",
  59438=>"011110111",
  59439=>"000110110",
  59440=>"011011010",
  59441=>"100100001",
  59442=>"111111110",
  59443=>"010010000",
  59444=>"111100001",
  59445=>"010000100",
  59446=>"101001111",
  59447=>"001010011",
  59448=>"010001000",
  59449=>"010100011",
  59450=>"100010010",
  59451=>"101101111",
  59452=>"101011100",
  59453=>"100101010",
  59454=>"001011000",
  59455=>"001001000",
  59456=>"110111000",
  59457=>"000010000",
  59458=>"111101001",
  59459=>"100101110",
  59460=>"101100000",
  59461=>"111100000",
  59462=>"011101001",
  59463=>"111100000",
  59464=>"001010101",
  59465=>"011111011",
  59466=>"010101100",
  59467=>"110011000",
  59468=>"011000010",
  59469=>"101101101",
  59470=>"110110111",
  59471=>"010100110",
  59472=>"110110100",
  59473=>"010100011",
  59474=>"011001000",
  59475=>"001111100",
  59476=>"110011110",
  59477=>"111100000",
  59478=>"101011111",
  59479=>"000010100",
  59480=>"111111001",
  59481=>"100111010",
  59482=>"101111101",
  59483=>"101111110",
  59484=>"011010111",
  59485=>"111100100",
  59486=>"011011101",
  59487=>"100010111",
  59488=>"001101111",
  59489=>"110111000",
  59490=>"101010111",
  59491=>"101001001",
  59492=>"001010000",
  59493=>"000110100",
  59494=>"111010101",
  59495=>"100110001",
  59496=>"100001100",
  59497=>"110001111",
  59498=>"001100110",
  59499=>"010110111",
  59500=>"000100100",
  59501=>"100001011",
  59502=>"110110001",
  59503=>"000001011",
  59504=>"000100110",
  59505=>"010101011",
  59506=>"000001101",
  59507=>"000011000",
  59508=>"101010001",
  59509=>"000110011",
  59510=>"100111011",
  59511=>"010000001",
  59512=>"001000000",
  59513=>"001100011",
  59514=>"110001110",
  59515=>"100011000",
  59516=>"001100000",
  59517=>"000000110",
  59518=>"111110010",
  59519=>"110000100",
  59520=>"000011000",
  59521=>"011001010",
  59522=>"011011010",
  59523=>"110111001",
  59524=>"011010111",
  59525=>"010110100",
  59526=>"010001101",
  59527=>"110111111",
  59528=>"010101011",
  59529=>"100111101",
  59530=>"110101101",
  59531=>"111010001",
  59532=>"011101001",
  59533=>"101101111",
  59534=>"110101000",
  59535=>"000111011",
  59536=>"110000010",
  59537=>"111110101",
  59538=>"001010011",
  59539=>"101100100",
  59540=>"110101100",
  59541=>"111001000",
  59542=>"101101010",
  59543=>"001100100",
  59544=>"100010100",
  59545=>"101111110",
  59546=>"011000011",
  59547=>"011010101",
  59548=>"110110000",
  59549=>"010101011",
  59550=>"101010011",
  59551=>"001011000",
  59552=>"001111100",
  59553=>"101000001",
  59554=>"000000001",
  59555=>"000110110",
  59556=>"011001010",
  59557=>"000001101",
  59558=>"010011011",
  59559=>"100000111",
  59560=>"100111000",
  59561=>"111110100",
  59562=>"111011100",
  59563=>"110010010",
  59564=>"111110100",
  59565=>"000010101",
  59566=>"111111111",
  59567=>"000011001",
  59568=>"000101001",
  59569=>"000000010",
  59570=>"011110111",
  59571=>"111001111",
  59572=>"100011001",
  59573=>"101111111",
  59574=>"110001011",
  59575=>"101111001",
  59576=>"001110100",
  59577=>"000010010",
  59578=>"001110100",
  59579=>"111011110",
  59580=>"111001101",
  59581=>"111111111",
  59582=>"001111110",
  59583=>"010101011",
  59584=>"000100011",
  59585=>"110001010",
  59586=>"100011110",
  59587=>"001011000",
  59588=>"011010011",
  59589=>"010111011",
  59590=>"100001101",
  59591=>"111100011",
  59592=>"101011000",
  59593=>"001100001",
  59594=>"111111111",
  59595=>"011010111",
  59596=>"001010000",
  59597=>"000110100",
  59598=>"101111101",
  59599=>"110001010",
  59600=>"101111000",
  59601=>"111101100",
  59602=>"010110011",
  59603=>"000111100",
  59604=>"101000100",
  59605=>"011100101",
  59606=>"101011100",
  59607=>"001110111",
  59608=>"011101100",
  59609=>"000001100",
  59610=>"100000100",
  59611=>"010111100",
  59612=>"011011011",
  59613=>"011110010",
  59614=>"110001111",
  59615=>"000011110",
  59616=>"100000011",
  59617=>"000011011",
  59618=>"001000111",
  59619=>"000110000",
  59620=>"000110010",
  59621=>"000011111",
  59622=>"100011100",
  59623=>"101000100",
  59624=>"010000101",
  59625=>"011011110",
  59626=>"001110001",
  59627=>"010111000",
  59628=>"110100000",
  59629=>"001010000",
  59630=>"010001000",
  59631=>"000000110",
  59632=>"000000010",
  59633=>"000010111",
  59634=>"011110000",
  59635=>"010100101",
  59636=>"000011100",
  59637=>"001101001",
  59638=>"000100000",
  59639=>"101000110",
  59640=>"000111100",
  59641=>"010101101",
  59642=>"110100000",
  59643=>"100001101",
  59644=>"110101010",
  59645=>"111110100",
  59646=>"101001100",
  59647=>"010110100",
  59648=>"110101100",
  59649=>"110011101",
  59650=>"111000101",
  59651=>"011000001",
  59652=>"001011011",
  59653=>"010001110",
  59654=>"100111101",
  59655=>"010100101",
  59656=>"101001000",
  59657=>"010111100",
  59658=>"111010011",
  59659=>"001000000",
  59660=>"001111000",
  59661=>"011101001",
  59662=>"110000000",
  59663=>"000100100",
  59664=>"000110000",
  59665=>"001101001",
  59666=>"000101000",
  59667=>"110100111",
  59668=>"101011001",
  59669=>"000001010",
  59670=>"010101100",
  59671=>"000000000",
  59672=>"110110100",
  59673=>"111101010",
  59674=>"001011101",
  59675=>"011010101",
  59676=>"110111011",
  59677=>"001101111",
  59678=>"001001011",
  59679=>"011011001",
  59680=>"111101001",
  59681=>"011111101",
  59682=>"000000011",
  59683=>"000101110",
  59684=>"000001111",
  59685=>"001010101",
  59686=>"101101101",
  59687=>"010001111",
  59688=>"100100100",
  59689=>"100110001",
  59690=>"011101011",
  59691=>"110001111",
  59692=>"010010000",
  59693=>"010010101",
  59694=>"000001000",
  59695=>"010111110",
  59696=>"000000111",
  59697=>"010111011",
  59698=>"000101101",
  59699=>"000100011",
  59700=>"001110100",
  59701=>"110000111",
  59702=>"001011010",
  59703=>"110111010",
  59704=>"111100111",
  59705=>"000001100",
  59706=>"100001001",
  59707=>"110100001",
  59708=>"100001010",
  59709=>"110011010",
  59710=>"000101010",
  59711=>"100011110",
  59712=>"111110000",
  59713=>"110000000",
  59714=>"000100110",
  59715=>"001101000",
  59716=>"011010111",
  59717=>"111000111",
  59718=>"101000111",
  59719=>"101000111",
  59720=>"110011000",
  59721=>"111010010",
  59722=>"001001100",
  59723=>"011011101",
  59724=>"101101110",
  59725=>"011001101",
  59726=>"101100010",
  59727=>"000101001",
  59728=>"010000000",
  59729=>"101010110",
  59730=>"000100000",
  59731=>"110110100",
  59732=>"001000000",
  59733=>"001110000",
  59734=>"011101010",
  59735=>"011100000",
  59736=>"110111111",
  59737=>"100001100",
  59738=>"000011100",
  59739=>"100010110",
  59740=>"011110111",
  59741=>"111100101",
  59742=>"100100000",
  59743=>"010100111",
  59744=>"110011100",
  59745=>"101100010",
  59746=>"001110101",
  59747=>"110000101",
  59748=>"100100010",
  59749=>"111101111",
  59750=>"011111001",
  59751=>"010000001",
  59752=>"100001111",
  59753=>"101011000",
  59754=>"111110110",
  59755=>"000101001",
  59756=>"101000000",
  59757=>"100001010",
  59758=>"000011000",
  59759=>"010001001",
  59760=>"100100101",
  59761=>"110001101",
  59762=>"010100011",
  59763=>"111101101",
  59764=>"000111001",
  59765=>"010101011",
  59766=>"010110011",
  59767=>"001011011",
  59768=>"111100101",
  59769=>"001001111",
  59770=>"100101011",
  59771=>"010110100",
  59772=>"000000111",
  59773=>"001001010",
  59774=>"000100101",
  59775=>"110000101",
  59776=>"110101001",
  59777=>"011111101",
  59778=>"010111111",
  59779=>"000101010",
  59780=>"100110011",
  59781=>"011011000",
  59782=>"000010000",
  59783=>"010010110",
  59784=>"101100111",
  59785=>"110101100",
  59786=>"011110111",
  59787=>"000001001",
  59788=>"110100111",
  59789=>"010111101",
  59790=>"100100010",
  59791=>"111000010",
  59792=>"010101111",
  59793=>"100100110",
  59794=>"000101010",
  59795=>"011000000",
  59796=>"010010010",
  59797=>"110011101",
  59798=>"000010000",
  59799=>"101111110",
  59800=>"001101101",
  59801=>"011000100",
  59802=>"111101110",
  59803=>"010010010",
  59804=>"101101001",
  59805=>"101001001",
  59806=>"111010000",
  59807=>"011001010",
  59808=>"101001010",
  59809=>"111111110",
  59810=>"001000101",
  59811=>"101001001",
  59812=>"110111110",
  59813=>"110111000",
  59814=>"110111001",
  59815=>"101000100",
  59816=>"110100011",
  59817=>"000001111",
  59818=>"010100000",
  59819=>"111010110",
  59820=>"010010000",
  59821=>"010011001",
  59822=>"000101010",
  59823=>"011000010",
  59824=>"100000011",
  59825=>"100110100",
  59826=>"011011100",
  59827=>"011000111",
  59828=>"000110111",
  59829=>"000001011",
  59830=>"000010001",
  59831=>"000101011",
  59832=>"110001011",
  59833=>"010101010",
  59834=>"111101101",
  59835=>"101001001",
  59836=>"111100011",
  59837=>"101011100",
  59838=>"101111101",
  59839=>"010010000",
  59840=>"101001011",
  59841=>"011100110",
  59842=>"100111110",
  59843=>"111110111",
  59844=>"100000010",
  59845=>"011000111",
  59846=>"011000010",
  59847=>"111000101",
  59848=>"100111100",
  59849=>"010101110",
  59850=>"010011011",
  59851=>"100001101",
  59852=>"101100000",
  59853=>"111101111",
  59854=>"100011011",
  59855=>"000110010",
  59856=>"011101101",
  59857=>"100001100",
  59858=>"010000010",
  59859=>"111000101",
  59860=>"000011101",
  59861=>"111101101",
  59862=>"011001111",
  59863=>"000110110",
  59864=>"110000000",
  59865=>"100101100",
  59866=>"001000001",
  59867=>"101111011",
  59868=>"011011011",
  59869=>"000111100",
  59870=>"010101011",
  59871=>"100000010",
  59872=>"000011100",
  59873=>"111000100",
  59874=>"110110000",
  59875=>"000110101",
  59876=>"100001110",
  59877=>"111001001",
  59878=>"111000010",
  59879=>"010100001",
  59880=>"001001000",
  59881=>"111000010",
  59882=>"000011111",
  59883=>"110110101",
  59884=>"000111000",
  59885=>"101101110",
  59886=>"110011111",
  59887=>"001101001",
  59888=>"001111100",
  59889=>"111001010",
  59890=>"000100100",
  59891=>"000000001",
  59892=>"101011100",
  59893=>"111011011",
  59894=>"101110100",
  59895=>"000100100",
  59896=>"100110010",
  59897=>"111000001",
  59898=>"111011010",
  59899=>"111101110",
  59900=>"001010101",
  59901=>"111111110",
  59902=>"100101111",
  59903=>"111111001",
  59904=>"110010011",
  59905=>"101011000",
  59906=>"100110001",
  59907=>"100111111",
  59908=>"100110111",
  59909=>"110010011",
  59910=>"001001011",
  59911=>"011011111",
  59912=>"101100001",
  59913=>"111011001",
  59914=>"011100001",
  59915=>"110010000",
  59916=>"011000110",
  59917=>"111110000",
  59918=>"110000010",
  59919=>"011011011",
  59920=>"110101000",
  59921=>"001110001",
  59922=>"111111100",
  59923=>"010100001",
  59924=>"111000111",
  59925=>"000111100",
  59926=>"001000111",
  59927=>"111000011",
  59928=>"000010010",
  59929=>"101001111",
  59930=>"100001000",
  59931=>"101000011",
  59932=>"110101001",
  59933=>"111011001",
  59934=>"100111000",
  59935=>"111011011",
  59936=>"110010100",
  59937=>"100101011",
  59938=>"001010010",
  59939=>"101110000",
  59940=>"101110110",
  59941=>"110011000",
  59942=>"010010001",
  59943=>"111100110",
  59944=>"111001011",
  59945=>"011001000",
  59946=>"111000000",
  59947=>"011000011",
  59948=>"111010001",
  59949=>"110001111",
  59950=>"110100011",
  59951=>"100110000",
  59952=>"110000100",
  59953=>"001111100",
  59954=>"010010110",
  59955=>"110010101",
  59956=>"010110111",
  59957=>"000111111",
  59958=>"000000100",
  59959=>"111000000",
  59960=>"111000011",
  59961=>"010010110",
  59962=>"110100010",
  59963=>"100110100",
  59964=>"000010011",
  59965=>"111000001",
  59966=>"101001111",
  59967=>"100000111",
  59968=>"111100100",
  59969=>"001010100",
  59970=>"110010100",
  59971=>"111110011",
  59972=>"100001010",
  59973=>"001101000",
  59974=>"010100000",
  59975=>"111100011",
  59976=>"111100010",
  59977=>"100010001",
  59978=>"111110011",
  59979=>"110011101",
  59980=>"011000111",
  59981=>"110100010",
  59982=>"101111000",
  59983=>"001100111",
  59984=>"100101010",
  59985=>"100111110",
  59986=>"010011111",
  59987=>"000100100",
  59988=>"110000000",
  59989=>"111011100",
  59990=>"010001111",
  59991=>"100001000",
  59992=>"111010101",
  59993=>"010101100",
  59994=>"001011010",
  59995=>"000100110",
  59996=>"100110110",
  59997=>"000110110",
  59998=>"110101010",
  59999=>"100000101",
  60000=>"010011101",
  60001=>"001010100",
  60002=>"010111011",
  60003=>"001111001",
  60004=>"011100110",
  60005=>"101111100",
  60006=>"000000001",
  60007=>"000011010",
  60008=>"001000000",
  60009=>"110110011",
  60010=>"011011010",
  60011=>"000000000",
  60012=>"000001100",
  60013=>"001101111",
  60014=>"011111100",
  60015=>"000111001",
  60016=>"011010010",
  60017=>"000011001",
  60018=>"100011010",
  60019=>"001000010",
  60020=>"000101110",
  60021=>"100100000",
  60022=>"111011101",
  60023=>"000111111",
  60024=>"011101101",
  60025=>"001001011",
  60026=>"111010101",
  60027=>"001100100",
  60028=>"001000001",
  60029=>"111010000",
  60030=>"111110111",
  60031=>"100110001",
  60032=>"111111101",
  60033=>"111100110",
  60034=>"100100100",
  60035=>"101000101",
  60036=>"100001001",
  60037=>"010111100",
  60038=>"000101110",
  60039=>"111111110",
  60040=>"000110011",
  60041=>"110010110",
  60042=>"000000111",
  60043=>"101111000",
  60044=>"010011010",
  60045=>"000111101",
  60046=>"101011111",
  60047=>"100111010",
  60048=>"000011000",
  60049=>"111101011",
  60050=>"110101100",
  60051=>"101110011",
  60052=>"110010101",
  60053=>"000100000",
  60054=>"110101100",
  60055=>"101001001",
  60056=>"100001100",
  60057=>"110001100",
  60058=>"010011000",
  60059=>"101101100",
  60060=>"000001110",
  60061=>"100100010",
  60062=>"110011100",
  60063=>"001100101",
  60064=>"110100001",
  60065=>"100111001",
  60066=>"110000111",
  60067=>"011101000",
  60068=>"110000000",
  60069=>"100100101",
  60070=>"001101101",
  60071=>"100111101",
  60072=>"001000110",
  60073=>"010111011",
  60074=>"101110100",
  60075=>"000001011",
  60076=>"011110001",
  60077=>"110000000",
  60078=>"111001010",
  60079=>"101110000",
  60080=>"000100011",
  60081=>"101101010",
  60082=>"011010100",
  60083=>"001010110",
  60084=>"110001000",
  60085=>"011011010",
  60086=>"111011100",
  60087=>"011111000",
  60088=>"000010110",
  60089=>"001111011",
  60090=>"101110011",
  60091=>"011010001",
  60092=>"101110101",
  60093=>"000000100",
  60094=>"011001001",
  60095=>"111011000",
  60096=>"111010101",
  60097=>"011101110",
  60098=>"000110101",
  60099=>"100011110",
  60100=>"111101111",
  60101=>"100101100",
  60102=>"011110011",
  60103=>"111110100",
  60104=>"010000001",
  60105=>"111000000",
  60106=>"000101011",
  60107=>"001010011",
  60108=>"001111000",
  60109=>"000000010",
  60110=>"011110010",
  60111=>"010100100",
  60112=>"110010001",
  60113=>"100110101",
  60114=>"010010110",
  60115=>"011011110",
  60116=>"010111010",
  60117=>"011010100",
  60118=>"101000110",
  60119=>"000110110",
  60120=>"110001000",
  60121=>"111101101",
  60122=>"001010100",
  60123=>"011011010",
  60124=>"111000101",
  60125=>"011010111",
  60126=>"011011010",
  60127=>"000000001",
  60128=>"011100000",
  60129=>"010011100",
  60130=>"100000010",
  60131=>"011000111",
  60132=>"101111111",
  60133=>"001100111",
  60134=>"110001100",
  60135=>"001110101",
  60136=>"000001110",
  60137=>"001100101",
  60138=>"111111110",
  60139=>"101111010",
  60140=>"000000001",
  60141=>"101001001",
  60142=>"110011000",
  60143=>"100011010",
  60144=>"101101110",
  60145=>"010010101",
  60146=>"011101111",
  60147=>"011100010",
  60148=>"011011110",
  60149=>"100011101",
  60150=>"010001110",
  60151=>"100001011",
  60152=>"111101000",
  60153=>"000010101",
  60154=>"000110001",
  60155=>"101110011",
  60156=>"110000110",
  60157=>"000111011",
  60158=>"101100010",
  60159=>"111011000",
  60160=>"101010101",
  60161=>"000101110",
  60162=>"111111110",
  60163=>"011011010",
  60164=>"001100000",
  60165=>"011011000",
  60166=>"100001110",
  60167=>"110010111",
  60168=>"000100001",
  60169=>"000101100",
  60170=>"101001001",
  60171=>"000000010",
  60172=>"001010111",
  60173=>"001010010",
  60174=>"110101000",
  60175=>"011100100",
  60176=>"101001100",
  60177=>"000001100",
  60178=>"101110100",
  60179=>"011001010",
  60180=>"011110101",
  60181=>"111001100",
  60182=>"111100101",
  60183=>"010100001",
  60184=>"111011010",
  60185=>"000001111",
  60186=>"001111010",
  60187=>"110010101",
  60188=>"101000110",
  60189=>"000101101",
  60190=>"110100101",
  60191=>"000100101",
  60192=>"010011110",
  60193=>"011000011",
  60194=>"110111111",
  60195=>"000100010",
  60196=>"110111100",
  60197=>"011111111",
  60198=>"010011111",
  60199=>"010010111",
  60200=>"000001001",
  60201=>"000111011",
  60202=>"010110000",
  60203=>"011000111",
  60204=>"001001001",
  60205=>"000000011",
  60206=>"011101000",
  60207=>"011100100",
  60208=>"100010110",
  60209=>"110111100",
  60210=>"000110010",
  60211=>"010111011",
  60212=>"110000001",
  60213=>"010001111",
  60214=>"100110101",
  60215=>"001000001",
  60216=>"100011111",
  60217=>"110001010",
  60218=>"010001000",
  60219=>"110101111",
  60220=>"111000100",
  60221=>"110000011",
  60222=>"101101010",
  60223=>"011101111",
  60224=>"110001110",
  60225=>"111010010",
  60226=>"010001000",
  60227=>"111000101",
  60228=>"110111100",
  60229=>"101101101",
  60230=>"111101011",
  60231=>"100010111",
  60232=>"001100111",
  60233=>"010001000",
  60234=>"100001101",
  60235=>"110100010",
  60236=>"110100011",
  60237=>"011011100",
  60238=>"100011000",
  60239=>"111000001",
  60240=>"110111011",
  60241=>"100010011",
  60242=>"001001000",
  60243=>"110011000",
  60244=>"010010010",
  60245=>"010111111",
  60246=>"001100010",
  60247=>"000010111",
  60248=>"010110111",
  60249=>"011100111",
  60250=>"001101001",
  60251=>"010101011",
  60252=>"001010010",
  60253=>"000100001",
  60254=>"001100100",
  60255=>"100100001",
  60256=>"010010101",
  60257=>"111110011",
  60258=>"000001010",
  60259=>"011000010",
  60260=>"011010100",
  60261=>"000011011",
  60262=>"011111010",
  60263=>"101111110",
  60264=>"110110000",
  60265=>"010011100",
  60266=>"111111010",
  60267=>"000011000",
  60268=>"111110110",
  60269=>"000100100",
  60270=>"001101001",
  60271=>"110001100",
  60272=>"010010100",
  60273=>"010000001",
  60274=>"000101110",
  60275=>"100010001",
  60276=>"100010010",
  60277=>"111100100",
  60278=>"101111011",
  60279=>"011101110",
  60280=>"100010011",
  60281=>"001101000",
  60282=>"010100010",
  60283=>"001000011",
  60284=>"000000000",
  60285=>"001100000",
  60286=>"010110101",
  60287=>"111101010",
  60288=>"010101000",
  60289=>"101010001",
  60290=>"100101011",
  60291=>"110000011",
  60292=>"001001100",
  60293=>"110110100",
  60294=>"010000100",
  60295=>"000101101",
  60296=>"100000011",
  60297=>"010101010",
  60298=>"111111111",
  60299=>"000000101",
  60300=>"110100101",
  60301=>"001100010",
  60302=>"001100111",
  60303=>"001100001",
  60304=>"111111000",
  60305=>"010010000",
  60306=>"101110100",
  60307=>"111000001",
  60308=>"110011100",
  60309=>"101110111",
  60310=>"010101011",
  60311=>"110111101",
  60312=>"011100100",
  60313=>"100001011",
  60314=>"111100110",
  60315=>"000000010",
  60316=>"111101100",
  60317=>"011001001",
  60318=>"111100010",
  60319=>"010000100",
  60320=>"100001110",
  60321=>"100111010",
  60322=>"011101000",
  60323=>"100000101",
  60324=>"001011100",
  60325=>"010100101",
  60326=>"100110101",
  60327=>"011110101",
  60328=>"110001010",
  60329=>"010101011",
  60330=>"011010010",
  60331=>"010000000",
  60332=>"000011111",
  60333=>"011101000",
  60334=>"110111010",
  60335=>"000101111",
  60336=>"011011000",
  60337=>"111010100",
  60338=>"000111000",
  60339=>"011011101",
  60340=>"110101100",
  60341=>"010001100",
  60342=>"000000010",
  60343=>"100001001",
  60344=>"010111001",
  60345=>"111011110",
  60346=>"011010010",
  60347=>"000000011",
  60348=>"010111110",
  60349=>"000000001",
  60350=>"111101011",
  60351=>"011001011",
  60352=>"101000111",
  60353=>"001011001",
  60354=>"000000110",
  60355=>"110000011",
  60356=>"000110000",
  60357=>"000001100",
  60358=>"101011000",
  60359=>"011110011",
  60360=>"100100011",
  60361=>"100000100",
  60362=>"000110010",
  60363=>"101010111",
  60364=>"011011010",
  60365=>"100101111",
  60366=>"001111011",
  60367=>"100010111",
  60368=>"100111011",
  60369=>"001111100",
  60370=>"000101010",
  60371=>"001100111",
  60372=>"101101000",
  60373=>"010010000",
  60374=>"011010000",
  60375=>"000010111",
  60376=>"001100010",
  60377=>"000010011",
  60378=>"001101111",
  60379=>"101001001",
  60380=>"101100010",
  60381=>"010110001",
  60382=>"110111000",
  60383=>"110111101",
  60384=>"110000010",
  60385=>"100100010",
  60386=>"111000101",
  60387=>"010001100",
  60388=>"010111101",
  60389=>"010110011",
  60390=>"001000111",
  60391=>"100101010",
  60392=>"011110000",
  60393=>"101110111",
  60394=>"000111000",
  60395=>"110001000",
  60396=>"010101101",
  60397=>"111000110",
  60398=>"001111101",
  60399=>"000000101",
  60400=>"011010010",
  60401=>"000110110",
  60402=>"001110001",
  60403=>"101000111",
  60404=>"011100010",
  60405=>"101000100",
  60406=>"101011100",
  60407=>"011001101",
  60408=>"000010001",
  60409=>"101010101",
  60410=>"101101110",
  60411=>"000110110",
  60412=>"100100000",
  60413=>"001011010",
  60414=>"001010011",
  60415=>"111011110",
  60416=>"000011011",
  60417=>"111000101",
  60418=>"010100011",
  60419=>"001001110",
  60420=>"110110100",
  60421=>"001100011",
  60422=>"000100011",
  60423=>"111000100",
  60424=>"100000101",
  60425=>"001101000",
  60426=>"010011110",
  60427=>"000101100",
  60428=>"000010011",
  60429=>"010100101",
  60430=>"100101011",
  60431=>"000001111",
  60432=>"000101111",
  60433=>"111101101",
  60434=>"011000111",
  60435=>"100010001",
  60436=>"000101000",
  60437=>"110111011",
  60438=>"110100011",
  60439=>"110011110",
  60440=>"100100011",
  60441=>"111101011",
  60442=>"010000010",
  60443=>"010010010",
  60444=>"010011101",
  60445=>"010110001",
  60446=>"000010010",
  60447=>"101011110",
  60448=>"111110110",
  60449=>"110011100",
  60450=>"101011110",
  60451=>"001111100",
  60452=>"111010100",
  60453=>"111011011",
  60454=>"111001001",
  60455=>"111111000",
  60456=>"111111010",
  60457=>"100001100",
  60458=>"100111111",
  60459=>"001001100",
  60460=>"001011101",
  60461=>"000010110",
  60462=>"000010011",
  60463=>"101110001",
  60464=>"010100110",
  60465=>"101011101",
  60466=>"101011001",
  60467=>"011000011",
  60468=>"000001100",
  60469=>"100110000",
  60470=>"101111011",
  60471=>"111111101",
  60472=>"010010101",
  60473=>"000100011",
  60474=>"101110001",
  60475=>"111111111",
  60476=>"101110111",
  60477=>"011001011",
  60478=>"110110100",
  60479=>"011010101",
  60480=>"010111110",
  60481=>"000100001",
  60482=>"111001000",
  60483=>"001000010",
  60484=>"010001000",
  60485=>"010011101",
  60486=>"000100111",
  60487=>"111101001",
  60488=>"110100101",
  60489=>"100100101",
  60490=>"000001100",
  60491=>"000000100",
  60492=>"110111101",
  60493=>"000110101",
  60494=>"110100011",
  60495=>"001111010",
  60496=>"101110100",
  60497=>"000010010",
  60498=>"000110100",
  60499=>"011110111",
  60500=>"100100000",
  60501=>"011110001",
  60502=>"100011101",
  60503=>"001011010",
  60504=>"100100110",
  60505=>"111101100",
  60506=>"101011111",
  60507=>"001001000",
  60508=>"000011001",
  60509=>"010100111",
  60510=>"110111000",
  60511=>"011011000",
  60512=>"111111111",
  60513=>"000010101",
  60514=>"001000010",
  60515=>"100000011",
  60516=>"110011100",
  60517=>"110000000",
  60518=>"101100000",
  60519=>"001001000",
  60520=>"001001100",
  60521=>"110111011",
  60522=>"010100101",
  60523=>"001101011",
  60524=>"010000011",
  60525=>"111101101",
  60526=>"000010101",
  60527=>"011001000",
  60528=>"011111100",
  60529=>"110001101",
  60530=>"110101111",
  60531=>"010001000",
  60532=>"001111110",
  60533=>"100010011",
  60534=>"000101110",
  60535=>"100001010",
  60536=>"001000011",
  60537=>"101011010",
  60538=>"000000100",
  60539=>"110001010",
  60540=>"011001110",
  60541=>"110100011",
  60542=>"010111010",
  60543=>"111110101",
  60544=>"011101000",
  60545=>"001110011",
  60546=>"111111101",
  60547=>"111001011",
  60548=>"000011011",
  60549=>"011100111",
  60550=>"000000111",
  60551=>"011001101",
  60552=>"000011110",
  60553=>"101100001",
  60554=>"111010000",
  60555=>"111100101",
  60556=>"100111101",
  60557=>"011001100",
  60558=>"011001011",
  60559=>"010110010",
  60560=>"011101100",
  60561=>"001000111",
  60562=>"100000100",
  60563=>"011011011",
  60564=>"011001001",
  60565=>"101011100",
  60566=>"111110010",
  60567=>"111111111",
  60568=>"000000100",
  60569=>"010100000",
  60570=>"111100001",
  60571=>"011110010",
  60572=>"011000101",
  60573=>"000010100",
  60574=>"001100000",
  60575=>"101111011",
  60576=>"001100100",
  60577=>"101001000",
  60578=>"010001000",
  60579=>"001001101",
  60580=>"000000010",
  60581=>"010010100",
  60582=>"010101000",
  60583=>"001000010",
  60584=>"111010000",
  60585=>"110111111",
  60586=>"100000110",
  60587=>"010000000",
  60588=>"110011011",
  60589=>"010010011",
  60590=>"010110100",
  60591=>"111001010",
  60592=>"011101011",
  60593=>"010000100",
  60594=>"100101100",
  60595=>"001001100",
  60596=>"001111011",
  60597=>"000110011",
  60598=>"000011110",
  60599=>"110100101",
  60600=>"010101011",
  60601=>"001101001",
  60602=>"000000111",
  60603=>"000101001",
  60604=>"011111110",
  60605=>"000011001",
  60606=>"111001010",
  60607=>"000101101",
  60608=>"111101001",
  60609=>"011111011",
  60610=>"001001101",
  60611=>"111111110",
  60612=>"100000101",
  60613=>"101011011",
  60614=>"101011100",
  60615=>"100110011",
  60616=>"111000011",
  60617=>"111011000",
  60618=>"100000000",
  60619=>"011101111",
  60620=>"010100010",
  60621=>"110110011",
  60622=>"100111110",
  60623=>"101000101",
  60624=>"001000011",
  60625=>"101110111",
  60626=>"000001000",
  60627=>"001010101",
  60628=>"010111101",
  60629=>"011000110",
  60630=>"101010100",
  60631=>"100010001",
  60632=>"101011001",
  60633=>"011110010",
  60634=>"100101000",
  60635=>"011011111",
  60636=>"001001010",
  60637=>"001010100",
  60638=>"110000100",
  60639=>"101011110",
  60640=>"011000010",
  60641=>"011001100",
  60642=>"100111010",
  60643=>"011111001",
  60644=>"111100111",
  60645=>"000001110",
  60646=>"010011001",
  60647=>"100110010",
  60648=>"111110110",
  60649=>"010110100",
  60650=>"100001011",
  60651=>"000011000",
  60652=>"000100010",
  60653=>"110101001",
  60654=>"100001111",
  60655=>"100010011",
  60656=>"110010101",
  60657=>"000000011",
  60658=>"111011010",
  60659=>"101001100",
  60660=>"101101110",
  60661=>"010110111",
  60662=>"001111111",
  60663=>"000100000",
  60664=>"000000001",
  60665=>"100111110",
  60666=>"111101110",
  60667=>"001100011",
  60668=>"010000111",
  60669=>"111001001",
  60670=>"101111100",
  60671=>"000001011",
  60672=>"011000111",
  60673=>"101111100",
  60674=>"010100111",
  60675=>"111110001",
  60676=>"010010100",
  60677=>"111101111",
  60678=>"111000110",
  60679=>"010100001",
  60680=>"010101000",
  60681=>"010000110",
  60682=>"100110100",
  60683=>"010100101",
  60684=>"110001100",
  60685=>"001000011",
  60686=>"010111010",
  60687=>"100100110",
  60688=>"100111110",
  60689=>"101011000",
  60690=>"001000010",
  60691=>"101101001",
  60692=>"010010001",
  60693=>"111010110",
  60694=>"100011111",
  60695=>"111111100",
  60696=>"111000011",
  60697=>"101111110",
  60698=>"110010000",
  60699=>"100011000",
  60700=>"000110010",
  60701=>"100110001",
  60702=>"000001110",
  60703=>"010111110",
  60704=>"010000110",
  60705=>"101110110",
  60706=>"010101111",
  60707=>"110110100",
  60708=>"000100110",
  60709=>"100011001",
  60710=>"101010110",
  60711=>"111001101",
  60712=>"010011010",
  60713=>"111111000",
  60714=>"100111000",
  60715=>"000110011",
  60716=>"010110011",
  60717=>"001010001",
  60718=>"110111111",
  60719=>"110000111",
  60720=>"001011011",
  60721=>"001010001",
  60722=>"010110100",
  60723=>"110100011",
  60724=>"000101010",
  60725=>"101100110",
  60726=>"000001010",
  60727=>"111011000",
  60728=>"110010100",
  60729=>"010011001",
  60730=>"001000001",
  60731=>"110001010",
  60732=>"001101011",
  60733=>"111110000",
  60734=>"100101100",
  60735=>"111011010",
  60736=>"111010000",
  60737=>"111011000",
  60738=>"100001111",
  60739=>"111100001",
  60740=>"010100001",
  60741=>"000000111",
  60742=>"101100101",
  60743=>"000011001",
  60744=>"001001000",
  60745=>"001111101",
  60746=>"001111110",
  60747=>"001111011",
  60748=>"000110001",
  60749=>"000000101",
  60750=>"011100011",
  60751=>"101001001",
  60752=>"100100101",
  60753=>"001010110",
  60754=>"110101010",
  60755=>"100001001",
  60756=>"110000100",
  60757=>"100110001",
  60758=>"111000000",
  60759=>"110000000",
  60760=>"001110011",
  60761=>"100001100",
  60762=>"100000000",
  60763=>"110011001",
  60764=>"110101111",
  60765=>"000001001",
  60766=>"010111111",
  60767=>"101011101",
  60768=>"001000100",
  60769=>"001111110",
  60770=>"100010011",
  60771=>"110111001",
  60772=>"011110001",
  60773=>"101001001",
  60774=>"110111101",
  60775=>"010000011",
  60776=>"000101111",
  60777=>"110001010",
  60778=>"011101001",
  60779=>"000010001",
  60780=>"101111101",
  60781=>"011101111",
  60782=>"000111011",
  60783=>"111011010",
  60784=>"110111111",
  60785=>"011001000",
  60786=>"101001111",
  60787=>"011000000",
  60788=>"010000000",
  60789=>"100011101",
  60790=>"010011000",
  60791=>"000110000",
  60792=>"000010110",
  60793=>"010000000",
  60794=>"100111011",
  60795=>"001011101",
  60796=>"101000000",
  60797=>"111001001",
  60798=>"011111010",
  60799=>"000100001",
  60800=>"111110011",
  60801=>"001100000",
  60802=>"110111111",
  60803=>"110101001",
  60804=>"000111000",
  60805=>"100100100",
  60806=>"011110101",
  60807=>"101100011",
  60808=>"100011110",
  60809=>"110111110",
  60810=>"011110111",
  60811=>"110110010",
  60812=>"100001001",
  60813=>"111111110",
  60814=>"101000010",
  60815=>"101000110",
  60816=>"000100110",
  60817=>"001101011",
  60818=>"000000010",
  60819=>"010100001",
  60820=>"010000010",
  60821=>"110111011",
  60822=>"110001011",
  60823=>"110001001",
  60824=>"010101010",
  60825=>"010001010",
  60826=>"001011011",
  60827=>"010111011",
  60828=>"001010000",
  60829=>"010100011",
  60830=>"010111111",
  60831=>"101000011",
  60832=>"000011000",
  60833=>"110000110",
  60834=>"101101111",
  60835=>"101010101",
  60836=>"100010000",
  60837=>"001000010",
  60838=>"011100110",
  60839=>"101111000",
  60840=>"010100010",
  60841=>"110101111",
  60842=>"001011001",
  60843=>"001100110",
  60844=>"001001001",
  60845=>"110000110",
  60846=>"011011111",
  60847=>"001101001",
  60848=>"010110010",
  60849=>"011100000",
  60850=>"001000100",
  60851=>"011011010",
  60852=>"101111011",
  60853=>"101100111",
  60854=>"001001001",
  60855=>"111101110",
  60856=>"011101100",
  60857=>"111011100",
  60858=>"001001001",
  60859=>"010010110",
  60860=>"110110010",
  60861=>"001110101",
  60862=>"011010101",
  60863=>"100010111",
  60864=>"000111001",
  60865=>"011000110",
  60866=>"111101010",
  60867=>"101100111",
  60868=>"011001000",
  60869=>"001110111",
  60870=>"001111111",
  60871=>"100100111",
  60872=>"001101101",
  60873=>"001111111",
  60874=>"000101011",
  60875=>"010100110",
  60876=>"001000001",
  60877=>"010001010",
  60878=>"010101111",
  60879=>"000110000",
  60880=>"000010110",
  60881=>"010010010",
  60882=>"110111100",
  60883=>"001010111",
  60884=>"110110000",
  60885=>"001001110",
  60886=>"001110001",
  60887=>"101010011",
  60888=>"101100110",
  60889=>"110001111",
  60890=>"100110100",
  60891=>"111001000",
  60892=>"100001001",
  60893=>"001000000",
  60894=>"110111101",
  60895=>"100101100",
  60896=>"100110110",
  60897=>"111000010",
  60898=>"000110011",
  60899=>"010010101",
  60900=>"101000101",
  60901=>"110111101",
  60902=>"010010101",
  60903=>"110110111",
  60904=>"011100111",
  60905=>"010011100",
  60906=>"110010000",
  60907=>"100001010",
  60908=>"010111111",
  60909=>"111011101",
  60910=>"010010001",
  60911=>"000110001",
  60912=>"001110110",
  60913=>"100110110",
  60914=>"001101010",
  60915=>"011110010",
  60916=>"111111100",
  60917=>"111010000",
  60918=>"100110101",
  60919=>"111100101",
  60920=>"011111110",
  60921=>"001110011",
  60922=>"010011010",
  60923=>"111100111",
  60924=>"000111010",
  60925=>"101010011",
  60926=>"010011101",
  60927=>"100110100",
  60928=>"110000111",
  60929=>"010010101",
  60930=>"011010100",
  60931=>"001010011",
  60932=>"110000100",
  60933=>"110111000",
  60934=>"101111111",
  60935=>"101010100",
  60936=>"110110001",
  60937=>"000101001",
  60938=>"110011101",
  60939=>"010000110",
  60940=>"110011010",
  60941=>"001010110",
  60942=>"010101000",
  60943=>"001001001",
  60944=>"110000101",
  60945=>"011001111",
  60946=>"000100110",
  60947=>"011110000",
  60948=>"111101011",
  60949=>"101101010",
  60950=>"000100001",
  60951=>"101011110",
  60952=>"011011000",
  60953=>"001000011",
  60954=>"110011011",
  60955=>"000111111",
  60956=>"001001010",
  60957=>"101011000",
  60958=>"000110100",
  60959=>"111100110",
  60960=>"101010101",
  60961=>"101000100",
  60962=>"110100101",
  60963=>"000011010",
  60964=>"011110101",
  60965=>"111110011",
  60966=>"111110001",
  60967=>"001111010",
  60968=>"001111010",
  60969=>"101100110",
  60970=>"100110001",
  60971=>"100010110",
  60972=>"100100111",
  60973=>"000011000",
  60974=>"100101001",
  60975=>"011111011",
  60976=>"111011101",
  60977=>"010000100",
  60978=>"101011011",
  60979=>"011000001",
  60980=>"100001111",
  60981=>"111010111",
  60982=>"100010110",
  60983=>"101110100",
  60984=>"000011101",
  60985=>"111110111",
  60986=>"011111111",
  60987=>"111001101",
  60988=>"011101110",
  60989=>"110011111",
  60990=>"100010000",
  60991=>"000111100",
  60992=>"010110110",
  60993=>"111011001",
  60994=>"001100101",
  60995=>"010100010",
  60996=>"011010110",
  60997=>"100001010",
  60998=>"000000111",
  60999=>"010110011",
  61000=>"011011110",
  61001=>"010011101",
  61002=>"111100010",
  61003=>"000111110",
  61004=>"001101110",
  61005=>"000000011",
  61006=>"111001100",
  61007=>"100101111",
  61008=>"011001010",
  61009=>"110001110",
  61010=>"110011101",
  61011=>"000011110",
  61012=>"101101001",
  61013=>"101100101",
  61014=>"000001000",
  61015=>"001111110",
  61016=>"010011110",
  61017=>"011001111",
  61018=>"010100010",
  61019=>"000000110",
  61020=>"110010101",
  61021=>"000000001",
  61022=>"110011100",
  61023=>"001100100",
  61024=>"001101010",
  61025=>"011010000",
  61026=>"000001011",
  61027=>"110010111",
  61028=>"110101001",
  61029=>"111101010",
  61030=>"110111010",
  61031=>"010101101",
  61032=>"110101100",
  61033=>"100100101",
  61034=>"101110010",
  61035=>"111100110",
  61036=>"110011011",
  61037=>"001010111",
  61038=>"110011110",
  61039=>"100001100",
  61040=>"010011011",
  61041=>"000100001",
  61042=>"001000100",
  61043=>"011100101",
  61044=>"001110001",
  61045=>"000010110",
  61046=>"100110101",
  61047=>"101000001",
  61048=>"100011110",
  61049=>"001110011",
  61050=>"100010000",
  61051=>"111000000",
  61052=>"010000010",
  61053=>"000011001",
  61054=>"001100001",
  61055=>"110011010",
  61056=>"100100110",
  61057=>"011100100",
  61058=>"011000000",
  61059=>"010000101",
  61060=>"101011111",
  61061=>"101101000",
  61062=>"111111000",
  61063=>"011010001",
  61064=>"111100100",
  61065=>"011100100",
  61066=>"100110110",
  61067=>"101110111",
  61068=>"101111011",
  61069=>"000011110",
  61070=>"011001010",
  61071=>"100111001",
  61072=>"010001011",
  61073=>"111111001",
  61074=>"010110011",
  61075=>"000101111",
  61076=>"011001101",
  61077=>"100000000",
  61078=>"101001100",
  61079=>"101101000",
  61080=>"011111010",
  61081=>"111000011",
  61082=>"010010001",
  61083=>"111101110",
  61084=>"101001111",
  61085=>"001100011",
  61086=>"110000000",
  61087=>"100100101",
  61088=>"100000001",
  61089=>"001010101",
  61090=>"100011011",
  61091=>"111001011",
  61092=>"011010111",
  61093=>"010000001",
  61094=>"100000001",
  61095=>"110100111",
  61096=>"111100100",
  61097=>"001100010",
  61098=>"111010011",
  61099=>"111010100",
  61100=>"100001100",
  61101=>"001111101",
  61102=>"011110011",
  61103=>"100101000",
  61104=>"001000001",
  61105=>"110011100",
  61106=>"010101011",
  61107=>"100000011",
  61108=>"001010111",
  61109=>"110011011",
  61110=>"111010101",
  61111=>"100011000",
  61112=>"010001001",
  61113=>"000100111",
  61114=>"000100010",
  61115=>"110011110",
  61116=>"000000100",
  61117=>"001001011",
  61118=>"011010100",
  61119=>"110000111",
  61120=>"011111010",
  61121=>"011101010",
  61122=>"101001001",
  61123=>"101100101",
  61124=>"101110001",
  61125=>"111001101",
  61126=>"000011111",
  61127=>"101110011",
  61128=>"011010001",
  61129=>"010000000",
  61130=>"111101100",
  61131=>"100100001",
  61132=>"111011110",
  61133=>"100000001",
  61134=>"110000011",
  61135=>"001010011",
  61136=>"111010101",
  61137=>"101100101",
  61138=>"000111011",
  61139=>"011011011",
  61140=>"001100010",
  61141=>"000101110",
  61142=>"000100111",
  61143=>"001000000",
  61144=>"001000100",
  61145=>"110100011",
  61146=>"011111100",
  61147=>"100110101",
  61148=>"110010010",
  61149=>"110000000",
  61150=>"011101101",
  61151=>"110011110",
  61152=>"000110111",
  61153=>"001110000",
  61154=>"110110111",
  61155=>"000110000",
  61156=>"010001000",
  61157=>"110100000",
  61158=>"100010111",
  61159=>"110110010",
  61160=>"101010000",
  61161=>"101011100",
  61162=>"111101100",
  61163=>"111011110",
  61164=>"000110010",
  61165=>"000001010",
  61166=>"111111110",
  61167=>"010111000",
  61168=>"011110100",
  61169=>"000101000",
  61170=>"110000100",
  61171=>"001010111",
  61172=>"100010001",
  61173=>"010110100",
  61174=>"110110111",
  61175=>"111110110",
  61176=>"001101011",
  61177=>"001001100",
  61178=>"000100111",
  61179=>"001000010",
  61180=>"101100100",
  61181=>"011110110",
  61182=>"011010111",
  61183=>"000001010",
  61184=>"000101011",
  61185=>"010111010",
  61186=>"111011011",
  61187=>"100111001",
  61188=>"011101011",
  61189=>"001101010",
  61190=>"110110101",
  61191=>"000011011",
  61192=>"110110001",
  61193=>"111010001",
  61194=>"100111101",
  61195=>"000001101",
  61196=>"100100001",
  61197=>"110111010",
  61198=>"011100101",
  61199=>"111111011",
  61200=>"000000010",
  61201=>"001001011",
  61202=>"011111010",
  61203=>"110100100",
  61204=>"010110111",
  61205=>"000101101",
  61206=>"011111011",
  61207=>"011111010",
  61208=>"001101001",
  61209=>"011111100",
  61210=>"001110110",
  61211=>"011101110",
  61212=>"101001101",
  61213=>"010111011",
  61214=>"011000010",
  61215=>"000000101",
  61216=>"001011000",
  61217=>"110011101",
  61218=>"000001110",
  61219=>"011110010",
  61220=>"001010101",
  61221=>"110010101",
  61222=>"101000110",
  61223=>"000011101",
  61224=>"101110100",
  61225=>"001011001",
  61226=>"000101101",
  61227=>"011111001",
  61228=>"101111101",
  61229=>"001111111",
  61230=>"000000111",
  61231=>"100001001",
  61232=>"110011010",
  61233=>"000011011",
  61234=>"110001010",
  61235=>"110111101",
  61236=>"011111001",
  61237=>"010100011",
  61238=>"011011111",
  61239=>"101000100",
  61240=>"111110010",
  61241=>"001000110",
  61242=>"011110000",
  61243=>"011110100",
  61244=>"101011110",
  61245=>"000011000",
  61246=>"001101010",
  61247=>"110101001",
  61248=>"000100110",
  61249=>"010010111",
  61250=>"011000100",
  61251=>"100001010",
  61252=>"111101011",
  61253=>"100100000",
  61254=>"001000000",
  61255=>"101000101",
  61256=>"100000011",
  61257=>"000101011",
  61258=>"101000101",
  61259=>"101011110",
  61260=>"011101010",
  61261=>"100010010",
  61262=>"100110000",
  61263=>"001000010",
  61264=>"110010010",
  61265=>"000000100",
  61266=>"011101010",
  61267=>"110011010",
  61268=>"110000011",
  61269=>"110000010",
  61270=>"010011010",
  61271=>"000100000",
  61272=>"110100110",
  61273=>"011101100",
  61274=>"010100000",
  61275=>"000101000",
  61276=>"101111111",
  61277=>"100110001",
  61278=>"011111011",
  61279=>"001010001",
  61280=>"010100001",
  61281=>"111011110",
  61282=>"111100111",
  61283=>"111011110",
  61284=>"100111001",
  61285=>"101001101",
  61286=>"100101011",
  61287=>"000001101",
  61288=>"100000100",
  61289=>"000100110",
  61290=>"101110001",
  61291=>"101110101",
  61292=>"000000101",
  61293=>"001000011",
  61294=>"011011000",
  61295=>"001001110",
  61296=>"111111011",
  61297=>"111000111",
  61298=>"011000110",
  61299=>"111010011",
  61300=>"111100001",
  61301=>"001010000",
  61302=>"001001101",
  61303=>"101101000",
  61304=>"100001111",
  61305=>"110110010",
  61306=>"011100101",
  61307=>"101111001",
  61308=>"010011011",
  61309=>"000101100",
  61310=>"100000010",
  61311=>"010010110",
  61312=>"000110101",
  61313=>"100110000",
  61314=>"101011101",
  61315=>"011001011",
  61316=>"110100111",
  61317=>"000111010",
  61318=>"011010110",
  61319=>"000001001",
  61320=>"011101101",
  61321=>"111011101",
  61322=>"010100110",
  61323=>"001011101",
  61324=>"110001111",
  61325=>"101010101",
  61326=>"111000101",
  61327=>"100110101",
  61328=>"010111000",
  61329=>"110110101",
  61330=>"101011000",
  61331=>"011001010",
  61332=>"011010101",
  61333=>"000110001",
  61334=>"011011111",
  61335=>"001110111",
  61336=>"010110100",
  61337=>"111001001",
  61338=>"110101010",
  61339=>"000101001",
  61340=>"010101001",
  61341=>"100101100",
  61342=>"101010111",
  61343=>"110010001",
  61344=>"011001111",
  61345=>"001001011",
  61346=>"000111101",
  61347=>"011110010",
  61348=>"100111011",
  61349=>"010111100",
  61350=>"000101101",
  61351=>"110011000",
  61352=>"101111001",
  61353=>"110011100",
  61354=>"111110010",
  61355=>"110101111",
  61356=>"111011111",
  61357=>"000110011",
  61358=>"100100100",
  61359=>"010000011",
  61360=>"111100100",
  61361=>"000100010",
  61362=>"011111010",
  61363=>"000011100",
  61364=>"000101100",
  61365=>"100111111",
  61366=>"111000101",
  61367=>"001000110",
  61368=>"000101011",
  61369=>"010110000",
  61370=>"110010100",
  61371=>"111011111",
  61372=>"111011111",
  61373=>"010100011",
  61374=>"001101100",
  61375=>"000000000",
  61376=>"101011000",
  61377=>"101010011",
  61378=>"100000111",
  61379=>"111110010",
  61380=>"011000011",
  61381=>"101001101",
  61382=>"001111110",
  61383=>"111001100",
  61384=>"111000000",
  61385=>"100101100",
  61386=>"000100000",
  61387=>"000011001",
  61388=>"000000100",
  61389=>"010001100",
  61390=>"001101101",
  61391=>"101010011",
  61392=>"001101001",
  61393=>"101111010",
  61394=>"010101100",
  61395=>"111000000",
  61396=>"101010011",
  61397=>"001001111",
  61398=>"000001010",
  61399=>"010100011",
  61400=>"001001001",
  61401=>"011101011",
  61402=>"101101000",
  61403=>"000010100",
  61404=>"000010010",
  61405=>"111001000",
  61406=>"100011011",
  61407=>"011000000",
  61408=>"101101001",
  61409=>"011011110",
  61410=>"110010010",
  61411=>"001011011",
  61412=>"000001010",
  61413=>"111000111",
  61414=>"101000010",
  61415=>"111001010",
  61416=>"010011001",
  61417=>"011010000",
  61418=>"001000001",
  61419=>"011111100",
  61420=>"000010101",
  61421=>"101011001",
  61422=>"111101011",
  61423=>"001100001",
  61424=>"000001000",
  61425=>"111001111",
  61426=>"111001011",
  61427=>"010001011",
  61428=>"110001001",
  61429=>"101110000",
  61430=>"100111010",
  61431=>"111111001",
  61432=>"100100010",
  61433=>"101101100",
  61434=>"101101011",
  61435=>"111011010",
  61436=>"011110000",
  61437=>"110100111",
  61438=>"110000110",
  61439=>"111111100",
  61440=>"000010110",
  61441=>"011001111",
  61442=>"011000101",
  61443=>"001001111",
  61444=>"111100101",
  61445=>"000001100",
  61446=>"011110000",
  61447=>"000110110",
  61448=>"011111000",
  61449=>"001101011",
  61450=>"011001111",
  61451=>"110011111",
  61452=>"010110100",
  61453=>"001101001",
  61454=>"011110010",
  61455=>"111111111",
  61456=>"110100111",
  61457=>"101001001",
  61458=>"101100011",
  61459=>"101101101",
  61460=>"000110011",
  61461=>"000110101",
  61462=>"100001011",
  61463=>"110110011",
  61464=>"111001111",
  61465=>"111000110",
  61466=>"010000001",
  61467=>"000110100",
  61468=>"011010010",
  61469=>"010011111",
  61470=>"001100101",
  61471=>"000011000",
  61472=>"000100111",
  61473=>"111111010",
  61474=>"010111110",
  61475=>"111001110",
  61476=>"110101100",
  61477=>"000001000",
  61478=>"100010100",
  61479=>"110010000",
  61480=>"011100101",
  61481=>"001100010",
  61482=>"010101101",
  61483=>"111001111",
  61484=>"000111100",
  61485=>"100110100",
  61486=>"101101111",
  61487=>"010011010",
  61488=>"001100110",
  61489=>"111011000",
  61490=>"001110110",
  61491=>"011001011",
  61492=>"101101111",
  61493=>"000000001",
  61494=>"111110001",
  61495=>"100100100",
  61496=>"011011100",
  61497=>"010101010",
  61498=>"111011010",
  61499=>"010101111",
  61500=>"100101101",
  61501=>"110100000",
  61502=>"011010110",
  61503=>"001010001",
  61504=>"101110011",
  61505=>"001001011",
  61506=>"110010110",
  61507=>"000011000",
  61508=>"000110100",
  61509=>"010000011",
  61510=>"111111010",
  61511=>"101000100",
  61512=>"111000001",
  61513=>"111000100",
  61514=>"000101101",
  61515=>"010011010",
  61516=>"111000011",
  61517=>"000111000",
  61518=>"101101110",
  61519=>"100110001",
  61520=>"000101001",
  61521=>"010111001",
  61522=>"111101000",
  61523=>"000111000",
  61524=>"011100101",
  61525=>"011001101",
  61526=>"001110011",
  61527=>"111010111",
  61528=>"010111110",
  61529=>"000111101",
  61530=>"010110110",
  61531=>"001110100",
  61532=>"010111010",
  61533=>"011111100",
  61534=>"101111100",
  61535=>"110010000",
  61536=>"100001101",
  61537=>"010110111",
  61538=>"001101010",
  61539=>"000100110",
  61540=>"100010000",
  61541=>"101001011",
  61542=>"110001100",
  61543=>"100011110",
  61544=>"000010001",
  61545=>"110110011",
  61546=>"000000011",
  61547=>"011100110",
  61548=>"111010101",
  61549=>"000111111",
  61550=>"001000011",
  61551=>"001001100",
  61552=>"100110100",
  61553=>"101001101",
  61554=>"101011011",
  61555=>"000100011",
  61556=>"010100111",
  61557=>"011011010",
  61558=>"110011101",
  61559=>"000111000",
  61560=>"001111011",
  61561=>"000000111",
  61562=>"101100001",
  61563=>"001101000",
  61564=>"000101010",
  61565=>"011100100",
  61566=>"111011010",
  61567=>"110001110",
  61568=>"010000111",
  61569=>"111101000",
  61570=>"101000010",
  61571=>"110110100",
  61572=>"010001011",
  61573=>"000100001",
  61574=>"111111110",
  61575=>"100110010",
  61576=>"000110110",
  61577=>"111011011",
  61578=>"000001101",
  61579=>"101001000",
  61580=>"011101010",
  61581=>"110000110",
  61582=>"110001000",
  61583=>"010110101",
  61584=>"000010100",
  61585=>"011100001",
  61586=>"111110001",
  61587=>"011110001",
  61588=>"011101110",
  61589=>"010111110",
  61590=>"110111110",
  61591=>"111011001",
  61592=>"101000000",
  61593=>"011010000",
  61594=>"010100011",
  61595=>"100100001",
  61596=>"101110011",
  61597=>"000100011",
  61598=>"101101101",
  61599=>"001100100",
  61600=>"000000001",
  61601=>"111000110",
  61602=>"010111111",
  61603=>"001000001",
  61604=>"011000000",
  61605=>"010010110",
  61606=>"100011010",
  61607=>"111000000",
  61608=>"110101111",
  61609=>"111000011",
  61610=>"100101010",
  61611=>"101101101",
  61612=>"110110001",
  61613=>"111001100",
  61614=>"010110000",
  61615=>"100101111",
  61616=>"101010101",
  61617=>"000100110",
  61618=>"000111101",
  61619=>"100001111",
  61620=>"011100011",
  61621=>"110010110",
  61622=>"001010110",
  61623=>"111000111",
  61624=>"001100000",
  61625=>"011100101",
  61626=>"101011001",
  61627=>"111111011",
  61628=>"110001000",
  61629=>"010011001",
  61630=>"011011100",
  61631=>"100001111",
  61632=>"011011101",
  61633=>"110010010",
  61634=>"110001001",
  61635=>"110001001",
  61636=>"010101111",
  61637=>"101110001",
  61638=>"101101110",
  61639=>"011111010",
  61640=>"111000001",
  61641=>"011110110",
  61642=>"101111111",
  61643=>"010010001",
  61644=>"000001001",
  61645=>"111100100",
  61646=>"100001110",
  61647=>"101111100",
  61648=>"011100111",
  61649=>"000000011",
  61650=>"000101000",
  61651=>"011010010",
  61652=>"111010110",
  61653=>"101100100",
  61654=>"101011101",
  61655=>"100110101",
  61656=>"001001010",
  61657=>"110101100",
  61658=>"000110010",
  61659=>"010011101",
  61660=>"110000001",
  61661=>"001011011",
  61662=>"010100010",
  61663=>"110100000",
  61664=>"000100101",
  61665=>"110100001",
  61666=>"110001100",
  61667=>"111011000",
  61668=>"101010100",
  61669=>"011111100",
  61670=>"110110000",
  61671=>"011001111",
  61672=>"111010100",
  61673=>"100111101",
  61674=>"011000100",
  61675=>"010000010",
  61676=>"111101110",
  61677=>"111010100",
  61678=>"010111110",
  61679=>"110001111",
  61680=>"100011100",
  61681=>"010000001",
  61682=>"010010100",
  61683=>"000111011",
  61684=>"101001111",
  61685=>"010010100",
  61686=>"110101100",
  61687=>"000100101",
  61688=>"010100000",
  61689=>"011011100",
  61690=>"000000000",
  61691=>"001101011",
  61692=>"010101111",
  61693=>"001111111",
  61694=>"011101010",
  61695=>"110000000",
  61696=>"111100010",
  61697=>"010100010",
  61698=>"000010010",
  61699=>"111111101",
  61700=>"000110000",
  61701=>"110111110",
  61702=>"001111011",
  61703=>"010001100",
  61704=>"011010011",
  61705=>"111110101",
  61706=>"110001100",
  61707=>"000001111",
  61708=>"111110110",
  61709=>"011000010",
  61710=>"011101001",
  61711=>"010110101",
  61712=>"111001111",
  61713=>"101010100",
  61714=>"000100100",
  61715=>"111111100",
  61716=>"001001001",
  61717=>"010000111",
  61718=>"011000011",
  61719=>"101011111",
  61720=>"110000110",
  61721=>"110011100",
  61722=>"001000000",
  61723=>"001001001",
  61724=>"110001001",
  61725=>"101110010",
  61726=>"001010010",
  61727=>"000101101",
  61728=>"110000000",
  61729=>"111000001",
  61730=>"001110001",
  61731=>"100000011",
  61732=>"101110010",
  61733=>"111101111",
  61734=>"010100101",
  61735=>"000001110",
  61736=>"001011101",
  61737=>"101100010",
  61738=>"000010100",
  61739=>"011111101",
  61740=>"000010100",
  61741=>"110001111",
  61742=>"101101101",
  61743=>"111000110",
  61744=>"100000001",
  61745=>"101110011",
  61746=>"101010000",
  61747=>"110100001",
  61748=>"110000110",
  61749=>"011110100",
  61750=>"110001010",
  61751=>"001111110",
  61752=>"011011000",
  61753=>"001000111",
  61754=>"001001110",
  61755=>"010111010",
  61756=>"010101001",
  61757=>"010100100",
  61758=>"110001011",
  61759=>"101100101",
  61760=>"010010010",
  61761=>"111100101",
  61762=>"101000111",
  61763=>"011001000",
  61764=>"110101001",
  61765=>"110111011",
  61766=>"111000011",
  61767=>"001000001",
  61768=>"010000001",
  61769=>"100000001",
  61770=>"001101100",
  61771=>"010011111",
  61772=>"101000110",
  61773=>"011000100",
  61774=>"001010101",
  61775=>"111001000",
  61776=>"101011010",
  61777=>"011101000",
  61778=>"100111011",
  61779=>"010110011",
  61780=>"011011111",
  61781=>"011001011",
  61782=>"011101100",
  61783=>"011110111",
  61784=>"000010001",
  61785=>"010110011",
  61786=>"000001100",
  61787=>"100110111",
  61788=>"110011101",
  61789=>"010110101",
  61790=>"100111010",
  61791=>"001001111",
  61792=>"100001111",
  61793=>"001001001",
  61794=>"101010100",
  61795=>"100001001",
  61796=>"001001001",
  61797=>"111100101",
  61798=>"101101001",
  61799=>"010000000",
  61800=>"101100001",
  61801=>"010011011",
  61802=>"111101101",
  61803=>"000110100",
  61804=>"100000011",
  61805=>"000101111",
  61806=>"010000010",
  61807=>"000100010",
  61808=>"000100101",
  61809=>"110100110",
  61810=>"000011000",
  61811=>"111110110",
  61812=>"001101011",
  61813=>"011011110",
  61814=>"001000111",
  61815=>"010001111",
  61816=>"011010100",
  61817=>"000110011",
  61818=>"111000111",
  61819=>"000010000",
  61820=>"000111100",
  61821=>"011110000",
  61822=>"010101001",
  61823=>"001011110",
  61824=>"001100100",
  61825=>"000110010",
  61826=>"101101011",
  61827=>"010110010",
  61828=>"110111001",
  61829=>"011101110",
  61830=>"001110100",
  61831=>"010010100",
  61832=>"111001110",
  61833=>"010110010",
  61834=>"100010011",
  61835=>"100110010",
  61836=>"011101111",
  61837=>"100100001",
  61838=>"000011111",
  61839=>"110010000",
  61840=>"110010010",
  61841=>"001011001",
  61842=>"110100100",
  61843=>"100000000",
  61844=>"101110011",
  61845=>"000011111",
  61846=>"010011011",
  61847=>"001100100",
  61848=>"111110101",
  61849=>"010010010",
  61850=>"101101000",
  61851=>"100111100",
  61852=>"111100001",
  61853=>"000001010",
  61854=>"001101101",
  61855=>"110010100",
  61856=>"000000001",
  61857=>"001010110",
  61858=>"111000010",
  61859=>"110111111",
  61860=>"110001000",
  61861=>"100011100",
  61862=>"110100100",
  61863=>"000011000",
  61864=>"010000100",
  61865=>"111111000",
  61866=>"000011010",
  61867=>"000001101",
  61868=>"110101101",
  61869=>"010000011",
  61870=>"101110011",
  61871=>"000010010",
  61872=>"001100111",
  61873=>"000010111",
  61874=>"111000100",
  61875=>"011111111",
  61876=>"001101111",
  61877=>"000101001",
  61878=>"001000001",
  61879=>"110111110",
  61880=>"011010010",
  61881=>"110001111",
  61882=>"011101000",
  61883=>"010101101",
  61884=>"110011110",
  61885=>"010011010",
  61886=>"100000000",
  61887=>"010110010",
  61888=>"001100111",
  61889=>"000101000",
  61890=>"101100001",
  61891=>"000111011",
  61892=>"110011110",
  61893=>"111001100",
  61894=>"111111010",
  61895=>"100111011",
  61896=>"111110010",
  61897=>"011011101",
  61898=>"111011001",
  61899=>"000100101",
  61900=>"111000100",
  61901=>"000010111",
  61902=>"011000110",
  61903=>"100100100",
  61904=>"011001110",
  61905=>"111001001",
  61906=>"001011101",
  61907=>"000001100",
  61908=>"011111110",
  61909=>"000001011",
  61910=>"001001010",
  61911=>"010110000",
  61912=>"010010101",
  61913=>"000101011",
  61914=>"111101011",
  61915=>"100100001",
  61916=>"011101010",
  61917=>"000010100",
  61918=>"111101101",
  61919=>"100110100",
  61920=>"100011001",
  61921=>"010011000",
  61922=>"100100001",
  61923=>"000111000",
  61924=>"100010000",
  61925=>"000001000",
  61926=>"111011110",
  61927=>"010011101",
  61928=>"010011100",
  61929=>"111100010",
  61930=>"001101010",
  61931=>"010110101",
  61932=>"011100000",
  61933=>"101100011",
  61934=>"100000101",
  61935=>"110100100",
  61936=>"001010000",
  61937=>"110000011",
  61938=>"111011101",
  61939=>"011010001",
  61940=>"010101110",
  61941=>"010101010",
  61942=>"000110100",
  61943=>"001001010",
  61944=>"011000101",
  61945=>"111111111",
  61946=>"111011110",
  61947=>"001101010",
  61948=>"010101101",
  61949=>"010000111",
  61950=>"111101010",
  61951=>"000000100",
  61952=>"111001101",
  61953=>"101110110",
  61954=>"111010111",
  61955=>"001111011",
  61956=>"110110110",
  61957=>"000000000",
  61958=>"101110111",
  61959=>"000110111",
  61960=>"101111101",
  61961=>"111110110",
  61962=>"101001001",
  61963=>"001000101",
  61964=>"000110111",
  61965=>"000010101",
  61966=>"000011010",
  61967=>"010011110",
  61968=>"101001111",
  61969=>"111111011",
  61970=>"100001011",
  61971=>"000011000",
  61972=>"100111000",
  61973=>"100000011",
  61974=>"000101000",
  61975=>"000101001",
  61976=>"001110111",
  61977=>"000000100",
  61978=>"011000110",
  61979=>"111111100",
  61980=>"110010101",
  61981=>"010011000",
  61982=>"010100000",
  61983=>"110000010",
  61984=>"110111101",
  61985=>"011011001",
  61986=>"001101010",
  61987=>"010101111",
  61988=>"111010101",
  61989=>"011000010",
  61990=>"101100010",
  61991=>"101111001",
  61992=>"011000100",
  61993=>"110010011",
  61994=>"010111011",
  61995=>"101111010",
  61996=>"010110100",
  61997=>"000100001",
  61998=>"110111000",
  61999=>"100111001",
  62000=>"110110001",
  62001=>"100001100",
  62002=>"011010001",
  62003=>"011011011",
  62004=>"010111111",
  62005=>"101000111",
  62006=>"001101110",
  62007=>"111011011",
  62008=>"110000011",
  62009=>"111011010",
  62010=>"101011011",
  62011=>"011110111",
  62012=>"000011100",
  62013=>"000100001",
  62014=>"110100001",
  62015=>"111111111",
  62016=>"101011001",
  62017=>"010101000",
  62018=>"110001011",
  62019=>"100011111",
  62020=>"110101100",
  62021=>"101100011",
  62022=>"000101011",
  62023=>"111111101",
  62024=>"111010000",
  62025=>"000000001",
  62026=>"011100011",
  62027=>"111011010",
  62028=>"011000010",
  62029=>"010111000",
  62030=>"110010100",
  62031=>"100110110",
  62032=>"111001001",
  62033=>"100010001",
  62034=>"011110011",
  62035=>"001110111",
  62036=>"111010100",
  62037=>"110100111",
  62038=>"100101001",
  62039=>"101100111",
  62040=>"110011001",
  62041=>"011011100",
  62042=>"101011111",
  62043=>"000011010",
  62044=>"000010000",
  62045=>"011001111",
  62046=>"110001000",
  62047=>"111111011",
  62048=>"100000111",
  62049=>"111001000",
  62050=>"110000111",
  62051=>"000101000",
  62052=>"101111100",
  62053=>"111000100",
  62054=>"100111001",
  62055=>"111101111",
  62056=>"000100011",
  62057=>"010110101",
  62058=>"111001101",
  62059=>"100111100",
  62060=>"000011100",
  62061=>"001100110",
  62062=>"000101000",
  62063=>"111101010",
  62064=>"111011010",
  62065=>"011000101",
  62066=>"111101000",
  62067=>"001010000",
  62068=>"000000010",
  62069=>"110101100",
  62070=>"000000010",
  62071=>"100001100",
  62072=>"110100001",
  62073=>"010001011",
  62074=>"111111110",
  62075=>"011000101",
  62076=>"110011010",
  62077=>"111111100",
  62078=>"011010001",
  62079=>"101010101",
  62080=>"101100010",
  62081=>"011110000",
  62082=>"100010110",
  62083=>"001101010",
  62084=>"101100001",
  62085=>"000011111",
  62086=>"010001001",
  62087=>"011011100",
  62088=>"110001011",
  62089=>"000010001",
  62090=>"001101110",
  62091=>"011101111",
  62092=>"011010011",
  62093=>"000001000",
  62094=>"011001010",
  62095=>"000111010",
  62096=>"110111100",
  62097=>"001001111",
  62098=>"101000001",
  62099=>"101101110",
  62100=>"110111111",
  62101=>"010010111",
  62102=>"111110101",
  62103=>"010011100",
  62104=>"110000001",
  62105=>"100010111",
  62106=>"101011010",
  62107=>"101011101",
  62108=>"110100110",
  62109=>"001101100",
  62110=>"010000100",
  62111=>"000011000",
  62112=>"101110100",
  62113=>"010111100",
  62114=>"001011101",
  62115=>"110101100",
  62116=>"110000011",
  62117=>"110110001",
  62118=>"011000100",
  62119=>"011000011",
  62120=>"000010000",
  62121=>"000010000",
  62122=>"000110111",
  62123=>"010111000",
  62124=>"101000011",
  62125=>"000110010",
  62126=>"000001101",
  62127=>"111011110",
  62128=>"001100000",
  62129=>"110011000",
  62130=>"101111010",
  62131=>"110110110",
  62132=>"110001001",
  62133=>"010010101",
  62134=>"010101110",
  62135=>"001000101",
  62136=>"110100101",
  62137=>"001011101",
  62138=>"000101010",
  62139=>"101000101",
  62140=>"111100001",
  62141=>"011100010",
  62142=>"000011100",
  62143=>"000000111",
  62144=>"001100100",
  62145=>"110001100",
  62146=>"111111010",
  62147=>"111010011",
  62148=>"100010100",
  62149=>"010101100",
  62150=>"110111100",
  62151=>"101110100",
  62152=>"100000000",
  62153=>"000111111",
  62154=>"101111111",
  62155=>"000101111",
  62156=>"100010000",
  62157=>"001011111",
  62158=>"000001000",
  62159=>"011101111",
  62160=>"110001100",
  62161=>"101110110",
  62162=>"110111000",
  62163=>"010010011",
  62164=>"110010101",
  62165=>"001010111",
  62166=>"101101011",
  62167=>"111100011",
  62168=>"010010000",
  62169=>"011001000",
  62170=>"111000001",
  62171=>"000000000",
  62172=>"101111100",
  62173=>"001101010",
  62174=>"111100110",
  62175=>"101100100",
  62176=>"010000000",
  62177=>"101111001",
  62178=>"001011011",
  62179=>"011001100",
  62180=>"100010010",
  62181=>"111101010",
  62182=>"110111100",
  62183=>"111111111",
  62184=>"011110001",
  62185=>"100001011",
  62186=>"011001110",
  62187=>"110111011",
  62188=>"001010001",
  62189=>"100100110",
  62190=>"001010001",
  62191=>"000100110",
  62192=>"110111111",
  62193=>"010010101",
  62194=>"000011010",
  62195=>"100000111",
  62196=>"010000100",
  62197=>"101000000",
  62198=>"001100001",
  62199=>"000000110",
  62200=>"101111000",
  62201=>"110110110",
  62202=>"101001110",
  62203=>"000110110",
  62204=>"001110101",
  62205=>"011001100",
  62206=>"101001001",
  62207=>"001011111",
  62208=>"010110100",
  62209=>"001100111",
  62210=>"111100010",
  62211=>"010111010",
  62212=>"010100101",
  62213=>"010000001",
  62214=>"000111011",
  62215=>"110011101",
  62216=>"111110000",
  62217=>"101011010",
  62218=>"011110110",
  62219=>"000000001",
  62220=>"111000000",
  62221=>"111011110",
  62222=>"100111000",
  62223=>"100101101",
  62224=>"110101101",
  62225=>"000000001",
  62226=>"011000010",
  62227=>"100111010",
  62228=>"001110110",
  62229=>"100100100",
  62230=>"110110010",
  62231=>"011010001",
  62232=>"001011010",
  62233=>"100000101",
  62234=>"010111111",
  62235=>"110000010",
  62236=>"001000110",
  62237=>"100011101",
  62238=>"110000011",
  62239=>"101101001",
  62240=>"010101110",
  62241=>"010000010",
  62242=>"110010010",
  62243=>"001011100",
  62244=>"101011001",
  62245=>"000110111",
  62246=>"101000111",
  62247=>"010000101",
  62248=>"110100001",
  62249=>"110011001",
  62250=>"100001010",
  62251=>"101100100",
  62252=>"101001111",
  62253=>"000001110",
  62254=>"011000010",
  62255=>"000111011",
  62256=>"110010111",
  62257=>"001111101",
  62258=>"000010110",
  62259=>"110001101",
  62260=>"100001001",
  62261=>"110111001",
  62262=>"101010010",
  62263=>"001101000",
  62264=>"011111011",
  62265=>"001110010",
  62266=>"101101111",
  62267=>"100000100",
  62268=>"010010011",
  62269=>"001101011",
  62270=>"101110001",
  62271=>"000100110",
  62272=>"101101000",
  62273=>"001010000",
  62274=>"000010000",
  62275=>"000000001",
  62276=>"011010001",
  62277=>"001010010",
  62278=>"111000010",
  62279=>"011110100",
  62280=>"100100010",
  62281=>"111111001",
  62282=>"011110010",
  62283=>"111111100",
  62284=>"010000110",
  62285=>"010001101",
  62286=>"000111000",
  62287=>"111111101",
  62288=>"000100001",
  62289=>"000101001",
  62290=>"001011011",
  62291=>"111011101",
  62292=>"101000100",
  62293=>"111011001",
  62294=>"001100100",
  62295=>"101100111",
  62296=>"111010000",
  62297=>"100101101",
  62298=>"010000101",
  62299=>"000100110",
  62300=>"010001001",
  62301=>"110110001",
  62302=>"001000000",
  62303=>"010111011",
  62304=>"100110110",
  62305=>"100000001",
  62306=>"000010110",
  62307=>"101011111",
  62308=>"100100010",
  62309=>"011100110",
  62310=>"111111101",
  62311=>"110011001",
  62312=>"011101001",
  62313=>"111111010",
  62314=>"000101010",
  62315=>"110101001",
  62316=>"001110000",
  62317=>"111111110",
  62318=>"101011011",
  62319=>"110111010",
  62320=>"111111001",
  62321=>"010000110",
  62322=>"111101111",
  62323=>"001111000",
  62324=>"111010101",
  62325=>"010111001",
  62326=>"011111000",
  62327=>"001100000",
  62328=>"111101110",
  62329=>"000001001",
  62330=>"101011010",
  62331=>"100111111",
  62332=>"010000001",
  62333=>"111000110",
  62334=>"001111001",
  62335=>"100110100",
  62336=>"011001000",
  62337=>"001110011",
  62338=>"000100010",
  62339=>"010000010",
  62340=>"001011001",
  62341=>"011000000",
  62342=>"101101111",
  62343=>"010011101",
  62344=>"100100000",
  62345=>"000000000",
  62346=>"010011110",
  62347=>"000100011",
  62348=>"000001010",
  62349=>"000110010",
  62350=>"100001001",
  62351=>"100100001",
  62352=>"111000011",
  62353=>"101110010",
  62354=>"101100100",
  62355=>"001001100",
  62356=>"011001011",
  62357=>"011111111",
  62358=>"110100100",
  62359=>"101110110",
  62360=>"110001110",
  62361=>"010001000",
  62362=>"000111110",
  62363=>"001101101",
  62364=>"100011111",
  62365=>"010100101",
  62366=>"010010011",
  62367=>"010110011",
  62368=>"100110101",
  62369=>"101110110",
  62370=>"001001000",
  62371=>"100101011",
  62372=>"001110011",
  62373=>"101111110",
  62374=>"100111010",
  62375=>"111010010",
  62376=>"111100101",
  62377=>"011001001",
  62378=>"110011011",
  62379=>"001001100",
  62380=>"000100010",
  62381=>"001000001",
  62382=>"001101000",
  62383=>"001101100",
  62384=>"101000100",
  62385=>"010000111",
  62386=>"000010001",
  62387=>"100110111",
  62388=>"110110100",
  62389=>"010100010",
  62390=>"101101101",
  62391=>"000111011",
  62392=>"000011010",
  62393=>"010000011",
  62394=>"111011011",
  62395=>"010011001",
  62396=>"110010001",
  62397=>"011100100",
  62398=>"000000011",
  62399=>"110011111",
  62400=>"100111111",
  62401=>"101110011",
  62402=>"011000010",
  62403=>"010011101",
  62404=>"010101111",
  62405=>"101100011",
  62406=>"101010101",
  62407=>"000010100",
  62408=>"000010111",
  62409=>"011010000",
  62410=>"111101101",
  62411=>"001101001",
  62412=>"110110100",
  62413=>"000000111",
  62414=>"101011010",
  62415=>"000010111",
  62416=>"000001110",
  62417=>"101001100",
  62418=>"100111011",
  62419=>"000001111",
  62420=>"000101111",
  62421=>"000101101",
  62422=>"111000011",
  62423=>"011100111",
  62424=>"000001010",
  62425=>"010110000",
  62426=>"000011111",
  62427=>"010100100",
  62428=>"110111000",
  62429=>"011010011",
  62430=>"110010010",
  62431=>"100000011",
  62432=>"010010101",
  62433=>"000100010",
  62434=>"000010000",
  62435=>"000000010",
  62436=>"000110011",
  62437=>"000000000",
  62438=>"001110011",
  62439=>"110111111",
  62440=>"010101010",
  62441=>"111001100",
  62442=>"000110101",
  62443=>"111000000",
  62444=>"000100110",
  62445=>"000111101",
  62446=>"101110111",
  62447=>"001010100",
  62448=>"010101010",
  62449=>"001001010",
  62450=>"110010000",
  62451=>"100110011",
  62452=>"010101001",
  62453=>"011001101",
  62454=>"010010100",
  62455=>"101111101",
  62456=>"010011001",
  62457=>"100111001",
  62458=>"011010001",
  62459=>"110000001",
  62460=>"011111001",
  62461=>"001100110",
  62462=>"110110010",
  62463=>"001101000",
  62464=>"010111100",
  62465=>"110010101",
  62466=>"101001000",
  62467=>"001000111",
  62468=>"001001100",
  62469=>"111111000",
  62470=>"111111000",
  62471=>"010010100",
  62472=>"111111001",
  62473=>"011101101",
  62474=>"111100101",
  62475=>"011101110",
  62476=>"001111111",
  62477=>"000000111",
  62478=>"010011111",
  62479=>"111110111",
  62480=>"010101010",
  62481=>"011110110",
  62482=>"110011101",
  62483=>"110110011",
  62484=>"000000010",
  62485=>"100011001",
  62486=>"101101011",
  62487=>"001011000",
  62488=>"001110110",
  62489=>"100001011",
  62490=>"111100101",
  62491=>"001100110",
  62492=>"000110100",
  62493=>"100001001",
  62494=>"011100110",
  62495=>"111100010",
  62496=>"010101111",
  62497=>"111000000",
  62498=>"100000000",
  62499=>"001000101",
  62500=>"010001100",
  62501=>"001101011",
  62502=>"011111100",
  62503=>"000100001",
  62504=>"101100101",
  62505=>"000110101",
  62506=>"100100111",
  62507=>"100011011",
  62508=>"101101000",
  62509=>"001011010",
  62510=>"000101110",
  62511=>"110010101",
  62512=>"000100100",
  62513=>"011011010",
  62514=>"011101101",
  62515=>"010001001",
  62516=>"010011011",
  62517=>"111010010",
  62518=>"011100101",
  62519=>"001010010",
  62520=>"010010111",
  62521=>"001101011",
  62522=>"001010101",
  62523=>"000010111",
  62524=>"011011011",
  62525=>"110000011",
  62526=>"110011011",
  62527=>"010010010",
  62528=>"011011100",
  62529=>"111100110",
  62530=>"010100010",
  62531=>"000100111",
  62532=>"000011000",
  62533=>"111101010",
  62534=>"000000011",
  62535=>"110110101",
  62536=>"100110110",
  62537=>"010110111",
  62538=>"001110001",
  62539=>"001010011",
  62540=>"000111101",
  62541=>"000100001",
  62542=>"000000111",
  62543=>"111101011",
  62544=>"111111100",
  62545=>"010100001",
  62546=>"011011111",
  62547=>"100000001",
  62548=>"110110010",
  62549=>"000110100",
  62550=>"011010011",
  62551=>"011011111",
  62552=>"111111111",
  62553=>"101111110",
  62554=>"101011001",
  62555=>"011100001",
  62556=>"011000010",
  62557=>"110101110",
  62558=>"100000010",
  62559=>"001000000",
  62560=>"100111100",
  62561=>"001110010",
  62562=>"000100011",
  62563=>"111100101",
  62564=>"100111100",
  62565=>"110111001",
  62566=>"100110111",
  62567=>"110100101",
  62568=>"010101000",
  62569=>"100001011",
  62570=>"011000010",
  62571=>"011001011",
  62572=>"110011110",
  62573=>"011010100",
  62574=>"101010110",
  62575=>"000100111",
  62576=>"101101001",
  62577=>"001000001",
  62578=>"001110001",
  62579=>"000010101",
  62580=>"110101111",
  62581=>"100111101",
  62582=>"011101001",
  62583=>"100000111",
  62584=>"101001100",
  62585=>"111011111",
  62586=>"111101001",
  62587=>"000010011",
  62588=>"101011011",
  62589=>"110010000",
  62590=>"011100100",
  62591=>"111001011",
  62592=>"111111000",
  62593=>"111101101",
  62594=>"110100011",
  62595=>"011110011",
  62596=>"011001000",
  62597=>"110011110",
  62598=>"011111111",
  62599=>"000001010",
  62600=>"010010101",
  62601=>"000011001",
  62602=>"010001000",
  62603=>"011001100",
  62604=>"111001010",
  62605=>"111111101",
  62606=>"000100011",
  62607=>"001101001",
  62608=>"001100010",
  62609=>"010011100",
  62610=>"010101111",
  62611=>"101100111",
  62612=>"101111110",
  62613=>"011011011",
  62614=>"101011000",
  62615=>"011100001",
  62616=>"100000111",
  62617=>"011011111",
  62618=>"110101101",
  62619=>"000010010",
  62620=>"001011110",
  62621=>"100010110",
  62622=>"001001011",
  62623=>"110110011",
  62624=>"001001011",
  62625=>"101111011",
  62626=>"010101110",
  62627=>"000001111",
  62628=>"100011110",
  62629=>"110000110",
  62630=>"010100111",
  62631=>"110001111",
  62632=>"010100100",
  62633=>"110001010",
  62634=>"101110000",
  62635=>"111000010",
  62636=>"101101011",
  62637=>"010011001",
  62638=>"001101111",
  62639=>"110111010",
  62640=>"111011100",
  62641=>"000101011",
  62642=>"000000111",
  62643=>"010010001",
  62644=>"000010111",
  62645=>"100001000",
  62646=>"111001111",
  62647=>"101100100",
  62648=>"101110000",
  62649=>"111001011",
  62650=>"100100010",
  62651=>"001100111",
  62652=>"110111110",
  62653=>"111010110",
  62654=>"111101111",
  62655=>"001010000",
  62656=>"010110001",
  62657=>"100100100",
  62658=>"001110001",
  62659=>"000111101",
  62660=>"110101110",
  62661=>"000111001",
  62662=>"111110110",
  62663=>"000000001",
  62664=>"010001110",
  62665=>"011001010",
  62666=>"110100101",
  62667=>"000101000",
  62668=>"000101010",
  62669=>"010101101",
  62670=>"011011111",
  62671=>"000100111",
  62672=>"100101100",
  62673=>"111110100",
  62674=>"000010011",
  62675=>"101111010",
  62676=>"000000000",
  62677=>"110001101",
  62678=>"101111000",
  62679=>"010011100",
  62680=>"011011011",
  62681=>"001101010",
  62682=>"001010100",
  62683=>"101101101",
  62684=>"010100010",
  62685=>"000101010",
  62686=>"100001000",
  62687=>"111000000",
  62688=>"000011100",
  62689=>"011011100",
  62690=>"101111101",
  62691=>"000000110",
  62692=>"011010000",
  62693=>"000111011",
  62694=>"111000011",
  62695=>"000011100",
  62696=>"010001001",
  62697=>"110001000",
  62698=>"011110101",
  62699=>"010011011",
  62700=>"101110000",
  62701=>"001000001",
  62702=>"010101011",
  62703=>"110010000",
  62704=>"001110011",
  62705=>"010010010",
  62706=>"010111011",
  62707=>"110001010",
  62708=>"011101010",
  62709=>"000001000",
  62710=>"000101110",
  62711=>"111101110",
  62712=>"101011110",
  62713=>"000101111",
  62714=>"110110101",
  62715=>"000011011",
  62716=>"011011101",
  62717=>"010101100",
  62718=>"111111000",
  62719=>"100001010",
  62720=>"101001000",
  62721=>"110011000",
  62722=>"011000010",
  62723=>"110000001",
  62724=>"100100101",
  62725=>"010011100",
  62726=>"100000011",
  62727=>"111110011",
  62728=>"001001101",
  62729=>"011010011",
  62730=>"100100100",
  62731=>"111100100",
  62732=>"010000001",
  62733=>"000001010",
  62734=>"000000111",
  62735=>"000001001",
  62736=>"110011001",
  62737=>"011001111",
  62738=>"010011000",
  62739=>"111100010",
  62740=>"100011100",
  62741=>"100010110",
  62742=>"110110011",
  62743=>"110111000",
  62744=>"111000011",
  62745=>"111111001",
  62746=>"111000001",
  62747=>"101001111",
  62748=>"110100111",
  62749=>"001010101",
  62750=>"101100100",
  62751=>"101001101",
  62752=>"111100110",
  62753=>"000111110",
  62754=>"100001101",
  62755=>"111111001",
  62756=>"110110111",
  62757=>"100101101",
  62758=>"000010101",
  62759=>"111000101",
  62760=>"010111110",
  62761=>"011001101",
  62762=>"101111000",
  62763=>"100010101",
  62764=>"100110110",
  62765=>"110101101",
  62766=>"110110100",
  62767=>"110101110",
  62768=>"110101010",
  62769=>"010000110",
  62770=>"010111101",
  62771=>"011010010",
  62772=>"010001010",
  62773=>"110001001",
  62774=>"011011110",
  62775=>"010110100",
  62776=>"011100011",
  62777=>"001110010",
  62778=>"011110100",
  62779=>"010001100",
  62780=>"001101010",
  62781=>"100101111",
  62782=>"010010000",
  62783=>"001000011",
  62784=>"101000010",
  62785=>"010011110",
  62786=>"001101110",
  62787=>"010110110",
  62788=>"110011000",
  62789=>"001110000",
  62790=>"001001100",
  62791=>"110001101",
  62792=>"000011001",
  62793=>"000000001",
  62794=>"111010101",
  62795=>"001110011",
  62796=>"011110101",
  62797=>"011111010",
  62798=>"101010011",
  62799=>"111001001",
  62800=>"111001011",
  62801=>"101010111",
  62802=>"110101010",
  62803=>"100000000",
  62804=>"001011000",
  62805=>"000111110",
  62806=>"110110010",
  62807=>"011101011",
  62808=>"011111111",
  62809=>"100100100",
  62810=>"001111000",
  62811=>"101001001",
  62812=>"100010010",
  62813=>"000010001",
  62814=>"001000001",
  62815=>"000100001",
  62816=>"001110110",
  62817=>"101000010",
  62818=>"100101100",
  62819=>"000010111",
  62820=>"110111100",
  62821=>"110100111",
  62822=>"111110111",
  62823=>"100111000",
  62824=>"010000001",
  62825=>"101011111",
  62826=>"100101000",
  62827=>"101101111",
  62828=>"010100000",
  62829=>"001000111",
  62830=>"000101110",
  62831=>"011011011",
  62832=>"110011011",
  62833=>"011000100",
  62834=>"110101001",
  62835=>"111100111",
  62836=>"001000001",
  62837=>"011101001",
  62838=>"010111110",
  62839=>"001000110",
  62840=>"111100101",
  62841=>"001000001",
  62842=>"000000111",
  62843=>"000110011",
  62844=>"010010111",
  62845=>"000000111",
  62846=>"001010100",
  62847=>"010111111",
  62848=>"010111100",
  62849=>"010011000",
  62850=>"111110010",
  62851=>"100010101",
  62852=>"100101011",
  62853=>"101011010",
  62854=>"110000010",
  62855=>"011011100",
  62856=>"100000010",
  62857=>"100010011",
  62858=>"101101110",
  62859=>"000101010",
  62860=>"111110001",
  62861=>"011011101",
  62862=>"110100001",
  62863=>"001000010",
  62864=>"000000100",
  62865=>"101011011",
  62866=>"110011101",
  62867=>"001101010",
  62868=>"000101001",
  62869=>"110100111",
  62870=>"110111111",
  62871=>"010101010",
  62872=>"101011111",
  62873=>"101100100",
  62874=>"111101010",
  62875=>"011001011",
  62876=>"100011000",
  62877=>"010010010",
  62878=>"110111101",
  62879=>"111100111",
  62880=>"111110101",
  62881=>"000101101",
  62882=>"010001010",
  62883=>"010001001",
  62884=>"100010000",
  62885=>"101010001",
  62886=>"001111000",
  62887=>"001011001",
  62888=>"111010110",
  62889=>"001100110",
  62890=>"000000100",
  62891=>"100000011",
  62892=>"101101011",
  62893=>"001101101",
  62894=>"001100011",
  62895=>"010001101",
  62896=>"010000011",
  62897=>"010111110",
  62898=>"111001100",
  62899=>"001010000",
  62900=>"100101001",
  62901=>"010011100",
  62902=>"010100000",
  62903=>"000000001",
  62904=>"110010000",
  62905=>"010110111",
  62906=>"000011001",
  62907=>"101000100",
  62908=>"010010001",
  62909=>"101011010",
  62910=>"001101110",
  62911=>"011010010",
  62912=>"101111000",
  62913=>"011100010",
  62914=>"000000110",
  62915=>"010001101",
  62916=>"000010010",
  62917=>"000101010",
  62918=>"000001000",
  62919=>"001000011",
  62920=>"101011000",
  62921=>"001011000",
  62922=>"011010101",
  62923=>"001111110",
  62924=>"100001100",
  62925=>"110101100",
  62926=>"100001001",
  62927=>"111111111",
  62928=>"111100110",
  62929=>"111001110",
  62930=>"010000001",
  62931=>"001010100",
  62932=>"100011110",
  62933=>"110100101",
  62934=>"101110001",
  62935=>"110010110",
  62936=>"000001111",
  62937=>"101100000",
  62938=>"110111111",
  62939=>"110101111",
  62940=>"101011100",
  62941=>"010001010",
  62942=>"100000000",
  62943=>"001011111",
  62944=>"111110101",
  62945=>"110001111",
  62946=>"110100101",
  62947=>"111000110",
  62948=>"010100111",
  62949=>"000000010",
  62950=>"011010110",
  62951=>"011001100",
  62952=>"000011111",
  62953=>"100000010",
  62954=>"110101111",
  62955=>"000000000",
  62956=>"011110011",
  62957=>"111101111",
  62958=>"111110111",
  62959=>"010010010",
  62960=>"001010110",
  62961=>"000100100",
  62962=>"010001111",
  62963=>"111001101",
  62964=>"000011101",
  62965=>"111001000",
  62966=>"101011011",
  62967=>"110011001",
  62968=>"110110111",
  62969=>"100110100",
  62970=>"000000110",
  62971=>"110010010",
  62972=>"111100001",
  62973=>"011100000",
  62974=>"100110010",
  62975=>"001010100",
  62976=>"010101111",
  62977=>"100010110",
  62978=>"110110000",
  62979=>"101101001",
  62980=>"010001001",
  62981=>"110100001",
  62982=>"100001100",
  62983=>"000000111",
  62984=>"000000111",
  62985=>"011100001",
  62986=>"101110000",
  62987=>"011101010",
  62988=>"110011100",
  62989=>"001000000",
  62990=>"100101110",
  62991=>"101100111",
  62992=>"101000101",
  62993=>"001011000",
  62994=>"011000101",
  62995=>"000101101",
  62996=>"000101100",
  62997=>"010010011",
  62998=>"110010100",
  62999=>"101001111",
  63000=>"000011000",
  63001=>"010001100",
  63002=>"000110000",
  63003=>"110100110",
  63004=>"000000011",
  63005=>"000111100",
  63006=>"000000010",
  63007=>"111101001",
  63008=>"011010111",
  63009=>"111111010",
  63010=>"001010001",
  63011=>"001101000",
  63012=>"011101101",
  63013=>"101100011",
  63014=>"100011001",
  63015=>"001010010",
  63016=>"100001010",
  63017=>"001101101",
  63018=>"110011101",
  63019=>"010111110",
  63020=>"110111000",
  63021=>"000001010",
  63022=>"110010101",
  63023=>"000011000",
  63024=>"011001000",
  63025=>"100001010",
  63026=>"001111000",
  63027=>"011011011",
  63028=>"000001000",
  63029=>"001111011",
  63030=>"001101110",
  63031=>"010010000",
  63032=>"010001011",
  63033=>"000110100",
  63034=>"111001100",
  63035=>"111010000",
  63036=>"100000101",
  63037=>"100000110",
  63038=>"000110001",
  63039=>"110111001",
  63040=>"111100111",
  63041=>"100110000",
  63042=>"011001000",
  63043=>"100010000",
  63044=>"101000101",
  63045=>"100011011",
  63046=>"101100010",
  63047=>"010101100",
  63048=>"110111000",
  63049=>"100111011",
  63050=>"010001010",
  63051=>"010011010",
  63052=>"111001101",
  63053=>"100010101",
  63054=>"000100011",
  63055=>"010010010",
  63056=>"001000111",
  63057=>"100001000",
  63058=>"011011101",
  63059=>"000010111",
  63060=>"000000010",
  63061=>"011100001",
  63062=>"010101011",
  63063=>"111010010",
  63064=>"100010100",
  63065=>"000010101",
  63066=>"000000011",
  63067=>"000110001",
  63068=>"001010111",
  63069=>"100010111",
  63070=>"110110010",
  63071=>"111011100",
  63072=>"001111101",
  63073=>"011001000",
  63074=>"111000100",
  63075=>"101111001",
  63076=>"001111010",
  63077=>"010011000",
  63078=>"100111110",
  63079=>"111100001",
  63080=>"110010110",
  63081=>"110100000",
  63082=>"011111110",
  63083=>"110111111",
  63084=>"110000011",
  63085=>"000000000",
  63086=>"100100000",
  63087=>"110011111",
  63088=>"001000010",
  63089=>"010100100",
  63090=>"100000010",
  63091=>"110111010",
  63092=>"101111110",
  63093=>"000010100",
  63094=>"000001010",
  63095=>"100110110",
  63096=>"001011001",
  63097=>"101001011",
  63098=>"011111111",
  63099=>"100010111",
  63100=>"001111000",
  63101=>"010010100",
  63102=>"101011010",
  63103=>"010010111",
  63104=>"100001001",
  63105=>"000010110",
  63106=>"100001011",
  63107=>"000001001",
  63108=>"100000000",
  63109=>"000000000",
  63110=>"011100001",
  63111=>"111101011",
  63112=>"110111000",
  63113=>"100110111",
  63114=>"111110010",
  63115=>"101101001",
  63116=>"001000111",
  63117=>"000000111",
  63118=>"010111111",
  63119=>"111000000",
  63120=>"110111001",
  63121=>"000100110",
  63122=>"110001001",
  63123=>"110000110",
  63124=>"010100011",
  63125=>"011010000",
  63126=>"010100110",
  63127=>"000000100",
  63128=>"010110001",
  63129=>"111100001",
  63130=>"001111111",
  63131=>"100010011",
  63132=>"100011011",
  63133=>"110000110",
  63134=>"011110011",
  63135=>"000010000",
  63136=>"000010100",
  63137=>"010011010",
  63138=>"010000100",
  63139=>"000111100",
  63140=>"100000011",
  63141=>"010001111",
  63142=>"000100010",
  63143=>"110000001",
  63144=>"010111001",
  63145=>"010000001",
  63146=>"001110011",
  63147=>"111101010",
  63148=>"101111010",
  63149=>"110011001",
  63150=>"100001110",
  63151=>"011110101",
  63152=>"100010101",
  63153=>"101011100",
  63154=>"101100101",
  63155=>"100110110",
  63156=>"000101010",
  63157=>"011101110",
  63158=>"000000010",
  63159=>"110010101",
  63160=>"011100000",
  63161=>"110011011",
  63162=>"111100111",
  63163=>"000001101",
  63164=>"100011011",
  63165=>"100111000",
  63166=>"000011110",
  63167=>"100010110",
  63168=>"100001100",
  63169=>"111100001",
  63170=>"000011101",
  63171=>"000011001",
  63172=>"010111111",
  63173=>"100110000",
  63174=>"111000101",
  63175=>"000000111",
  63176=>"000111000",
  63177=>"111001111",
  63178=>"101110100",
  63179=>"110101010",
  63180=>"110111011",
  63181=>"000000110",
  63182=>"011010000",
  63183=>"000100011",
  63184=>"110101001",
  63185=>"111111011",
  63186=>"010001111",
  63187=>"100110111",
  63188=>"010011010",
  63189=>"001101110",
  63190=>"001101001",
  63191=>"011001110",
  63192=>"111010000",
  63193=>"111100111",
  63194=>"001111000",
  63195=>"010000011",
  63196=>"000111010",
  63197=>"000110001",
  63198=>"011011010",
  63199=>"000001011",
  63200=>"010000000",
  63201=>"110111010",
  63202=>"010000011",
  63203=>"111100101",
  63204=>"001001000",
  63205=>"010111100",
  63206=>"001011111",
  63207=>"010011110",
  63208=>"000110101",
  63209=>"001101011",
  63210=>"011110111",
  63211=>"111001110",
  63212=>"101101110",
  63213=>"001000100",
  63214=>"101011001",
  63215=>"010010010",
  63216=>"101111110",
  63217=>"100000000",
  63218=>"101001010",
  63219=>"011111010",
  63220=>"001001101",
  63221=>"001010001",
  63222=>"110110110",
  63223=>"010010001",
  63224=>"111101111",
  63225=>"110001110",
  63226=>"111110001",
  63227=>"001101001",
  63228=>"111010010",
  63229=>"101100001",
  63230=>"011010011",
  63231=>"100111000",
  63232=>"000011010",
  63233=>"111101010",
  63234=>"110010100",
  63235=>"110010100",
  63236=>"011001010",
  63237=>"001110100",
  63238=>"001010000",
  63239=>"111101111",
  63240=>"000111010",
  63241=>"101001111",
  63242=>"001011111",
  63243=>"110101101",
  63244=>"110111110",
  63245=>"110010011",
  63246=>"111000011",
  63247=>"011101000",
  63248=>"010000000",
  63249=>"110100011",
  63250=>"100000000",
  63251=>"001011110",
  63252=>"001000111",
  63253=>"000110001",
  63254=>"011010100",
  63255=>"110110111",
  63256=>"000101000",
  63257=>"110000001",
  63258=>"000011001",
  63259=>"011111100",
  63260=>"001000111",
  63261=>"111100111",
  63262=>"111011001",
  63263=>"100100100",
  63264=>"001001010",
  63265=>"010111101",
  63266=>"110100001",
  63267=>"011111111",
  63268=>"011010010",
  63269=>"000000110",
  63270=>"001011110",
  63271=>"101111011",
  63272=>"000100010",
  63273=>"010100101",
  63274=>"011000011",
  63275=>"001100101",
  63276=>"001110111",
  63277=>"001001010",
  63278=>"010000011",
  63279=>"011000011",
  63280=>"110000101",
  63281=>"111110110",
  63282=>"110100000",
  63283=>"110000100",
  63284=>"001010001",
  63285=>"101001100",
  63286=>"101000100",
  63287=>"110001110",
  63288=>"101101110",
  63289=>"111101111",
  63290=>"100000111",
  63291=>"000000001",
  63292=>"001011011",
  63293=>"100100101",
  63294=>"010110000",
  63295=>"111000011",
  63296=>"110111001",
  63297=>"101001100",
  63298=>"011000101",
  63299=>"001100000",
  63300=>"110011001",
  63301=>"110011011",
  63302=>"010010111",
  63303=>"110101010",
  63304=>"110110100",
  63305=>"101111010",
  63306=>"010011010",
  63307=>"110000111",
  63308=>"111110101",
  63309=>"010000001",
  63310=>"000100111",
  63311=>"000100101",
  63312=>"000111011",
  63313=>"010010110",
  63314=>"111010100",
  63315=>"001101101",
  63316=>"111011001",
  63317=>"110011100",
  63318=>"001000010",
  63319=>"011110000",
  63320=>"010111111",
  63321=>"011110000",
  63322=>"010110101",
  63323=>"101101000",
  63324=>"111100010",
  63325=>"101110010",
  63326=>"000111011",
  63327=>"010010100",
  63328=>"000110110",
  63329=>"010001111",
  63330=>"100000000",
  63331=>"011101011",
  63332=>"000100010",
  63333=>"100111011",
  63334=>"101011001",
  63335=>"110101010",
  63336=>"011111110",
  63337=>"010010000",
  63338=>"001000110",
  63339=>"101111101",
  63340=>"001110000",
  63341=>"100000000",
  63342=>"111101000",
  63343=>"000000000",
  63344=>"110101110",
  63345=>"000001000",
  63346=>"110010001",
  63347=>"100100010",
  63348=>"110000101",
  63349=>"111111101",
  63350=>"011010100",
  63351=>"100000110",
  63352=>"010100111",
  63353=>"110011100",
  63354=>"110000011",
  63355=>"101101000",
  63356=>"000011111",
  63357=>"001001001",
  63358=>"110000001",
  63359=>"001011110",
  63360=>"001110111",
  63361=>"110000101",
  63362=>"011011100",
  63363=>"110111110",
  63364=>"010111001",
  63365=>"001110110",
  63366=>"000110001",
  63367=>"100000110",
  63368=>"011001101",
  63369=>"110010101",
  63370=>"111110010",
  63371=>"001000101",
  63372=>"110010101",
  63373=>"010111000",
  63374=>"110011101",
  63375=>"100010001",
  63376=>"000101100",
  63377=>"101000110",
  63378=>"010000100",
  63379=>"000010110",
  63380=>"110001110",
  63381=>"000111010",
  63382=>"100010001",
  63383=>"111001111",
  63384=>"100010010",
  63385=>"011011111",
  63386=>"101101111",
  63387=>"101000100",
  63388=>"011010010",
  63389=>"111010111",
  63390=>"001111100",
  63391=>"000001111",
  63392=>"010000000",
  63393=>"110000100",
  63394=>"100100111",
  63395=>"100111101",
  63396=>"110101111",
  63397=>"101101010",
  63398=>"111010010",
  63399=>"000100110",
  63400=>"111111111",
  63401=>"010111010",
  63402=>"001010111",
  63403=>"100110101",
  63404=>"110101110",
  63405=>"010100010",
  63406=>"100001111",
  63407=>"100100110",
  63408=>"001101101",
  63409=>"001110110",
  63410=>"111110000",
  63411=>"011001010",
  63412=>"110111100",
  63413=>"100011111",
  63414=>"111110100",
  63415=>"000100001",
  63416=>"010110111",
  63417=>"111101100",
  63418=>"001110101",
  63419=>"010111011",
  63420=>"100111110",
  63421=>"001101111",
  63422=>"111001000",
  63423=>"000110001",
  63424=>"011110000",
  63425=>"010100110",
  63426=>"000100101",
  63427=>"010011100",
  63428=>"001001000",
  63429=>"110010111",
  63430=>"101110110",
  63431=>"100101100",
  63432=>"111101111",
  63433=>"000111010",
  63434=>"101110011",
  63435=>"001000001",
  63436=>"001101110",
  63437=>"000101101",
  63438=>"100001011",
  63439=>"011000000",
  63440=>"110001011",
  63441=>"101000011",
  63442=>"011001111",
  63443=>"110011010",
  63444=>"011010001",
  63445=>"010001100",
  63446=>"001001000",
  63447=>"011001110",
  63448=>"011101001",
  63449=>"001011011",
  63450=>"110111010",
  63451=>"110000100",
  63452=>"101001111",
  63453=>"111101001",
  63454=>"100000000",
  63455=>"001111111",
  63456=>"010000010",
  63457=>"010110011",
  63458=>"100000110",
  63459=>"000110000",
  63460=>"101001000",
  63461=>"000010010",
  63462=>"001110110",
  63463=>"010011110",
  63464=>"100111011",
  63465=>"111011111",
  63466=>"110111011",
  63467=>"111101000",
  63468=>"010110010",
  63469=>"110001111",
  63470=>"011010110",
  63471=>"110000000",
  63472=>"010110111",
  63473=>"000110110",
  63474=>"011011111",
  63475=>"111000110",
  63476=>"000110010",
  63477=>"001001001",
  63478=>"110010100",
  63479=>"011000101",
  63480=>"000011011",
  63481=>"111001111",
  63482=>"011010011",
  63483=>"001001111",
  63484=>"100101110",
  63485=>"010011101",
  63486=>"010110010",
  63487=>"000100110",
  63488=>"110100000",
  63489=>"100001001",
  63490=>"011101011",
  63491=>"111101101",
  63492=>"100110001",
  63493=>"100111100",
  63494=>"010001000",
  63495=>"011101001",
  63496=>"101000010",
  63497=>"010000011",
  63498=>"000000101",
  63499=>"001011011",
  63500=>"000100010",
  63501=>"010111101",
  63502=>"111100001",
  63503=>"110111000",
  63504=>"100010110",
  63505=>"001100111",
  63506=>"011110001",
  63507=>"110100000",
  63508=>"011011011",
  63509=>"111010101",
  63510=>"100101101",
  63511=>"010010001",
  63512=>"011000101",
  63513=>"100101010",
  63514=>"110100011",
  63515=>"010001100",
  63516=>"010010011",
  63517=>"010010101",
  63518=>"000010100",
  63519=>"111000000",
  63520=>"010111010",
  63521=>"011100010",
  63522=>"010100010",
  63523=>"110111101",
  63524=>"101010010",
  63525=>"111111001",
  63526=>"010000100",
  63527=>"101000100",
  63528=>"011010010",
  63529=>"101111000",
  63530=>"110111111",
  63531=>"110011101",
  63532=>"010000001",
  63533=>"100110011",
  63534=>"101101100",
  63535=>"111001101",
  63536=>"110111101",
  63537=>"110110001",
  63538=>"101011001",
  63539=>"110100111",
  63540=>"110011000",
  63541=>"100101000",
  63542=>"010100010",
  63543=>"010001000",
  63544=>"110011100",
  63545=>"011110011",
  63546=>"000110011",
  63547=>"110010100",
  63548=>"011101010",
  63549=>"000011010",
  63550=>"110100110",
  63551=>"000011101",
  63552=>"011100001",
  63553=>"110010111",
  63554=>"110011001",
  63555=>"000101101",
  63556=>"110110100",
  63557=>"111110010",
  63558=>"110110111",
  63559=>"100101110",
  63560=>"000001100",
  63561=>"000001011",
  63562=>"100001011",
  63563=>"000011111",
  63564=>"001110110",
  63565=>"101010100",
  63566=>"011110111",
  63567=>"010011010",
  63568=>"010101011",
  63569=>"010110011",
  63570=>"101110010",
  63571=>"111100111",
  63572=>"010100011",
  63573=>"000000011",
  63574=>"011011001",
  63575=>"000010000",
  63576=>"001011110",
  63577=>"110001111",
  63578=>"010000000",
  63579=>"101001110",
  63580=>"010110111",
  63581=>"100100101",
  63582=>"011000011",
  63583=>"000000100",
  63584=>"011101111",
  63585=>"111010101",
  63586=>"010110001",
  63587=>"001000011",
  63588=>"011110100",
  63589=>"001100000",
  63590=>"010011111",
  63591=>"100010100",
  63592=>"001001001",
  63593=>"001110000",
  63594=>"110110100",
  63595=>"000101010",
  63596=>"111100101",
  63597=>"001101101",
  63598=>"001000101",
  63599=>"000100111",
  63600=>"111000001",
  63601=>"100000011",
  63602=>"111011111",
  63603=>"010111101",
  63604=>"000111100",
  63605=>"010101100",
  63606=>"010011010",
  63607=>"100011010",
  63608=>"011010000",
  63609=>"100000100",
  63610=>"001000100",
  63611=>"101000110",
  63612=>"000101001",
  63613=>"011100100",
  63614=>"000011000",
  63615=>"111100011",
  63616=>"101011111",
  63617=>"100010000",
  63618=>"010000010",
  63619=>"010110011",
  63620=>"010000111",
  63621=>"000001000",
  63622=>"100000001",
  63623=>"100110001",
  63624=>"010001101",
  63625=>"011100101",
  63626=>"111000100",
  63627=>"001100010",
  63628=>"001111101",
  63629=>"110000011",
  63630=>"111111110",
  63631=>"010101000",
  63632=>"000000010",
  63633=>"110000011",
  63634=>"011100110",
  63635=>"100010111",
  63636=>"100001010",
  63637=>"010011101",
  63638=>"001001100",
  63639=>"111011110",
  63640=>"101100110",
  63641=>"111111110",
  63642=>"000000111",
  63643=>"101101000",
  63644=>"010011001",
  63645=>"100110001",
  63646=>"000001111",
  63647=>"101111111",
  63648=>"101101111",
  63649=>"101110110",
  63650=>"110001100",
  63651=>"000100100",
  63652=>"000101110",
  63653=>"001001110",
  63654=>"010111011",
  63655=>"100110011",
  63656=>"110011011",
  63657=>"100110000",
  63658=>"110100100",
  63659=>"001100000",
  63660=>"110101001",
  63661=>"110011011",
  63662=>"111110111",
  63663=>"010011010",
  63664=>"000111110",
  63665=>"000011011",
  63666=>"100110110",
  63667=>"101001001",
  63668=>"111001001",
  63669=>"110000111",
  63670=>"011001110",
  63671=>"100010010",
  63672=>"100011000",
  63673=>"110101000",
  63674=>"000010100",
  63675=>"011110001",
  63676=>"011011100",
  63677=>"000000010",
  63678=>"111111100",
  63679=>"111100011",
  63680=>"100101110",
  63681=>"000101110",
  63682=>"011011000",
  63683=>"011001011",
  63684=>"010111110",
  63685=>"001001110",
  63686=>"110101110",
  63687=>"001100010",
  63688=>"111100101",
  63689=>"100100001",
  63690=>"010010000",
  63691=>"000100110",
  63692=>"110000000",
  63693=>"100001111",
  63694=>"110000101",
  63695=>"111010111",
  63696=>"001010000",
  63697=>"010010010",
  63698=>"101000010",
  63699=>"101001001",
  63700=>"010001000",
  63701=>"011100011",
  63702=>"101111000",
  63703=>"000010011",
  63704=>"101001000",
  63705=>"011100101",
  63706=>"110110000",
  63707=>"100010101",
  63708=>"001000001",
  63709=>"101100110",
  63710=>"100001001",
  63711=>"101011000",
  63712=>"110000010",
  63713=>"000111000",
  63714=>"110110001",
  63715=>"011001100",
  63716=>"010100011",
  63717=>"010000101",
  63718=>"000100110",
  63719=>"001100110",
  63720=>"100111110",
  63721=>"110111100",
  63722=>"101101101",
  63723=>"001110111",
  63724=>"111100110",
  63725=>"100100001",
  63726=>"110010000",
  63727=>"000111011",
  63728=>"111000010",
  63729=>"010010101",
  63730=>"010000100",
  63731=>"111101101",
  63732=>"101011000",
  63733=>"011100011",
  63734=>"111111101",
  63735=>"000011100",
  63736=>"111100010",
  63737=>"110100001",
  63738=>"100010100",
  63739=>"110001100",
  63740=>"010010010",
  63741=>"011110001",
  63742=>"001011101",
  63743=>"101101111",
  63744=>"110000000",
  63745=>"100010010",
  63746=>"010110011",
  63747=>"000000001",
  63748=>"111101100",
  63749=>"100111011",
  63750=>"010101001",
  63751=>"010101010",
  63752=>"110000000",
  63753=>"000100001",
  63754=>"110011011",
  63755=>"101101100",
  63756=>"010011100",
  63757=>"011101111",
  63758=>"101010001",
  63759=>"101000011",
  63760=>"100000100",
  63761=>"101010100",
  63762=>"010111110",
  63763=>"111111110",
  63764=>"001101000",
  63765=>"100100001",
  63766=>"110110100",
  63767=>"010111001",
  63768=>"011011100",
  63769=>"011101000",
  63770=>"011001111",
  63771=>"001001010",
  63772=>"011010011",
  63773=>"111000110",
  63774=>"001111010",
  63775=>"000000010",
  63776=>"010001011",
  63777=>"011101010",
  63778=>"001101010",
  63779=>"111101111",
  63780=>"111101101",
  63781=>"000011110",
  63782=>"011000000",
  63783=>"001001101",
  63784=>"001110100",
  63785=>"011001110",
  63786=>"000001011",
  63787=>"101010110",
  63788=>"000001011",
  63789=>"001001010",
  63790=>"110100100",
  63791=>"000000011",
  63792=>"000001110",
  63793=>"011111101",
  63794=>"001101101",
  63795=>"010101001",
  63796=>"011001100",
  63797=>"000011111",
  63798=>"000011001",
  63799=>"010010011",
  63800=>"001100011",
  63801=>"011000101",
  63802=>"010011001",
  63803=>"100010000",
  63804=>"000001101",
  63805=>"111100110",
  63806=>"101011001",
  63807=>"100110101",
  63808=>"000000111",
  63809=>"110100010",
  63810=>"010010000",
  63811=>"101111110",
  63812=>"011101111",
  63813=>"001011010",
  63814=>"111001010",
  63815=>"100011101",
  63816=>"001110011",
  63817=>"000001111",
  63818=>"110010011",
  63819=>"110011011",
  63820=>"000001100",
  63821=>"101011011",
  63822=>"010111011",
  63823=>"110000111",
  63824=>"111000111",
  63825=>"111011001",
  63826=>"000100011",
  63827=>"000101101",
  63828=>"111100111",
  63829=>"010101000",
  63830=>"001101000",
  63831=>"100011100",
  63832=>"010100010",
  63833=>"000001000",
  63834=>"101101011",
  63835=>"011001101",
  63836=>"111011000",
  63837=>"011110000",
  63838=>"101000011",
  63839=>"000000110",
  63840=>"101110101",
  63841=>"101101111",
  63842=>"001000101",
  63843=>"000011010",
  63844=>"000000100",
  63845=>"010000001",
  63846=>"000000111",
  63847=>"011001011",
  63848=>"111001001",
  63849=>"100100100",
  63850=>"111111010",
  63851=>"101100111",
  63852=>"001011111",
  63853=>"000111101",
  63854=>"100101100",
  63855=>"111011011",
  63856=>"010000000",
  63857=>"010101110",
  63858=>"000000001",
  63859=>"001010101",
  63860=>"111111011",
  63861=>"101100101",
  63862=>"001101011",
  63863=>"111010010",
  63864=>"001001001",
  63865=>"010110010",
  63866=>"101110000",
  63867=>"101111000",
  63868=>"000100101",
  63869=>"100100010",
  63870=>"100011100",
  63871=>"100001100",
  63872=>"000011100",
  63873=>"011011111",
  63874=>"111111010",
  63875=>"001010100",
  63876=>"111100001",
  63877=>"001100100",
  63878=>"010010000",
  63879=>"000010000",
  63880=>"000000100",
  63881=>"110000111",
  63882=>"100100011",
  63883=>"010101011",
  63884=>"000000110",
  63885=>"000010110",
  63886=>"111001110",
  63887=>"101100100",
  63888=>"110001011",
  63889=>"000101110",
  63890=>"101110111",
  63891=>"101111100",
  63892=>"001100111",
  63893=>"100101101",
  63894=>"011110100",
  63895=>"100111110",
  63896=>"011001001",
  63897=>"101011001",
  63898=>"010110100",
  63899=>"011010100",
  63900=>"111011010",
  63901=>"010100011",
  63902=>"110101001",
  63903=>"001110101",
  63904=>"101100000",
  63905=>"111001111",
  63906=>"010001100",
  63907=>"010100100",
  63908=>"011000000",
  63909=>"011101010",
  63910=>"111110000",
  63911=>"100110111",
  63912=>"101100100",
  63913=>"100111010",
  63914=>"100111100",
  63915=>"000001110",
  63916=>"100000010",
  63917=>"101100101",
  63918=>"111000100",
  63919=>"010010110",
  63920=>"001011110",
  63921=>"111100111",
  63922=>"101111100",
  63923=>"000001111",
  63924=>"100010110",
  63925=>"000111010",
  63926=>"111000010",
  63927=>"101010010",
  63928=>"101000000",
  63929=>"001101110",
  63930=>"111001000",
  63931=>"111100101",
  63932=>"101110111",
  63933=>"110011111",
  63934=>"100011111",
  63935=>"110100001",
  63936=>"101000001",
  63937=>"010101010",
  63938=>"011010001",
  63939=>"111110010",
  63940=>"000010001",
  63941=>"111000000",
  63942=>"010000011",
  63943=>"010000101",
  63944=>"010110100",
  63945=>"101011111",
  63946=>"111101110",
  63947=>"011010110",
  63948=>"100000000",
  63949=>"110111001",
  63950=>"011000110",
  63951=>"000101110",
  63952=>"111111100",
  63953=>"110110011",
  63954=>"110101010",
  63955=>"111101000",
  63956=>"000011111",
  63957=>"110110010",
  63958=>"011010001",
  63959=>"001001001",
  63960=>"010110010",
  63961=>"011111100",
  63962=>"011110100",
  63963=>"100111101",
  63964=>"010010010",
  63965=>"100100110",
  63966=>"110001110",
  63967=>"010101111",
  63968=>"100100000",
  63969=>"000110101",
  63970=>"010010100",
  63971=>"101011111",
  63972=>"110000110",
  63973=>"100001001",
  63974=>"101010001",
  63975=>"111100111",
  63976=>"011001101",
  63977=>"110000011",
  63978=>"010011000",
  63979=>"100000101",
  63980=>"000000011",
  63981=>"100000011",
  63982=>"010000110",
  63983=>"000111000",
  63984=>"111011000",
  63985=>"110001010",
  63986=>"101110100",
  63987=>"100101101",
  63988=>"110100010",
  63989=>"111011010",
  63990=>"001100000",
  63991=>"011011000",
  63992=>"111111010",
  63993=>"010111011",
  63994=>"101001100",
  63995=>"111100111",
  63996=>"010101111",
  63997=>"000110101",
  63998=>"010111111",
  63999=>"101000100",
  64000=>"011101001",
  64001=>"010100100",
  64002=>"111000111",
  64003=>"001111111",
  64004=>"101101100",
  64005=>"010110101",
  64006=>"100000011",
  64007=>"111001000",
  64008=>"110000101",
  64009=>"101101010",
  64010=>"010001111",
  64011=>"111110001",
  64012=>"000101111",
  64013=>"110111100",
  64014=>"110010100",
  64015=>"001001101",
  64016=>"000011011",
  64017=>"011111100",
  64018=>"100001010",
  64019=>"111111111",
  64020=>"000100100",
  64021=>"000000101",
  64022=>"100101110",
  64023=>"110000111",
  64024=>"001001111",
  64025=>"000101000",
  64026=>"001110100",
  64027=>"010101111",
  64028=>"011010000",
  64029=>"000001001",
  64030=>"001101110",
  64031=>"000011110",
  64032=>"100110011",
  64033=>"000100110",
  64034=>"100000010",
  64035=>"111000000",
  64036=>"100001001",
  64037=>"101100001",
  64038=>"111100110",
  64039=>"000011100",
  64040=>"011000100",
  64041=>"111101100",
  64042=>"101001111",
  64043=>"101111001",
  64044=>"110011011",
  64045=>"000100111",
  64046=>"000110100",
  64047=>"000000001",
  64048=>"101110000",
  64049=>"010100101",
  64050=>"011010101",
  64051=>"101100000",
  64052=>"000100001",
  64053=>"001100110",
  64054=>"011101110",
  64055=>"100100111",
  64056=>"111111011",
  64057=>"111110010",
  64058=>"100100101",
  64059=>"010011000",
  64060=>"000101011",
  64061=>"010010011",
  64062=>"110011000",
  64063=>"000101011",
  64064=>"011101000",
  64065=>"110001010",
  64066=>"000010001",
  64067=>"111111001",
  64068=>"000100000",
  64069=>"000001110",
  64070=>"011110010",
  64071=>"000101100",
  64072=>"011101010",
  64073=>"101001110",
  64074=>"011010101",
  64075=>"101101001",
  64076=>"000100000",
  64077=>"100011010",
  64078=>"111000111",
  64079=>"001111101",
  64080=>"110011011",
  64081=>"001110011",
  64082=>"100011110",
  64083=>"000000101",
  64084=>"001000111",
  64085=>"000101000",
  64086=>"101010101",
  64087=>"100100110",
  64088=>"100011111",
  64089=>"111010101",
  64090=>"000110110",
  64091=>"101000110",
  64092=>"011001000",
  64093=>"000101111",
  64094=>"000101101",
  64095=>"110000000",
  64096=>"101101010",
  64097=>"111010101",
  64098=>"011011111",
  64099=>"111001100",
  64100=>"111101101",
  64101=>"011101110",
  64102=>"010011010",
  64103=>"011000111",
  64104=>"111010000",
  64105=>"101001010",
  64106=>"111011100",
  64107=>"000111000",
  64108=>"101101100",
  64109=>"000100110",
  64110=>"100010001",
  64111=>"011100010",
  64112=>"011010001",
  64113=>"000001000",
  64114=>"111110001",
  64115=>"101000110",
  64116=>"111110100",
  64117=>"011001110",
  64118=>"001110010",
  64119=>"100010100",
  64120=>"010100100",
  64121=>"001001001",
  64122=>"101000001",
  64123=>"001101001",
  64124=>"000010001",
  64125=>"011110010",
  64126=>"100011000",
  64127=>"110111011",
  64128=>"110000110",
  64129=>"110000111",
  64130=>"111110010",
  64131=>"011101001",
  64132=>"000001101",
  64133=>"101100000",
  64134=>"101101101",
  64135=>"101001111",
  64136=>"110000000",
  64137=>"000000011",
  64138=>"000100011",
  64139=>"111010000",
  64140=>"000011100",
  64141=>"011000011",
  64142=>"101011101",
  64143=>"110001100",
  64144=>"100100110",
  64145=>"010110010",
  64146=>"111011010",
  64147=>"111101110",
  64148=>"101101100",
  64149=>"110011111",
  64150=>"101110111",
  64151=>"010001010",
  64152=>"011010010",
  64153=>"001110010",
  64154=>"101010101",
  64155=>"001110111",
  64156=>"000000000",
  64157=>"000010101",
  64158=>"110001011",
  64159=>"001101010",
  64160=>"111010101",
  64161=>"010110000",
  64162=>"101100110",
  64163=>"011111110",
  64164=>"110110001",
  64165=>"010101011",
  64166=>"000001101",
  64167=>"010100001",
  64168=>"000011010",
  64169=>"100100011",
  64170=>"011101011",
  64171=>"001110011",
  64172=>"011000011",
  64173=>"100001011",
  64174=>"011101110",
  64175=>"000001100",
  64176=>"011110010",
  64177=>"111110110",
  64178=>"111011111",
  64179=>"111111110",
  64180=>"110111100",
  64181=>"000011101",
  64182=>"001110100",
  64183=>"001011010",
  64184=>"001010110",
  64185=>"100011000",
  64186=>"001101010",
  64187=>"000111001",
  64188=>"010111100",
  64189=>"000010001",
  64190=>"110010001",
  64191=>"011001110",
  64192=>"010000101",
  64193=>"010100000",
  64194=>"110000100",
  64195=>"001101111",
  64196=>"100111110",
  64197=>"011001111",
  64198=>"110100111",
  64199=>"000111010",
  64200=>"110000110",
  64201=>"001001101",
  64202=>"111101101",
  64203=>"110101111",
  64204=>"110101111",
  64205=>"100001110",
  64206=>"111000010",
  64207=>"001110011",
  64208=>"010000001",
  64209=>"100010110",
  64210=>"100010000",
  64211=>"010010011",
  64212=>"011110000",
  64213=>"000110101",
  64214=>"000100111",
  64215=>"101001001",
  64216=>"111000011",
  64217=>"010011111",
  64218=>"110100100",
  64219=>"001000000",
  64220=>"000011001",
  64221=>"110101110",
  64222=>"001111110",
  64223=>"010101100",
  64224=>"100000100",
  64225=>"100011001",
  64226=>"101011011",
  64227=>"111001111",
  64228=>"011111000",
  64229=>"001100000",
  64230=>"010101010",
  64231=>"010101101",
  64232=>"010010011",
  64233=>"000101110",
  64234=>"101111000",
  64235=>"111110100",
  64236=>"000111001",
  64237=>"111100101",
  64238=>"011111001",
  64239=>"001010011",
  64240=>"110111110",
  64241=>"001100111",
  64242=>"001011111",
  64243=>"000000001",
  64244=>"010110011",
  64245=>"101101111",
  64246=>"011101000",
  64247=>"010010000",
  64248=>"111110011",
  64249=>"011000110",
  64250=>"101100100",
  64251=>"011000000",
  64252=>"001010010",
  64253=>"110000111",
  64254=>"110100001",
  64255=>"111110000",
  64256=>"101001001",
  64257=>"101111101",
  64258=>"000101101",
  64259=>"010001011",
  64260=>"110011000",
  64261=>"100101100",
  64262=>"100101100",
  64263=>"101010100",
  64264=>"100100011",
  64265=>"011010000",
  64266=>"101010101",
  64267=>"010010001",
  64268=>"110010011",
  64269=>"001111001",
  64270=>"011010010",
  64271=>"111110110",
  64272=>"100110000",
  64273=>"000111100",
  64274=>"010011101",
  64275=>"000011000",
  64276=>"010011011",
  64277=>"001110110",
  64278=>"110010000",
  64279=>"011011111",
  64280=>"010000110",
  64281=>"000011111",
  64282=>"001110011",
  64283=>"101000011",
  64284=>"010001010",
  64285=>"011000011",
  64286=>"100110100",
  64287=>"001000011",
  64288=>"100010010",
  64289=>"011001001",
  64290=>"111100101",
  64291=>"110011110",
  64292=>"111101101",
  64293=>"010010100",
  64294=>"101011001",
  64295=>"110110110",
  64296=>"001000001",
  64297=>"000110100",
  64298=>"101001111",
  64299=>"111011011",
  64300=>"011000111",
  64301=>"011100110",
  64302=>"000110101",
  64303=>"100011101",
  64304=>"101101100",
  64305=>"111011010",
  64306=>"000011001",
  64307=>"101101110",
  64308=>"000001111",
  64309=>"010101101",
  64310=>"101011001",
  64311=>"000000111",
  64312=>"111011111",
  64313=>"000110101",
  64314=>"001000111",
  64315=>"100011010",
  64316=>"111010001",
  64317=>"101000000",
  64318=>"000100000",
  64319=>"111010011",
  64320=>"000010101",
  64321=>"000100101",
  64322=>"001001011",
  64323=>"010011010",
  64324=>"110010001",
  64325=>"000100101",
  64326=>"000111110",
  64327=>"000001111",
  64328=>"000000010",
  64329=>"101110110",
  64330=>"000101111",
  64331=>"111101100",
  64332=>"010101100",
  64333=>"010000100",
  64334=>"010011111",
  64335=>"100011111",
  64336=>"110011011",
  64337=>"000100011",
  64338=>"000111000",
  64339=>"011101000",
  64340=>"101101100",
  64341=>"100100100",
  64342=>"110110110",
  64343=>"011011010",
  64344=>"011000001",
  64345=>"000110010",
  64346=>"001111001",
  64347=>"110001001",
  64348=>"000000111",
  64349=>"110111000",
  64350=>"000101111",
  64351=>"001001110",
  64352=>"101011110",
  64353=>"000011100",
  64354=>"001111111",
  64355=>"110100110",
  64356=>"100100010",
  64357=>"000011000",
  64358=>"100111010",
  64359=>"001100111",
  64360=>"000000100",
  64361=>"111010000",
  64362=>"101010000",
  64363=>"000101100",
  64364=>"001110110",
  64365=>"111110101",
  64366=>"000111100",
  64367=>"101111010",
  64368=>"001011111",
  64369=>"001111000",
  64370=>"001010111",
  64371=>"101101100",
  64372=>"100001101",
  64373=>"111110000",
  64374=>"011000100",
  64375=>"011100011",
  64376=>"010101101",
  64377=>"100010001",
  64378=>"011110001",
  64379=>"110111100",
  64380=>"010010010",
  64381=>"100100011",
  64382=>"100000001",
  64383=>"000110011",
  64384=>"111011110",
  64385=>"110111011",
  64386=>"000010001",
  64387=>"011010010",
  64388=>"111001000",
  64389=>"110000000",
  64390=>"001100101",
  64391=>"101100001",
  64392=>"001001111",
  64393=>"010001001",
  64394=>"010000101",
  64395=>"001100101",
  64396=>"110010001",
  64397=>"001110110",
  64398=>"010111011",
  64399=>"101011110",
  64400=>"100000010",
  64401=>"011110000",
  64402=>"011010100",
  64403=>"010010100",
  64404=>"000010010",
  64405=>"101100100",
  64406=>"000001001",
  64407=>"001110110",
  64408=>"011001100",
  64409=>"111110000",
  64410=>"000110011",
  64411=>"011011111",
  64412=>"000101101",
  64413=>"001100010",
  64414=>"001010101",
  64415=>"000001001",
  64416=>"010100010",
  64417=>"101101100",
  64418=>"100111010",
  64419=>"110110111",
  64420=>"000100001",
  64421=>"111010011",
  64422=>"011011010",
  64423=>"110011111",
  64424=>"001101000",
  64425=>"110111011",
  64426=>"101101110",
  64427=>"100000000",
  64428=>"101000011",
  64429=>"001000110",
  64430=>"000100101",
  64431=>"111010010",
  64432=>"101111001",
  64433=>"001111101",
  64434=>"000011111",
  64435=>"011101111",
  64436=>"100111110",
  64437=>"011000001",
  64438=>"001110000",
  64439=>"000010001",
  64440=>"101011011",
  64441=>"000111110",
  64442=>"001101101",
  64443=>"010100000",
  64444=>"011110011",
  64445=>"001011000",
  64446=>"111110111",
  64447=>"100001000",
  64448=>"011010101",
  64449=>"101101011",
  64450=>"110001100",
  64451=>"110110101",
  64452=>"101110110",
  64453=>"101011100",
  64454=>"101110100",
  64455=>"000100010",
  64456=>"100100110",
  64457=>"001110001",
  64458=>"100100000",
  64459=>"110001101",
  64460=>"010100010",
  64461=>"111000100",
  64462=>"000011101",
  64463=>"111011111",
  64464=>"001110001",
  64465=>"011000001",
  64466=>"100111101",
  64467=>"110000011",
  64468=>"100000000",
  64469=>"001001111",
  64470=>"001101100",
  64471=>"111101110",
  64472=>"110100010",
  64473=>"000101101",
  64474=>"100101010",
  64475=>"101001011",
  64476=>"001001100",
  64477=>"011111001",
  64478=>"001011100",
  64479=>"010110011",
  64480=>"001101000",
  64481=>"100111010",
  64482=>"011101111",
  64483=>"010000000",
  64484=>"101100101",
  64485=>"001110111",
  64486=>"001001011",
  64487=>"000111110",
  64488=>"100110111",
  64489=>"000010111",
  64490=>"111001101",
  64491=>"010011001",
  64492=>"001101100",
  64493=>"011100111",
  64494=>"001001110",
  64495=>"001010001",
  64496=>"100001101",
  64497=>"010001010",
  64498=>"100001010",
  64499=>"011001101",
  64500=>"001111100",
  64501=>"001000100",
  64502=>"111110001",
  64503=>"110110010",
  64504=>"000001001",
  64505=>"010001111",
  64506=>"001100110",
  64507=>"000010111",
  64508=>"110101101",
  64509=>"101000010",
  64510=>"111010001",
  64511=>"001000110",
  64512=>"011011000",
  64513=>"000011011",
  64514=>"000110101",
  64515=>"110000000",
  64516=>"101111011",
  64517=>"111101101",
  64518=>"011001011",
  64519=>"000111111",
  64520=>"010011101",
  64521=>"111000001",
  64522=>"111101001",
  64523=>"011101000",
  64524=>"101100001",
  64525=>"110111011",
  64526=>"011000001",
  64527=>"111000110",
  64528=>"001110101",
  64529=>"010000010",
  64530=>"100110101",
  64531=>"110110000",
  64532=>"101001110",
  64533=>"010000100",
  64534=>"110011111",
  64535=>"010000001",
  64536=>"111100100",
  64537=>"001000110",
  64538=>"111011100",
  64539=>"100110010",
  64540=>"111000100",
  64541=>"110001110",
  64542=>"001001101",
  64543=>"111001101",
  64544=>"010011110",
  64545=>"110011001",
  64546=>"000101101",
  64547=>"000000010",
  64548=>"010101111",
  64549=>"001010010",
  64550=>"000111011",
  64551=>"010000010",
  64552=>"011111100",
  64553=>"100011111",
  64554=>"010000111",
  64555=>"100001001",
  64556=>"101110001",
  64557=>"111100000",
  64558=>"100010001",
  64559=>"001111001",
  64560=>"101101011",
  64561=>"110010100",
  64562=>"110110000",
  64563=>"010010010",
  64564=>"101111100",
  64565=>"011010001",
  64566=>"110010000",
  64567=>"001101111",
  64568=>"000111011",
  64569=>"001000000",
  64570=>"100110001",
  64571=>"011001010",
  64572=>"100001010",
  64573=>"001010010",
  64574=>"101100100",
  64575=>"010100010",
  64576=>"111001111",
  64577=>"010110001",
  64578=>"110001110",
  64579=>"000010000",
  64580=>"010101010",
  64581=>"101111001",
  64582=>"011001111",
  64583=>"111101110",
  64584=>"101001111",
  64585=>"101001000",
  64586=>"000011011",
  64587=>"011000000",
  64588=>"000110100",
  64589=>"111111101",
  64590=>"110111110",
  64591=>"111111110",
  64592=>"101010110",
  64593=>"111110111",
  64594=>"100011110",
  64595=>"011110110",
  64596=>"100110111",
  64597=>"001101001",
  64598=>"110001010",
  64599=>"100101101",
  64600=>"000000100",
  64601=>"001000000",
  64602=>"111001010",
  64603=>"010100001",
  64604=>"010001101",
  64605=>"110100000",
  64606=>"010010000",
  64607=>"001111001",
  64608=>"100110001",
  64609=>"000101111",
  64610=>"000000000",
  64611=>"101100011",
  64612=>"110101100",
  64613=>"110111101",
  64614=>"100000110",
  64615=>"100110000",
  64616=>"001010001",
  64617=>"011110000",
  64618=>"011110001",
  64619=>"000010110",
  64620=>"100100000",
  64621=>"111110110",
  64622=>"100001000",
  64623=>"100101000",
  64624=>"111101110",
  64625=>"100110001",
  64626=>"111101001",
  64627=>"100010000",
  64628=>"111110000",
  64629=>"110010111",
  64630=>"111000111",
  64631=>"000010011",
  64632=>"110110110",
  64633=>"111110011",
  64634=>"011011000",
  64635=>"101111010",
  64636=>"001011010",
  64637=>"010001111",
  64638=>"010110000",
  64639=>"000010000",
  64640=>"101011100",
  64641=>"101011000",
  64642=>"110011001",
  64643=>"101100000",
  64644=>"011001110",
  64645=>"011010111",
  64646=>"100011011",
  64647=>"110011000",
  64648=>"101001011",
  64649=>"111001111",
  64650=>"101110000",
  64651=>"000100111",
  64652=>"111000111",
  64653=>"101111101",
  64654=>"111110000",
  64655=>"001110001",
  64656=>"101001111",
  64657=>"111011010",
  64658=>"011001001",
  64659=>"101001101",
  64660=>"001011000",
  64661=>"011000000",
  64662=>"001110000",
  64663=>"011011011",
  64664=>"100100110",
  64665=>"011111001",
  64666=>"010001110",
  64667=>"010101001",
  64668=>"110110000",
  64669=>"011001101",
  64670=>"010101010",
  64671=>"101011110",
  64672=>"111001001",
  64673=>"110001110",
  64674=>"110000101",
  64675=>"010100101",
  64676=>"001011001",
  64677=>"001010011",
  64678=>"110010100",
  64679=>"001001011",
  64680=>"010110100",
  64681=>"010111111",
  64682=>"100000111",
  64683=>"100100111",
  64684=>"010011111",
  64685=>"001100010",
  64686=>"110100100",
  64687=>"110101100",
  64688=>"011101100",
  64689=>"101010000",
  64690=>"000110100",
  64691=>"101111100",
  64692=>"100111101",
  64693=>"100010110",
  64694=>"000101101",
  64695=>"011100001",
  64696=>"110001001",
  64697=>"100101011",
  64698=>"000111110",
  64699=>"111111111",
  64700=>"001011011",
  64701=>"010011011",
  64702=>"000100000",
  64703=>"100111011",
  64704=>"110100000",
  64705=>"001010101",
  64706=>"101001100",
  64707=>"011011001",
  64708=>"010110010",
  64709=>"100111000",
  64710=>"010110001",
  64711=>"001000110",
  64712=>"101100010",
  64713=>"100101011",
  64714=>"000111111",
  64715=>"001111111",
  64716=>"111001001",
  64717=>"101111110",
  64718=>"010110010",
  64719=>"101101000",
  64720=>"110101000",
  64721=>"100001010",
  64722=>"100110100",
  64723=>"011100110",
  64724=>"111011011",
  64725=>"101011011",
  64726=>"101111101",
  64727=>"000110011",
  64728=>"101111011",
  64729=>"100011011",
  64730=>"100110100",
  64731=>"110110001",
  64732=>"111011101",
  64733=>"100001010",
  64734=>"111111100",
  64735=>"001100111",
  64736=>"100001101",
  64737=>"111011100",
  64738=>"101001100",
  64739=>"000001001",
  64740=>"100010111",
  64741=>"111111010",
  64742=>"000001101",
  64743=>"111001101",
  64744=>"111010010",
  64745=>"011000101",
  64746=>"001010101",
  64747=>"000101111",
  64748=>"010000110",
  64749=>"101001001",
  64750=>"100000001",
  64751=>"010000100",
  64752=>"101011100",
  64753=>"101101110",
  64754=>"000100011",
  64755=>"011111111",
  64756=>"001100001",
  64757=>"010001101",
  64758=>"001111000",
  64759=>"011100101",
  64760=>"001111011",
  64761=>"011110111",
  64762=>"101101110",
  64763=>"011110111",
  64764=>"101001001",
  64765=>"000010010",
  64766=>"100011101",
  64767=>"101111100",
  64768=>"010110100",
  64769=>"001000101",
  64770=>"100000110",
  64771=>"110111011",
  64772=>"111110100",
  64773=>"111001110",
  64774=>"001000100",
  64775=>"000111101",
  64776=>"011111000",
  64777=>"011010011",
  64778=>"101011011",
  64779=>"010111100",
  64780=>"111100001",
  64781=>"101100000",
  64782=>"111010010",
  64783=>"010101000",
  64784=>"011010001",
  64785=>"010101001",
  64786=>"101101010",
  64787=>"000010101",
  64788=>"100011011",
  64789=>"101110110",
  64790=>"100000111",
  64791=>"100111000",
  64792=>"000000110",
  64793=>"111011000",
  64794=>"100100111",
  64795=>"101110100",
  64796=>"100100100",
  64797=>"000111100",
  64798=>"101001110",
  64799=>"011011101",
  64800=>"010001101",
  64801=>"100110100",
  64802=>"011101110",
  64803=>"101100110",
  64804=>"001111111",
  64805=>"101001111",
  64806=>"110100001",
  64807=>"000101011",
  64808=>"010101111",
  64809=>"001010010",
  64810=>"110010110",
  64811=>"000101000",
  64812=>"111010011",
  64813=>"001100011",
  64814=>"000110011",
  64815=>"011110010",
  64816=>"000110011",
  64817=>"011100010",
  64818=>"001000101",
  64819=>"101001011",
  64820=>"010001011",
  64821=>"011101000",
  64822=>"100101100",
  64823=>"111100111",
  64824=>"000000110",
  64825=>"100010101",
  64826=>"100111001",
  64827=>"110001100",
  64828=>"101000101",
  64829=>"000110110",
  64830=>"110010110",
  64831=>"001001011",
  64832=>"100100101",
  64833=>"100000001",
  64834=>"111110001",
  64835=>"110110101",
  64836=>"001001001",
  64837=>"101010000",
  64838=>"000000000",
  64839=>"000000011",
  64840=>"001111001",
  64841=>"100101000",
  64842=>"111110001",
  64843=>"100000100",
  64844=>"101100111",
  64845=>"111000110",
  64846=>"010011011",
  64847=>"110011101",
  64848=>"000111110",
  64849=>"011000101",
  64850=>"011011011",
  64851=>"111000001",
  64852=>"100010100",
  64853=>"011000011",
  64854=>"111111001",
  64855=>"001001100",
  64856=>"000101110",
  64857=>"110110101",
  64858=>"010100100",
  64859=>"001010001",
  64860=>"101100000",
  64861=>"011010010",
  64862=>"111010111",
  64863=>"000111101",
  64864=>"101010110",
  64865=>"101010010",
  64866=>"000110010",
  64867=>"100101101",
  64868=>"000011101",
  64869=>"100000100",
  64870=>"101100001",
  64871=>"010110011",
  64872=>"011110010",
  64873=>"000001010",
  64874=>"100011011",
  64875=>"000000001",
  64876=>"001010110",
  64877=>"101010101",
  64878=>"000010111",
  64879=>"001101010",
  64880=>"010011111",
  64881=>"111111110",
  64882=>"011101110",
  64883=>"111111001",
  64884=>"011100011",
  64885=>"111011111",
  64886=>"000000001",
  64887=>"000001110",
  64888=>"111111101",
  64889=>"001010101",
  64890=>"010101101",
  64891=>"110111101",
  64892=>"101011111",
  64893=>"101101001",
  64894=>"000100001",
  64895=>"010111101",
  64896=>"011111110",
  64897=>"001000010",
  64898=>"100100111",
  64899=>"001001101",
  64900=>"111001111",
  64901=>"111001010",
  64902=>"001011000",
  64903=>"000010010",
  64904=>"010010011",
  64905=>"001011101",
  64906=>"100110010",
  64907=>"001111010",
  64908=>"100000011",
  64909=>"111111101",
  64910=>"011001010",
  64911=>"100111100",
  64912=>"010101110",
  64913=>"101100001",
  64914=>"011000001",
  64915=>"001001001",
  64916=>"010010011",
  64917=>"100111010",
  64918=>"101011010",
  64919=>"100110001",
  64920=>"101000001",
  64921=>"111110001",
  64922=>"001000101",
  64923=>"110111101",
  64924=>"000010011",
  64925=>"111011001",
  64926=>"011000010",
  64927=>"110111011",
  64928=>"011101111",
  64929=>"100110000",
  64930=>"110000101",
  64931=>"000101001",
  64932=>"101000111",
  64933=>"100000001",
  64934=>"100110001",
  64935=>"000100000",
  64936=>"111010111",
  64937=>"011010011",
  64938=>"000000001",
  64939=>"001111000",
  64940=>"111011011",
  64941=>"000010010",
  64942=>"110001011",
  64943=>"001011100",
  64944=>"100010011",
  64945=>"110101011",
  64946=>"001101101",
  64947=>"001110001",
  64948=>"011111010",
  64949=>"100100000",
  64950=>"101010100",
  64951=>"000111110",
  64952=>"011011010",
  64953=>"011111110",
  64954=>"010000111",
  64955=>"000011011",
  64956=>"010111011",
  64957=>"101111110",
  64958=>"100001010",
  64959=>"010100111",
  64960=>"110001001",
  64961=>"010001111",
  64962=>"101010001",
  64963=>"110011000",
  64964=>"011010101",
  64965=>"001011110",
  64966=>"001101101",
  64967=>"111011110",
  64968=>"001101011",
  64969=>"011011100",
  64970=>"101000001",
  64971=>"011110011",
  64972=>"000010100",
  64973=>"000011001",
  64974=>"011001110",
  64975=>"000011100",
  64976=>"011000110",
  64977=>"001011111",
  64978=>"011010011",
  64979=>"010111011",
  64980=>"100111111",
  64981=>"000001101",
  64982=>"101110101",
  64983=>"101100001",
  64984=>"010101001",
  64985=>"001110010",
  64986=>"101101010",
  64987=>"010111001",
  64988=>"010110100",
  64989=>"010001111",
  64990=>"101100101",
  64991=>"110111100",
  64992=>"000000111",
  64993=>"100101001",
  64994=>"110011100",
  64995=>"111110010",
  64996=>"110101001",
  64997=>"111111011",
  64998=>"100011110",
  64999=>"101100110",
  65000=>"001000001",
  65001=>"000110010",
  65002=>"111011100",
  65003=>"111110000",
  65004=>"000000100",
  65005=>"100000111",
  65006=>"110111101",
  65007=>"101000101",
  65008=>"111001010",
  65009=>"111101010",
  65010=>"010100111",
  65011=>"001110001",
  65012=>"011001011",
  65013=>"101111110",
  65014=>"101001011",
  65015=>"101100000",
  65016=>"110100101",
  65017=>"010011110",
  65018=>"111011100",
  65019=>"001100100",
  65020=>"011000001",
  65021=>"000010011",
  65022=>"010011111",
  65023=>"110010000",
  65024=>"011011011",
  65025=>"001000100",
  65026=>"000001011",
  65027=>"010000101",
  65028=>"101011001",
  65029=>"110100000",
  65030=>"101011111",
  65031=>"111010000",
  65032=>"101101001",
  65033=>"001110110",
  65034=>"000110100",
  65035=>"000001001",
  65036=>"101000101",
  65037=>"110001110",
  65038=>"111001000",
  65039=>"100100101",
  65040=>"101101111",
  65041=>"011100011",
  65042=>"011010000",
  65043=>"100101001",
  65044=>"011000010",
  65045=>"101000011",
  65046=>"010010101",
  65047=>"010011101",
  65048=>"101000000",
  65049=>"001001100",
  65050=>"001000001",
  65051=>"000000000",
  65052=>"001110000",
  65053=>"100000101",
  65054=>"100101111",
  65055=>"011110101",
  65056=>"101001010",
  65057=>"111100010",
  65058=>"000011111",
  65059=>"100101010",
  65060=>"001100110",
  65061=>"110011010",
  65062=>"010001001",
  65063=>"000011011",
  65064=>"111001000",
  65065=>"111001011",
  65066=>"001101000",
  65067=>"000101101",
  65068=>"100100101",
  65069=>"010011010",
  65070=>"100001001",
  65071=>"110100100",
  65072=>"111011101",
  65073=>"000001001",
  65074=>"100000111",
  65075=>"010110010",
  65076=>"000101001",
  65077=>"111110100",
  65078=>"101100110",
  65079=>"100001010",
  65080=>"101011010",
  65081=>"001001001",
  65082=>"111010110",
  65083=>"110110001",
  65084=>"101001110",
  65085=>"100010001",
  65086=>"010010100",
  65087=>"110100001",
  65088=>"010000100",
  65089=>"111111100",
  65090=>"011001100",
  65091=>"101000101",
  65092=>"000000011",
  65093=>"000011100",
  65094=>"010101010",
  65095=>"110010110",
  65096=>"011100100",
  65097=>"111100011",
  65098=>"101110100",
  65099=>"100000100",
  65100=>"000010111",
  65101=>"000101110",
  65102=>"000001001",
  65103=>"001101001",
  65104=>"010001110",
  65105=>"001011101",
  65106=>"111101001",
  65107=>"001010010",
  65108=>"000011000",
  65109=>"101110001",
  65110=>"111101001",
  65111=>"111010101",
  65112=>"101000011",
  65113=>"110011101",
  65114=>"101000100",
  65115=>"001111110",
  65116=>"101110000",
  65117=>"000011001",
  65118=>"100000100",
  65119=>"011110000",
  65120=>"111101001",
  65121=>"100100101",
  65122=>"010100011",
  65123=>"101101011",
  65124=>"110011001",
  65125=>"101100001",
  65126=>"011100110",
  65127=>"000011001",
  65128=>"000000100",
  65129=>"010011110",
  65130=>"100010000",
  65131=>"000111001",
  65132=>"011100100",
  65133=>"100001000",
  65134=>"100111000",
  65135=>"011100111",
  65136=>"011011011",
  65137=>"000000010",
  65138=>"100010000",
  65139=>"001000111",
  65140=>"101100110",
  65141=>"010011100",
  65142=>"101111001",
  65143=>"111000010",
  65144=>"010111111",
  65145=>"001001111",
  65146=>"000011000",
  65147=>"010111101",
  65148=>"010000000",
  65149=>"001111101",
  65150=>"100011000",
  65151=>"011100011",
  65152=>"010010000",
  65153=>"000000001",
  65154=>"011011010",
  65155=>"111001001",
  65156=>"100101001",
  65157=>"110101001",
  65158=>"100110101",
  65159=>"110010001",
  65160=>"100110100",
  65161=>"111101001",
  65162=>"100101010",
  65163=>"011011001",
  65164=>"000001100",
  65165=>"001101011",
  65166=>"111100111",
  65167=>"100000101",
  65168=>"110101010",
  65169=>"101101011",
  65170=>"111001011",
  65171=>"101001100",
  65172=>"101100100",
  65173=>"001011100",
  65174=>"011100110",
  65175=>"100101111",
  65176=>"010010010",
  65177=>"110101100",
  65178=>"101110010",
  65179=>"010110000",
  65180=>"010000000",
  65181=>"000110110",
  65182=>"110110111",
  65183=>"010000110",
  65184=>"100010010",
  65185=>"101001011",
  65186=>"011001000",
  65187=>"001000100",
  65188=>"010000001",
  65189=>"000010101",
  65190=>"100101111",
  65191=>"000001010",
  65192=>"010011011",
  65193=>"111010001",
  65194=>"000001011",
  65195=>"010010011",
  65196=>"001011100",
  65197=>"011110110",
  65198=>"001001000",
  65199=>"010000000",
  65200=>"100001000",
  65201=>"000100100",
  65202=>"011110101",
  65203=>"101100011",
  65204=>"111001110",
  65205=>"101010100",
  65206=>"110011000",
  65207=>"110010000",
  65208=>"110010110",
  65209=>"100000111",
  65210=>"010110111",
  65211=>"101001000",
  65212=>"110111111",
  65213=>"001110001",
  65214=>"001100100",
  65215=>"010110111",
  65216=>"001001101",
  65217=>"101100001",
  65218=>"110110001",
  65219=>"000011010",
  65220=>"000111100",
  65221=>"110110001",
  65222=>"010011110",
  65223=>"100010100",
  65224=>"111010101",
  65225=>"100111100",
  65226=>"000010011",
  65227=>"101111010",
  65228=>"001000100",
  65229=>"111111000",
  65230=>"010000011",
  65231=>"011101111",
  65232=>"110011111",
  65233=>"101111111",
  65234=>"000000011",
  65235=>"111101011",
  65236=>"011001011",
  65237=>"110001110",
  65238=>"010000011",
  65239=>"001010010",
  65240=>"000110010",
  65241=>"111000001",
  65242=>"010001111",
  65243=>"001001100",
  65244=>"101101101",
  65245=>"000110000",
  65246=>"000001010",
  65247=>"100011110",
  65248=>"011111001",
  65249=>"010100001",
  65250=>"101101011",
  65251=>"111000000",
  65252=>"001001011",
  65253=>"110010001",
  65254=>"011010010",
  65255=>"101001011",
  65256=>"110100111",
  65257=>"000101011",
  65258=>"110011111",
  65259=>"010100000",
  65260=>"111001110",
  65261=>"001001000",
  65262=>"011000011",
  65263=>"101010111",
  65264=>"001011000",
  65265=>"110110010",
  65266=>"100010111",
  65267=>"001001011",
  65268=>"001010110",
  65269=>"001111100",
  65270=>"000010111",
  65271=>"101011001",
  65272=>"011001010",
  65273=>"010001000",
  65274=>"101111100",
  65275=>"001010101",
  65276=>"001101011",
  65277=>"000000100",
  65278=>"110000101",
  65279=>"000110000",
  65280=>"000101001",
  65281=>"001100100",
  65282=>"001001011",
  65283=>"000100000",
  65284=>"111110110",
  65285=>"100111011",
  65286=>"001111010",
  65287=>"011111101",
  65288=>"100100010",
  65289=>"001100001",
  65290=>"001110100",
  65291=>"010001000",
  65292=>"100110101",
  65293=>"111110001",
  65294=>"110100100",
  65295=>"111100101",
  65296=>"010111001",
  65297=>"100101101",
  65298=>"001111011",
  65299=>"010011001",
  65300=>"111111101",
  65301=>"000000010",
  65302=>"110101101",
  65303=>"101101110",
  65304=>"001000000",
  65305=>"100000011",
  65306=>"101000010",
  65307=>"000111101",
  65308=>"111000100",
  65309=>"101000001",
  65310=>"001110110",
  65311=>"010010101",
  65312=>"010011000",
  65313=>"010011111",
  65314=>"001111000",
  65315=>"000000000",
  65316=>"001011111",
  65317=>"111101011",
  65318=>"111001100",
  65319=>"000011000",
  65320=>"010101001",
  65321=>"001000010",
  65322=>"011011111",
  65323=>"100100001",
  65324=>"110111000",
  65325=>"101000111",
  65326=>"101010111",
  65327=>"011010010",
  65328=>"101010001",
  65329=>"110001111",
  65330=>"000100100",
  65331=>"010100100",
  65332=>"101000101",
  65333=>"100000001",
  65334=>"111000001",
  65335=>"111110010",
  65336=>"001111100",
  65337=>"000000000",
  65338=>"111001010",
  65339=>"111000110",
  65340=>"110110100",
  65341=>"010010100",
  65342=>"101001100",
  65343=>"010001000",
  65344=>"011111001",
  65345=>"000111001",
  65346=>"010000111",
  65347=>"011110100",
  65348=>"111111001",
  65349=>"011001011",
  65350=>"101110110",
  65351=>"101010010",
  65352=>"100000011",
  65353=>"000011111",
  65354=>"000100000",
  65355=>"001000011",
  65356=>"000000110",
  65357=>"101011001",
  65358=>"100101111",
  65359=>"010101000",
  65360=>"101110111",
  65361=>"001111010",
  65362=>"111011111",
  65363=>"010000000",
  65364=>"010011011",
  65365=>"110000000",
  65366=>"001011100",
  65367=>"100011000",
  65368=>"001111011",
  65369=>"011010010",
  65370=>"110111010",
  65371=>"111100101",
  65372=>"000110111",
  65373=>"001110011",
  65374=>"010010110",
  65375=>"100001010",
  65376=>"000010110",
  65377=>"100101101",
  65378=>"111000111",
  65379=>"001111011",
  65380=>"111111000",
  65381=>"000100101",
  65382=>"110100001",
  65383=>"011000100",
  65384=>"000101111",
  65385=>"101001011",
  65386=>"100101001",
  65387=>"100110000",
  65388=>"100001110",
  65389=>"001000111",
  65390=>"000000000",
  65391=>"111001101",
  65392=>"011001000",
  65393=>"011000011",
  65394=>"011010111",
  65395=>"101111001",
  65396=>"000010011",
  65397=>"110000001",
  65398=>"111000101",
  65399=>"101110101",
  65400=>"001000001",
  65401=>"110100000",
  65402=>"100011001",
  65403=>"000000100",
  65404=>"011000001",
  65405=>"110001010",
  65406=>"011101110",
  65407=>"001111000",
  65408=>"101100101",
  65409=>"110110111",
  65410=>"000110000",
  65411=>"000100000",
  65412=>"100010110",
  65413=>"001110101",
  65414=>"110100011",
  65415=>"011100010",
  65416=>"000000000",
  65417=>"000110110",
  65418=>"000000001",
  65419=>"100001111",
  65420=>"110110011",
  65421=>"010100001",
  65422=>"010100101",
  65423=>"010000010",
  65424=>"110001001",
  65425=>"100000101",
  65426=>"100001011",
  65427=>"101110111",
  65428=>"111110001",
  65429=>"101001010",
  65430=>"001110010",
  65431=>"110000001",
  65432=>"101010110",
  65433=>"101101101",
  65434=>"110001000",
  65435=>"110000101",
  65436=>"001110011",
  65437=>"111000001",
  65438=>"100111110",
  65439=>"011001011",
  65440=>"001110100",
  65441=>"001000011",
  65442=>"011011101",
  65443=>"101001101",
  65444=>"101000010",
  65445=>"000000110",
  65446=>"110100011",
  65447=>"010010011",
  65448=>"001101000",
  65449=>"000011101",
  65450=>"110110101",
  65451=>"000001100",
  65452=>"100001011",
  65453=>"111111001",
  65454=>"001101100",
  65455=>"000011110",
  65456=>"000101110",
  65457=>"001111101",
  65458=>"011110001",
  65459=>"111010010",
  65460=>"100010111",
  65461=>"111101111",
  65462=>"111100010",
  65463=>"010110111",
  65464=>"000100010",
  65465=>"101010001",
  65466=>"110111110",
  65467=>"010010000",
  65468=>"111110101",
  65469=>"000110000",
  65470=>"100011010",
  65471=>"000100101",
  65472=>"101100101",
  65473=>"000101111",
  65474=>"110100000",
  65475=>"001000001",
  65476=>"011000100",
  65477=>"000010001",
  65478=>"111000100",
  65479=>"100010011",
  65480=>"000101110",
  65481=>"111010010",
  65482=>"111110001",
  65483=>"001111010",
  65484=>"001001011",
  65485=>"101100100",
  65486=>"000110010",
  65487=>"011110101",
  65488=>"001101000",
  65489=>"101000000",
  65490=>"100010100",
  65491=>"011100000",
  65492=>"101001011",
  65493=>"000001001",
  65494=>"101001111",
  65495=>"011110001",
  65496=>"100010000",
  65497=>"001101101",
  65498=>"001101100",
  65499=>"100101010",
  65500=>"101010000",
  65501=>"010001101",
  65502=>"010111110",
  65503=>"011111001",
  65504=>"101101000",
  65505=>"000110110",
  65506=>"101101101",
  65507=>"111000011",
  65508=>"100000001",
  65509=>"101111110",
  65510=>"001110000",
  65511=>"100001000",
  65512=>"000000010",
  65513=>"101000010",
  65514=>"000110110",
  65515=>"111100010",
  65516=>"010110101",
  65517=>"101111101",
  65518=>"000010011",
  65519=>"000000011",
  65520=>"101000111",
  65521=>"111000111",
  65522=>"000010100",
  65523=>"100111101",
  65524=>"111011011",
  65525=>"010001101",
  65526=>"101111011",
  65527=>"101111000",
  65528=>"100000100",
  65529=>"111011000",
  65530=>"000100111",
  65531=>"111010001",
  65532=>"111111101",
  65533=>"001000001",
  65534=>"100010010",
  65535=>"000110111");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;