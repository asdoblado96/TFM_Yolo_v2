LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_2_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(5 DOWNTO 0));
END L8_2_BNROM;

ARCHITECTURE RTL OF L8_2_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 63) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"0010010001001101"&"0010001001110110",
  1=>"0001000101000110"&"0001111110101000",
  2=>"0010010001000111"&"0010001110111010",
  3=>"0001011111000111"&"0001011011100110",
  4=>"0001111000101011"&"0010000111000001",
  5=>"0011001110001101"&"0010001101100000",
  6=>"0001010111000111"&"0010010101110101",
  7=>"0000110001001111"&"0010010111010101",
  8=>"0000101101000010"&"0010010110000101",
  9=>"0001011111010001"&"0010010101001000",
  10=>"0001000000001100"&"0010001010110000",
  11=>"0001101110100010"&"0001111101010111",
  12=>"0001010001001111"&"0010011001111100",
  13=>"0000010100101001"&"0010011000111100",
  14=>"0001101011100001"&"0010001101100011",
  15=>"0010001001100111"&"0001110001101010",
  16=>"0010011100101011"&"0010011010011000",
  17=>"0001110100110101"&"0010001010010110",
  18=>"0000000101010010"&"0010001111000010",
  19=>"0000101001100110"&"0010010000110001",
  20=>"0000111110011011"&"0010011110011000",
  21=>"0001010110100100"&"0010001101110010",
  22=>"0001000111100111"&"0010011011011100",
  23=>"0010000111001010"&"0001111010111001",
  24=>"0001010001100001"&"0010010010111110",
  25=>"0001010101010101"&"0010001110101001",
  26=>"0000111011001011"&"0010000010101001",
  27=>"0001001001111001"&"0010001000001001",
  28=>"0010000001110001"&"0010010010011111",
  29=>"0010001000001110"&"0010001011111010",
  30=>"0000101111001000"&"0010001000010110",
  31=>"1111111101011001"&"0010011101111111",
  32=>"0000101001101100"&"0010011101110111",
  33=>"0000110110010010"&"0010010001110011",
  34=>"0001100111000000"&"0010010100111011",
  35=>"0001010001110101"&"0010010111100110",
  36=>"0001011101010110"&"0010011100101100",
  37=>"0001000101000001"&"0010000001101000",
  38=>"0000111111011011"&"0010000110101010",
  39=>"0010011111001101"&"0010000110010001",
  40=>"0001101101001010"&"0010001000000110",
  41=>"0001001110001101"&"0010010110110111",
  42=>"0010000011010010"&"0010000111100011",
  43=>"0011011001000011"&"0010001010110111",
  44=>"0000111110110100"&"0010011110101010",
  45=>"0001000110011001"&"0010011101001100",
  46=>"0001110100010010"&"0010000111101010",
  47=>"0000011000000101"&"0010000011010110",
  48=>"0010001111101110"&"0010010010001011",
  49=>"0010000010100101"&"0010000000001001",
  50=>"0010010110011111"&"0010010000001111",
  51=>"0000010000111100"&"0010001111011111",
  52=>"0000111000100101"&"0001111100111001",
  53=>"0000010100111100"&"0010001011001111",
  54=>"0001111011011000"&"0010011010111110",
  55=>"0000000110100100"&"0010001101001010",
  56=>"0000010111101010"&"0010011011100110",
  57=>"0010110111101110"&"0010000101101100",
  58=>"0010001111000001"&"0010010000000000",
  59=>"1111111010010110"&"0010001000111000",
  60=>"0001011101001011"&"0010000110111100",
  61=>"0000100010111010"&"0001110011110010",
  62=>"0001111110100001"&"0001111001001111",
  63=>"0000100101100011"&"0010001010110001");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;