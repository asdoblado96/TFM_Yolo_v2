LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L4_2_BNROM IS
    PORT (
        coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        address : IN unsigned(5 DOWNTO 0));
END L4_2_BNROM;

ARCHITECTURE RTL OF L4_2_BNROM IS

    TYPE ROM_mem IS ARRAY (0 TO 63) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

    CONSTANT ROM_content : ROM_mem :=
    (0=>"0000001010001111"&"0000111001100111",
    1=>"1111100011111101"&"0001011100001001",
    2=>"1111111000010011"&"0001001110100111",
    3=>"1110101001100011"&"0001101101110110",
    4=>"1111101111011111"&"0001010011011011",
    5=>"0000000001110100"&"0001100001110011",
    6=>"1110001100101110"&"0001101000011001",
    7=>"0000010101110111"&"0001000110011001",
    8=>"0000011001111010"&"0000110111001110",
    9=>"0000011011011001"&"0000111100111111",
    10=>"1111111010110000"&"0001000111101001",
    11=>"1101111001001011"&"0000101110110111",
    12=>"0000010101110110"&"0001001001110100",
    13=>"1111111010100100"&"0000110111101110",
    14=>"1111011100011100"&"0001001001100100",
    15=>"0000110111101100"&"0000111000001101",
    16=>"1111111001110110"&"0001001111110001",
    17=>"0000100101011111"&"0001010100101000",
    18=>"1111000100100101"&"0000110011000111",
    19=>"1111101101001001"&"0001010000110111",
    20=>"0000010000001001"&"0001100010001100",
    21=>"0001110011011000"&"0001011111000011",
    22=>"1111100001111011"&"0001101011101000",
    23=>"1111001010111000"&"0010000001110010",
    24=>"0000010001101100"&"0001010111111010",
    25=>"1111101001000111"&"0001011010000111",
    26=>"1111100110100000"&"0001110001001110",
    27=>"1111101111001110"&"0001010001101010",
    28=>"0000000010011000"&"0001001001010101",
    29=>"0001010111111111"&"0001000011010101",
    30=>"0000101100110010"&"0001011000111100",
    31=>"1111010011010101"&"0001010110100110",
    32=>"1111101101011010"&"0001011000100010",
    33=>"1111000100100010"&"0001100100011110",
    34=>"0001010011000001"&"0000111100100001",
    35=>"0000101100100111"&"0000101111110010",
    36=>"0000001110011100"&"0001010111100101",
    37=>"1101100000101011"&"0001001000100100",
    38=>"1111100111100000"&"0001010110101100",
    39=>"1111100110000001"&"0001010100001000",
    40=>"0000111010111100"&"0001001011100000",
    41=>"0001010011111001"&"0001011001101100",
    42=>"0000011101010110"&"0001010110010100",
    43=>"0000010010010010"&"0001100000001100",
    44=>"0000011100101010"&"0001001000101100",
    45=>"1111001000100000"&"0001101011100010",
    46=>"1111110000111001"&"0001001101011111",
    47=>"0000010100001011"&"0001011011101100",
    48=>"0000101001001110"&"0000111010011010",
    49=>"1111100001101010"&"0001011010101111",
    50=>"0000010010101011"&"0000111011010111",
    51=>"0000100001111110"&"0000101101111100",
    52=>"1111100010110110"&"0001001101110001",
    53=>"1100101011010100"&"0001011010101101",
    54=>"0000000011111100"&"0001001110111000",
    55=>"1111111110110000"&"0001010111001111",
    56=>"0000000111111000"&"0001000001000100",
    57=>"0000011111010111"&"0001010011011011",
    58=>"0000111011010011"&"0001000111001010",
    59=>"0000101100110101"&"0000101101100000",
    60=>"1111111000111101"&"0001100110110101",
    61=>"0000100000100100"&"0001001101001110",
    62=>"0001000001010110"&"0001011001111110",
    63=>"0001010011111100"&"0001001101110100");
    
BEGIN
    coefs <= ROM_content(to_integer(address));
END RTL;