LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_10_BNROM IS
  PORT (
    coefs : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    address : IN unsigned(5 DOWNTO 0));
END L8_10_BNROM;

ARCHITECTURE RTL OF L8_10_BNROM IS

  TYPE ROM_mem IS ARRAY (0 TO 63) OF STD_LOGIC_VECTOR(31 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem :=

  --Contenido bias || scale
  (0=>"0010000011000110"&"0010001111011101",
  1=>"0000011111000001"&"0010001100011101",
  2=>"0010011001000010"&"0010001110000000",
  3=>"0010000101010111"&"0010001011010110",
  4=>"0001011101000111"&"0010001011001110",
  5=>"0000101010010010"&"0010010100110100",
  6=>"0000101000100011"&"0010010011010111",
  7=>"0001010001010110"&"0010011000010010",
  8=>"0001101100001111"&"0010011100011010",
  9=>"1101010101001011"&"0001001011111001",
  10=>"0000101000010011"&"0010001100000011",
  11=>"0000110101101111"&"0010011010100011",
  12=>"1101110000011010"&"0001110111111010",
  13=>"0001000110101010"&"0010010100100011",
  14=>"0001011111100001"&"0010010000110011",
  15=>"0000111110110010"&"0010010111001000",
  16=>"1110111001011010"&"0001110111111011",
  17=>"0001001111100100"&"0010010111010010",
  18=>"0001001111111110"&"0010000111101000",
  19=>"0001011010110101"&"0001110101101111",
  20=>"0001111110000000"&"0010001010000110",
  21=>"0001001101100101"&"0010000111111001",
  22=>"0010101110110111"&"0010001111100111",
  23=>"1110101011110001"&"0001101110000111",
  24=>"0000110110001111"&"0010011011110101",
  25=>"0010011010011100"&"0010010100011011",
  26=>"0010100111010001"&"0001111001101011",
  27=>"0000011010111001"&"0010010111101111",
  28=>"0000110101110001"&"0010011111001011",
  29=>"1110010101101100"&"0001010101101010",
  30=>"0000100100001010"&"0010011000010101",
  31=>"0000011101000101"&"0001110101001111",
  32=>"0000101101101110"&"0010001111001010",
  33=>"0001110001101111"&"0010010011001111",
  34=>"0001000100000001"&"0010001110100100",
  35=>"0000101100101100"&"0010100001110011",
  36=>"0010001111000001"&"0010010101111111",
  37=>"0001001110011011"&"0010001000110001",
  38=>"0010100101101100"&"0001101110111100",
  39=>"0001100001110001"&"0010010110000101",
  40=>"0001001001100000"&"0010010101000011",
  41=>"0001011000010001"&"0010010001000101",
  42=>"0001100110111011"&"0001101110110100",
  43=>"0001010011101101"&"0010010000011100",
  44=>"0010001111010001"&"0010001111100101",
  45=>"0001010111110000"&"0010010101001010",
  46=>"0001001010011011"&"0010010111101101",
  47=>"0000101100110001"&"0010100000100111",
  48=>"0010001010111000"&"0010010011101100",
  49=>"0001111110110110"&"0010000001111011",
  50=>"0001011011001000"&"0010000100110100",
  51=>"0000100101000011"&"0010000011011101",
  52=>"0001011101011010"&"0001101110110110",
  53=>"0000010011100110"&"0001111100000000",
  54=>"0000101011010100"&"0010001001001100",
  55=>"0000101111110111"&"0010011110110101",
  56=>"0001100010000000"&"0010001111101110",
  57=>"0000011110001111"&"0001110010111000",
  58=>"0010001101110011"&"0010010101110000",
  59=>"0001101000111110"&"0010001000001100",
  60=>"0010000111000010"&"0001110010100010",
  61=>"0011001110110110"&"0010001000100111",
  62=>"0000100001001110"&"0010011001000010",
  63=>"0000110010100000"&"0001111001010100");

BEGIN
  coefs <= ROM_content(to_integer(address));
END RTL;