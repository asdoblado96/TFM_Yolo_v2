LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_5_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(8)-1 DOWNTO 0));
END L8_5_WROM;

ARCHITECTURE RTL OF L8_5_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"100010111",
  1=>"110101000",
  2=>"010010111",
  3=>"010000110",
  4=>"111110101",
  5=>"111111001",
  6=>"001011111",
  7=>"101011100",
  8=>"100010010",
  9=>"111101000",
  10=>"111010100",
  11=>"111101010",
  12=>"100100010",
  13=>"011101011",
  14=>"100010011",
  15=>"111011011",
  16=>"001101011",
  17=>"000111001",
  18=>"000101101",
  19=>"000011001",
  20=>"101010100",
  21=>"100011011",
  22=>"001110101",
  23=>"001010001",
  24=>"000010110",
  25=>"100000010",
  26=>"010000001",
  27=>"001011000",
  28=>"110001011",
  29=>"011011111",
  30=>"011010101",
  31=>"101101000",
  32=>"101111100",
  33=>"001110110",
  34=>"101111011",
  35=>"001010101",
  36=>"011010010",
  37=>"101000110",
  38=>"111111001",
  39=>"110111001",
  40=>"011100010",
  41=>"000001110",
  42=>"101111100",
  43=>"110111000",
  44=>"001100100",
  45=>"100001110",
  46=>"011000100",
  47=>"000110000",
  48=>"101011000",
  49=>"111010011",
  50=>"001010100",
  51=>"110001011",
  52=>"001000010",
  53=>"110101100",
  54=>"101100011",
  55=>"011101111",
  56=>"110011001",
  57=>"110000101",
  58=>"011010101",
  59=>"010010011",
  60=>"110110111",
  61=>"010001100",
  62=>"001101011",
  63=>"000001100",
  64=>"111101011",
  65=>"111001000",
  66=>"001111011",
  67=>"101101100",
  68=>"101000011",
  69=>"010100111",
  70=>"001100110",
  71=>"110000110",
  72=>"011001011",
  73=>"101101001",
  74=>"001011100",
  75=>"011101101",
  76=>"001101110",
  77=>"001001001",
  78=>"111101111",
  79=>"100001001",
  80=>"010000100",
  81=>"100000000",
  82=>"100110101",
  83=>"100000111",
  84=>"010011010",
  85=>"110111100",
  86=>"000010111",
  87=>"000101010",
  88=>"010011101",
  89=>"010000001",
  90=>"100001000",
  91=>"101111111",
  92=>"110010000",
  93=>"000100101",
  94=>"101000011",
  95=>"011010101",
  96=>"011100100",
  97=>"001110010",
  98=>"100000101",
  99=>"101101100",
  100=>"010010000",
  101=>"010110110",
  102=>"111111100",
  103=>"000001111",
  104=>"010000011",
  105=>"010001110",
  106=>"001001101",
  107=>"110010110",
  108=>"101000111",
  109=>"101000111",
  110=>"101000110",
  111=>"000000111",
  112=>"100001011",
  113=>"100000010",
  114=>"100010001",
  115=>"110110100",
  116=>"011000110",
  117=>"111110110",
  118=>"000000110",
  119=>"000100111",
  120=>"000110111",
  121=>"001110010",
  122=>"000110011",
  123=>"111100000",
  124=>"011000111",
  125=>"001101011",
  126=>"101111011",
  127=>"010111010",
  128=>"010010000",
  129=>"100101000",
  130=>"101111101",
  131=>"101011011",
  132=>"110000000",
  133=>"111011010",
  134=>"111110111",
  135=>"001110110",
  136=>"001101001",
  137=>"000000011",
  138=>"111001101",
  139=>"101000110",
  140=>"111111111",
  141=>"111100000",
  142=>"101111001",
  143=>"001110101",
  144=>"000000010",
  145=>"001111001",
  146=>"011001011",
  147=>"001110101",
  148=>"001001001",
  149=>"100110010",
  150=>"001100100",
  151=>"010011110",
  152=>"101101011",
  153=>"001011000",
  154=>"001000101",
  155=>"101110010",
  156=>"011111000",
  157=>"011011111",
  158=>"111101011",
  159=>"101100010",
  160=>"001100101",
  161=>"111010000",
  162=>"010000101",
  163=>"010101010",
  164=>"000010101",
  165=>"110110110",
  166=>"011000100",
  167=>"110101000",
  168=>"101000111",
  169=>"111111111",
  170=>"111001011",
  171=>"010100011",
  172=>"100011011",
  173=>"101100110",
  174=>"011101011",
  175=>"110000111",
  176=>"001011111",
  177=>"100100110",
  178=>"000110000",
  179=>"110100010",
  180=>"110110000",
  181=>"000110101",
  182=>"110001100",
  183=>"000101100",
  184=>"101011000",
  185=>"001110101",
  186=>"001100101",
  187=>"111111110",
  188=>"001011100",
  189=>"011101111",
  190=>"110101101",
  191=>"011111001",
  192=>"101000110",
  193=>"000011010",
  194=>"000110111",
  195=>"010111110",
  196=>"101000001",
  197=>"011010010",
  198=>"001010011",
  199=>"100100111",
  200=>"100011001",
  201=>"001000001",
  202=>"011000101",
  203=>"111100111",
  204=>"011000011",
  205=>"011001100",
  206=>"100000011",
  207=>"000111101",
  208=>"100001001",
  209=>"100011111",
  210=>"000101011",
  211=>"111000111",
  212=>"111010101",
  213=>"011111010",
  214=>"100011000",
  215=>"011101101",
  216=>"110110001",
  217=>"011001010",
  218=>"000000100",
  219=>"101011110",
  220=>"101001010",
  221=>"111000111",
  222=>"010100000",
  223=>"111011000",
  224=>"001100101",
  225=>"101000001",
  226=>"110100111",
  227=>"000000010",
  228=>"001001111",
  229=>"000011011",
  230=>"000001111",
  231=>"111000000",
  232=>"000010010",
  233=>"101110111",
  234=>"000000100",
  235=>"111011011",
  236=>"100110101",
  237=>"110010110",
  238=>"110110101",
  239=>"011101100",
  240=>"011110110",
  241=>"000011010",
  242=>"101000100",
  243=>"101000001",
  244=>"110101111",
  245=>"110101000",
  246=>"101011100",
  247=>"000111000",
  248=>"011101011",
  249=>"101101001",
  250=>"101100001",
  251=>"011010111",
  252=>"001010110",
  253=>"100011011",
  254=>"111010010",
  255=>"110100000",
  256=>"101111001",
  257=>"101000000",
  258=>"110110110",
  259=>"011001000",
  260=>"010110100",
  261=>"011101100",
  262=>"011001101",
  263=>"111111000",
  264=>"001100011",
  265=>"110010000",
  266=>"101010111",
  267=>"000110001",
  268=>"110010000",
  269=>"001111000",
  270=>"110101001",
  271=>"000001110",
  272=>"110000010",
  273=>"100100011",
  274=>"011000110",
  275=>"001101101",
  276=>"010010111",
  277=>"100100011",
  278=>"010111001",
  279=>"000111111",
  280=>"010010001",
  281=>"111010000",
  282=>"001001010",
  283=>"010101000",
  284=>"110101011",
  285=>"000111011",
  286=>"010000001",
  287=>"101011111",
  288=>"011111100",
  289=>"010111010",
  290=>"100111001",
  291=>"110111000",
  292=>"011110111",
  293=>"111111011",
  294=>"101100101",
  295=>"001111100",
  296=>"111101100",
  297=>"100001011",
  298=>"111010011",
  299=>"100001000",
  300=>"111001011",
  301=>"110100010",
  302=>"101101100",
  303=>"110011100",
  304=>"111001001",
  305=>"000100011",
  306=>"001000001",
  307=>"010001010",
  308=>"110101010",
  309=>"111000000",
  310=>"100011100",
  311=>"111000000",
  312=>"000010000",
  313=>"011001110",
  314=>"101110010",
  315=>"100010110",
  316=>"011000100",
  317=>"110000100",
  318=>"100001110",
  319=>"010100100",
  320=>"011111100",
  321=>"010111111",
  322=>"010100100",
  323=>"010001011",
  324=>"101101011",
  325=>"101011010",
  326=>"110110100",
  327=>"101100000",
  328=>"100010000",
  329=>"001000111",
  330=>"110110101",
  331=>"111010000",
  332=>"110011001",
  333=>"011000000",
  334=>"110010001",
  335=>"000001010",
  336=>"111100011",
  337=>"100110101",
  338=>"101110111",
  339=>"001000111",
  340=>"000010010",
  341=>"000000010",
  342=>"000000101",
  343=>"011001101",
  344=>"000011011",
  345=>"000100000",
  346=>"101000010",
  347=>"110000111",
  348=>"001010011",
  349=>"010100111",
  350=>"110011101",
  351=>"010000110",
  352=>"011101100",
  353=>"101001101",
  354=>"011011000",
  355=>"011000001",
  356=>"101010100",
  357=>"101011100",
  358=>"001101010",
  359=>"111111010",
  360=>"111000101",
  361=>"000100010",
  362=>"101101111",
  363=>"100011010",
  364=>"000010000",
  365=>"010100100",
  366=>"000100111",
  367=>"010001101",
  368=>"001000001",
  369=>"100011001",
  370=>"011000110",
  371=>"110001011",
  372=>"110111110",
  373=>"000010010",
  374=>"100111111",
  375=>"010110001",
  376=>"000111100",
  377=>"100010110",
  378=>"110110111",
  379=>"010110000",
  380=>"100001001",
  381=>"100111110",
  382=>"110010101",
  383=>"110000100",
  384=>"011100011",
  385=>"100001110",
  386=>"000101100",
  387=>"110010010",
  388=>"011010000",
  389=>"000000001",
  390=>"001001101",
  391=>"101100100",
  392=>"111000100",
  393=>"001111111",
  394=>"100010101",
  395=>"000011010",
  396=>"000101000",
  397=>"100110110",
  398=>"011110110",
  399=>"100101010",
  400=>"110011010",
  401=>"111001011",
  402=>"010000101",
  403=>"000000110",
  404=>"010011001",
  405=>"000101010",
  406=>"100001001",
  407=>"100010010",
  408=>"100001100",
  409=>"101000001",
  410=>"011011010",
  411=>"100001101",
  412=>"010011011",
  413=>"010100001",
  414=>"011110010",
  415=>"100100111",
  416=>"110100111",
  417=>"111011010",
  418=>"001000110",
  419=>"111000110",
  420=>"010100110",
  421=>"001110100",
  422=>"110100111",
  423=>"011111010",
  424=>"011001010",
  425=>"000100010",
  426=>"010101010",
  427=>"001000010",
  428=>"100000000",
  429=>"110010000",
  430=>"110000111",
  431=>"011111010",
  432=>"101010110",
  433=>"111111011",
  434=>"111100001",
  435=>"101001001",
  436=>"110100101",
  437=>"001010100",
  438=>"001001010",
  439=>"111001101",
  440=>"010001101",
  441=>"011111001",
  442=>"000010001",
  443=>"001111111",
  444=>"100011100",
  445=>"000011110",
  446=>"111000000",
  447=>"111000101",
  448=>"000110011",
  449=>"101000010",
  450=>"010100010",
  451=>"111110101",
  452=>"011010010",
  453=>"110101111",
  454=>"100001010",
  455=>"110001000",
  456=>"111001011",
  457=>"010110101",
  458=>"101110110",
  459=>"101111110",
  460=>"011001011",
  461=>"100001111",
  462=>"010010001",
  463=>"101010110",
  464=>"101011111",
  465=>"100010100",
  466=>"000001100",
  467=>"100010010",
  468=>"010000011",
  469=>"011011101",
  470=>"010110111",
  471=>"111011110",
  472=>"100001010",
  473=>"100110101",
  474=>"101101110",
  475=>"001110111",
  476=>"000001100",
  477=>"001100001",
  478=>"111100110",
  479=>"100011101",
  480=>"001100010",
  481=>"100000000",
  482=>"001010101",
  483=>"111000010",
  484=>"000000101",
  485=>"011010001",
  486=>"000010100",
  487=>"100000010",
  488=>"111111111",
  489=>"101101101",
  490=>"001101100",
  491=>"000111111",
  492=>"000101111",
  493=>"000010110",
  494=>"111110110",
  495=>"100001101",
  496=>"010111111",
  497=>"010101001",
  498=>"101110001",
  499=>"011110011",
  500=>"011001111",
  501=>"110100000",
  502=>"000101001",
  503=>"111111011",
  504=>"110100111",
  505=>"010011011",
  506=>"000101110",
  507=>"000111011",
  508=>"000100010",
  509=>"101100100",
  510=>"100110010",
  511=>"011100001",
  512=>"001001001",
  513=>"101111110",
  514=>"101101111",
  515=>"100101111",
  516=>"010010010",
  517=>"100000100",
  518=>"111111100",
  519=>"011100000",
  520=>"011100100",
  521=>"100010001",
  522=>"111011111",
  523=>"000010010",
  524=>"001100011",
  525=>"000000110",
  526=>"101000011",
  527=>"010111001",
  528=>"011001100",
  529=>"101110111",
  530=>"111011100",
  531=>"000011010",
  532=>"000010000",
  533=>"101110101",
  534=>"011011111",
  535=>"100111001",
  536=>"010110010",
  537=>"010100111",
  538=>"101010110",
  539=>"111000111",
  540=>"110100010",
  541=>"010011001",
  542=>"010000100",
  543=>"001011011",
  544=>"100001001",
  545=>"110011100",
  546=>"001101101",
  547=>"001111001",
  548=>"010011011",
  549=>"111000001",
  550=>"110110010",
  551=>"110101000",
  552=>"100101101",
  553=>"101101100",
  554=>"000001001",
  555=>"001000010",
  556=>"011000011",
  557=>"101010011",
  558=>"101100111",
  559=>"000111110",
  560=>"110111011",
  561=>"110011110",
  562=>"110110101",
  563=>"101000010",
  564=>"101011110",
  565=>"111100111",
  566=>"011110110",
  567=>"010010011",
  568=>"101110101",
  569=>"101101000",
  570=>"011111100",
  571=>"001110010",
  572=>"000011101",
  573=>"001011011",
  574=>"101111111",
  575=>"111100101",
  576=>"001010101",
  577=>"100100111",
  578=>"110001010",
  579=>"001110001",
  580=>"101010110",
  581=>"100111100",
  582=>"101110110",
  583=>"001111101",
  584=>"100101111",
  585=>"101100111",
  586=>"111011011",
  587=>"100100010",
  588=>"110101001",
  589=>"101100000",
  590=>"011100100",
  591=>"000011101",
  592=>"110110000",
  593=>"111111110",
  594=>"000010000",
  595=>"111101100",
  596=>"011000101",
  597=>"010001101",
  598=>"111011001",
  599=>"101000111",
  600=>"101111001",
  601=>"010101010",
  602=>"101100001",
  603=>"000000110",
  604=>"100001110",
  605=>"000010000",
  606=>"001001011",
  607=>"111101011",
  608=>"101111100",
  609=>"011000111",
  610=>"010000100",
  611=>"000010111",
  612=>"010011110",
  613=>"011000100",
  614=>"100000010",
  615=>"110101100",
  616=>"010100110",
  617=>"001101110",
  618=>"011101111",
  619=>"001100101",
  620=>"101010111",
  621=>"001111101",
  622=>"000100001",
  623=>"110110000",
  624=>"100011000",
  625=>"001001110",
  626=>"100101110",
  627=>"001011100",
  628=>"001111101",
  629=>"101000110",
  630=>"111000101",
  631=>"111100000",
  632=>"101101111",
  633=>"101100111",
  634=>"101111110",
  635=>"110111011",
  636=>"000100011",
  637=>"111000110",
  638=>"111100100",
  639=>"111110100",
  640=>"010101100",
  641=>"100111000",
  642=>"111010001",
  643=>"000000000",
  644=>"101000001",
  645=>"001010110",
  646=>"010000010",
  647=>"010111111",
  648=>"001111110",
  649=>"110100001",
  650=>"100110010",
  651=>"110110111",
  652=>"001011111",
  653=>"111000000",
  654=>"110101100",
  655=>"011010000",
  656=>"011000010",
  657=>"001110111",
  658=>"011110000",
  659=>"100110101",
  660=>"000000000",
  661=>"011110100",
  662=>"110101000",
  663=>"010111000",
  664=>"100111011",
  665=>"101101000",
  666=>"100010111",
  667=>"010001010",
  668=>"011000010",
  669=>"010011110",
  670=>"100101011",
  671=>"101100111",
  672=>"100000111",
  673=>"111111100",
  674=>"101111011",
  675=>"000101000",
  676=>"111001100",
  677=>"100110000",
  678=>"001100101",
  679=>"011000001",
  680=>"101011011",
  681=>"111010111",
  682=>"000111101",
  683=>"111011010",
  684=>"011110011",
  685=>"000010111",
  686=>"010001000",
  687=>"111011101",
  688=>"010011111",
  689=>"111010111",
  690=>"001110110",
  691=>"010100011",
  692=>"101110001",
  693=>"101001001",
  694=>"111101111",
  695=>"010110000",
  696=>"011010011",
  697=>"111100000",
  698=>"100100000",
  699=>"100010000",
  700=>"101001110",
  701=>"100001001",
  702=>"100000010",
  703=>"010001001",
  704=>"000101000",
  705=>"110100111",
  706=>"010110101",
  707=>"111111011",
  708=>"110011010",
  709=>"101011101",
  710=>"101010100",
  711=>"101100001",
  712=>"000010000",
  713=>"010100001",
  714=>"101100000",
  715=>"100001001",
  716=>"110110000",
  717=>"011001010",
  718=>"000011011",
  719=>"110011100",
  720=>"111010101",
  721=>"100111000",
  722=>"111011111",
  723=>"010001000",
  724=>"101000111",
  725=>"000011011",
  726=>"000100111",
  727=>"001110110",
  728=>"100100111",
  729=>"111001100",
  730=>"010000100",
  731=>"101111000",
  732=>"011111101",
  733=>"111011010",
  734=>"101111011",
  735=>"011001000",
  736=>"110100100",
  737=>"111010001",
  738=>"001100111",
  739=>"001100111",
  740=>"110001010",
  741=>"011001010",
  742=>"000010011",
  743=>"101000101",
  744=>"101011111",
  745=>"111110110",
  746=>"001100010",
  747=>"100111111",
  748=>"010010000",
  749=>"010000010",
  750=>"011010100",
  751=>"000111000",
  752=>"101001011",
  753=>"101100111",
  754=>"000010000",
  755=>"000110101",
  756=>"101011110",
  757=>"001100011",
  758=>"001001111",
  759=>"101110011",
  760=>"010011010",
  761=>"110111010",
  762=>"011111100",
  763=>"111101111",
  764=>"110110001",
  765=>"111110111",
  766=>"000011001",
  767=>"000100110",
  768=>"010111011",
  769=>"100000011",
  770=>"000000111",
  771=>"101011000",
  772=>"010111111",
  773=>"100100000",
  774=>"111010110",
  775=>"101111001",
  776=>"001001010",
  777=>"010000011",
  778=>"111011110",
  779=>"011001101",
  780=>"111111000",
  781=>"011011111",
  782=>"100001111",
  783=>"000000011",
  784=>"110101000",
  785=>"010000001",
  786=>"000011011",
  787=>"001011101",
  788=>"111111000",
  789=>"010011000",
  790=>"010010000",
  791=>"111100000",
  792=>"011010101",
  793=>"110011100",
  794=>"001111111",
  795=>"010101011",
  796=>"001000000",
  797=>"100001111",
  798=>"100110100",
  799=>"100011110",
  800=>"010001111",
  801=>"000100111",
  802=>"111101100",
  803=>"111111111",
  804=>"000011101",
  805=>"110111100",
  806=>"111101100",
  807=>"001011010",
  808=>"000100001",
  809=>"000011100",
  810=>"101111011",
  811=>"100001011",
  812=>"000101100",
  813=>"101010101",
  814=>"100000001",
  815=>"000011011",
  816=>"110000011",
  817=>"001111011",
  818=>"101110111",
  819=>"011010001",
  820=>"001100101",
  821=>"111010011",
  822=>"110100000",
  823=>"000100101",
  824=>"111111010",
  825=>"001011111",
  826=>"110110001",
  827=>"100010001",
  828=>"110101100",
  829=>"111011110",
  830=>"111101000",
  831=>"011011101",
  832=>"001111001",
  833=>"010010011",
  834=>"111000001",
  835=>"110010001",
  836=>"011110001",
  837=>"100100100",
  838=>"000101100",
  839=>"011110110",
  840=>"111111001",
  841=>"000101101",
  842=>"000101010",
  843=>"100001100",
  844=>"111101011",
  845=>"100110110",
  846=>"100101010",
  847=>"100000100",
  848=>"110001101",
  849=>"110100100",
  850=>"001100011",
  851=>"011000110",
  852=>"101110111",
  853=>"100001110",
  854=>"111000011",
  855=>"011011011",
  856=>"110011111",
  857=>"011010110",
  858=>"010001111",
  859=>"010100001",
  860=>"111110001",
  861=>"110010010",
  862=>"001111011",
  863=>"011010111",
  864=>"110010011",
  865=>"111000001",
  866=>"001010010",
  867=>"100000110",
  868=>"100100001",
  869=>"010001100",
  870=>"000000101",
  871=>"010011001",
  872=>"111000000",
  873=>"001101110",
  874=>"000101010",
  875=>"010100011",
  876=>"110010101",
  877=>"111110111",
  878=>"010110000",
  879=>"110011110",
  880=>"000111111",
  881=>"101011110",
  882=>"110010101",
  883=>"110011011",
  884=>"000001111",
  885=>"000100101",
  886=>"010111011",
  887=>"001001110",
  888=>"011101010",
  889=>"000010010",
  890=>"110001100",
  891=>"111100011",
  892=>"010000100",
  893=>"111100111",
  894=>"000011001",
  895=>"111111100",
  896=>"010100011",
  897=>"110001111",
  898=>"011000000",
  899=>"000010100",
  900=>"000010100",
  901=>"111101101",
  902=>"011011000",
  903=>"010100000",
  904=>"000110110",
  905=>"000110011",
  906=>"001111111",
  907=>"010100010",
  908=>"000010100",
  909=>"110100110",
  910=>"001101111",
  911=>"011110101",
  912=>"110110100",
  913=>"000011101",
  914=>"001000011",
  915=>"001010000",
  916=>"001101101",
  917=>"111110101",
  918=>"000010111",
  919=>"000000001",
  920=>"110101110",
  921=>"101111010",
  922=>"000010001",
  923=>"101100101",
  924=>"010101000",
  925=>"110011101",
  926=>"110111000",
  927=>"110001110",
  928=>"010111101",
  929=>"111110001",
  930=>"100000010",
  931=>"001011100",
  932=>"000000011",
  933=>"111110111",
  934=>"100001110",
  935=>"101001101",
  936=>"111101100",
  937=>"110010101",
  938=>"010111011",
  939=>"000101110",
  940=>"010100010",
  941=>"100010111",
  942=>"010110111",
  943=>"001110010",
  944=>"000011101",
  945=>"110111101",
  946=>"000101001",
  947=>"001111011",
  948=>"011100111",
  949=>"110010111",
  950=>"111010111",
  951=>"101000111",
  952=>"011100010",
  953=>"001110100",
  954=>"100010000",
  955=>"111011011",
  956=>"010001111",
  957=>"010010000",
  958=>"000010001",
  959=>"101110001",
  960=>"000100101",
  961=>"011000010",
  962=>"001011011",
  963=>"101001100",
  964=>"100100010",
  965=>"011100001",
  966=>"001101000",
  967=>"010111000",
  968=>"000110100",
  969=>"111110011",
  970=>"001111101",
  971=>"001111100",
  972=>"111010000",
  973=>"011000011",
  974=>"100010110",
  975=>"101001111",
  976=>"010101001",
  977=>"011010111",
  978=>"010011110",
  979=>"001000011",
  980=>"010101110",
  981=>"100101010",
  982=>"001011011",
  983=>"110110010",
  984=>"110000001",
  985=>"110001011",
  986=>"100000010",
  987=>"010111111",
  988=>"101111101",
  989=>"100010100",
  990=>"000010101",
  991=>"101001111",
  992=>"011000101",
  993=>"100000110",
  994=>"101111010",
  995=>"011001110",
  996=>"000100111",
  997=>"001011001",
  998=>"111111000",
  999=>"011110111",
  1000=>"010000110",
  1001=>"000000010",
  1002=>"000000010",
  1003=>"111011001",
  1004=>"111101010",
  1005=>"000111111",
  1006=>"101110111",
  1007=>"001011010",
  1008=>"000000101",
  1009=>"111011100",
  1010=>"110101111",
  1011=>"110110101",
  1012=>"011001110",
  1013=>"010010011",
  1014=>"010101111",
  1015=>"111111000",
  1016=>"111100010",
  1017=>"101000010",
  1018=>"001000110",
  1019=>"000110011",
  1020=>"110001100",
  1021=>"011000101",
  1022=>"001011111",
  1023=>"100010111",
  1024=>"010100001",
  1025=>"100100001",
  1026=>"001011101",
  1027=>"101011101",
  1028=>"110100100",
  1029=>"010100010",
  1030=>"001111000",
  1031=>"111110100",
  1032=>"100000101",
  1033=>"010000010",
  1034=>"000100011",
  1035=>"110100011",
  1036=>"100010010",
  1037=>"100000011",
  1038=>"100000101",
  1039=>"100100111",
  1040=>"110011011",
  1041=>"101000100",
  1042=>"111010001",
  1043=>"110010110",
  1044=>"010100011",
  1045=>"000100001",
  1046=>"111111011",
  1047=>"010010011",
  1048=>"101110010",
  1049=>"001001100",
  1050=>"101000110",
  1051=>"101100010",
  1052=>"011100001",
  1053=>"101111100",
  1054=>"010110110",
  1055=>"111101110",
  1056=>"100010010",
  1057=>"011100111",
  1058=>"101110110",
  1059=>"100100110",
  1060=>"010101010",
  1061=>"101010110",
  1062=>"101000110",
  1063=>"111101101",
  1064=>"100111101",
  1065=>"010001000",
  1066=>"011001100",
  1067=>"000010110",
  1068=>"000000111",
  1069=>"100101100",
  1070=>"000110100",
  1071=>"011001110",
  1072=>"110110101",
  1073=>"010110110",
  1074=>"110010000",
  1075=>"111110111",
  1076=>"101011000",
  1077=>"110111111",
  1078=>"010110011",
  1079=>"011101110",
  1080=>"000000101",
  1081=>"011010111",
  1082=>"110110011",
  1083=>"000111000",
  1084=>"101010100",
  1085=>"010111111",
  1086=>"011100010",
  1087=>"001000101",
  1088=>"100101111",
  1089=>"110110011",
  1090=>"110111101",
  1091=>"100110111",
  1092=>"111000110",
  1093=>"101111010",
  1094=>"001111100",
  1095=>"000111100",
  1096=>"111000011",
  1097=>"100011101",
  1098=>"000110010",
  1099=>"000001000",
  1100=>"010001101",
  1101=>"101000100",
  1102=>"001011110",
  1103=>"000111100",
  1104=>"100010001",
  1105=>"011110001",
  1106=>"011011101",
  1107=>"101001000",
  1108=>"100110100",
  1109=>"100011101",
  1110=>"110010110",
  1111=>"101001101",
  1112=>"111000011",
  1113=>"011101101",
  1114=>"001100100",
  1115=>"010010100",
  1116=>"100111111",
  1117=>"111110010",
  1118=>"001001111",
  1119=>"001010111",
  1120=>"101010100",
  1121=>"000100000",
  1122=>"000001110",
  1123=>"101101001",
  1124=>"100000011",
  1125=>"110000110",
  1126=>"111100100",
  1127=>"101111111",
  1128=>"100111101",
  1129=>"101110111",
  1130=>"100110011",
  1131=>"001100011",
  1132=>"000101011",
  1133=>"000100000",
  1134=>"000000001",
  1135=>"010010111",
  1136=>"010100000",
  1137=>"101001110",
  1138=>"100010110",
  1139=>"011111100",
  1140=>"100001100",
  1141=>"011010000",
  1142=>"000101001",
  1143=>"010011100",
  1144=>"011000000",
  1145=>"111101010",
  1146=>"010000000",
  1147=>"000010100",
  1148=>"001100000",
  1149=>"000110000",
  1150=>"001001010",
  1151=>"111101111",
  1152=>"101010010",
  1153=>"010111011",
  1154=>"011101101",
  1155=>"001110101",
  1156=>"001010100",
  1157=>"011010110",
  1158=>"101110111",
  1159=>"100001000",
  1160=>"111111000",
  1161=>"110101100",
  1162=>"111000011",
  1163=>"010111101",
  1164=>"000001101",
  1165=>"011110111",
  1166=>"101001100",
  1167=>"111111111",
  1168=>"001100111",
  1169=>"011111100",
  1170=>"010001111",
  1171=>"000111110",
  1172=>"010001100",
  1173=>"000010010",
  1174=>"010110010",
  1175=>"001000000",
  1176=>"111001110",
  1177=>"010001110",
  1178=>"111111100",
  1179=>"100100110",
  1180=>"001001110",
  1181=>"001101101",
  1182=>"110111000",
  1183=>"010101110",
  1184=>"100010110",
  1185=>"111100000",
  1186=>"011001101",
  1187=>"100011011",
  1188=>"111010101",
  1189=>"100101010",
  1190=>"110000100",
  1191=>"010000101",
  1192=>"100010110",
  1193=>"111100111",
  1194=>"010001000",
  1195=>"011011001",
  1196=>"001010001",
  1197=>"001000111",
  1198=>"100111111",
  1199=>"100000000",
  1200=>"010101010",
  1201=>"101011000",
  1202=>"000011100",
  1203=>"101001101",
  1204=>"100000100",
  1205=>"111000100",
  1206=>"100100100",
  1207=>"000111010",
  1208=>"010110101",
  1209=>"000010010",
  1210=>"001111000",
  1211=>"110011111",
  1212=>"000110010",
  1213=>"110101100",
  1214=>"100011011",
  1215=>"011011010",
  1216=>"000001000",
  1217=>"010010100",
  1218=>"100111011",
  1219=>"011101100",
  1220=>"101111010",
  1221=>"010010001",
  1222=>"011010100",
  1223=>"001011000",
  1224=>"110010101",
  1225=>"100110010",
  1226=>"011011010",
  1227=>"011010100",
  1228=>"100101111",
  1229=>"011000101",
  1230=>"111011100",
  1231=>"110010000",
  1232=>"010110100",
  1233=>"101110111",
  1234=>"011111100",
  1235=>"001110100",
  1236=>"110011110",
  1237=>"100111100",
  1238=>"011100011",
  1239=>"111111011",
  1240=>"111000101",
  1241=>"011001001",
  1242=>"000100101",
  1243=>"100100001",
  1244=>"011011100",
  1245=>"110101000",
  1246=>"010011101",
  1247=>"111111011",
  1248=>"011011000",
  1249=>"000100101",
  1250=>"000101101",
  1251=>"001101110",
  1252=>"000010111",
  1253=>"100111111",
  1254=>"010010101",
  1255=>"000101110",
  1256=>"001000010",
  1257=>"110101111",
  1258=>"000110011",
  1259=>"110010011",
  1260=>"100001000",
  1261=>"000111011",
  1262=>"010010001",
  1263=>"001100000",
  1264=>"101110010",
  1265=>"011011111",
  1266=>"010001011",
  1267=>"110111110",
  1268=>"101011111",
  1269=>"101000100",
  1270=>"110100101",
  1271=>"000010011",
  1272=>"110101010",
  1273=>"101000101",
  1274=>"111000010",
  1275=>"010111000",
  1276=>"111001100",
  1277=>"010100100",
  1278=>"001111010",
  1279=>"101001101",
  1280=>"100101001",
  1281=>"011100001",
  1282=>"001101100",
  1283=>"010100001",
  1284=>"001001001",
  1285=>"001011110",
  1286=>"000001100",
  1287=>"101101000",
  1288=>"110100011",
  1289=>"100111101",
  1290=>"011110001",
  1291=>"011111110",
  1292=>"100110000",
  1293=>"110101010",
  1294=>"101000011",
  1295=>"100011001",
  1296=>"111101111",
  1297=>"101001001",
  1298=>"101000101",
  1299=>"111001011",
  1300=>"111110000",
  1301=>"001010111",
  1302=>"101010011",
  1303=>"011011000",
  1304=>"101011010",
  1305=>"101011001",
  1306=>"100010000",
  1307=>"110000100",
  1308=>"000011001",
  1309=>"111101011",
  1310=>"100101110",
  1311=>"010001001",
  1312=>"001100001",
  1313=>"001100110",
  1314=>"100110010",
  1315=>"101100001",
  1316=>"110110111",
  1317=>"110101001",
  1318=>"000101111",
  1319=>"001100001",
  1320=>"011110011",
  1321=>"011010111",
  1322=>"001000100",
  1323=>"011010110",
  1324=>"101100010",
  1325=>"001000000",
  1326=>"001000110",
  1327=>"000000110",
  1328=>"001000111",
  1329=>"000111110",
  1330=>"010011101",
  1331=>"001100000",
  1332=>"110110100",
  1333=>"000101111",
  1334=>"000010011",
  1335=>"110101111",
  1336=>"000010110",
  1337=>"111011001",
  1338=>"100010100",
  1339=>"110010000",
  1340=>"010101010",
  1341=>"001111100",
  1342=>"001110101",
  1343=>"110010001",
  1344=>"110000100",
  1345=>"000010010",
  1346=>"000000000",
  1347=>"100000100",
  1348=>"010011111",
  1349=>"010011101",
  1350=>"001000110",
  1351=>"010010100",
  1352=>"111011010",
  1353=>"011101101",
  1354=>"000011101",
  1355=>"010010110",
  1356=>"001101001",
  1357=>"001101011",
  1358=>"011111000",
  1359=>"110111101",
  1360=>"010111111",
  1361=>"111011000",
  1362=>"010010000",
  1363=>"011101010",
  1364=>"010001011",
  1365=>"100000111",
  1366=>"100110111",
  1367=>"000111100",
  1368=>"101111000",
  1369=>"111010101",
  1370=>"110001101",
  1371=>"111110100",
  1372=>"110100111",
  1373=>"110110000",
  1374=>"110010000",
  1375=>"111100001",
  1376=>"001010011",
  1377=>"011110001",
  1378=>"010110001",
  1379=>"100110010",
  1380=>"101010100",
  1381=>"100011001",
  1382=>"010011001",
  1383=>"111111110",
  1384=>"010011100",
  1385=>"000001000",
  1386=>"011100000",
  1387=>"010001111",
  1388=>"001010110",
  1389=>"101110111",
  1390=>"001101111",
  1391=>"100001010",
  1392=>"110101110",
  1393=>"010100100",
  1394=>"111010111",
  1395=>"101110110",
  1396=>"000111010",
  1397=>"000110111",
  1398=>"101111010",
  1399=>"001010111",
  1400=>"111100101",
  1401=>"001110100",
  1402=>"011011000",
  1403=>"010001000",
  1404=>"011011111",
  1405=>"000011110",
  1406=>"111101110",
  1407=>"110101001",
  1408=>"001001001",
  1409=>"000110111",
  1410=>"000000010",
  1411=>"101110010",
  1412=>"011100001",
  1413=>"110011111",
  1414=>"111011001",
  1415=>"011110111",
  1416=>"111101100",
  1417=>"001111100",
  1418=>"001100001",
  1419=>"000000100",
  1420=>"001101001",
  1421=>"100100101",
  1422=>"101010110",
  1423=>"110100011",
  1424=>"011011010",
  1425=>"010000000",
  1426=>"001001011",
  1427=>"000010101",
  1428=>"110100110",
  1429=>"110001001",
  1430=>"000010100",
  1431=>"111011111",
  1432=>"001111101",
  1433=>"000001111",
  1434=>"001011010",
  1435=>"000111000",
  1436=>"101110000",
  1437=>"101001000",
  1438=>"100111000",
  1439=>"111110000",
  1440=>"000000101",
  1441=>"110100011",
  1442=>"110011101",
  1443=>"000101111",
  1444=>"010101100",
  1445=>"101100100",
  1446=>"100100110",
  1447=>"001011010",
  1448=>"110111001",
  1449=>"101101010",
  1450=>"101101100",
  1451=>"000011010",
  1452=>"110111001",
  1453=>"101111110",
  1454=>"101010010",
  1455=>"000000001",
  1456=>"110000100",
  1457=>"110100101",
  1458=>"111001111",
  1459=>"110000111",
  1460=>"001000111",
  1461=>"110001111",
  1462=>"001000111",
  1463=>"011111101",
  1464=>"011010001",
  1465=>"001010110",
  1466=>"000110011",
  1467=>"000110110",
  1468=>"100111010",
  1469=>"111110011",
  1470=>"001000011",
  1471=>"111111001",
  1472=>"110010010",
  1473=>"011011111",
  1474=>"001111110",
  1475=>"111010110",
  1476=>"110100100",
  1477=>"001001001",
  1478=>"010010111",
  1479=>"101100000",
  1480=>"111100111",
  1481=>"000010001",
  1482=>"010010110",
  1483=>"000100100",
  1484=>"010101100",
  1485=>"111101110",
  1486=>"110011011",
  1487=>"110011010",
  1488=>"100010110",
  1489=>"011001100",
  1490=>"010011011",
  1491=>"110110000",
  1492=>"000111100",
  1493=>"010010111",
  1494=>"111111010",
  1495=>"000111011",
  1496=>"001000100",
  1497=>"101110110",
  1498=>"011101110",
  1499=>"010010011",
  1500=>"101001001",
  1501=>"111110110",
  1502=>"100011101",
  1503=>"001001000",
  1504=>"010110010",
  1505=>"001101101",
  1506=>"111000100",
  1507=>"111100000",
  1508=>"111110000",
  1509=>"101011111",
  1510=>"010100001",
  1511=>"010100101",
  1512=>"010100100",
  1513=>"000001010",
  1514=>"111000001",
  1515=>"101111000",
  1516=>"011101110",
  1517=>"111011110",
  1518=>"010111100",
  1519=>"011110011",
  1520=>"000011110",
  1521=>"101111000",
  1522=>"111010100",
  1523=>"011111000",
  1524=>"110001000",
  1525=>"000100011",
  1526=>"101110010",
  1527=>"110010010",
  1528=>"001001011",
  1529=>"010001100",
  1530=>"011101110",
  1531=>"000100000",
  1532=>"011110101",
  1533=>"010001110",
  1534=>"001000100",
  1535=>"111011111",
  1536=>"011101010",
  1537=>"001000001",
  1538=>"110111000",
  1539=>"001101100",
  1540=>"111111101",
  1541=>"000000101",
  1542=>"000110111",
  1543=>"001000010",
  1544=>"000110000",
  1545=>"010001011",
  1546=>"100000010",
  1547=>"100100000",
  1548=>"000110010",
  1549=>"000110101",
  1550=>"011111100",
  1551=>"000000001",
  1552=>"001101111",
  1553=>"000110101",
  1554=>"011010011",
  1555=>"101111010",
  1556=>"100011110",
  1557=>"110001001",
  1558=>"011011101",
  1559=>"100110101",
  1560=>"110100110",
  1561=>"000000000",
  1562=>"000101101",
  1563=>"011001000",
  1564=>"010111000",
  1565=>"001000100",
  1566=>"110000001",
  1567=>"011111111",
  1568=>"011101111",
  1569=>"100110100",
  1570=>"001101111",
  1571=>"100010110",
  1572=>"101011011",
  1573=>"111110011",
  1574=>"000011010",
  1575=>"111011111",
  1576=>"110101000",
  1577=>"000011010",
  1578=>"000111000",
  1579=>"011111101",
  1580=>"001110001",
  1581=>"101011101",
  1582=>"111110100",
  1583=>"000011000",
  1584=>"010001000",
  1585=>"101011111",
  1586=>"000101101",
  1587=>"001100000",
  1588=>"010100000",
  1589=>"000111011",
  1590=>"100000001",
  1591=>"111011010",
  1592=>"111000000",
  1593=>"001001011",
  1594=>"011100100",
  1595=>"111001111",
  1596=>"001000100",
  1597=>"100010110",
  1598=>"011001100",
  1599=>"101001010",
  1600=>"001100011",
  1601=>"110011100",
  1602=>"010011011",
  1603=>"001010011",
  1604=>"010110011",
  1605=>"011011100",
  1606=>"010011100",
  1607=>"101001110",
  1608=>"100101111",
  1609=>"100001000",
  1610=>"010110000",
  1611=>"000000011",
  1612=>"010100100",
  1613=>"101100110",
  1614=>"000010010",
  1615=>"100001100",
  1616=>"101010100",
  1617=>"000000010",
  1618=>"100100111",
  1619=>"110111110",
  1620=>"111011010",
  1621=>"101011000",
  1622=>"110101101",
  1623=>"000101101",
  1624=>"111110000",
  1625=>"111100101",
  1626=>"100010101",
  1627=>"000011011",
  1628=>"001000001",
  1629=>"100100101",
  1630=>"001111101",
  1631=>"100010001",
  1632=>"000000000",
  1633=>"111101110",
  1634=>"110001110",
  1635=>"001110001",
  1636=>"000000111",
  1637=>"100000101",
  1638=>"011001100",
  1639=>"101011100",
  1640=>"010111011",
  1641=>"111011111",
  1642=>"010111100",
  1643=>"100000001",
  1644=>"111111101",
  1645=>"001010000",
  1646=>"100100000",
  1647=>"001000110",
  1648=>"100111101",
  1649=>"110100100",
  1650=>"101010000",
  1651=>"010011100",
  1652=>"111100111",
  1653=>"101000100",
  1654=>"000010100",
  1655=>"000011001",
  1656=>"111101111",
  1657=>"010111001",
  1658=>"111100110",
  1659=>"010001100",
  1660=>"111000111",
  1661=>"010001101",
  1662=>"001010101",
  1663=>"001111100",
  1664=>"011101100",
  1665=>"100100010",
  1666=>"001111111",
  1667=>"111110001",
  1668=>"000000101",
  1669=>"110011011",
  1670=>"100011110",
  1671=>"011011000",
  1672=>"010010111",
  1673=>"001000110",
  1674=>"001010110",
  1675=>"111100000",
  1676=>"001000110",
  1677=>"101100111",
  1678=>"101000001",
  1679=>"000110111",
  1680=>"111111110",
  1681=>"001001100",
  1682=>"000110011",
  1683=>"001000011",
  1684=>"001011100",
  1685=>"110110111",
  1686=>"010000010",
  1687=>"110011011",
  1688=>"110010010",
  1689=>"111011000",
  1690=>"101010000",
  1691=>"000110001",
  1692=>"000111101",
  1693=>"111101000",
  1694=>"110011000",
  1695=>"001011011",
  1696=>"101010100",
  1697=>"111100011",
  1698=>"110001100",
  1699=>"100000010",
  1700=>"011000101",
  1701=>"111100110",
  1702=>"011110010",
  1703=>"110001110",
  1704=>"010011100",
  1705=>"010100001",
  1706=>"001111111",
  1707=>"110101000",
  1708=>"000101010",
  1709=>"010000010",
  1710=>"100001101",
  1711=>"100110101",
  1712=>"110110111",
  1713=>"010011001",
  1714=>"011000000",
  1715=>"110010101",
  1716=>"001111100",
  1717=>"111110111",
  1718=>"111111110",
  1719=>"111110110",
  1720=>"000101010",
  1721=>"011101001",
  1722=>"110010110",
  1723=>"101100100",
  1724=>"100001000",
  1725=>"101000000",
  1726=>"100100001",
  1727=>"101111010",
  1728=>"110111001",
  1729=>"111011010",
  1730=>"010000100",
  1731=>"100101000",
  1732=>"101000000",
  1733=>"101000111",
  1734=>"110101101",
  1735=>"101011010",
  1736=>"010111100",
  1737=>"000011000",
  1738=>"110010000",
  1739=>"001001111",
  1740=>"011000010",
  1741=>"001101111",
  1742=>"011010000",
  1743=>"010100111",
  1744=>"110000000",
  1745=>"100011111",
  1746=>"101001000",
  1747=>"001001101",
  1748=>"101000001",
  1749=>"011011111",
  1750=>"111011101",
  1751=>"100111000",
  1752=>"010000001",
  1753=>"001101101",
  1754=>"001011101",
  1755=>"110110100",
  1756=>"011000100",
  1757=>"010011011",
  1758=>"001010011",
  1759=>"100010110",
  1760=>"110000100",
  1761=>"000111110",
  1762=>"000011010",
  1763=>"001000011",
  1764=>"001111010",
  1765=>"100010011",
  1766=>"101100100",
  1767=>"101000110",
  1768=>"001000010",
  1769=>"101111111",
  1770=>"100100101",
  1771=>"000011000",
  1772=>"000001011",
  1773=>"001000101",
  1774=>"010001111",
  1775=>"000011000",
  1776=>"010110110",
  1777=>"001011011",
  1778=>"100001011",
  1779=>"000101101",
  1780=>"110011000",
  1781=>"100000001",
  1782=>"011101011",
  1783=>"111101011",
  1784=>"111000010",
  1785=>"111110111",
  1786=>"010011000",
  1787=>"000101010",
  1788=>"001100000",
  1789=>"101010100",
  1790=>"110010010",
  1791=>"001011010",
  1792=>"110100100",
  1793=>"100011001",
  1794=>"111111101",
  1795=>"110011111",
  1796=>"010011111",
  1797=>"011000110",
  1798=>"000100101",
  1799=>"110000100",
  1800=>"010101001",
  1801=>"101010101",
  1802=>"001101001",
  1803=>"100101110",
  1804=>"000001100",
  1805=>"010111111",
  1806=>"010000011",
  1807=>"000010000",
  1808=>"000000110",
  1809=>"000011100",
  1810=>"000011101",
  1811=>"111010100",
  1812=>"010000010",
  1813=>"000001111",
  1814=>"101000000",
  1815=>"101100011",
  1816=>"111010101",
  1817=>"101011100",
  1818=>"000011111",
  1819=>"110001101",
  1820=>"010100101",
  1821=>"011001010",
  1822=>"100101100",
  1823=>"100000101",
  1824=>"011001001",
  1825=>"010111101",
  1826=>"111101011",
  1827=>"100001011",
  1828=>"001110001",
  1829=>"000001011",
  1830=>"101010101",
  1831=>"111110111",
  1832=>"011000001",
  1833=>"000001111",
  1834=>"000111100",
  1835=>"111001101",
  1836=>"110010011",
  1837=>"110010011",
  1838=>"000011011",
  1839=>"000001010",
  1840=>"110111000",
  1841=>"011011001",
  1842=>"010011010",
  1843=>"000010111",
  1844=>"010101100",
  1845=>"111000100",
  1846=>"101010000",
  1847=>"010001011",
  1848=>"010100010",
  1849=>"110100111",
  1850=>"111100111",
  1851=>"101100001",
  1852=>"011010101",
  1853=>"101010011",
  1854=>"101111010",
  1855=>"110111000",
  1856=>"101111011",
  1857=>"111010100",
  1858=>"111110100",
  1859=>"110000100",
  1860=>"001011001",
  1861=>"100110001",
  1862=>"101001000",
  1863=>"110010000",
  1864=>"111001110",
  1865=>"101001000",
  1866=>"110000011",
  1867=>"100010100",
  1868=>"100100010",
  1869=>"001000100",
  1870=>"101100000",
  1871=>"000010100",
  1872=>"011100010",
  1873=>"100101111",
  1874=>"100100010",
  1875=>"010010001",
  1876=>"011010001",
  1877=>"000101000",
  1878=>"010011110",
  1879=>"001000111",
  1880=>"000011001",
  1881=>"100011000",
  1882=>"000100010",
  1883=>"100000111",
  1884=>"110010010",
  1885=>"110010101",
  1886=>"100011100",
  1887=>"101101111",
  1888=>"000000101",
  1889=>"111110100",
  1890=>"011011000",
  1891=>"100000110",
  1892=>"000100110",
  1893=>"110010101",
  1894=>"000111100",
  1895=>"110101100",
  1896=>"111011111",
  1897=>"111100011",
  1898=>"011101101",
  1899=>"011001011",
  1900=>"100000100",
  1901=>"001100111",
  1902=>"001010001",
  1903=>"000000001",
  1904=>"001000001",
  1905=>"010100111",
  1906=>"101111111",
  1907=>"100000000",
  1908=>"101000001",
  1909=>"011111110",
  1910=>"110010000",
  1911=>"011100111",
  1912=>"010111110",
  1913=>"110011010",
  1914=>"101000100",
  1915=>"010111111",
  1916=>"110101101",
  1917=>"011101010",
  1918=>"000110010",
  1919=>"011000100",
  1920=>"100100101",
  1921=>"110111011",
  1922=>"111111111",
  1923=>"001111010",
  1924=>"000110010",
  1925=>"101011000",
  1926=>"001001011",
  1927=>"101100100",
  1928=>"001000011",
  1929=>"000101111",
  1930=>"111111010",
  1931=>"000011010",
  1932=>"000010001",
  1933=>"110100010",
  1934=>"101010111",
  1935=>"001111111",
  1936=>"111000101",
  1937=>"001001100",
  1938=>"101011000",
  1939=>"110010101",
  1940=>"011010111",
  1941=>"110010100",
  1942=>"000100101",
  1943=>"101111111",
  1944=>"101110001",
  1945=>"111101011",
  1946=>"000101101",
  1947=>"110011111",
  1948=>"111000000",
  1949=>"100101000",
  1950=>"000010011",
  1951=>"100101000",
  1952=>"100101000",
  1953=>"100011001",
  1954=>"000000000",
  1955=>"010101001",
  1956=>"111000001",
  1957=>"110011111",
  1958=>"101110001",
  1959=>"101100101",
  1960=>"011001101",
  1961=>"010110000",
  1962=>"100111110",
  1963=>"100010000",
  1964=>"011111111",
  1965=>"010000110",
  1966=>"111110111",
  1967=>"001000001",
  1968=>"000001111",
  1969=>"111100111",
  1970=>"011110101",
  1971=>"100010101",
  1972=>"101111011",
  1973=>"111010010",
  1974=>"001001001",
  1975=>"110010100",
  1976=>"011010110",
  1977=>"001010100",
  1978=>"111110010",
  1979=>"001110011",
  1980=>"001100010",
  1981=>"010100000",
  1982=>"111110001",
  1983=>"100100011",
  1984=>"000000101",
  1985=>"111000011",
  1986=>"000111000",
  1987=>"101101000",
  1988=>"000101100",
  1989=>"101100000",
  1990=>"001011100",
  1991=>"000110011",
  1992=>"001000000",
  1993=>"001000110",
  1994=>"000110011",
  1995=>"111001000",
  1996=>"110011000",
  1997=>"101011111",
  1998=>"111101011",
  1999=>"100011001",
  2000=>"001011100",
  2001=>"101000011",
  2002=>"110111110",
  2003=>"001000010",
  2004=>"110011001",
  2005=>"000000011",
  2006=>"011100001",
  2007=>"011001110",
  2008=>"100001000",
  2009=>"111011011",
  2010=>"100111010",
  2011=>"010010000",
  2012=>"001011001",
  2013=>"100010100",
  2014=>"010110110",
  2015=>"110010000",
  2016=>"000101111",
  2017=>"010100110",
  2018=>"101000000",
  2019=>"000011101",
  2020=>"101000000",
  2021=>"000100000",
  2022=>"100100111",
  2023=>"000010001",
  2024=>"111101101",
  2025=>"111111001",
  2026=>"001010010",
  2027=>"101011000",
  2028=>"101100101",
  2029=>"000010101",
  2030=>"001001110",
  2031=>"110111011",
  2032=>"101000111",
  2033=>"000001011",
  2034=>"111100001",
  2035=>"111001000",
  2036=>"011100000",
  2037=>"110111101",
  2038=>"010010110",
  2039=>"011100110",
  2040=>"111010001",
  2041=>"001101000",
  2042=>"100110110",
  2043=>"110010011",
  2044=>"111111101",
  2045=>"010010101",
  2046=>"000110100",
  2047=>"110001010",
  2048=>"110110000",
  2049=>"011010101",
  2050=>"100010110",
  2051=>"010111111",
  2052=>"110001010",
  2053=>"000011001",
  2054=>"111111000",
  2055=>"011001010",
  2056=>"111000101",
  2057=>"001110001",
  2058=>"111101100",
  2059=>"001101001",
  2060=>"101000011",
  2061=>"111111011",
  2062=>"100010100",
  2063=>"010010000",
  2064=>"100110001",
  2065=>"111001111",
  2066=>"011111011",
  2067=>"011100000",
  2068=>"000001111",
  2069=>"100010010",
  2070=>"000011101",
  2071=>"101110010",
  2072=>"010100001",
  2073=>"000001000",
  2074=>"111110000",
  2075=>"111000111",
  2076=>"111110000",
  2077=>"100000011",
  2078=>"111100000",
  2079=>"010001101",
  2080=>"101110100",
  2081=>"011000110",
  2082=>"001010101",
  2083=>"101111011",
  2084=>"010111101",
  2085=>"011111101",
  2086=>"000110000",
  2087=>"110011001",
  2088=>"101100010",
  2089=>"111111000",
  2090=>"001110110",
  2091=>"011010100",
  2092=>"010110011",
  2093=>"100000100",
  2094=>"011001000",
  2095=>"011100011",
  2096=>"011101000",
  2097=>"100101110",
  2098=>"110101111",
  2099=>"111100011",
  2100=>"001000110",
  2101=>"100111101",
  2102=>"111111101",
  2103=>"000101110",
  2104=>"101000001",
  2105=>"010100101",
  2106=>"001110010",
  2107=>"000000010",
  2108=>"100100101",
  2109=>"010101110",
  2110=>"000001110",
  2111=>"000000000",
  2112=>"000000000",
  2113=>"000100011",
  2114=>"111010100",
  2115=>"101111010",
  2116=>"001010011",
  2117=>"111111000",
  2118=>"011101001",
  2119=>"010010110",
  2120=>"001111001",
  2121=>"111001101",
  2122=>"100001010",
  2123=>"110010010",
  2124=>"001100000",
  2125=>"011011011",
  2126=>"101000000",
  2127=>"110110101",
  2128=>"001101000",
  2129=>"111110010",
  2130=>"111100101",
  2131=>"010100111",
  2132=>"010011000",
  2133=>"111101100",
  2134=>"110100010",
  2135=>"101111011",
  2136=>"111011001",
  2137=>"111111011",
  2138=>"101100100",
  2139=>"100001000",
  2140=>"101000000",
  2141=>"100111110",
  2142=>"100100111",
  2143=>"100000010",
  2144=>"010011111",
  2145=>"100111111",
  2146=>"010010001",
  2147=>"100010000",
  2148=>"011110010",
  2149=>"111111011",
  2150=>"101111011",
  2151=>"010110010",
  2152=>"111100100",
  2153=>"110000111",
  2154=>"111001111",
  2155=>"000110001",
  2156=>"101110010",
  2157=>"110111011",
  2158=>"011101000",
  2159=>"001001000",
  2160=>"000101100",
  2161=>"000110100",
  2162=>"111101110",
  2163=>"110010110",
  2164=>"100101000",
  2165=>"010100100",
  2166=>"111111111",
  2167=>"010011110",
  2168=>"101010111",
  2169=>"000011000",
  2170=>"110101011",
  2171=>"101101001",
  2172=>"100111100",
  2173=>"100011110",
  2174=>"000010100",
  2175=>"111010111",
  2176=>"001001011",
  2177=>"001000101",
  2178=>"100011111",
  2179=>"000011010",
  2180=>"110110011",
  2181=>"110100110",
  2182=>"101000101",
  2183=>"000110011",
  2184=>"111111101",
  2185=>"011001010",
  2186=>"111100011",
  2187=>"110010101",
  2188=>"101011000",
  2189=>"010101000",
  2190=>"100100111",
  2191=>"110011000",
  2192=>"110111100",
  2193=>"111000010",
  2194=>"111110101",
  2195=>"111000011",
  2196=>"000001110",
  2197=>"101010011",
  2198=>"111101101",
  2199=>"110101111",
  2200=>"100001100",
  2201=>"010110101",
  2202=>"110011100",
  2203=>"101000111",
  2204=>"110001000",
  2205=>"110010101",
  2206=>"010101011",
  2207=>"011110101",
  2208=>"101000110",
  2209=>"100000110",
  2210=>"101001101",
  2211=>"001100110",
  2212=>"010011101",
  2213=>"100010100",
  2214=>"101100010",
  2215=>"100011011",
  2216=>"100001100",
  2217=>"100000111",
  2218=>"100010001",
  2219=>"111001111",
  2220=>"010100000",
  2221=>"100010010",
  2222=>"110111111",
  2223=>"000010000",
  2224=>"101011001",
  2225=>"000101110",
  2226=>"000011110",
  2227=>"110001011",
  2228=>"011000111",
  2229=>"001011010",
  2230=>"111001101",
  2231=>"101110110",
  2232=>"001100011",
  2233=>"001100100",
  2234=>"001001011",
  2235=>"111111100",
  2236=>"000110001",
  2237=>"101111011",
  2238=>"001111010",
  2239=>"111111111",
  2240=>"110111110",
  2241=>"100011101",
  2242=>"000001010",
  2243=>"110011100",
  2244=>"000110000",
  2245=>"111011011",
  2246=>"101110100",
  2247=>"111101101",
  2248=>"111100000",
  2249=>"110101010",
  2250=>"110010001",
  2251=>"001110111",
  2252=>"111110011",
  2253=>"011111000",
  2254=>"110010000",
  2255=>"101000000",
  2256=>"101011011",
  2257=>"110101000",
  2258=>"010101111",
  2259=>"010100010",
  2260=>"010000010",
  2261=>"011001101",
  2262=>"110110101",
  2263=>"010000110",
  2264=>"001100000",
  2265=>"101010100",
  2266=>"000100100",
  2267=>"000000010",
  2268=>"101011110",
  2269=>"001010100",
  2270=>"001000010",
  2271=>"010110110",
  2272=>"100010001",
  2273=>"010000000",
  2274=>"000100110",
  2275=>"110111010",
  2276=>"100100110",
  2277=>"001001110",
  2278=>"010000001",
  2279=>"101011100",
  2280=>"101001110",
  2281=>"000111010",
  2282=>"111111011",
  2283=>"101101110",
  2284=>"001010111",
  2285=>"010101111",
  2286=>"111001000",
  2287=>"001001000",
  2288=>"010000001",
  2289=>"110110111",
  2290=>"000100111",
  2291=>"010100100",
  2292=>"111011110",
  2293=>"101000110",
  2294=>"100011110",
  2295=>"101100010",
  2296=>"110000110",
  2297=>"100010010",
  2298=>"000001010",
  2299=>"010101111",
  2300=>"101001000",
  2301=>"100111001",
  2302=>"000110111",
  2303=>"001001101",
  2304=>"110001010",
  2305=>"100001101",
  2306=>"110000111",
  2307=>"111100100",
  2308=>"101001100",
  2309=>"010010010",
  2310=>"110001110",
  2311=>"110101111",
  2312=>"000110001",
  2313=>"000100100",
  2314=>"100101000",
  2315=>"111100001",
  2316=>"001000010",
  2317=>"011101001",
  2318=>"101001001",
  2319=>"001111100",
  2320=>"000011010",
  2321=>"110111101",
  2322=>"001000100",
  2323=>"100101011",
  2324=>"111011101",
  2325=>"011000000",
  2326=>"010111000",
  2327=>"001101110",
  2328=>"000110100",
  2329=>"100010101",
  2330=>"100101100",
  2331=>"101100100",
  2332=>"000011110",
  2333=>"111100101",
  2334=>"011000100",
  2335=>"100001010",
  2336=>"001001101",
  2337=>"101011001",
  2338=>"010111110",
  2339=>"001000110",
  2340=>"011111100",
  2341=>"000010011",
  2342=>"001010001",
  2343=>"001110000",
  2344=>"100000000",
  2345=>"111101000",
  2346=>"111011000",
  2347=>"000000001",
  2348=>"000010000",
  2349=>"101111101",
  2350=>"001011000",
  2351=>"011111001",
  2352=>"010000000",
  2353=>"110010000",
  2354=>"111010110",
  2355=>"010000011",
  2356=>"011111101",
  2357=>"001101001",
  2358=>"010100001",
  2359=>"010100100",
  2360=>"110000000",
  2361=>"001111110",
  2362=>"010100111",
  2363=>"011001010",
  2364=>"100101110",
  2365=>"011011111",
  2366=>"101011011",
  2367=>"101101101",
  2368=>"011100100",
  2369=>"010011101",
  2370=>"100001111",
  2371=>"010000110",
  2372=>"111110101",
  2373=>"010100100",
  2374=>"000010000",
  2375=>"100111001",
  2376=>"111101111",
  2377=>"010000100",
  2378=>"010000101",
  2379=>"110110100",
  2380=>"010000111",
  2381=>"111011110",
  2382=>"111101110",
  2383=>"100010010",
  2384=>"100011000",
  2385=>"000001000",
  2386=>"011110011",
  2387=>"111111011",
  2388=>"101000010",
  2389=>"011000000",
  2390=>"100111010",
  2391=>"110110110",
  2392=>"011000001",
  2393=>"101100111",
  2394=>"110110111",
  2395=>"100010010",
  2396=>"001100101",
  2397=>"100110111",
  2398=>"111100010",
  2399=>"101100100",
  2400=>"110101111",
  2401=>"110000101",
  2402=>"001011010",
  2403=>"000100010",
  2404=>"000111100",
  2405=>"000001111",
  2406=>"010001100",
  2407=>"011110100",
  2408=>"110010111",
  2409=>"111001001",
  2410=>"010001000",
  2411=>"101110100",
  2412=>"100011111",
  2413=>"001001110",
  2414=>"111001010",
  2415=>"100111011",
  2416=>"110010001",
  2417=>"000000110",
  2418=>"001100110",
  2419=>"110011101",
  2420=>"111111001",
  2421=>"001111011",
  2422=>"101111011",
  2423=>"000101101",
  2424=>"001001101",
  2425=>"100000000",
  2426=>"000001001",
  2427=>"110000101",
  2428=>"101110010",
  2429=>"111101001",
  2430=>"111111110",
  2431=>"011101101",
  2432=>"001010110",
  2433=>"111111100",
  2434=>"001001101",
  2435=>"011001000",
  2436=>"100010001",
  2437=>"110000010",
  2438=>"010001110",
  2439=>"101000000",
  2440=>"000010011",
  2441=>"111000000",
  2442=>"110001001",
  2443=>"100111000",
  2444=>"000000110",
  2445=>"011111000",
  2446=>"111111100",
  2447=>"001011101",
  2448=>"000110101",
  2449=>"010100010",
  2450=>"100001011",
  2451=>"000011000",
  2452=>"100101110",
  2453=>"111011010",
  2454=>"011000011",
  2455=>"110101111",
  2456=>"000001000",
  2457=>"110000101",
  2458=>"000001100",
  2459=>"001110100",
  2460=>"101101001",
  2461=>"010100001",
  2462=>"101110011",
  2463=>"010100101",
  2464=>"001011011",
  2465=>"001100111",
  2466=>"100101110",
  2467=>"000101101",
  2468=>"110011010",
  2469=>"100000100",
  2470=>"000100000",
  2471=>"000111001",
  2472=>"110000001",
  2473=>"001111110",
  2474=>"000011110",
  2475=>"001010010",
  2476=>"011001010",
  2477=>"100111001",
  2478=>"111100110",
  2479=>"011111111",
  2480=>"100010000",
  2481=>"101101011",
  2482=>"110000001",
  2483=>"111101000",
  2484=>"100100000",
  2485=>"000000001",
  2486=>"001001101",
  2487=>"000110100",
  2488=>"000011011",
  2489=>"100111111",
  2490=>"001001001",
  2491=>"101001111",
  2492=>"101101101",
  2493=>"010000101",
  2494=>"100010010",
  2495=>"110001111",
  2496=>"111001001",
  2497=>"001011001",
  2498=>"100101010",
  2499=>"100101101",
  2500=>"011100111",
  2501=>"101010111",
  2502=>"110111001",
  2503=>"110101100",
  2504=>"111101110",
  2505=>"101001000",
  2506=>"001011010",
  2507=>"000010101",
  2508=>"010111100",
  2509=>"110000100",
  2510=>"110110010",
  2511=>"001111010",
  2512=>"010100100",
  2513=>"000100100",
  2514=>"001011101",
  2515=>"011000110",
  2516=>"111110000",
  2517=>"100000011",
  2518=>"000101011",
  2519=>"000111010",
  2520=>"111100100",
  2521=>"111010011",
  2522=>"110100000",
  2523=>"100001110",
  2524=>"010001010",
  2525=>"010100001",
  2526=>"100101001",
  2527=>"101000111",
  2528=>"010001100",
  2529=>"100111111",
  2530=>"111110101",
  2531=>"011101101",
  2532=>"000110000",
  2533=>"111101100",
  2534=>"101011000",
  2535=>"111110111",
  2536=>"011011001",
  2537=>"110011001",
  2538=>"001001011",
  2539=>"111000110",
  2540=>"100100100",
  2541=>"011001100",
  2542=>"110000000",
  2543=>"111111001",
  2544=>"100011011",
  2545=>"110000111",
  2546=>"000110011",
  2547=>"010011010",
  2548=>"000011100",
  2549=>"001010001",
  2550=>"110100011",
  2551=>"011101101",
  2552=>"100101010",
  2553=>"101001111",
  2554=>"010010101",
  2555=>"001010011",
  2556=>"000011101",
  2557=>"100100101",
  2558=>"000000010",
  2559=>"101111011",
  2560=>"011100000",
  2561=>"111101110",
  2562=>"000100010",
  2563=>"000001001",
  2564=>"011011001",
  2565=>"010010100",
  2566=>"100011011",
  2567=>"010100010",
  2568=>"011110000",
  2569=>"101001100",
  2570=>"100111101",
  2571=>"100010110",
  2572=>"011011100",
  2573=>"111101100",
  2574=>"100101000",
  2575=>"110011101",
  2576=>"111110001",
  2577=>"000001101",
  2578=>"011001011",
  2579=>"101011000",
  2580=>"011010101",
  2581=>"010100000",
  2582=>"100000010",
  2583=>"010000011",
  2584=>"000011000",
  2585=>"111001010",
  2586=>"111101110",
  2587=>"101100101",
  2588=>"100101110",
  2589=>"010110110",
  2590=>"000001100",
  2591=>"110010000",
  2592=>"110001010",
  2593=>"000011000",
  2594=>"111000101",
  2595=>"010010101",
  2596=>"111100001",
  2597=>"100001111",
  2598=>"111010111",
  2599=>"000110010",
  2600=>"001000010",
  2601=>"001101010",
  2602=>"100000000",
  2603=>"111001001",
  2604=>"111110000",
  2605=>"011000011",
  2606=>"100011111",
  2607=>"111101110",
  2608=>"101001101",
  2609=>"011111011",
  2610=>"110000000",
  2611=>"100001010",
  2612=>"101001000",
  2613=>"000100010",
  2614=>"010010111",
  2615=>"010101011",
  2616=>"110001001",
  2617=>"001100111",
  2618=>"011110001",
  2619=>"100100111",
  2620=>"110111111",
  2621=>"010010110",
  2622=>"000111010",
  2623=>"010100011",
  2624=>"110001101",
  2625=>"011011111",
  2626=>"111100000",
  2627=>"110011111",
  2628=>"010001001",
  2629=>"001110000",
  2630=>"001100100",
  2631=>"110100110",
  2632=>"101111111",
  2633=>"101010010",
  2634=>"001110110",
  2635=>"111101000",
  2636=>"000101110",
  2637=>"110101011",
  2638=>"010111110",
  2639=>"100011001",
  2640=>"010010110",
  2641=>"010011000",
  2642=>"010010101",
  2643=>"000010111",
  2644=>"110001001",
  2645=>"011111100",
  2646=>"011100001",
  2647=>"011010010",
  2648=>"011111110",
  2649=>"101001101",
  2650=>"010100001",
  2651=>"000000000",
  2652=>"000010101",
  2653=>"010001001",
  2654=>"110001000",
  2655=>"100010010",
  2656=>"110000100",
  2657=>"111110111",
  2658=>"001010000",
  2659=>"000001111",
  2660=>"100011100",
  2661=>"111101101",
  2662=>"111010000",
  2663=>"011111111",
  2664=>"111111001",
  2665=>"110001011",
  2666=>"000101001",
  2667=>"011010001",
  2668=>"101101110",
  2669=>"100110100",
  2670=>"110011101",
  2671=>"101100111",
  2672=>"010011100",
  2673=>"100011011",
  2674=>"001101011",
  2675=>"101011100",
  2676=>"011011100",
  2677=>"110001000",
  2678=>"011000101",
  2679=>"111100110",
  2680=>"010000111",
  2681=>"001101001",
  2682=>"100110010",
  2683=>"001000111",
  2684=>"001001100",
  2685=>"111011101",
  2686=>"111111000",
  2687=>"101101001",
  2688=>"101011010",
  2689=>"011000000",
  2690=>"100110001",
  2691=>"000000101",
  2692=>"101110101",
  2693=>"101100000",
  2694=>"111001001",
  2695=>"100110011",
  2696=>"101010010",
  2697=>"100100000",
  2698=>"111101111",
  2699=>"011011111",
  2700=>"010010101",
  2701=>"111011111",
  2702=>"000001000",
  2703=>"010010101",
  2704=>"010111111",
  2705=>"000111100",
  2706=>"111000110",
  2707=>"000000000",
  2708=>"011110110",
  2709=>"010111100",
  2710=>"011001100",
  2711=>"110110100",
  2712=>"010001001",
  2713=>"011110000",
  2714=>"011100101",
  2715=>"000000010",
  2716=>"001110010",
  2717=>"100000011",
  2718=>"010010001",
  2719=>"111111111",
  2720=>"000100001",
  2721=>"000010110",
  2722=>"101000100",
  2723=>"101001111",
  2724=>"000011110",
  2725=>"001000010",
  2726=>"011000010",
  2727=>"000000000",
  2728=>"001100010",
  2729=>"000111110",
  2730=>"110011001",
  2731=>"000010101",
  2732=>"001011110",
  2733=>"011111110",
  2734=>"101110111",
  2735=>"010111110",
  2736=>"000011100",
  2737=>"000110111",
  2738=>"001001001",
  2739=>"110010011",
  2740=>"100000011",
  2741=>"110100010",
  2742=>"000100100",
  2743=>"001100110",
  2744=>"100100101",
  2745=>"011001111",
  2746=>"110011011",
  2747=>"001101011",
  2748=>"011011101",
  2749=>"010110010",
  2750=>"111101100",
  2751=>"001011111",
  2752=>"001001110",
  2753=>"001101011",
  2754=>"001000110",
  2755=>"001001000",
  2756=>"011110000",
  2757=>"100101010",
  2758=>"001100100",
  2759=>"001110101",
  2760=>"000010011",
  2761=>"001010110",
  2762=>"101000010",
  2763=>"011011001",
  2764=>"000010010",
  2765=>"011101011",
  2766=>"111101101",
  2767=>"111000111",
  2768=>"001011110",
  2769=>"001000000",
  2770=>"001011001",
  2771=>"000011111",
  2772=>"110001100",
  2773=>"000001111",
  2774=>"011001111",
  2775=>"101000000",
  2776=>"000100101",
  2777=>"011111111",
  2778=>"110100001",
  2779=>"110011000",
  2780=>"100101111",
  2781=>"001010110",
  2782=>"001001100",
  2783=>"010111101",
  2784=>"011011101",
  2785=>"001111110",
  2786=>"111110000",
  2787=>"011100001",
  2788=>"000110001",
  2789=>"001011011",
  2790=>"011110100",
  2791=>"111111110",
  2792=>"001011001",
  2793=>"100001101",
  2794=>"010011101",
  2795=>"000100000",
  2796=>"010110111",
  2797=>"111111111",
  2798=>"010000000",
  2799=>"011000011",
  2800=>"111100111",
  2801=>"011000000",
  2802=>"011110110",
  2803=>"000000101",
  2804=>"101101000",
  2805=>"111100000",
  2806=>"111100111",
  2807=>"001011100",
  2808=>"110111110",
  2809=>"100011000",
  2810=>"010000000",
  2811=>"000011001",
  2812=>"100000000",
  2813=>"000000010",
  2814=>"101001101",
  2815=>"100010101",
  2816=>"111000100",
  2817=>"001111001",
  2818=>"001100000",
  2819=>"111110110",
  2820=>"111001100",
  2821=>"001010011",
  2822=>"111100101",
  2823=>"011010001",
  2824=>"111000000",
  2825=>"011100101",
  2826=>"000110101",
  2827=>"001101110",
  2828=>"001000100",
  2829=>"000100001",
  2830=>"011000000",
  2831=>"111001110",
  2832=>"100000101",
  2833=>"101011111",
  2834=>"111011111",
  2835=>"000000100",
  2836=>"010111110",
  2837=>"111111110",
  2838=>"001011000",
  2839=>"100100001",
  2840=>"001100000",
  2841=>"000000110",
  2842=>"100110011",
  2843=>"110101101",
  2844=>"100101000",
  2845=>"111111011",
  2846=>"110000001",
  2847=>"100100100",
  2848=>"001010101",
  2849=>"110000111",
  2850=>"110101111",
  2851=>"101011100",
  2852=>"001011001",
  2853=>"101111110",
  2854=>"101101001",
  2855=>"001111111",
  2856=>"001111111",
  2857=>"011001011",
  2858=>"111101010",
  2859=>"000110110",
  2860=>"001000100",
  2861=>"100010110",
  2862=>"100011000",
  2863=>"100011001",
  2864=>"010000100",
  2865=>"000101100",
  2866=>"010111111",
  2867=>"000010010",
  2868=>"101111111",
  2869=>"001001010",
  2870=>"001100001",
  2871=>"011011000",
  2872=>"001001010",
  2873=>"100100010",
  2874=>"010000010",
  2875=>"000101111",
  2876=>"100110000",
  2877=>"000010000",
  2878=>"101101000",
  2879=>"111110111",
  2880=>"000110000",
  2881=>"011001010",
  2882=>"001010001",
  2883=>"010101001",
  2884=>"100101001",
  2885=>"111101010",
  2886=>"110110011",
  2887=>"000011010",
  2888=>"100011110",
  2889=>"010110011",
  2890=>"011101001",
  2891=>"000011100",
  2892=>"011011001",
  2893=>"110000110",
  2894=>"000100001",
  2895=>"101001100",
  2896=>"101011000",
  2897=>"110111001",
  2898=>"111001100",
  2899=>"100011001",
  2900=>"111110101",
  2901=>"010111111",
  2902=>"111001111",
  2903=>"010010110",
  2904=>"000111010",
  2905=>"100001010",
  2906=>"100110001",
  2907=>"010010100",
  2908=>"010000100",
  2909=>"101100110",
  2910=>"100100011",
  2911=>"101101111",
  2912=>"100010111",
  2913=>"000001000",
  2914=>"000001011",
  2915=>"000100000",
  2916=>"101000111",
  2917=>"011000000",
  2918=>"100100011",
  2919=>"101101010",
  2920=>"111010111",
  2921=>"110111011",
  2922=>"111011010",
  2923=>"110101011",
  2924=>"110001000",
  2925=>"000100101",
  2926=>"001110100",
  2927=>"111011001",
  2928=>"010111101",
  2929=>"111001001",
  2930=>"001010010",
  2931=>"000001011",
  2932=>"000100111",
  2933=>"001010101",
  2934=>"001011011",
  2935=>"111110000",
  2936=>"011001000",
  2937=>"000100110",
  2938=>"010001100",
  2939=>"000010011",
  2940=>"101010111",
  2941=>"000001111",
  2942=>"011111110",
  2943=>"011101111",
  2944=>"000100011",
  2945=>"000111000",
  2946=>"100000001",
  2947=>"111010010",
  2948=>"110101010",
  2949=>"011001110",
  2950=>"110101000",
  2951=>"111110000",
  2952=>"101001010",
  2953=>"101000011",
  2954=>"101101000",
  2955=>"010111100",
  2956=>"101000000",
  2957=>"100000001",
  2958=>"100001001",
  2959=>"001010000",
  2960=>"011101110",
  2961=>"010110010",
  2962=>"000000000",
  2963=>"110100010",
  2964=>"111110111",
  2965=>"110110001",
  2966=>"010010111",
  2967=>"110010001",
  2968=>"110000101",
  2969=>"000110001",
  2970=>"111110111",
  2971=>"010100001",
  2972=>"001000110",
  2973=>"110111000",
  2974=>"001001010",
  2975=>"111111111",
  2976=>"001111010",
  2977=>"010000001",
  2978=>"111011010",
  2979=>"100011101",
  2980=>"000110110",
  2981=>"010100100",
  2982=>"000001010",
  2983=>"111110110",
  2984=>"100000000",
  2985=>"010000010",
  2986=>"011111101",
  2987=>"000010101",
  2988=>"101001100",
  2989=>"101011101",
  2990=>"101001111",
  2991=>"101010000",
  2992=>"010110100",
  2993=>"110000111",
  2994=>"100110000",
  2995=>"101100010",
  2996=>"100110011",
  2997=>"110000110",
  2998=>"101101110",
  2999=>"001010110",
  3000=>"110001110",
  3001=>"000010011",
  3002=>"010011001",
  3003=>"010011100",
  3004=>"100101000",
  3005=>"110111010",
  3006=>"110000010",
  3007=>"000101110",
  3008=>"100011000",
  3009=>"110011100",
  3010=>"011010111",
  3011=>"111100010",
  3012=>"110011010",
  3013=>"011011001",
  3014=>"101010111",
  3015=>"010111110",
  3016=>"101000000",
  3017=>"110110010",
  3018=>"001101001",
  3019=>"010110011",
  3020=>"000010101",
  3021=>"100101110",
  3022=>"010111000",
  3023=>"101011001",
  3024=>"111001000",
  3025=>"000000001",
  3026=>"110100100",
  3027=>"100011110",
  3028=>"001111000",
  3029=>"011000011",
  3030=>"001000100",
  3031=>"010011000",
  3032=>"101000110",
  3033=>"010101111",
  3034=>"000000000",
  3035=>"001010011",
  3036=>"010100101",
  3037=>"001001110",
  3038=>"000000000",
  3039=>"000010101",
  3040=>"011111011",
  3041=>"100000111",
  3042=>"001011110",
  3043=>"111010001",
  3044=>"110101000",
  3045=>"111100111",
  3046=>"000110001",
  3047=>"110101010",
  3048=>"001110100",
  3049=>"101001111",
  3050=>"000000011",
  3051=>"001100100",
  3052=>"111011101",
  3053=>"101100100",
  3054=>"010000000",
  3055=>"111110110",
  3056=>"001101111",
  3057=>"111011001",
  3058=>"011111110",
  3059=>"110111010",
  3060=>"111111101",
  3061=>"011110100",
  3062=>"011010111",
  3063=>"100110101",
  3064=>"011010000",
  3065=>"001001010",
  3066=>"010100000",
  3067=>"010011000",
  3068=>"001111100",
  3069=>"100011110",
  3070=>"111100111",
  3071=>"100000010",
  3072=>"110000000",
  3073=>"000110100",
  3074=>"001100001",
  3075=>"000100011",
  3076=>"100010110",
  3077=>"111011000",
  3078=>"001110010",
  3079=>"111001001",
  3080=>"100111010",
  3081=>"001010110",
  3082=>"110010110",
  3083=>"010010001",
  3084=>"001001110",
  3085=>"011001100",
  3086=>"111001000",
  3087=>"011011011",
  3088=>"110001001",
  3089=>"010000000",
  3090=>"011110000",
  3091=>"100110000",
  3092=>"110111100",
  3093=>"010101011",
  3094=>"111011010",
  3095=>"011010010",
  3096=>"000101110",
  3097=>"001001000",
  3098=>"000110110",
  3099=>"101011001",
  3100=>"000001001",
  3101=>"100101100",
  3102=>"110010001",
  3103=>"100010011",
  3104=>"000101100",
  3105=>"100101101",
  3106=>"011101010",
  3107=>"010010110",
  3108=>"010100011",
  3109=>"111011110",
  3110=>"011001001",
  3111=>"001110100",
  3112=>"000100101",
  3113=>"101011101",
  3114=>"110010101",
  3115=>"100001101",
  3116=>"100111111",
  3117=>"101100111",
  3118=>"100100110",
  3119=>"000000101",
  3120=>"111000100",
  3121=>"110111001",
  3122=>"101100011",
  3123=>"001111000",
  3124=>"010110011",
  3125=>"010010011",
  3126=>"000001011",
  3127=>"101111010",
  3128=>"111001101",
  3129=>"111001100",
  3130=>"110100011",
  3131=>"101010011",
  3132=>"001100011",
  3133=>"110101110",
  3134=>"011010111",
  3135=>"000110111",
  3136=>"010010100",
  3137=>"000000011",
  3138=>"001010110",
  3139=>"100011000",
  3140=>"111000011",
  3141=>"001110111",
  3142=>"100001010",
  3143=>"100010010",
  3144=>"010001100",
  3145=>"110111110",
  3146=>"001000101",
  3147=>"001011101",
  3148=>"010101110",
  3149=>"100110101",
  3150=>"100101010",
  3151=>"001110011",
  3152=>"100001110",
  3153=>"100101101",
  3154=>"011111010",
  3155=>"111010010",
  3156=>"000001111",
  3157=>"000010001",
  3158=>"001010011",
  3159=>"001101110",
  3160=>"011000100",
  3161=>"001001101",
  3162=>"011111110",
  3163=>"001000000",
  3164=>"100100101",
  3165=>"100001101",
  3166=>"110101111",
  3167=>"010110111",
  3168=>"000010101",
  3169=>"001110011",
  3170=>"110100111",
  3171=>"100000110",
  3172=>"100001001",
  3173=>"100001101",
  3174=>"010011000",
  3175=>"101001111",
  3176=>"010000011",
  3177=>"010110011",
  3178=>"100110001",
  3179=>"111110001",
  3180=>"101110110",
  3181=>"111001101",
  3182=>"001101100",
  3183=>"100111101",
  3184=>"000010000",
  3185=>"000001001",
  3186=>"110010011",
  3187=>"010111000",
  3188=>"001111111",
  3189=>"100110110",
  3190=>"100101011",
  3191=>"011010001",
  3192=>"101011101",
  3193=>"000011000",
  3194=>"001100010",
  3195=>"111001011",
  3196=>"000110000",
  3197=>"001010100",
  3198=>"010110011",
  3199=>"010110011",
  3200=>"111110110",
  3201=>"000111100",
  3202=>"001001101",
  3203=>"100100101",
  3204=>"011010110",
  3205=>"000111100",
  3206=>"000111011",
  3207=>"110111001",
  3208=>"010100011",
  3209=>"101101001",
  3210=>"101110101",
  3211=>"101111011",
  3212=>"011011110",
  3213=>"111111001",
  3214=>"001010010",
  3215=>"110000101",
  3216=>"101111010",
  3217=>"011101111",
  3218=>"010110100",
  3219=>"100010010",
  3220=>"001001000",
  3221=>"111101111",
  3222=>"100001010",
  3223=>"110000000",
  3224=>"100000010",
  3225=>"001100100",
  3226=>"111101100",
  3227=>"100000000",
  3228=>"110111101",
  3229=>"000010010",
  3230=>"101100011",
  3231=>"100011011",
  3232=>"001100111",
  3233=>"110011010",
  3234=>"011100011",
  3235=>"110001000",
  3236=>"010110000",
  3237=>"001111110",
  3238=>"110011101",
  3239=>"100001101",
  3240=>"011011010",
  3241=>"100010100",
  3242=>"000001011",
  3243=>"000101101",
  3244=>"000100110",
  3245=>"111001100",
  3246=>"111111100",
  3247=>"000111010",
  3248=>"001101001",
  3249=>"010010110",
  3250=>"111010110",
  3251=>"111100010",
  3252=>"011111100",
  3253=>"010101010",
  3254=>"000110010",
  3255=>"101001011",
  3256=>"111001011",
  3257=>"010000111",
  3258=>"100000000",
  3259=>"100101001",
  3260=>"010100010",
  3261=>"111001101",
  3262=>"110000000",
  3263=>"111110111",
  3264=>"000111110",
  3265=>"101000001",
  3266=>"100001001",
  3267=>"100100111",
  3268=>"111001001",
  3269=>"110101111",
  3270=>"111111110",
  3271=>"111001110",
  3272=>"110101110",
  3273=>"011011011",
  3274=>"001011011",
  3275=>"110010001",
  3276=>"011000010",
  3277=>"010010001",
  3278=>"101101011",
  3279=>"100101100",
  3280=>"000100110",
  3281=>"001110111",
  3282=>"101001001",
  3283=>"000111010",
  3284=>"111001111",
  3285=>"000101111",
  3286=>"000100010",
  3287=>"000001100",
  3288=>"101100101",
  3289=>"110011110",
  3290=>"001100100",
  3291=>"111011101",
  3292=>"011011010",
  3293=>"110110011",
  3294=>"001101010",
  3295=>"011110111",
  3296=>"001100100",
  3297=>"011100100",
  3298=>"010111011",
  3299=>"100000001",
  3300=>"000001010",
  3301=>"100111001",
  3302=>"010101010",
  3303=>"100110111",
  3304=>"101110101",
  3305=>"100111111",
  3306=>"000001101",
  3307=>"101101100",
  3308=>"001000001",
  3309=>"010001110",
  3310=>"111111100",
  3311=>"101111110",
  3312=>"101101101",
  3313=>"000011101",
  3314=>"100110010",
  3315=>"100100111",
  3316=>"100011101",
  3317=>"001110110",
  3318=>"111100111",
  3319=>"000101011",
  3320=>"110010000",
  3321=>"010001001",
  3322=>"111001110",
  3323=>"111010010",
  3324=>"110001000",
  3325=>"110000010",
  3326=>"110110011",
  3327=>"001101101",
  3328=>"111101110",
  3329=>"111000001",
  3330=>"011000110",
  3331=>"111011011",
  3332=>"000000111",
  3333=>"110001001",
  3334=>"011011100",
  3335=>"111110010",
  3336=>"000001010",
  3337=>"111110100",
  3338=>"010010101",
  3339=>"110001110",
  3340=>"010000101",
  3341=>"110000000",
  3342=>"101000101",
  3343=>"110001010",
  3344=>"011011111",
  3345=>"101101001",
  3346=>"100010101",
  3347=>"011010111",
  3348=>"001110010",
  3349=>"011101010",
  3350=>"001000000",
  3351=>"000001010",
  3352=>"101000001",
  3353=>"100011111",
  3354=>"100100100",
  3355=>"010010100",
  3356=>"001101101",
  3357=>"010001000",
  3358=>"111001011",
  3359=>"000101000",
  3360=>"000110111",
  3361=>"101111111",
  3362=>"110111101",
  3363=>"000000101",
  3364=>"011101010",
  3365=>"111001100",
  3366=>"010011000",
  3367=>"100000110",
  3368=>"000101110",
  3369=>"000001011",
  3370=>"111101001",
  3371=>"101000101",
  3372=>"110101110",
  3373=>"110000010",
  3374=>"000001000",
  3375=>"100000100",
  3376=>"000010001",
  3377=>"111011110",
  3378=>"111100001",
  3379=>"011100001",
  3380=>"011011110",
  3381=>"100110110",
  3382=>"010100110",
  3383=>"110100110",
  3384=>"110110101",
  3385=>"011000010",
  3386=>"010100000",
  3387=>"111100011",
  3388=>"001011010",
  3389=>"101010001",
  3390=>"001011001",
  3391=>"110000101",
  3392=>"011010010",
  3393=>"111110011",
  3394=>"110100000",
  3395=>"000011010",
  3396=>"011101111",
  3397=>"110111000",
  3398=>"000010101",
  3399=>"100101100",
  3400=>"111001000",
  3401=>"000000001",
  3402=>"000100101",
  3403=>"101001000",
  3404=>"011011101",
  3405=>"010111011",
  3406=>"000100111",
  3407=>"100001110",
  3408=>"011010000",
  3409=>"010100101",
  3410=>"000111110",
  3411=>"101011110",
  3412=>"010000010",
  3413=>"011110010",
  3414=>"111111101",
  3415=>"001101011",
  3416=>"001100110",
  3417=>"011010001",
  3418=>"100110011",
  3419=>"110000011",
  3420=>"110110100",
  3421=>"011000101",
  3422=>"100000111",
  3423=>"111010100",
  3424=>"010110000",
  3425=>"011011110",
  3426=>"101101000",
  3427=>"000111111",
  3428=>"101011110",
  3429=>"100101011",
  3430=>"000001111",
  3431=>"011010001",
  3432=>"110001011",
  3433=>"111101100",
  3434=>"010101111",
  3435=>"101101100",
  3436=>"111100110",
  3437=>"001000001",
  3438=>"000101011",
  3439=>"011110000",
  3440=>"000101010",
  3441=>"111111110",
  3442=>"000110001",
  3443=>"001110101",
  3444=>"000100000",
  3445=>"011010101",
  3446=>"111100111",
  3447=>"010001110",
  3448=>"100001110",
  3449=>"001000100",
  3450=>"111100101",
  3451=>"110100001",
  3452=>"110111011",
  3453=>"010011000",
  3454=>"100110111",
  3455=>"110011111",
  3456=>"100111100",
  3457=>"101001111",
  3458=>"110101100",
  3459=>"011110010",
  3460=>"100001100",
  3461=>"110001110",
  3462=>"010010011",
  3463=>"110110111",
  3464=>"011101000",
  3465=>"111000000",
  3466=>"011001000",
  3467=>"110110011",
  3468=>"111111111",
  3469=>"000001110",
  3470=>"000100011",
  3471=>"000111110",
  3472=>"110010011",
  3473=>"100000001",
  3474=>"001001101",
  3475=>"101010011",
  3476=>"111110000",
  3477=>"000101010",
  3478=>"101110011",
  3479=>"001011011",
  3480=>"011100010",
  3481=>"101000101",
  3482=>"110101001",
  3483=>"000111000",
  3484=>"111011010",
  3485=>"011100000",
  3486=>"010111111",
  3487=>"100100101",
  3488=>"000011000",
  3489=>"001100000",
  3490=>"001110010",
  3491=>"000100011",
  3492=>"010100001",
  3493=>"100100100",
  3494=>"010010011",
  3495=>"001000001",
  3496=>"111101100",
  3497=>"011010000",
  3498=>"111100000",
  3499=>"101011100",
  3500=>"100000110",
  3501=>"110100110",
  3502=>"100000100",
  3503=>"111100100",
  3504=>"101110111",
  3505=>"111001010",
  3506=>"110001010",
  3507=>"010000101",
  3508=>"000000101",
  3509=>"100011001",
  3510=>"001010101",
  3511=>"111111110",
  3512=>"110010110",
  3513=>"010001101",
  3514=>"001001101",
  3515=>"111011010",
  3516=>"111011111",
  3517=>"111000101",
  3518=>"101001000",
  3519=>"110101001",
  3520=>"011000101",
  3521=>"011001010",
  3522=>"110111100",
  3523=>"100110011",
  3524=>"111110001",
  3525=>"001001111",
  3526=>"110110111",
  3527=>"000001001",
  3528=>"100110111",
  3529=>"101010011",
  3530=>"111001101",
  3531=>"110100101",
  3532=>"001011100",
  3533=>"100100000",
  3534=>"000111010",
  3535=>"000011110",
  3536=>"001100010",
  3537=>"001101001",
  3538=>"001001100",
  3539=>"100110111",
  3540=>"111110111",
  3541=>"001100001",
  3542=>"010101000",
  3543=>"100001101",
  3544=>"001011101",
  3545=>"000111000",
  3546=>"110011000",
  3547=>"111010110",
  3548=>"011110010",
  3549=>"010000110",
  3550=>"000010111",
  3551=>"011011000",
  3552=>"010100000",
  3553=>"111000011",
  3554=>"101001010",
  3555=>"110000110",
  3556=>"100101100",
  3557=>"010100011",
  3558=>"100111101",
  3559=>"111100100",
  3560=>"101000011",
  3561=>"100000000",
  3562=>"000010000",
  3563=>"001001100",
  3564=>"000110010",
  3565=>"000111110",
  3566=>"111000100",
  3567=>"110111111",
  3568=>"100011100",
  3569=>"000100000",
  3570=>"001011110",
  3571=>"011101100",
  3572=>"111101011",
  3573=>"000111000",
  3574=>"010000111",
  3575=>"000100000",
  3576=>"100100011",
  3577=>"111011011",
  3578=>"100001011",
  3579=>"101101100",
  3580=>"000111110",
  3581=>"000110101",
  3582=>"011011110",
  3583=>"100000100",
  3584=>"010110001",
  3585=>"001000001",
  3586=>"000000011",
  3587=>"000111011",
  3588=>"110000111",
  3589=>"010111111",
  3590=>"011000000",
  3591=>"011100000",
  3592=>"100001000",
  3593=>"000110010",
  3594=>"101101000",
  3595=>"001010001",
  3596=>"010011110",
  3597=>"111010101",
  3598=>"011100000",
  3599=>"010010001",
  3600=>"111010110",
  3601=>"111101111",
  3602=>"100010011",
  3603=>"100100010",
  3604=>"111111111",
  3605=>"010101011",
  3606=>"101111100",
  3607=>"111101100",
  3608=>"010111010",
  3609=>"111001110",
  3610=>"100000101",
  3611=>"101101011",
  3612=>"110011111",
  3613=>"111001000",
  3614=>"011101101",
  3615=>"100110110",
  3616=>"110000011",
  3617=>"100101000",
  3618=>"110000100",
  3619=>"100000101",
  3620=>"111001010",
  3621=>"011001110",
  3622=>"000000100",
  3623=>"111111011",
  3624=>"100011100",
  3625=>"111100111",
  3626=>"001101010",
  3627=>"110010011",
  3628=>"010001011",
  3629=>"100011001",
  3630=>"010001010",
  3631=>"011110101",
  3632=>"110101100",
  3633=>"001101010",
  3634=>"010100010",
  3635=>"000000010",
  3636=>"010111010",
  3637=>"110111111",
  3638=>"010101000",
  3639=>"011111001",
  3640=>"110011111",
  3641=>"110010110",
  3642=>"001100110",
  3643=>"001110101",
  3644=>"110001011",
  3645=>"001101100",
  3646=>"111000100",
  3647=>"000010111",
  3648=>"000011110",
  3649=>"001101101",
  3650=>"010101100",
  3651=>"001110001",
  3652=>"001111101",
  3653=>"011001101",
  3654=>"001001111",
  3655=>"111001101",
  3656=>"011001010",
  3657=>"000111101",
  3658=>"000110000",
  3659=>"000110111",
  3660=>"110010110",
  3661=>"000010011",
  3662=>"001111000",
  3663=>"100011101",
  3664=>"011000001",
  3665=>"011011110",
  3666=>"110011010",
  3667=>"001100010",
  3668=>"001000110",
  3669=>"100000000",
  3670=>"100010111",
  3671=>"001111001",
  3672=>"100110001",
  3673=>"101100100",
  3674=>"000011000",
  3675=>"101011110",
  3676=>"111100100",
  3677=>"000000100",
  3678=>"101010111",
  3679=>"101110001",
  3680=>"001001000",
  3681=>"101011000",
  3682=>"011001001",
  3683=>"001010110",
  3684=>"101101100",
  3685=>"111111011",
  3686=>"001110001",
  3687=>"001100000",
  3688=>"010000111",
  3689=>"010110011",
  3690=>"011010010",
  3691=>"010000010",
  3692=>"010110101",
  3693=>"010000111",
  3694=>"110000010",
  3695=>"111010011",
  3696=>"110110101",
  3697=>"110001100",
  3698=>"111011111",
  3699=>"000001011",
  3700=>"101100110",
  3701=>"100000010",
  3702=>"111110110",
  3703=>"100010010",
  3704=>"110110111",
  3705=>"110111100",
  3706=>"111111111",
  3707=>"100000101",
  3708=>"101100001",
  3709=>"001110000",
  3710=>"010100010",
  3711=>"101011010",
  3712=>"100000000",
  3713=>"011110111",
  3714=>"010000110",
  3715=>"110100111",
  3716=>"000111001",
  3717=>"100000011",
  3718=>"110110011",
  3719=>"110001011",
  3720=>"101110111",
  3721=>"010000101",
  3722=>"010010010",
  3723=>"110010111",
  3724=>"000000000",
  3725=>"100001100",
  3726=>"010100100",
  3727=>"110011100",
  3728=>"110001011",
  3729=>"100010000",
  3730=>"101111000",
  3731=>"111111111",
  3732=>"000000001",
  3733=>"110000111",
  3734=>"010110011",
  3735=>"000101110",
  3736=>"101111100",
  3737=>"110100101",
  3738=>"010100111",
  3739=>"001101111",
  3740=>"101100110",
  3741=>"110111011",
  3742=>"001010111",
  3743=>"010111001",
  3744=>"101001001",
  3745=>"000001000",
  3746=>"010000101",
  3747=>"111110101",
  3748=>"011101011",
  3749=>"110010101",
  3750=>"111011010",
  3751=>"001100011",
  3752=>"110100110",
  3753=>"001101000",
  3754=>"000010011",
  3755=>"010100100",
  3756=>"101001110",
  3757=>"000000101",
  3758=>"101100001",
  3759=>"001111000",
  3760=>"011001000",
  3761=>"010010111",
  3762=>"100100000",
  3763=>"010000010",
  3764=>"110100100",
  3765=>"000100110",
  3766=>"001000110",
  3767=>"101101011",
  3768=>"110010011",
  3769=>"011110111",
  3770=>"101001100",
  3771=>"111100011",
  3772=>"110101011",
  3773=>"000110110",
  3774=>"111010001",
  3775=>"110000000",
  3776=>"000110110",
  3777=>"000110001",
  3778=>"010111000",
  3779=>"010111110",
  3780=>"011000111",
  3781=>"110100101",
  3782=>"000101000",
  3783=>"110000010",
  3784=>"010011000",
  3785=>"010000001",
  3786=>"001111000",
  3787=>"000101100",
  3788=>"110000000",
  3789=>"110111111",
  3790=>"111111101",
  3791=>"000010100",
  3792=>"100001011",
  3793=>"111111011",
  3794=>"101100010",
  3795=>"000001101",
  3796=>"101100010",
  3797=>"100001110",
  3798=>"110101111",
  3799=>"010000110",
  3800=>"100110000",
  3801=>"100010000",
  3802=>"010001001",
  3803=>"011111011",
  3804=>"111100111",
  3805=>"100001010",
  3806=>"100110001",
  3807=>"111011110",
  3808=>"111111111",
  3809=>"111111001",
  3810=>"001010110",
  3811=>"001110011",
  3812=>"111000101",
  3813=>"101000101",
  3814=>"001001111",
  3815=>"100110000",
  3816=>"101010111",
  3817=>"010000111",
  3818=>"101111110",
  3819=>"010011110",
  3820=>"000101101",
  3821=>"000111101",
  3822=>"000101010",
  3823=>"100100010",
  3824=>"010001101",
  3825=>"111100010",
  3826=>"011000011",
  3827=>"010010110",
  3828=>"001110010",
  3829=>"111010111",
  3830=>"010001111",
  3831=>"011111011",
  3832=>"101010010",
  3833=>"011101110",
  3834=>"101000100",
  3835=>"111110010",
  3836=>"110100110",
  3837=>"011000010",
  3838=>"011111000",
  3839=>"111011001",
  3840=>"010000011",
  3841=>"000000000",
  3842=>"110110110",
  3843=>"000000011",
  3844=>"100110111",
  3845=>"010010101",
  3846=>"111000101",
  3847=>"011001010",
  3848=>"110010101",
  3849=>"111111010",
  3850=>"011010111",
  3851=>"101100011",
  3852=>"001111110",
  3853=>"111110110",
  3854=>"100101110",
  3855=>"001100100",
  3856=>"000010111",
  3857=>"001111000",
  3858=>"001000101",
  3859=>"001011101",
  3860=>"000000111",
  3861=>"100100100",
  3862=>"100001110",
  3863=>"101001111",
  3864=>"101101110",
  3865=>"001101100",
  3866=>"011111100",
  3867=>"101000000",
  3868=>"001100010",
  3869=>"011101011",
  3870=>"001111010",
  3871=>"001111111",
  3872=>"100011000",
  3873=>"010110100",
  3874=>"111100011",
  3875=>"011000010",
  3876=>"101101101",
  3877=>"000001000",
  3878=>"010111100",
  3879=>"010100100",
  3880=>"111100101",
  3881=>"110101101",
  3882=>"101101100",
  3883=>"010010110",
  3884=>"011011101",
  3885=>"001111100",
  3886=>"000000110",
  3887=>"110111010",
  3888=>"000000100",
  3889=>"100111100",
  3890=>"011110101",
  3891=>"111111111",
  3892=>"011000000",
  3893=>"010000001",
  3894=>"000010000",
  3895=>"101000010",
  3896=>"000110001",
  3897=>"000110000",
  3898=>"001101000",
  3899=>"011010001",
  3900=>"110110110",
  3901=>"000100000",
  3902=>"111010101",
  3903=>"001000010",
  3904=>"010110111",
  3905=>"111001100",
  3906=>"100101111",
  3907=>"111000010",
  3908=>"100000111",
  3909=>"101001100",
  3910=>"011000110",
  3911=>"110110001",
  3912=>"001111100",
  3913=>"110101110",
  3914=>"110011010",
  3915=>"001111001",
  3916=>"001011100",
  3917=>"111111000",
  3918=>"110010111",
  3919=>"100000011",
  3920=>"000110110",
  3921=>"100010000",
  3922=>"011000011",
  3923=>"100111110",
  3924=>"010010010",
  3925=>"110011001",
  3926=>"001101011",
  3927=>"100010011",
  3928=>"111111100",
  3929=>"110001101",
  3930=>"101001101",
  3931=>"111101010",
  3932=>"111101111",
  3933=>"001110001",
  3934=>"010101000",
  3935=>"100011010",
  3936=>"101000000",
  3937=>"100001010",
  3938=>"000011101",
  3939=>"000111111",
  3940=>"110010000",
  3941=>"010111100",
  3942=>"101011101",
  3943=>"010100111",
  3944=>"111000100",
  3945=>"011101010",
  3946=>"000000001",
  3947=>"010010111",
  3948=>"000011100",
  3949=>"000101010",
  3950=>"000100110",
  3951=>"101000000",
  3952=>"001011110",
  3953=>"111101010",
  3954=>"101000010",
  3955=>"101001001",
  3956=>"000010010",
  3957=>"011001000",
  3958=>"001011000",
  3959=>"011011000",
  3960=>"101101111",
  3961=>"011100110",
  3962=>"101100000",
  3963=>"110111100",
  3964=>"011101001",
  3965=>"111101010",
  3966=>"010010100",
  3967=>"111110111",
  3968=>"001001011",
  3969=>"100000111",
  3970=>"001101001",
  3971=>"110001001",
  3972=>"010111010",
  3973=>"011000001",
  3974=>"111011011",
  3975=>"000001010",
  3976=>"001001110",
  3977=>"000110111",
  3978=>"000010111",
  3979=>"000100111",
  3980=>"110111011",
  3981=>"111001010",
  3982=>"101000111",
  3983=>"011100000",
  3984=>"110001100",
  3985=>"111000101",
  3986=>"110110011",
  3987=>"011111101",
  3988=>"000111101",
  3989=>"110011011",
  3990=>"100010001",
  3991=>"110100010",
  3992=>"100110000",
  3993=>"001100011",
  3994=>"010000000",
  3995=>"010011111",
  3996=>"110111001",
  3997=>"000011110",
  3998=>"101011000",
  3999=>"111000101",
  4000=>"111101110",
  4001=>"100011001",
  4002=>"110111010",
  4003=>"111110100",
  4004=>"101100000",
  4005=>"100001110",
  4006=>"100111101",
  4007=>"001110110",
  4008=>"111100010",
  4009=>"100010010",
  4010=>"001111100",
  4011=>"110110010",
  4012=>"010110110",
  4013=>"001000101",
  4014=>"011011000",
  4015=>"100010001",
  4016=>"101100111",
  4017=>"111011010",
  4018=>"101011110",
  4019=>"101100101",
  4020=>"111011101",
  4021=>"000100000",
  4022=>"110011001",
  4023=>"011101000",
  4024=>"100000111",
  4025=>"011011101",
  4026=>"001001000",
  4027=>"111101010",
  4028=>"111110100",
  4029=>"000111110",
  4030=>"111101001",
  4031=>"111110111",
  4032=>"001110111",
  4033=>"000010001",
  4034=>"110111010",
  4035=>"111010011",
  4036=>"010100110",
  4037=>"001000010",
  4038=>"001011110",
  4039=>"001000000",
  4040=>"110000101",
  4041=>"011101001",
  4042=>"111001100",
  4043=>"011110011",
  4044=>"100011100",
  4045=>"110000110",
  4046=>"100110001",
  4047=>"110001011",
  4048=>"011001110",
  4049=>"000011010",
  4050=>"000111010",
  4051=>"001000101",
  4052=>"011100110",
  4053=>"100110001",
  4054=>"101100110",
  4055=>"101111111",
  4056=>"101101100",
  4057=>"000000001",
  4058=>"000001011",
  4059=>"100010011",
  4060=>"011010110",
  4061=>"100100011",
  4062=>"001101101",
  4063=>"011100010",
  4064=>"001000011",
  4065=>"010110011",
  4066=>"000011010",
  4067=>"111000110",
  4068=>"010010011",
  4069=>"010001000",
  4070=>"001100101",
  4071=>"110000010",
  4072=>"000001000",
  4073=>"011110000",
  4074=>"110000110",
  4075=>"010000100",
  4076=>"100100111",
  4077=>"001111100",
  4078=>"001101100",
  4079=>"001010111",
  4080=>"100101111",
  4081=>"010100010",
  4082=>"010011101",
  4083=>"111111000",
  4084=>"000000010",
  4085=>"100101001",
  4086=>"010010111",
  4087=>"111001100",
  4088=>"111010101",
  4089=>"111111100",
  4090=>"111101011",
  4091=>"100101110",
  4092=>"110001111",
  4093=>"001111001",
  4094=>"100100110",
  4095=>"101100001",
  4096=>"010110101",
  4097=>"100001101",
  4098=>"101010111",
  4099=>"000100001",
  4100=>"111010111",
  4101=>"011101011",
  4102=>"010101111",
  4103=>"001101110",
  4104=>"100001101",
  4105=>"110010110",
  4106=>"000010011",
  4107=>"000010000",
  4108=>"010100110",
  4109=>"010001010",
  4110=>"011111101",
  4111=>"011011100",
  4112=>"100010010",
  4113=>"100001101",
  4114=>"100101110",
  4115=>"001100111",
  4116=>"010010011",
  4117=>"110111101",
  4118=>"010101111",
  4119=>"100010011",
  4120=>"111110100",
  4121=>"000000100",
  4122=>"011010101",
  4123=>"011101110",
  4124=>"011001100",
  4125=>"111000010",
  4126=>"011110101",
  4127=>"001100100",
  4128=>"101101100",
  4129=>"001000000",
  4130=>"101101100",
  4131=>"011101001",
  4132=>"011010001",
  4133=>"101101000",
  4134=>"010010101",
  4135=>"110011101",
  4136=>"100011010",
  4137=>"000010110",
  4138=>"011100100",
  4139=>"100100110",
  4140=>"110110001",
  4141=>"001101011",
  4142=>"101110010",
  4143=>"101110010",
  4144=>"011111001",
  4145=>"110101101",
  4146=>"100111100",
  4147=>"010000011",
  4148=>"101100011",
  4149=>"111101100",
  4150=>"111010001",
  4151=>"000101111",
  4152=>"111100001",
  4153=>"101011011",
  4154=>"101000101",
  4155=>"010011000",
  4156=>"001101110",
  4157=>"110000001",
  4158=>"000110101",
  4159=>"100011000",
  4160=>"100111001",
  4161=>"000000000",
  4162=>"001001110",
  4163=>"011110100",
  4164=>"100101000",
  4165=>"111000011",
  4166=>"100010010",
  4167=>"010010100",
  4168=>"001100001",
  4169=>"100001011",
  4170=>"011101010",
  4171=>"000001101",
  4172=>"001010111",
  4173=>"101010000",
  4174=>"111111011",
  4175=>"111001001",
  4176=>"111101111",
  4177=>"111000101",
  4178=>"111001101",
  4179=>"110001010",
  4180=>"101111010",
  4181=>"000101100",
  4182=>"001110001",
  4183=>"000111110",
  4184=>"001000100",
  4185=>"111101001",
  4186=>"101000101",
  4187=>"111111101",
  4188=>"110000110",
  4189=>"000111100",
  4190=>"010101001",
  4191=>"001010001",
  4192=>"010101100",
  4193=>"010100111",
  4194=>"100110110",
  4195=>"010101000",
  4196=>"010000100",
  4197=>"010111000",
  4198=>"011011010",
  4199=>"000000011",
  4200=>"000110111",
  4201=>"010110011",
  4202=>"000001101",
  4203=>"100011001",
  4204=>"000000101",
  4205=>"101110010",
  4206=>"011101001",
  4207=>"010100011",
  4208=>"011000001",
  4209=>"001100001",
  4210=>"000101000",
  4211=>"110111101",
  4212=>"101110101",
  4213=>"111110111",
  4214=>"100111101",
  4215=>"011010000",
  4216=>"001010010",
  4217=>"100001110",
  4218=>"111001001",
  4219=>"000000000",
  4220=>"001100010",
  4221=>"001001001",
  4222=>"001110100",
  4223=>"101110010",
  4224=>"011010000",
  4225=>"010111111",
  4226=>"001101110",
  4227=>"101001101",
  4228=>"010010001",
  4229=>"101111000",
  4230=>"010110110",
  4231=>"010010101",
  4232=>"000101000",
  4233=>"000000001",
  4234=>"111100000",
  4235=>"111110001",
  4236=>"101110011",
  4237=>"001001111",
  4238=>"001111110",
  4239=>"011100001",
  4240=>"101111111",
  4241=>"011110110",
  4242=>"001000101",
  4243=>"111010101",
  4244=>"100101101",
  4245=>"110001101",
  4246=>"011011000",
  4247=>"000011110",
  4248=>"100001100",
  4249=>"001101100",
  4250=>"000110110",
  4251=>"011110111",
  4252=>"000110001",
  4253=>"000010100",
  4254=>"010101000",
  4255=>"111100011",
  4256=>"101001111",
  4257=>"010111100",
  4258=>"010100110",
  4259=>"100110001",
  4260=>"010110111",
  4261=>"100111000",
  4262=>"010000100",
  4263=>"000101001",
  4264=>"010010010",
  4265=>"110100111",
  4266=>"101100001",
  4267=>"000110010",
  4268=>"101111111",
  4269=>"101000001",
  4270=>"001100001",
  4271=>"011111000",
  4272=>"110101111",
  4273=>"100000001",
  4274=>"011000001",
  4275=>"000011100",
  4276=>"001011000",
  4277=>"100011001",
  4278=>"100001010",
  4279=>"001011001",
  4280=>"110011001",
  4281=>"001001110",
  4282=>"101100010",
  4283=>"111111110",
  4284=>"010111001",
  4285=>"010000001",
  4286=>"110011001",
  4287=>"111100000",
  4288=>"110110101",
  4289=>"011010000",
  4290=>"001111011",
  4291=>"110111001",
  4292=>"101011000",
  4293=>"110101111",
  4294=>"010000001",
  4295=>"000010001",
  4296=>"100010110",
  4297=>"001111110",
  4298=>"110110110",
  4299=>"110110110",
  4300=>"100111110",
  4301=>"010011000",
  4302=>"100101110",
  4303=>"010100101",
  4304=>"110001011",
  4305=>"001010110",
  4306=>"110001011",
  4307=>"010110100",
  4308=>"110010000",
  4309=>"011101101",
  4310=>"000010001",
  4311=>"100001000",
  4312=>"010000010",
  4313=>"110010100",
  4314=>"010101100",
  4315=>"100010110",
  4316=>"101010000",
  4317=>"111001111",
  4318=>"110111010",
  4319=>"000000010",
  4320=>"100000100",
  4321=>"000010011",
  4322=>"010001101",
  4323=>"010011000",
  4324=>"010101000",
  4325=>"010110011",
  4326=>"011011101",
  4327=>"101111011",
  4328=>"110010110",
  4329=>"100100100",
  4330=>"110001011",
  4331=>"101110010",
  4332=>"000110010",
  4333=>"011100001",
  4334=>"001001100",
  4335=>"000010100",
  4336=>"000111010",
  4337=>"110101001",
  4338=>"011010101",
  4339=>"000101001",
  4340=>"000000110",
  4341=>"101101010",
  4342=>"101110011",
  4343=>"111100011",
  4344=>"101001110",
  4345=>"001101111",
  4346=>"010110100",
  4347=>"001010110",
  4348=>"100111111",
  4349=>"000110001",
  4350=>"001100101",
  4351=>"101010110",
  4352=>"111010111",
  4353=>"110101111",
  4354=>"101000011",
  4355=>"010100100",
  4356=>"111100011",
  4357=>"000111100",
  4358=>"000011101",
  4359=>"111101100",
  4360=>"100011111",
  4361=>"111010010",
  4362=>"101100101",
  4363=>"000000100",
  4364=>"010110111",
  4365=>"001010000",
  4366=>"110101100",
  4367=>"010001110",
  4368=>"010010101",
  4369=>"110110000",
  4370=>"001101001",
  4371=>"101000000",
  4372=>"010000101",
  4373=>"110010100",
  4374=>"010011111",
  4375=>"011001100",
  4376=>"011110010",
  4377=>"011101000",
  4378=>"100100110",
  4379=>"001101000",
  4380=>"000011001",
  4381=>"110000001",
  4382=>"010101011",
  4383=>"100100110",
  4384=>"101010000",
  4385=>"100010110",
  4386=>"010010111",
  4387=>"011101011",
  4388=>"111110000",
  4389=>"011101110",
  4390=>"001110001",
  4391=>"010110001",
  4392=>"001111000",
  4393=>"100000100",
  4394=>"001000001",
  4395=>"011000011",
  4396=>"110010011",
  4397=>"110000101",
  4398=>"110101101",
  4399=>"101101010",
  4400=>"010001010",
  4401=>"101100111",
  4402=>"000001100",
  4403=>"000110111",
  4404=>"100101000",
  4405=>"011000001",
  4406=>"010001110",
  4407=>"110111010",
  4408=>"100011100",
  4409=>"011010110",
  4410=>"000000111",
  4411=>"001001001",
  4412=>"001100010",
  4413=>"101000010",
  4414=>"100010010",
  4415=>"100010101",
  4416=>"000101100",
  4417=>"111100010",
  4418=>"010001110",
  4419=>"010101011",
  4420=>"000011010",
  4421=>"011111000",
  4422=>"011010010",
  4423=>"000000001",
  4424=>"000011110",
  4425=>"000000011",
  4426=>"000110101",
  4427=>"100000110",
  4428=>"101110110",
  4429=>"000101011",
  4430=>"101000011",
  4431=>"111011001",
  4432=>"010100011",
  4433=>"000111110",
  4434=>"010011110",
  4435=>"000001001",
  4436=>"101011011",
  4437=>"000110111",
  4438=>"001011110",
  4439=>"100011010",
  4440=>"001000000",
  4441=>"000001111",
  4442=>"101111001",
  4443=>"011100101",
  4444=>"011000100",
  4445=>"001000101",
  4446=>"110110000",
  4447=>"001101111",
  4448=>"100001111",
  4449=>"100101010",
  4450=>"000110010",
  4451=>"000100001",
  4452=>"000011010",
  4453=>"100010000",
  4454=>"111010010",
  4455=>"100000100",
  4456=>"101100010",
  4457=>"001111010",
  4458=>"010000110",
  4459=>"100001100",
  4460=>"001111100",
  4461=>"010010111",
  4462=>"100001100",
  4463=>"000111010",
  4464=>"100000011",
  4465=>"010111010",
  4466=>"101010001",
  4467=>"110000100",
  4468=>"011111000",
  4469=>"000111010",
  4470=>"101101101",
  4471=>"000100101",
  4472=>"110001010",
  4473=>"100000011",
  4474=>"101110010",
  4475=>"001110011",
  4476=>"000101100",
  4477=>"011100100",
  4478=>"101000000",
  4479=>"001000100",
  4480=>"101110011",
  4481=>"101101010",
  4482=>"110100101",
  4483=>"000010101",
  4484=>"111110001",
  4485=>"000000001",
  4486=>"110010101",
  4487=>"110110001",
  4488=>"010110000",
  4489=>"100000110",
  4490=>"000010010",
  4491=>"000010010",
  4492=>"010101011",
  4493=>"000110010",
  4494=>"010000101",
  4495=>"110111010",
  4496=>"010101010",
  4497=>"111001000",
  4498=>"100111111",
  4499=>"100001001",
  4500=>"100000100",
  4501=>"011111101",
  4502=>"100101101",
  4503=>"111110000",
  4504=>"110010001",
  4505=>"100000111",
  4506=>"011010110",
  4507=>"001000100",
  4508=>"101100010",
  4509=>"000110000",
  4510=>"111000000",
  4511=>"011111010",
  4512=>"011101001",
  4513=>"111101101",
  4514=>"100110000",
  4515=>"001001101",
  4516=>"111101001",
  4517=>"110100100",
  4518=>"101101110",
  4519=>"011011000",
  4520=>"110010100",
  4521=>"001001000",
  4522=>"011100100",
  4523=>"111100011",
  4524=>"100100100",
  4525=>"101011111",
  4526=>"000011010",
  4527=>"010111000",
  4528=>"000001100",
  4529=>"000000010",
  4530=>"011001100",
  4531=>"001010110",
  4532=>"001111010",
  4533=>"000101010",
  4534=>"100011100",
  4535=>"010001000",
  4536=>"111110101",
  4537=>"100101000",
  4538=>"001000011",
  4539=>"110111101",
  4540=>"001000100",
  4541=>"101001100",
  4542=>"010000101",
  4543=>"100001111",
  4544=>"010000001",
  4545=>"100001110",
  4546=>"001011010",
  4547=>"000011011",
  4548=>"110110001",
  4549=>"101000101",
  4550=>"010101100",
  4551=>"011011000",
  4552=>"111010010",
  4553=>"001110010",
  4554=>"100100111",
  4555=>"100011101",
  4556=>"111011111",
  4557=>"111011100",
  4558=>"100100110",
  4559=>"111110011",
  4560=>"100100001",
  4561=>"000010101",
  4562=>"000001110",
  4563=>"011110010",
  4564=>"111110101",
  4565=>"110101100",
  4566=>"100000000",
  4567=>"001100111",
  4568=>"101101001",
  4569=>"100011010",
  4570=>"010001000",
  4571=>"001000010",
  4572=>"111111011",
  4573=>"101001011",
  4574=>"010100000",
  4575=>"100000001",
  4576=>"101001000",
  4577=>"111101110",
  4578=>"000011000",
  4579=>"100110000",
  4580=>"100010010",
  4581=>"101011101",
  4582=>"011011000",
  4583=>"101101001",
  4584=>"000101100",
  4585=>"100010111",
  4586=>"000110111",
  4587=>"100011010",
  4588=>"111011110",
  4589=>"011001000",
  4590=>"110001110",
  4591=>"010011000",
  4592=>"000001010",
  4593=>"010111010",
  4594=>"100100010",
  4595=>"000100101",
  4596=>"110100101",
  4597=>"000111010",
  4598=>"000000010",
  4599=>"011101011",
  4600=>"111010110",
  4601=>"111111010",
  4602=>"000001000",
  4603=>"110110101",
  4604=>"111110110",
  4605=>"110110001",
  4606=>"110010011",
  4607=>"001101110",
  4608=>"001101100",
  4609=>"000001101",
  4610=>"110000110",
  4611=>"010101111",
  4612=>"001111011",
  4613=>"101011100",
  4614=>"011101100",
  4615=>"011000000",
  4616=>"001010000",
  4617=>"000001010",
  4618=>"010000010",
  4619=>"010010010",
  4620=>"001000010",
  4621=>"010101100",
  4622=>"111101001",
  4623=>"111011000",
  4624=>"000100110",
  4625=>"000100100",
  4626=>"000100001",
  4627=>"100010001",
  4628=>"000001101",
  4629=>"111010010",
  4630=>"011010000",
  4631=>"110010101",
  4632=>"000000100",
  4633=>"011001111",
  4634=>"011010010",
  4635=>"111111000",
  4636=>"000000100",
  4637=>"101001010",
  4638=>"000111011",
  4639=>"011000100",
  4640=>"101010011",
  4641=>"110100110",
  4642=>"110111101",
  4643=>"110100101",
  4644=>"111010011",
  4645=>"010110100",
  4646=>"100111110",
  4647=>"101110011",
  4648=>"001100000",
  4649=>"011101100",
  4650=>"110110101",
  4651=>"101001010",
  4652=>"100110100",
  4653=>"001110110",
  4654=>"100101101",
  4655=>"001100001",
  4656=>"010110010",
  4657=>"100101101",
  4658=>"110101101",
  4659=>"100101101",
  4660=>"110001111",
  4661=>"111100001",
  4662=>"010010001",
  4663=>"011110000",
  4664=>"111001101",
  4665=>"110100111",
  4666=>"100100001",
  4667=>"000111110",
  4668=>"010000010",
  4669=>"000000110",
  4670=>"111001000",
  4671=>"010110011",
  4672=>"001110000",
  4673=>"010100110",
  4674=>"001000100",
  4675=>"001111110",
  4676=>"111000001",
  4677=>"010101000",
  4678=>"100001000",
  4679=>"010101010",
  4680=>"110110011",
  4681=>"011011111",
  4682=>"101011000",
  4683=>"101101000",
  4684=>"110110101",
  4685=>"010000010",
  4686=>"011000011",
  4687=>"110001010",
  4688=>"010000111",
  4689=>"100000001",
  4690=>"000001000",
  4691=>"010100001",
  4692=>"010000111",
  4693=>"010101101",
  4694=>"101000010",
  4695=>"000000010",
  4696=>"110111111",
  4697=>"100111101",
  4698=>"101011000",
  4699=>"000101100",
  4700=>"111100010",
  4701=>"000001000",
  4702=>"011100101",
  4703=>"010110111",
  4704=>"110001000",
  4705=>"011111000",
  4706=>"000100001",
  4707=>"010111010",
  4708=>"101000000",
  4709=>"001001001",
  4710=>"000111000",
  4711=>"000000011",
  4712=>"001100001",
  4713=>"001001000",
  4714=>"111011010",
  4715=>"111101010",
  4716=>"000100101",
  4717=>"100011010",
  4718=>"101110101",
  4719=>"110100100",
  4720=>"010001000",
  4721=>"000101010",
  4722=>"101000010",
  4723=>"100010110",
  4724=>"001100010",
  4725=>"000101001",
  4726=>"101110000",
  4727=>"011101110",
  4728=>"001110100",
  4729=>"101111011",
  4730=>"101111011",
  4731=>"101101111",
  4732=>"110100000",
  4733=>"001111001",
  4734=>"111100000",
  4735=>"000010011",
  4736=>"001000011",
  4737=>"000101101",
  4738=>"111001000",
  4739=>"001111100",
  4740=>"100111001",
  4741=>"000001000",
  4742=>"000001000",
  4743=>"011000101",
  4744=>"000111011",
  4745=>"101100010",
  4746=>"110010101",
  4747=>"110110011",
  4748=>"111001100",
  4749=>"001110010",
  4750=>"010101100",
  4751=>"001010111",
  4752=>"111100010",
  4753=>"100101000",
  4754=>"000010011",
  4755=>"111011101",
  4756=>"100101000",
  4757=>"100001010",
  4758=>"100111001",
  4759=>"101100000",
  4760=>"100001000",
  4761=>"110000011",
  4762=>"010010001",
  4763=>"011111011",
  4764=>"000011000",
  4765=>"101101111",
  4766=>"001100000",
  4767=>"001001111",
  4768=>"101110011",
  4769=>"011111110",
  4770=>"000010000",
  4771=>"011101111",
  4772=>"100011111",
  4773=>"000101111",
  4774=>"111001011",
  4775=>"011101000",
  4776=>"110111001",
  4777=>"110010000",
  4778=>"110111001",
  4779=>"011101110",
  4780=>"000000000",
  4781=>"011010101",
  4782=>"110010101",
  4783=>"001011101",
  4784=>"011110000",
  4785=>"011010011",
  4786=>"010000001",
  4787=>"010111011",
  4788=>"111001111",
  4789=>"010001011",
  4790=>"011110111",
  4791=>"010010010",
  4792=>"111000100",
  4793=>"101110011",
  4794=>"000010110",
  4795=>"010110000",
  4796=>"110000001",
  4797=>"001010100",
  4798=>"011000010",
  4799=>"000000001",
  4800=>"101010001",
  4801=>"111111000",
  4802=>"101010000",
  4803=>"001100110",
  4804=>"100110111",
  4805=>"010011010",
  4806=>"000101001",
  4807=>"101111100",
  4808=>"101100100",
  4809=>"110100011",
  4810=>"100110010",
  4811=>"001101000",
  4812=>"101010000",
  4813=>"110001100",
  4814=>"110011100",
  4815=>"000100000",
  4816=>"111010010",
  4817=>"000101100",
  4818=>"001011110",
  4819=>"100101100",
  4820=>"110011100",
  4821=>"000111000",
  4822=>"011000110",
  4823=>"000100100",
  4824=>"110101000",
  4825=>"110110100",
  4826=>"100001111",
  4827=>"111111001",
  4828=>"101101011",
  4829=>"011011010",
  4830=>"011001000",
  4831=>"100101111",
  4832=>"001001010",
  4833=>"000011000",
  4834=>"100100010",
  4835=>"000111111",
  4836=>"001100000",
  4837=>"100111011",
  4838=>"000101000",
  4839=>"110100000",
  4840=>"000000001",
  4841=>"100110101",
  4842=>"111101010",
  4843=>"010010101",
  4844=>"001100011",
  4845=>"011000101",
  4846=>"110111101",
  4847=>"001010011",
  4848=>"010100001",
  4849=>"000111100",
  4850=>"111110000",
  4851=>"101101011",
  4852=>"000110001",
  4853=>"101011111",
  4854=>"100101111",
  4855=>"011000101",
  4856=>"101101001",
  4857=>"100010110",
  4858=>"010001110",
  4859=>"100000010",
  4860=>"101111101",
  4861=>"011001101",
  4862=>"001010100",
  4863=>"010100100",
  4864=>"010010000",
  4865=>"111101011",
  4866=>"110101010",
  4867=>"000111011",
  4868=>"111001100",
  4869=>"010001001",
  4870=>"011100100",
  4871=>"111110110",
  4872=>"000111110",
  4873=>"010000001",
  4874=>"101110001",
  4875=>"111111001",
  4876=>"010000011",
  4877=>"000010101",
  4878=>"011000110",
  4879=>"110000110",
  4880=>"110101100",
  4881=>"101000000",
  4882=>"100101011",
  4883=>"001100110",
  4884=>"100101110",
  4885=>"010011110",
  4886=>"110110000",
  4887=>"000011111",
  4888=>"110110000",
  4889=>"001010100",
  4890=>"000100110",
  4891=>"111101000",
  4892=>"111111100",
  4893=>"010111000",
  4894=>"000011000",
  4895=>"110011110",
  4896=>"000110001",
  4897=>"100011001",
  4898=>"000001111",
  4899=>"000111110",
  4900=>"110111110",
  4901=>"001101100",
  4902=>"111101111",
  4903=>"010110101",
  4904=>"101001101",
  4905=>"100110000",
  4906=>"111001110",
  4907=>"110101010",
  4908=>"100110101",
  4909=>"101001011",
  4910=>"111110001",
  4911=>"100100011",
  4912=>"000100001",
  4913=>"001001110",
  4914=>"010100100",
  4915=>"100011111",
  4916=>"000101111",
  4917=>"011010101",
  4918=>"000111100",
  4919=>"000000011",
  4920=>"010111000",
  4921=>"111011111",
  4922=>"000110110",
  4923=>"110111011",
  4924=>"110000110",
  4925=>"101001000",
  4926=>"011111101",
  4927=>"100110011",
  4928=>"010001000",
  4929=>"110100111",
  4930=>"111010110",
  4931=>"101010100",
  4932=>"001001101",
  4933=>"111101000",
  4934=>"011110100",
  4935=>"010011001",
  4936=>"111110111",
  4937=>"011011010",
  4938=>"101100110",
  4939=>"000110000",
  4940=>"001101111",
  4941=>"010001111",
  4942=>"010000100",
  4943=>"110110100",
  4944=>"000011010",
  4945=>"100111110",
  4946=>"010100110",
  4947=>"010000100",
  4948=>"001100011",
  4949=>"000001101",
  4950=>"011000111",
  4951=>"011101001",
  4952=>"100011111",
  4953=>"110110010",
  4954=>"111010111",
  4955=>"101010101",
  4956=>"000011001",
  4957=>"100101101",
  4958=>"000111000",
  4959=>"001010001",
  4960=>"011100000",
  4961=>"001001101",
  4962=>"000100100",
  4963=>"111010011",
  4964=>"100000111",
  4965=>"101110100",
  4966=>"011100010",
  4967=>"101111100",
  4968=>"000110101",
  4969=>"000101000",
  4970=>"100100010",
  4971=>"010101100",
  4972=>"011000010",
  4973=>"000111100",
  4974=>"011001101",
  4975=>"011101111",
  4976=>"111001101",
  4977=>"101101111",
  4978=>"011001000",
  4979=>"111111011",
  4980=>"010000100",
  4981=>"010100000",
  4982=>"010100010",
  4983=>"100101110",
  4984=>"100001110",
  4985=>"011110011",
  4986=>"011010000",
  4987=>"001101110",
  4988=>"001100000",
  4989=>"011111110",
  4990=>"100011001",
  4991=>"010011001",
  4992=>"101000010",
  4993=>"110111010",
  4994=>"010010101",
  4995=>"000110110",
  4996=>"000011010",
  4997=>"100001101",
  4998=>"001101101",
  4999=>"001001011",
  5000=>"010111100",
  5001=>"111011100",
  5002=>"111110010",
  5003=>"000110001",
  5004=>"100010001",
  5005=>"001110001",
  5006=>"110001010",
  5007=>"011011001",
  5008=>"001001111",
  5009=>"001111011",
  5010=>"000000100",
  5011=>"110111000",
  5012=>"000000100",
  5013=>"100000100",
  5014=>"101000010",
  5015=>"101111100",
  5016=>"000010111",
  5017=>"101000110",
  5018=>"100100110",
  5019=>"000000111",
  5020=>"001110000",
  5021=>"111100100",
  5022=>"011000111",
  5023=>"000001111",
  5024=>"100011110",
  5025=>"110000000",
  5026=>"001100100",
  5027=>"000100000",
  5028=>"001000000",
  5029=>"100111111",
  5030=>"101000000",
  5031=>"110010000",
  5032=>"111001000",
  5033=>"011111110",
  5034=>"100101101",
  5035=>"001110001",
  5036=>"101000001",
  5037=>"101111011",
  5038=>"100111000",
  5039=>"111001110",
  5040=>"001000101",
  5041=>"111110111",
  5042=>"000100011",
  5043=>"000000001",
  5044=>"100111010",
  5045=>"001110101",
  5046=>"110011010",
  5047=>"001110000",
  5048=>"101100101",
  5049=>"100010100",
  5050=>"001001001",
  5051=>"101111010",
  5052=>"110001110",
  5053=>"100010101",
  5054=>"110001010",
  5055=>"000000010",
  5056=>"011010110",
  5057=>"010001011",
  5058=>"010111100",
  5059=>"010001011",
  5060=>"100101011",
  5061=>"010100100",
  5062=>"000110100",
  5063=>"111010101",
  5064=>"100000000",
  5065=>"101100100",
  5066=>"100000011",
  5067=>"010001011",
  5068=>"100100101",
  5069=>"001001011",
  5070=>"110000100",
  5071=>"110000000",
  5072=>"110011000",
  5073=>"011000111",
  5074=>"110001011",
  5075=>"011100000",
  5076=>"011010001",
  5077=>"100000110",
  5078=>"011000001",
  5079=>"110110000",
  5080=>"100010101",
  5081=>"010000110",
  5082=>"011000100",
  5083=>"100000010",
  5084=>"110010001",
  5085=>"100111110",
  5086=>"100101100",
  5087=>"001011101",
  5088=>"011101010",
  5089=>"000101111",
  5090=>"110001010",
  5091=>"100011001",
  5092=>"001010100",
  5093=>"000010110",
  5094=>"011110000",
  5095=>"001000100",
  5096=>"000100100",
  5097=>"010100100",
  5098=>"100101110",
  5099=>"000101010",
  5100=>"110000111",
  5101=>"101000001",
  5102=>"111010101",
  5103=>"010000110",
  5104=>"000100101",
  5105=>"010111100",
  5106=>"101011100",
  5107=>"000111110",
  5108=>"001001000",
  5109=>"011010000",
  5110=>"001110101",
  5111=>"100110111",
  5112=>"001101011",
  5113=>"110100011",
  5114=>"100010111",
  5115=>"101111101",
  5116=>"001000010",
  5117=>"000001011",
  5118=>"110011000",
  5119=>"110101001",
  5120=>"101110100",
  5121=>"001101000",
  5122=>"100101100",
  5123=>"110111001",
  5124=>"010001011",
  5125=>"010001001",
  5126=>"000011100",
  5127=>"111100110",
  5128=>"100001000",
  5129=>"111111001",
  5130=>"010111101",
  5131=>"001011011",
  5132=>"000101101",
  5133=>"111011100",
  5134=>"011001101",
  5135=>"011001100",
  5136=>"011000111",
  5137=>"000101101",
  5138=>"000100010",
  5139=>"000010011",
  5140=>"111111100",
  5141=>"010000001",
  5142=>"000111001",
  5143=>"101110001",
  5144=>"110110011",
  5145=>"110000010",
  5146=>"101001000",
  5147=>"011001101",
  5148=>"100001111",
  5149=>"011010100",
  5150=>"101011100",
  5151=>"010011010",
  5152=>"111101000",
  5153=>"110111110",
  5154=>"110110011",
  5155=>"001000110",
  5156=>"010000100",
  5157=>"110011000",
  5158=>"001001101",
  5159=>"000001010",
  5160=>"000110110",
  5161=>"001111100",
  5162=>"001111010",
  5163=>"111001001",
  5164=>"101000100",
  5165=>"110001110",
  5166=>"001110000",
  5167=>"010000001",
  5168=>"110100100",
  5169=>"010101010",
  5170=>"100001001",
  5171=>"000010000",
  5172=>"000000110",
  5173=>"000000110",
  5174=>"001000110",
  5175=>"110101011",
  5176=>"001111011",
  5177=>"000111000",
  5178=>"111100001",
  5179=>"100000000",
  5180=>"001011100",
  5181=>"001000101",
  5182=>"011101101",
  5183=>"111101000",
  5184=>"010111010",
  5185=>"100000100",
  5186=>"000111111",
  5187=>"001100010",
  5188=>"001001110",
  5189=>"001011001",
  5190=>"111001001",
  5191=>"101100100",
  5192=>"110100111",
  5193=>"110011000",
  5194=>"110110001",
  5195=>"010000100",
  5196=>"111100100",
  5197=>"010111100",
  5198=>"011100111",
  5199=>"001001011",
  5200=>"000010111",
  5201=>"100010100",
  5202=>"001111011",
  5203=>"110101111",
  5204=>"100101000",
  5205=>"000010111",
  5206=>"110010101",
  5207=>"100001000",
  5208=>"010010110",
  5209=>"011101101",
  5210=>"001110111",
  5211=>"101100011",
  5212=>"011010000",
  5213=>"101001010",
  5214=>"011001100",
  5215=>"000000011",
  5216=>"010111100",
  5217=>"110011100",
  5218=>"100000001",
  5219=>"000010110",
  5220=>"001000000",
  5221=>"000111111",
  5222=>"000111011",
  5223=>"110011111",
  5224=>"100100010",
  5225=>"100000000",
  5226=>"001100100",
  5227=>"110010111",
  5228=>"100010001",
  5229=>"011110111",
  5230=>"001001000",
  5231=>"111011000",
  5232=>"001110111",
  5233=>"000101111",
  5234=>"001110000",
  5235=>"100010110",
  5236=>"111110001",
  5237=>"000101000",
  5238=>"011101110",
  5239=>"011100000",
  5240=>"101111100",
  5241=>"001100111",
  5242=>"011010000",
  5243=>"111101100",
  5244=>"100010110",
  5245=>"001110111",
  5246=>"011101001",
  5247=>"000000100",
  5248=>"111110110",
  5249=>"100000011",
  5250=>"000101100",
  5251=>"001101001",
  5252=>"010001100",
  5253=>"010110011",
  5254=>"011110101",
  5255=>"011110001",
  5256=>"001000000",
  5257=>"111111111",
  5258=>"100001000",
  5259=>"011000110",
  5260=>"101101100",
  5261=>"010110101",
  5262=>"001101001",
  5263=>"101011010",
  5264=>"010011011",
  5265=>"011001110",
  5266=>"111100000",
  5267=>"000011100",
  5268=>"100011110",
  5269=>"111101111",
  5270=>"101010001",
  5271=>"111000011",
  5272=>"000001001",
  5273=>"111010011",
  5274=>"011001011",
  5275=>"011110110",
  5276=>"110111010",
  5277=>"111011000",
  5278=>"101000100",
  5279=>"000010101",
  5280=>"111100000",
  5281=>"000001011",
  5282=>"011111110",
  5283=>"001110111",
  5284=>"101010111",
  5285=>"010101000",
  5286=>"000100000",
  5287=>"011111110",
  5288=>"010110101",
  5289=>"100110000",
  5290=>"101010101",
  5291=>"111000111",
  5292=>"001100101",
  5293=>"100000001",
  5294=>"110110000",
  5295=>"011011111",
  5296=>"101100110",
  5297=>"010010000",
  5298=>"000110101",
  5299=>"010101100",
  5300=>"001101000",
  5301=>"111101011",
  5302=>"111011111",
  5303=>"011000011",
  5304=>"000011110",
  5305=>"110101111",
  5306=>"100000010",
  5307=>"010010101",
  5308=>"001001001",
  5309=>"010100010",
  5310=>"111001001",
  5311=>"111100010",
  5312=>"110100001",
  5313=>"100101101",
  5314=>"110101101",
  5315=>"100000100",
  5316=>"001000000",
  5317=>"001111011",
  5318=>"000000001",
  5319=>"100000100",
  5320=>"101011100",
  5321=>"011011010",
  5322=>"100001100",
  5323=>"000101000",
  5324=>"001100010",
  5325=>"000000100",
  5326=>"001001111",
  5327=>"100100111",
  5328=>"100000011",
  5329=>"010101010",
  5330=>"011000100",
  5331=>"110011010",
  5332=>"110101101",
  5333=>"011001010",
  5334=>"000100011",
  5335=>"110010001",
  5336=>"111100100",
  5337=>"010011011",
  5338=>"111011100",
  5339=>"011110111",
  5340=>"100101111",
  5341=>"100000011",
  5342=>"110111011",
  5343=>"110010001",
  5344=>"000110001",
  5345=>"001110010",
  5346=>"111110111",
  5347=>"000100010",
  5348=>"111001110",
  5349=>"011011000",
  5350=>"100010100",
  5351=>"010100000",
  5352=>"110011111",
  5353=>"100011000",
  5354=>"011100000",
  5355=>"011000001",
  5356=>"011001001",
  5357=>"000010111",
  5358=>"001000111",
  5359=>"100011001",
  5360=>"001110010",
  5361=>"110010011",
  5362=>"001010111",
  5363=>"011100111",
  5364=>"001110100",
  5365=>"101111011",
  5366=>"000001000",
  5367=>"110110110",
  5368=>"100100010",
  5369=>"000110111",
  5370=>"110000000",
  5371=>"111001001",
  5372=>"111011010",
  5373=>"001101000",
  5374=>"110111110",
  5375=>"100001001",
  5376=>"100011110",
  5377=>"101110010",
  5378=>"011010000",
  5379=>"011001100",
  5380=>"100110010",
  5381=>"111111110",
  5382=>"110011100",
  5383=>"000011000",
  5384=>"110000000",
  5385=>"111111010",
  5386=>"011011100",
  5387=>"101101111",
  5388=>"011001010",
  5389=>"110110111",
  5390=>"111000000",
  5391=>"100000001",
  5392=>"111001000",
  5393=>"110011110",
  5394=>"110110101",
  5395=>"000000101",
  5396=>"111100001",
  5397=>"010000101",
  5398=>"000111111",
  5399=>"000011010",
  5400=>"010100001",
  5401=>"101100101",
  5402=>"001000010",
  5403=>"001001101",
  5404=>"110111001",
  5405=>"000000001",
  5406=>"011001010",
  5407=>"000000110",
  5408=>"000010001",
  5409=>"101101010",
  5410=>"110110001",
  5411=>"111011101",
  5412=>"111001011",
  5413=>"110010010",
  5414=>"010011101",
  5415=>"111000110",
  5416=>"000011110",
  5417=>"100110111",
  5418=>"110011011",
  5419=>"010101110",
  5420=>"100000011",
  5421=>"001100110",
  5422=>"010111000",
  5423=>"100010001",
  5424=>"110100110",
  5425=>"000000100",
  5426=>"001111001",
  5427=>"011000001",
  5428=>"000110111",
  5429=>"001110010",
  5430=>"110001000",
  5431=>"111001000",
  5432=>"100100110",
  5433=>"100100110",
  5434=>"111011111",
  5435=>"001100010",
  5436=>"110000011",
  5437=>"110010111",
  5438=>"001001001",
  5439=>"001010000",
  5440=>"011101100",
  5441=>"001010100",
  5442=>"000011000",
  5443=>"101010100",
  5444=>"100100100",
  5445=>"110001111",
  5446=>"001110011",
  5447=>"000000101",
  5448=>"111111110",
  5449=>"011110101",
  5450=>"010011001",
  5451=>"001011001",
  5452=>"111010111",
  5453=>"100111011",
  5454=>"100111110",
  5455=>"000011111",
  5456=>"111110011",
  5457=>"110101110",
  5458=>"010000100",
  5459=>"010000101",
  5460=>"001110010",
  5461=>"010010100",
  5462=>"110001000",
  5463=>"010010100",
  5464=>"101010100",
  5465=>"111110110",
  5466=>"010001000",
  5467=>"101101100",
  5468=>"010111001",
  5469=>"010000011",
  5470=>"000110010",
  5471=>"101101010",
  5472=>"010100001",
  5473=>"010000000",
  5474=>"111000001",
  5475=>"000110001",
  5476=>"100000100",
  5477=>"011101100",
  5478=>"100100001",
  5479=>"000001001",
  5480=>"101111101",
  5481=>"010011101",
  5482=>"010101010",
  5483=>"111000010",
  5484=>"111111100",
  5485=>"001001001",
  5486=>"100001111",
  5487=>"101110000",
  5488=>"100001010",
  5489=>"100100010",
  5490=>"010110100",
  5491=>"011011111",
  5492=>"101101000",
  5493=>"100011011",
  5494=>"000100001",
  5495=>"100101010",
  5496=>"000110011",
  5497=>"100110000",
  5498=>"111011111",
  5499=>"010100110",
  5500=>"110110100",
  5501=>"111000001",
  5502=>"100011101",
  5503=>"011011110",
  5504=>"001000111",
  5505=>"000011000",
  5506=>"011001111",
  5507=>"000100011",
  5508=>"110111010",
  5509=>"100100100",
  5510=>"010101110",
  5511=>"011100101",
  5512=>"000010011",
  5513=>"100001111",
  5514=>"011010101",
  5515=>"111111101",
  5516=>"000000100",
  5517=>"111000001",
  5518=>"010110101",
  5519=>"100011001",
  5520=>"110100111",
  5521=>"111111110",
  5522=>"011010011",
  5523=>"011001101",
  5524=>"110011001",
  5525=>"111011111",
  5526=>"100100101",
  5527=>"011111000",
  5528=>"100110011",
  5529=>"011101111",
  5530=>"100100111",
  5531=>"011010101",
  5532=>"111101000",
  5533=>"011001010",
  5534=>"000010001",
  5535=>"101100010",
  5536=>"100010010",
  5537=>"000010001",
  5538=>"001000100",
  5539=>"110110101",
  5540=>"000111110",
  5541=>"000111100",
  5542=>"001010010",
  5543=>"100111110",
  5544=>"110101100",
  5545=>"101111110",
  5546=>"010110110",
  5547=>"011101100",
  5548=>"011010111",
  5549=>"000010000",
  5550=>"010000111",
  5551=>"100011101",
  5552=>"000111110",
  5553=>"100010010",
  5554=>"110111101",
  5555=>"000000111",
  5556=>"110010101",
  5557=>"101001110",
  5558=>"000011001",
  5559=>"001010100",
  5560=>"110001011",
  5561=>"100011101",
  5562=>"001001111",
  5563=>"001000110",
  5564=>"100101011",
  5565=>"011101010",
  5566=>"000111100",
  5567=>"000001011",
  5568=>"101000000",
  5569=>"100010010",
  5570=>"000000000",
  5571=>"110110011",
  5572=>"011100110",
  5573=>"101101110",
  5574=>"011111101",
  5575=>"000110111",
  5576=>"010001111",
  5577=>"100110100",
  5578=>"111110011",
  5579=>"011010110",
  5580=>"111010101",
  5581=>"001010110",
  5582=>"110101001",
  5583=>"001111111",
  5584=>"110010010",
  5585=>"111001000",
  5586=>"000011101",
  5587=>"000001100",
  5588=>"010101000",
  5589=>"000001100",
  5590=>"100011001",
  5591=>"010111000",
  5592=>"011000000",
  5593=>"101011110",
  5594=>"000000100",
  5595=>"000100010",
  5596=>"111011111",
  5597=>"111101001",
  5598=>"011000101",
  5599=>"011011011",
  5600=>"010100110",
  5601=>"101001110",
  5602=>"000000000",
  5603=>"101000101",
  5604=>"011001101",
  5605=>"000011010",
  5606=>"011011000",
  5607=>"100000010",
  5608=>"100011101",
  5609=>"100011100",
  5610=>"111101101",
  5611=>"011100010",
  5612=>"010111001",
  5613=>"111010100",
  5614=>"101001111",
  5615=>"011010100",
  5616=>"111010001",
  5617=>"001111110",
  5618=>"111110001",
  5619=>"000101010",
  5620=>"011101110",
  5621=>"010100001",
  5622=>"101100111",
  5623=>"000001000",
  5624=>"100011001",
  5625=>"110001011",
  5626=>"111011100",
  5627=>"110100100",
  5628=>"110110101",
  5629=>"111100010",
  5630=>"100011011",
  5631=>"110100010",
  5632=>"011110000",
  5633=>"011000100",
  5634=>"011010101",
  5635=>"001011100",
  5636=>"010111100",
  5637=>"101011110",
  5638=>"011011110",
  5639=>"111100010",
  5640=>"010111110",
  5641=>"010110100",
  5642=>"100111101",
  5643=>"011011010",
  5644=>"101100110",
  5645=>"010110101",
  5646=>"100101011",
  5647=>"110110111",
  5648=>"101010011",
  5649=>"100111011",
  5650=>"101011110",
  5651=>"011110011",
  5652=>"010011111",
  5653=>"110110000",
  5654=>"000001111",
  5655=>"000100010",
  5656=>"011101010",
  5657=>"001101100",
  5658=>"000000000",
  5659=>"100001010",
  5660=>"101011111",
  5661=>"100110111",
  5662=>"000100011",
  5663=>"011101101",
  5664=>"001000111",
  5665=>"111100010",
  5666=>"101000000",
  5667=>"100010010",
  5668=>"111110000",
  5669=>"000000011",
  5670=>"100011000",
  5671=>"110001100",
  5672=>"001000111",
  5673=>"101011101",
  5674=>"011111101",
  5675=>"010011100",
  5676=>"011110001",
  5677=>"110000001",
  5678=>"001111011",
  5679=>"111101111",
  5680=>"011101111",
  5681=>"111111110",
  5682=>"010111100",
  5683=>"101011110",
  5684=>"111111001",
  5685=>"110001010",
  5686=>"011001101",
  5687=>"001100111",
  5688=>"100001101",
  5689=>"101110011",
  5690=>"011100100",
  5691=>"010100010",
  5692=>"110101000",
  5693=>"111010011",
  5694=>"001000101",
  5695=>"001100011",
  5696=>"101110000",
  5697=>"101000010",
  5698=>"001000011",
  5699=>"111001100",
  5700=>"001001000",
  5701=>"000111101",
  5702=>"000100101",
  5703=>"001101010",
  5704=>"011101011",
  5705=>"110011111",
  5706=>"000101000",
  5707=>"011011101",
  5708=>"111010101",
  5709=>"011011110",
  5710=>"001010010",
  5711=>"010100110",
  5712=>"110110110",
  5713=>"011111000",
  5714=>"000000100",
  5715=>"000001000",
  5716=>"010001011",
  5717=>"001010110",
  5718=>"111011110",
  5719=>"100001101",
  5720=>"111101111",
  5721=>"110101011",
  5722=>"110001010",
  5723=>"000101101",
  5724=>"001100001",
  5725=>"111010100",
  5726=>"111100011",
  5727=>"011010101",
  5728=>"001000110",
  5729=>"001010110",
  5730=>"101000100",
  5731=>"001100000",
  5732=>"101000111",
  5733=>"111110001",
  5734=>"000100001",
  5735=>"010100011",
  5736=>"010001101",
  5737=>"000100110",
  5738=>"001100101",
  5739=>"001001111",
  5740=>"111110101",
  5741=>"101101110",
  5742=>"010001101",
  5743=>"000110100",
  5744=>"110000101",
  5745=>"001001111",
  5746=>"000010001",
  5747=>"101100001",
  5748=>"100011000",
  5749=>"100010110",
  5750=>"111111101",
  5751=>"110101111",
  5752=>"010100111",
  5753=>"011001100",
  5754=>"111100001",
  5755=>"110111100",
  5756=>"011010100",
  5757=>"000100011",
  5758=>"111111111",
  5759=>"000111111",
  5760=>"101010100",
  5761=>"110011000",
  5762=>"100010010",
  5763=>"101010001",
  5764=>"010100010",
  5765=>"011101101",
  5766=>"110001100",
  5767=>"011010001",
  5768=>"110000101",
  5769=>"010010111",
  5770=>"111111000",
  5771=>"001001111",
  5772=>"101011000",
  5773=>"010101110",
  5774=>"001110011",
  5775=>"010010010",
  5776=>"110000000",
  5777=>"000100000",
  5778=>"100011000",
  5779=>"100100011",
  5780=>"011101110",
  5781=>"000111110",
  5782=>"000101111",
  5783=>"100000110",
  5784=>"100010000",
  5785=>"110010110",
  5786=>"000001111",
  5787=>"111000001",
  5788=>"011010010",
  5789=>"101010111",
  5790=>"101011110",
  5791=>"111101111",
  5792=>"101000011",
  5793=>"011001011",
  5794=>"000110101",
  5795=>"110001001",
  5796=>"011000100",
  5797=>"011000000",
  5798=>"010110010",
  5799=>"101101111",
  5800=>"110001101",
  5801=>"010101011",
  5802=>"000000001",
  5803=>"010111111",
  5804=>"110111100",
  5805=>"100001001",
  5806=>"100110011",
  5807=>"100101010",
  5808=>"000000000",
  5809=>"110110001",
  5810=>"000101101",
  5811=>"101000100",
  5812=>"111000101",
  5813=>"101100100",
  5814=>"000011001",
  5815=>"110010101",
  5816=>"101100010",
  5817=>"110000110",
  5818=>"000110000",
  5819=>"110010000",
  5820=>"000111010",
  5821=>"110110110",
  5822=>"010001011",
  5823=>"110100111",
  5824=>"111000000",
  5825=>"011010101",
  5826=>"000000111",
  5827=>"111111111",
  5828=>"001001011",
  5829=>"111000011",
  5830=>"101010110",
  5831=>"001000001",
  5832=>"010101110",
  5833=>"011001100",
  5834=>"101100100",
  5835=>"101011111",
  5836=>"111110010",
  5837=>"101001001",
  5838=>"000101100",
  5839=>"000111111",
  5840=>"101100100",
  5841=>"011001111",
  5842=>"010010010",
  5843=>"100110010",
  5844=>"000001000",
  5845=>"101010110",
  5846=>"010111110",
  5847=>"010100011",
  5848=>"010010000",
  5849=>"001111111",
  5850=>"110111001",
  5851=>"011000011",
  5852=>"000000011",
  5853=>"010100101",
  5854=>"100010011",
  5855=>"000010111",
  5856=>"000100011",
  5857=>"010001000",
  5858=>"100100001",
  5859=>"111011101",
  5860=>"011101100",
  5861=>"010100101",
  5862=>"001011010",
  5863=>"010011001",
  5864=>"110011010",
  5865=>"110110010",
  5866=>"000101111",
  5867=>"010000100",
  5868=>"011100111",
  5869=>"001001001",
  5870=>"111101110",
  5871=>"011000011",
  5872=>"101001110",
  5873=>"000010010",
  5874=>"111101110",
  5875=>"011110111",
  5876=>"000110011",
  5877=>"001110110",
  5878=>"101001101",
  5879=>"010000111",
  5880=>"101100001",
  5881=>"000010011",
  5882=>"011000100",
  5883=>"100110101",
  5884=>"101110011",
  5885=>"001001100",
  5886=>"110011100",
  5887=>"001100101",
  5888=>"100111010",
  5889=>"000000111",
  5890=>"010001000",
  5891=>"010111000",
  5892=>"010111100",
  5893=>"110111101",
  5894=>"001001100",
  5895=>"001100110",
  5896=>"100000001",
  5897=>"110101111",
  5898=>"101110100",
  5899=>"100000001",
  5900=>"110000100",
  5901=>"011100101",
  5902=>"111011001",
  5903=>"110100110",
  5904=>"110010111",
  5905=>"001101011",
  5906=>"101101111",
  5907=>"111000011",
  5908=>"010011100",
  5909=>"100010000",
  5910=>"010011110",
  5911=>"011110001",
  5912=>"010100110",
  5913=>"100001000",
  5914=>"110000111",
  5915=>"100101011",
  5916=>"100100000",
  5917=>"111111111",
  5918=>"111001100",
  5919=>"011110110",
  5920=>"111100101",
  5921=>"111000011",
  5922=>"000001001",
  5923=>"010011110",
  5924=>"001010101",
  5925=>"001101110",
  5926=>"111111111",
  5927=>"010101000",
  5928=>"100100011",
  5929=>"110111010",
  5930=>"000010110",
  5931=>"100110000",
  5932=>"100000111",
  5933=>"000111111",
  5934=>"110100010",
  5935=>"001010101",
  5936=>"110001110",
  5937=>"110111011",
  5938=>"110001101",
  5939=>"111001110",
  5940=>"111111110",
  5941=>"011100001",
  5942=>"000101110",
  5943=>"000010010",
  5944=>"101011110",
  5945=>"100001011",
  5946=>"000000100",
  5947=>"001000001",
  5948=>"101110011",
  5949=>"100100110",
  5950=>"111110111",
  5951=>"101110001",
  5952=>"111001001",
  5953=>"110001110",
  5954=>"101001110",
  5955=>"111100001",
  5956=>"011101001",
  5957=>"001111001",
  5958=>"111110011",
  5959=>"100100111",
  5960=>"100011001",
  5961=>"100100100",
  5962=>"010110000",
  5963=>"110000111",
  5964=>"010011111",
  5965=>"001100100",
  5966=>"110010010",
  5967=>"110100101",
  5968=>"001000001",
  5969=>"000011000",
  5970=>"000100011",
  5971=>"010000100",
  5972=>"111011011",
  5973=>"101010011",
  5974=>"010001000",
  5975=>"100000111",
  5976=>"101101100",
  5977=>"111001011",
  5978=>"100110011",
  5979=>"000000110",
  5980=>"000100111",
  5981=>"110100101",
  5982=>"100011000",
  5983=>"010000110",
  5984=>"101000011",
  5985=>"001000110",
  5986=>"100110000",
  5987=>"010111111",
  5988=>"001111101",
  5989=>"110100100",
  5990=>"110010010",
  5991=>"010011110",
  5992=>"010110011",
  5993=>"010001111",
  5994=>"000010010",
  5995=>"101111011",
  5996=>"010000000",
  5997=>"011100000",
  5998=>"001000101",
  5999=>"100000101",
  6000=>"011011111",
  6001=>"100111110",
  6002=>"110010101",
  6003=>"010011101",
  6004=>"110100110",
  6005=>"000111100",
  6006=>"001100101",
  6007=>"101000010",
  6008=>"110000000",
  6009=>"101011100",
  6010=>"101110111",
  6011=>"101000001",
  6012=>"101000001",
  6013=>"100010010",
  6014=>"100000100",
  6015=>"011111101",
  6016=>"000100110",
  6017=>"010110110",
  6018=>"110000010",
  6019=>"110111111",
  6020=>"010111101",
  6021=>"010010000",
  6022=>"100111001",
  6023=>"000111101",
  6024=>"101000001",
  6025=>"101101000",
  6026=>"011110001",
  6027=>"010100011",
  6028=>"000100100",
  6029=>"000101101",
  6030=>"000100001",
  6031=>"101010110",
  6032=>"100100001",
  6033=>"001100000",
  6034=>"100110000",
  6035=>"011010101",
  6036=>"010100001",
  6037=>"101010000",
  6038=>"010010101",
  6039=>"010000110",
  6040=>"011101101",
  6041=>"010011000",
  6042=>"111001100",
  6043=>"111011011",
  6044=>"010111011",
  6045=>"001111111",
  6046=>"110101111",
  6047=>"011111110",
  6048=>"110110011",
  6049=>"001000011",
  6050=>"000000101",
  6051=>"001100110",
  6052=>"110100110",
  6053=>"010101001",
  6054=>"010111101",
  6055=>"100000000",
  6056=>"111001010",
  6057=>"011010110",
  6058=>"001111101",
  6059=>"101011111",
  6060=>"110110101",
  6061=>"111001111",
  6062=>"011000011",
  6063=>"000000000",
  6064=>"000000000",
  6065=>"000011000",
  6066=>"011101001",
  6067=>"110001011",
  6068=>"011010000",
  6069=>"101100101",
  6070=>"011011001",
  6071=>"110100010",
  6072=>"100100010",
  6073=>"100010111",
  6074=>"000011110",
  6075=>"110101001",
  6076=>"111100001",
  6077=>"001111001",
  6078=>"111101111",
  6079=>"000011101",
  6080=>"000111000",
  6081=>"110000100",
  6082=>"011100101",
  6083=>"111001111",
  6084=>"101110111",
  6085=>"110010000",
  6086=>"010100110",
  6087=>"000100110",
  6088=>"110000111",
  6089=>"010010001",
  6090=>"110101010",
  6091=>"110100111",
  6092=>"110011101",
  6093=>"010001100",
  6094=>"001110000",
  6095=>"001110100",
  6096=>"000100100",
  6097=>"101110100",
  6098=>"111111000",
  6099=>"101101111",
  6100=>"101100101",
  6101=>"110101001",
  6102=>"000110110",
  6103=>"000101011",
  6104=>"001000011",
  6105=>"011110110",
  6106=>"001111100",
  6107=>"011100110",
  6108=>"110111011",
  6109=>"110111110",
  6110=>"100110101",
  6111=>"011000101",
  6112=>"100011011",
  6113=>"110000100",
  6114=>"100101010",
  6115=>"001110110",
  6116=>"101000000",
  6117=>"111111100",
  6118=>"111010100",
  6119=>"000011111",
  6120=>"101110000",
  6121=>"001000001",
  6122=>"100000000",
  6123=>"100100110",
  6124=>"011111011",
  6125=>"100110110",
  6126=>"001000010",
  6127=>"101100111",
  6128=>"000111110",
  6129=>"011111001",
  6130=>"100110011",
  6131=>"001100100",
  6132=>"001000110",
  6133=>"000010111",
  6134=>"010000010",
  6135=>"011011001",
  6136=>"011100000",
  6137=>"101110110",
  6138=>"110001001",
  6139=>"101010000",
  6140=>"001010101",
  6141=>"010010100",
  6142=>"100110101",
  6143=>"110010000",
  6144=>"101001111",
  6145=>"101110000",
  6146=>"011010100",
  6147=>"010110110",
  6148=>"000100100",
  6149=>"101011101",
  6150=>"011001110",
  6151=>"110001011",
  6152=>"001110010",
  6153=>"000010110",
  6154=>"101101001",
  6155=>"111100101",
  6156=>"110101000",
  6157=>"100101111",
  6158=>"100011000",
  6159=>"111111011",
  6160=>"100011100",
  6161=>"001111111",
  6162=>"111001100",
  6163=>"100001010",
  6164=>"101101011",
  6165=>"110111111",
  6166=>"000110000",
  6167=>"111100010",
  6168=>"000110101",
  6169=>"000101001",
  6170=>"111110111",
  6171=>"011111100",
  6172=>"001110010",
  6173=>"101100110",
  6174=>"011011100",
  6175=>"101000011",
  6176=>"001101111",
  6177=>"110010011",
  6178=>"111010110",
  6179=>"000100000",
  6180=>"110001010",
  6181=>"111111011",
  6182=>"111011111",
  6183=>"101011111",
  6184=>"001100100",
  6185=>"001011110",
  6186=>"100000101",
  6187=>"001101001",
  6188=>"010111000",
  6189=>"110011011",
  6190=>"100111001",
  6191=>"001001110",
  6192=>"101100000",
  6193=>"111100001",
  6194=>"111101110",
  6195=>"000100001",
  6196=>"100101100",
  6197=>"001110111",
  6198=>"100001001",
  6199=>"101100100",
  6200=>"100101101",
  6201=>"000110111",
  6202=>"101011000",
  6203=>"101111101",
  6204=>"111011010",
  6205=>"111101011",
  6206=>"010010111",
  6207=>"110001101",
  6208=>"000011101",
  6209=>"100101001",
  6210=>"110001001",
  6211=>"011100101",
  6212=>"101000111",
  6213=>"010001101",
  6214=>"111111011",
  6215=>"111000000",
  6216=>"100100110",
  6217=>"110001111",
  6218=>"100001001",
  6219=>"000000100",
  6220=>"110001010",
  6221=>"111100000",
  6222=>"111111000",
  6223=>"100111110",
  6224=>"100101111",
  6225=>"110011011",
  6226=>"011011111",
  6227=>"111101001",
  6228=>"011001010",
  6229=>"011111010",
  6230=>"011001101",
  6231=>"101111000",
  6232=>"111001111",
  6233=>"001101011",
  6234=>"100100110",
  6235=>"001001001",
  6236=>"110100111",
  6237=>"100111111",
  6238=>"011100110",
  6239=>"110110110",
  6240=>"011001011",
  6241=>"000000110",
  6242=>"101001011",
  6243=>"000011000",
  6244=>"001111110",
  6245=>"111011011",
  6246=>"110000010",
  6247=>"101001000",
  6248=>"111110111",
  6249=>"111010111",
  6250=>"000010101",
  6251=>"001010110",
  6252=>"000010101",
  6253=>"001101011",
  6254=>"101100000",
  6255=>"111010110",
  6256=>"110111001",
  6257=>"010010111",
  6258=>"010001111",
  6259=>"000100000",
  6260=>"001011111",
  6261=>"011111010",
  6262=>"011110000",
  6263=>"111100101",
  6264=>"010111110",
  6265=>"000001001",
  6266=>"010101001",
  6267=>"111001011",
  6268=>"001111101",
  6269=>"100011010",
  6270=>"101101111",
  6271=>"000010111",
  6272=>"000010000",
  6273=>"011111100",
  6274=>"010010111",
  6275=>"010100100",
  6276=>"111100011",
  6277=>"111100010",
  6278=>"000001101",
  6279=>"000110000",
  6280=>"000001111",
  6281=>"110101111",
  6282=>"100101110",
  6283=>"110001000",
  6284=>"001111001",
  6285=>"101011011",
  6286=>"100110010",
  6287=>"101000101",
  6288=>"101101011",
  6289=>"101101010",
  6290=>"001101100",
  6291=>"000010101",
  6292=>"011101111",
  6293=>"001001001",
  6294=>"011000001",
  6295=>"100101000",
  6296=>"011111100",
  6297=>"000001010",
  6298=>"001011000",
  6299=>"110110111",
  6300=>"100010011",
  6301=>"000101100",
  6302=>"011100100",
  6303=>"101111110",
  6304=>"001110011",
  6305=>"100001110",
  6306=>"110010100",
  6307=>"100101100",
  6308=>"010000111",
  6309=>"011010011",
  6310=>"110010000",
  6311=>"001110101",
  6312=>"110011100",
  6313=>"010110110",
  6314=>"001101011",
  6315=>"101111001",
  6316=>"001101000",
  6317=>"000110001",
  6318=>"010101101",
  6319=>"000100010",
  6320=>"011101101",
  6321=>"000111010",
  6322=>"000111111",
  6323=>"011111101",
  6324=>"001101000",
  6325=>"011000110",
  6326=>"110111110",
  6327=>"011001000",
  6328=>"101110100",
  6329=>"100010000",
  6330=>"101000101",
  6331=>"111000111",
  6332=>"001000101",
  6333=>"111101100",
  6334=>"001000100",
  6335=>"010001101",
  6336=>"100100011",
  6337=>"011110011",
  6338=>"111001101",
  6339=>"000010010",
  6340=>"100001001",
  6341=>"010100010",
  6342=>"011110110",
  6343=>"011000111",
  6344=>"111000001",
  6345=>"100111000",
  6346=>"010100100",
  6347=>"101110010",
  6348=>"100011110",
  6349=>"010000010",
  6350=>"111001111",
  6351=>"100000111",
  6352=>"101100011",
  6353=>"011100101",
  6354=>"011100110",
  6355=>"001110111",
  6356=>"001100110",
  6357=>"011111110",
  6358=>"100011011",
  6359=>"000101000",
  6360=>"010101110",
  6361=>"000101000",
  6362=>"101000100",
  6363=>"101111111",
  6364=>"001110100",
  6365=>"001100011",
  6366=>"001100000",
  6367=>"001101000",
  6368=>"110101011",
  6369=>"011000010",
  6370=>"000001001",
  6371=>"101111001",
  6372=>"100110010",
  6373=>"000101010",
  6374=>"100111110",
  6375=>"110001010",
  6376=>"100000111",
  6377=>"001011111",
  6378=>"001011100",
  6379=>"010100000",
  6380=>"010000100",
  6381=>"110101011",
  6382=>"001000011",
  6383=>"010100011",
  6384=>"001101111",
  6385=>"010100100",
  6386=>"010100001",
  6387=>"100011011",
  6388=>"101111011",
  6389=>"110000100",
  6390=>"010001000",
  6391=>"000000100",
  6392=>"110001111",
  6393=>"110101000",
  6394=>"110011000",
  6395=>"110001010",
  6396=>"100111001",
  6397=>"101100000",
  6398=>"000000101",
  6399=>"111101000",
  6400=>"101110111",
  6401=>"000101001",
  6402=>"000010111",
  6403=>"010110100",
  6404=>"110000110",
  6405=>"011100101",
  6406=>"000000001",
  6407=>"111111101",
  6408=>"111010011",
  6409=>"000010001",
  6410=>"000010110",
  6411=>"000001010",
  6412=>"010001000",
  6413=>"111111111",
  6414=>"010000111",
  6415=>"100011110",
  6416=>"000111111",
  6417=>"101011110",
  6418=>"100010111",
  6419=>"111111010",
  6420=>"000111101",
  6421=>"011111100",
  6422=>"110100000",
  6423=>"111111010",
  6424=>"000010111",
  6425=>"110000101",
  6426=>"010011010",
  6427=>"011111010",
  6428=>"001000111",
  6429=>"111110110",
  6430=>"010100110",
  6431=>"000001010",
  6432=>"111000010",
  6433=>"111111011",
  6434=>"001111110",
  6435=>"000011100",
  6436=>"000011010",
  6437=>"110100001",
  6438=>"101101001",
  6439=>"101011001",
  6440=>"101101111",
  6441=>"010100101",
  6442=>"110011110",
  6443=>"110110111",
  6444=>"010001100",
  6445=>"011100000",
  6446=>"101111101",
  6447=>"011101101",
  6448=>"110001100",
  6449=>"000011000",
  6450=>"101011011",
  6451=>"111101111",
  6452=>"100110001",
  6453=>"100010110",
  6454=>"011110111",
  6455=>"100100110",
  6456=>"100000001",
  6457=>"111101111",
  6458=>"110100010",
  6459=>"000001011",
  6460=>"001011011",
  6461=>"101010101",
  6462=>"100100000",
  6463=>"100111010",
  6464=>"011111001",
  6465=>"110000100",
  6466=>"100001110",
  6467=>"100010001",
  6468=>"011101010",
  6469=>"000000110",
  6470=>"010110101",
  6471=>"100100100",
  6472=>"000001011",
  6473=>"001101010",
  6474=>"111111101",
  6475=>"111001000",
  6476=>"110100101",
  6477=>"000111110",
  6478=>"000100000",
  6479=>"011110011",
  6480=>"100110011",
  6481=>"110001010",
  6482=>"101111110",
  6483=>"100111011",
  6484=>"001011110",
  6485=>"100111011",
  6486=>"000111111",
  6487=>"000101000",
  6488=>"010000000",
  6489=>"100001100",
  6490=>"010000011",
  6491=>"101011100",
  6492=>"000001110",
  6493=>"111000100",
  6494=>"110001010",
  6495=>"000101111",
  6496=>"111000110",
  6497=>"000011100",
  6498=>"010000111",
  6499=>"111000010",
  6500=>"011111001",
  6501=>"000010100",
  6502=>"111101011",
  6503=>"010100101",
  6504=>"110010101",
  6505=>"111111110",
  6506=>"101011000",
  6507=>"010001011",
  6508=>"101100011",
  6509=>"000101010",
  6510=>"101010111",
  6511=>"010001101",
  6512=>"011110000",
  6513=>"111011110",
  6514=>"001101010",
  6515=>"001001001",
  6516=>"000101000",
  6517=>"101001100",
  6518=>"111111000",
  6519=>"101100101",
  6520=>"111100010",
  6521=>"100101001",
  6522=>"101100011",
  6523=>"011100111",
  6524=>"110111001",
  6525=>"010110100",
  6526=>"111110011",
  6527=>"100000100",
  6528=>"001100000",
  6529=>"011010100",
  6530=>"101000001",
  6531=>"000001100",
  6532=>"100111010",
  6533=>"100101001",
  6534=>"100010111",
  6535=>"100101000",
  6536=>"110101010",
  6537=>"101101111",
  6538=>"000000110",
  6539=>"111100100",
  6540=>"101000011",
  6541=>"010101111",
  6542=>"001110011",
  6543=>"011000000",
  6544=>"110000001",
  6545=>"110011001",
  6546=>"100001010",
  6547=>"011110011",
  6548=>"010110001",
  6549=>"000110001",
  6550=>"000001000",
  6551=>"001111010",
  6552=>"011000110",
  6553=>"110101000",
  6554=>"010011001",
  6555=>"101010110",
  6556=>"000010111",
  6557=>"011000101",
  6558=>"001100001",
  6559=>"101100010",
  6560=>"101101111",
  6561=>"001110100",
  6562=>"110000001",
  6563=>"001101100",
  6564=>"001010011",
  6565=>"110001010",
  6566=>"101011000",
  6567=>"000001010",
  6568=>"011000001",
  6569=>"000011000",
  6570=>"101001100",
  6571=>"110001001",
  6572=>"111110110",
  6573=>"000101010",
  6574=>"010100110",
  6575=>"110001001",
  6576=>"110110001",
  6577=>"111100101",
  6578=>"000010000",
  6579=>"000101111",
  6580=>"010010101",
  6581=>"001000101",
  6582=>"101010111",
  6583=>"100010111",
  6584=>"101011001",
  6585=>"100001001",
  6586=>"110001110",
  6587=>"111010011",
  6588=>"100110111",
  6589=>"101111100",
  6590=>"010101110",
  6591=>"110000000",
  6592=>"100110011",
  6593=>"110011111",
  6594=>"011100111",
  6595=>"000100101",
  6596=>"101100100",
  6597=>"000000111",
  6598=>"010110001",
  6599=>"011010100",
  6600=>"110011100",
  6601=>"000101001",
  6602=>"100101111",
  6603=>"100001001",
  6604=>"100100010",
  6605=>"110000101",
  6606=>"111111010",
  6607=>"001101101",
  6608=>"100010000",
  6609=>"111101000",
  6610=>"100001101",
  6611=>"101000101",
  6612=>"100000011",
  6613=>"111110101",
  6614=>"000110110",
  6615=>"111110000",
  6616=>"100011001",
  6617=>"001011111",
  6618=>"001110010",
  6619=>"010101100",
  6620=>"110111100",
  6621=>"011000110",
  6622=>"011001011",
  6623=>"100111001",
  6624=>"011101111",
  6625=>"100100110",
  6626=>"111010000",
  6627=>"111001010",
  6628=>"101001101",
  6629=>"110000001",
  6630=>"010110010",
  6631=>"110100011",
  6632=>"000010011",
  6633=>"001011010",
  6634=>"101101100",
  6635=>"011110011",
  6636=>"000010110",
  6637=>"101110111",
  6638=>"111110101",
  6639=>"101111011",
  6640=>"010111111",
  6641=>"010000010",
  6642=>"000001101",
  6643=>"000010100",
  6644=>"101000010",
  6645=>"110101000",
  6646=>"100011111",
  6647=>"001001100",
  6648=>"011101101",
  6649=>"101111001",
  6650=>"000100000",
  6651=>"000111000",
  6652=>"100111111",
  6653=>"101001110",
  6654=>"111010110",
  6655=>"110110010",
  6656=>"100010111",
  6657=>"111100100",
  6658=>"101111001",
  6659=>"100000100",
  6660=>"001100101",
  6661=>"111111010",
  6662=>"001100101",
  6663=>"110101001",
  6664=>"111101011",
  6665=>"100000011",
  6666=>"110000111",
  6667=>"000001100",
  6668=>"111110111",
  6669=>"101010001",
  6670=>"111101000",
  6671=>"000011000",
  6672=>"100110010",
  6673=>"110000010",
  6674=>"111011101",
  6675=>"011100101",
  6676=>"000000011",
  6677=>"101010110",
  6678=>"000110100",
  6679=>"000011110",
  6680=>"010000100",
  6681=>"010011110",
  6682=>"111100011",
  6683=>"100011011",
  6684=>"001001010",
  6685=>"101101110",
  6686=>"110011110",
  6687=>"101000011",
  6688=>"111010000",
  6689=>"000010101",
  6690=>"011001000",
  6691=>"110110000",
  6692=>"011010001",
  6693=>"010011100",
  6694=>"111101011",
  6695=>"111100101",
  6696=>"110111101",
  6697=>"101110101",
  6698=>"010000000",
  6699=>"011000000",
  6700=>"010100111",
  6701=>"110101110",
  6702=>"010000111",
  6703=>"000010000",
  6704=>"110111100",
  6705=>"110110001",
  6706=>"000001010",
  6707=>"011100100",
  6708=>"100010110",
  6709=>"110010101",
  6710=>"010110001",
  6711=>"110100010",
  6712=>"001010100",
  6713=>"011100011",
  6714=>"000001000",
  6715=>"101111001",
  6716=>"110101010",
  6717=>"000100000",
  6718=>"011001001",
  6719=>"101111101",
  6720=>"101101000",
  6721=>"111111101",
  6722=>"111000101",
  6723=>"010011100",
  6724=>"010000011",
  6725=>"001000111",
  6726=>"100110011",
  6727=>"110101011",
  6728=>"000111101",
  6729=>"110011101",
  6730=>"101110110",
  6731=>"111000000",
  6732=>"101110101",
  6733=>"100000110",
  6734=>"011101110",
  6735=>"010001110",
  6736=>"111001001",
  6737=>"101011111",
  6738=>"110110010",
  6739=>"111000111",
  6740=>"101100000",
  6741=>"101010111",
  6742=>"001110110",
  6743=>"110001011",
  6744=>"101111001",
  6745=>"001101111",
  6746=>"111000011",
  6747=>"110001100",
  6748=>"110001101",
  6749=>"111000101",
  6750=>"011101100",
  6751=>"000010101",
  6752=>"001010101",
  6753=>"000001111",
  6754=>"010011100",
  6755=>"011011001",
  6756=>"010100001",
  6757=>"100100100",
  6758=>"000100010",
  6759=>"000010110",
  6760=>"111111000",
  6761=>"010000111",
  6762=>"101111000",
  6763=>"010011100",
  6764=>"000111010",
  6765=>"100001000",
  6766=>"000100100",
  6767=>"000010011",
  6768=>"011010100",
  6769=>"111111001",
  6770=>"010100010",
  6771=>"011101110",
  6772=>"000101011",
  6773=>"110001000",
  6774=>"100100001",
  6775=>"011001100",
  6776=>"100110101",
  6777=>"110101000",
  6778=>"111111011",
  6779=>"001011101",
  6780=>"010111001",
  6781=>"111001110",
  6782=>"000101010",
  6783=>"010000001",
  6784=>"000001000",
  6785=>"000100111",
  6786=>"101101110",
  6787=>"100101110",
  6788=>"101110110",
  6789=>"110000011",
  6790=>"000001101",
  6791=>"101110101",
  6792=>"100011000",
  6793=>"001000111",
  6794=>"110000000",
  6795=>"011011010",
  6796=>"011101001",
  6797=>"100011011",
  6798=>"110101000",
  6799=>"111011101",
  6800=>"111000001",
  6801=>"001001011",
  6802=>"011010011",
  6803=>"110001101",
  6804=>"100111111",
  6805=>"001101000",
  6806=>"011000001",
  6807=>"001100010",
  6808=>"110110010",
  6809=>"100010011",
  6810=>"101000100",
  6811=>"001000010",
  6812=>"101001100",
  6813=>"000100101",
  6814=>"100111111",
  6815=>"011101101",
  6816=>"000111101",
  6817=>"000000101",
  6818=>"011000111",
  6819=>"101110101",
  6820=>"000001011",
  6821=>"101111101",
  6822=>"101111100",
  6823=>"111101001",
  6824=>"110111001",
  6825=>"010110010",
  6826=>"000000110",
  6827=>"111011000",
  6828=>"111101101",
  6829=>"000010111",
  6830=>"110010000",
  6831=>"100000001",
  6832=>"101000111",
  6833=>"001101100",
  6834=>"100101011",
  6835=>"111000011",
  6836=>"110001001",
  6837=>"111100000",
  6838=>"001100101",
  6839=>"101010111",
  6840=>"001110111",
  6841=>"101000000",
  6842=>"000011100",
  6843=>"010111100",
  6844=>"100000001",
  6845=>"011101001",
  6846=>"100001101",
  6847=>"110010000",
  6848=>"101110011",
  6849=>"011010001",
  6850=>"001111010",
  6851=>"000111101",
  6852=>"011100100",
  6853=>"100011111",
  6854=>"110000110",
  6855=>"101100000",
  6856=>"111100010",
  6857=>"101001101",
  6858=>"101010101",
  6859=>"011100000",
  6860=>"100100001",
  6861=>"110110101",
  6862=>"010011100",
  6863=>"010001001",
  6864=>"111001011",
  6865=>"101111111",
  6866=>"110001011",
  6867=>"101011000",
  6868=>"000000101",
  6869=>"111001001",
  6870=>"010100010",
  6871=>"000001001",
  6872=>"100101000",
  6873=>"111100101",
  6874=>"101111111",
  6875=>"100001110",
  6876=>"111101111",
  6877=>"011110001",
  6878=>"101101000",
  6879=>"100100000",
  6880=>"000001111",
  6881=>"001110010",
  6882=>"011001010",
  6883=>"100000001",
  6884=>"000101000",
  6885=>"000101011",
  6886=>"001011100",
  6887=>"111111010",
  6888=>"010101000",
  6889=>"101110010",
  6890=>"010011101",
  6891=>"110000011",
  6892=>"101001010",
  6893=>"001001101",
  6894=>"100110110",
  6895=>"100000000",
  6896=>"000010001",
  6897=>"010110100",
  6898=>"110010001",
  6899=>"000100110",
  6900=>"110100111",
  6901=>"110011011",
  6902=>"111100110",
  6903=>"001001000",
  6904=>"101101000",
  6905=>"001111100",
  6906=>"100000010",
  6907=>"010010010",
  6908=>"000100100",
  6909=>"001110100",
  6910=>"001001000",
  6911=>"111001111",
  6912=>"100010000",
  6913=>"010100111",
  6914=>"000000001",
  6915=>"000001100",
  6916=>"101011011",
  6917=>"100011011",
  6918=>"000111001",
  6919=>"011110011",
  6920=>"001111001",
  6921=>"011110011",
  6922=>"010110011",
  6923=>"001000101",
  6924=>"100101001",
  6925=>"111111101",
  6926=>"110100101",
  6927=>"101100011",
  6928=>"101101010",
  6929=>"001101001",
  6930=>"000101101",
  6931=>"101100110",
  6932=>"001110001",
  6933=>"000111011",
  6934=>"101110110",
  6935=>"100010010",
  6936=>"011011001",
  6937=>"010110101",
  6938=>"110010010",
  6939=>"111101011",
  6940=>"001111110",
  6941=>"100110100",
  6942=>"000101100",
  6943=>"010011111",
  6944=>"111011111",
  6945=>"100011000",
  6946=>"101010011",
  6947=>"101101000",
  6948=>"010111011",
  6949=>"110110111",
  6950=>"000001101",
  6951=>"101111110",
  6952=>"101000011",
  6953=>"011011110",
  6954=>"000101111",
  6955=>"010111010",
  6956=>"000010011",
  6957=>"001000110",
  6958=>"000110001",
  6959=>"111001010",
  6960=>"001000010",
  6961=>"100001101",
  6962=>"000000011",
  6963=>"011111101",
  6964=>"111101000",
  6965=>"100101000",
  6966=>"001011100",
  6967=>"010000011",
  6968=>"000010011",
  6969=>"111001000",
  6970=>"011001000",
  6971=>"011111011",
  6972=>"010010011",
  6973=>"100010100",
  6974=>"110111100",
  6975=>"100010010",
  6976=>"111011000",
  6977=>"101110101",
  6978=>"100010100",
  6979=>"100100100",
  6980=>"000110000",
  6981=>"000101110",
  6982=>"001110100",
  6983=>"101100011",
  6984=>"000101101",
  6985=>"100100000",
  6986=>"111011000",
  6987=>"000010001",
  6988=>"001111010",
  6989=>"100001101",
  6990=>"101110111",
  6991=>"000000000",
  6992=>"110100000",
  6993=>"011000001",
  6994=>"011011000",
  6995=>"000100101",
  6996=>"000101110",
  6997=>"110010000",
  6998=>"001011100",
  6999=>"100000110",
  7000=>"100101011",
  7001=>"011010101",
  7002=>"110110100",
  7003=>"011111110",
  7004=>"011001001",
  7005=>"001011000",
  7006=>"100000111",
  7007=>"111101101",
  7008=>"010000001",
  7009=>"110001001",
  7010=>"000110010",
  7011=>"101011001",
  7012=>"101000101",
  7013=>"100101010",
  7014=>"100001010",
  7015=>"100011001",
  7016=>"111110001",
  7017=>"011101100",
  7018=>"011101101",
  7019=>"010000001",
  7020=>"110010011",
  7021=>"000010000",
  7022=>"100111110",
  7023=>"100111011",
  7024=>"010111101",
  7025=>"000000010",
  7026=>"010010000",
  7027=>"000110011",
  7028=>"010001001",
  7029=>"101000011",
  7030=>"110111110",
  7031=>"101101011",
  7032=>"101010011",
  7033=>"000011101",
  7034=>"101001100",
  7035=>"001011111",
  7036=>"001001100",
  7037=>"101011111",
  7038=>"111100100",
  7039=>"101000111",
  7040=>"110000110",
  7041=>"000000010",
  7042=>"000101001",
  7043=>"000110011",
  7044=>"000110101",
  7045=>"011110100",
  7046=>"111011111",
  7047=>"001010001",
  7048=>"000101110",
  7049=>"111100000",
  7050=>"000100001",
  7051=>"110010111",
  7052=>"100010010",
  7053=>"101100000",
  7054=>"000010011",
  7055=>"100001110",
  7056=>"101111101",
  7057=>"110001010",
  7058=>"000011101",
  7059=>"111011111",
  7060=>"100101111",
  7061=>"010110000",
  7062=>"101111100",
  7063=>"011111100",
  7064=>"100010010",
  7065=>"111101010",
  7066=>"101110100",
  7067=>"010011111",
  7068=>"000011100",
  7069=>"001110001",
  7070=>"001011100",
  7071=>"010000001",
  7072=>"010010010",
  7073=>"001110001",
  7074=>"001011111",
  7075=>"011010000",
  7076=>"100100001",
  7077=>"000000111",
  7078=>"010010110",
  7079=>"110110111",
  7080=>"011110100",
  7081=>"110100101",
  7082=>"101101101",
  7083=>"011110100",
  7084=>"100000110",
  7085=>"111000101",
  7086=>"101111100",
  7087=>"101010110",
  7088=>"100111000",
  7089=>"101011100",
  7090=>"111111100",
  7091=>"110001000",
  7092=>"001011110",
  7093=>"001111000",
  7094=>"011000100",
  7095=>"110011101",
  7096=>"011101111",
  7097=>"001100011",
  7098=>"010100001",
  7099=>"101111011",
  7100=>"001001101",
  7101=>"000010100",
  7102=>"111111100",
  7103=>"001011110",
  7104=>"010000111",
  7105=>"100111010",
  7106=>"001010111",
  7107=>"101110101",
  7108=>"010000100",
  7109=>"110111101",
  7110=>"101110011",
  7111=>"111111101",
  7112=>"010001001",
  7113=>"101111111",
  7114=>"100111111",
  7115=>"101110101",
  7116=>"010010010",
  7117=>"101101111",
  7118=>"110011100",
  7119=>"010001101",
  7120=>"100100110",
  7121=>"010001001",
  7122=>"000011000",
  7123=>"011000000",
  7124=>"111000100",
  7125=>"011010011",
  7126=>"001001111",
  7127=>"101001111",
  7128=>"101111110",
  7129=>"111110101",
  7130=>"000111000",
  7131=>"011100100",
  7132=>"010111111",
  7133=>"000010110",
  7134=>"100100100",
  7135=>"110011000",
  7136=>"100010111",
  7137=>"110101101",
  7138=>"110111011",
  7139=>"100010001",
  7140=>"111101101",
  7141=>"101101101",
  7142=>"110001100",
  7143=>"100100011",
  7144=>"100000000",
  7145=>"001010111",
  7146=>"101100011",
  7147=>"100000000",
  7148=>"110010101",
  7149=>"001100100",
  7150=>"010101111",
  7151=>"001111000",
  7152=>"111000111",
  7153=>"011111111",
  7154=>"111101111",
  7155=>"101011111",
  7156=>"001110000",
  7157=>"000111001",
  7158=>"111101010",
  7159=>"101100001",
  7160=>"110010010",
  7161=>"010111010",
  7162=>"011011111",
  7163=>"100100100",
  7164=>"111011001",
  7165=>"010110101",
  7166=>"110110010",
  7167=>"001101000",
  7168=>"001100001",
  7169=>"110110001",
  7170=>"000110100",
  7171=>"000001101",
  7172=>"101111110",
  7173=>"011101001",
  7174=>"011011101",
  7175=>"100100101",
  7176=>"110000000",
  7177=>"001110000",
  7178=>"111101110",
  7179=>"010110110",
  7180=>"101011101",
  7181=>"001000100",
  7182=>"001000101",
  7183=>"011001000",
  7184=>"001101010",
  7185=>"110000101",
  7186=>"111110001",
  7187=>"000010101",
  7188=>"111100111",
  7189=>"001001110",
  7190=>"001100011",
  7191=>"000001100",
  7192=>"000101111",
  7193=>"101000100",
  7194=>"011101101",
  7195=>"101101010",
  7196=>"101001011",
  7197=>"011111111",
  7198=>"010101101",
  7199=>"100111100",
  7200=>"101010001",
  7201=>"110011001",
  7202=>"101011110",
  7203=>"101100001",
  7204=>"011001010",
  7205=>"110110000",
  7206=>"000111010",
  7207=>"111010000",
  7208=>"100000010",
  7209=>"100110000",
  7210=>"110100010",
  7211=>"100111001",
  7212=>"011001010",
  7213=>"111111010",
  7214=>"001110111",
  7215=>"000111001",
  7216=>"101101101",
  7217=>"000011001",
  7218=>"010011000",
  7219=>"110100000",
  7220=>"011101101",
  7221=>"101000010",
  7222=>"000110011",
  7223=>"010111010",
  7224=>"010101011",
  7225=>"100101010",
  7226=>"010001001",
  7227=>"101010000",
  7228=>"011101101",
  7229=>"101011011",
  7230=>"011010111",
  7231=>"100010000",
  7232=>"111110010",
  7233=>"111001001",
  7234=>"111010001",
  7235=>"110111100",
  7236=>"110110110",
  7237=>"101010110",
  7238=>"100110111",
  7239=>"100011010",
  7240=>"000110101",
  7241=>"101111111",
  7242=>"100110010",
  7243=>"000010101",
  7244=>"101101011",
  7245=>"110011110",
  7246=>"110010001",
  7247=>"100110101",
  7248=>"010010011",
  7249=>"000100000",
  7250=>"101111110",
  7251=>"101010110",
  7252=>"110111111",
  7253=>"011000111",
  7254=>"000111100",
  7255=>"011011010",
  7256=>"101010001",
  7257=>"100100000",
  7258=>"010001001",
  7259=>"110001110",
  7260=>"000110111",
  7261=>"111101101",
  7262=>"110110011",
  7263=>"110111000",
  7264=>"001001101",
  7265=>"100101011",
  7266=>"010111011",
  7267=>"011000001",
  7268=>"111010000",
  7269=>"011111000",
  7270=>"001111001",
  7271=>"101111110",
  7272=>"001011100",
  7273=>"110110101",
  7274=>"000001100",
  7275=>"000101000",
  7276=>"001000111",
  7277=>"110001001",
  7278=>"101100110",
  7279=>"111001111",
  7280=>"101011100",
  7281=>"101011011",
  7282=>"001000001",
  7283=>"001111111",
  7284=>"111000000",
  7285=>"010010000",
  7286=>"100100001",
  7287=>"100101001",
  7288=>"110101000",
  7289=>"111101010",
  7290=>"100101011",
  7291=>"100010000",
  7292=>"011110101",
  7293=>"010001100",
  7294=>"101101111",
  7295=>"000000001",
  7296=>"001110100",
  7297=>"010011011",
  7298=>"010111001",
  7299=>"010111110",
  7300=>"011000101",
  7301=>"011111011",
  7302=>"111000001",
  7303=>"001110011",
  7304=>"100011001",
  7305=>"111001011",
  7306=>"110000111",
  7307=>"000101101",
  7308=>"100100000",
  7309=>"111101111",
  7310=>"010100010",
  7311=>"110100000",
  7312=>"000100111",
  7313=>"010010110",
  7314=>"110011110",
  7315=>"101001000",
  7316=>"111000001",
  7317=>"101100010",
  7318=>"101001100",
  7319=>"110110111",
  7320=>"101111010",
  7321=>"111110010",
  7322=>"111111001",
  7323=>"010010000",
  7324=>"011111000",
  7325=>"010101110",
  7326=>"010101111",
  7327=>"010001011",
  7328=>"111011011",
  7329=>"001011001",
  7330=>"001110100",
  7331=>"100001011",
  7332=>"110110101",
  7333=>"000011111",
  7334=>"001000000",
  7335=>"011101101",
  7336=>"011010100",
  7337=>"001011110",
  7338=>"110010010",
  7339=>"100011001",
  7340=>"011001100",
  7341=>"101110000",
  7342=>"001100000",
  7343=>"110111000",
  7344=>"000010010",
  7345=>"101010000",
  7346=>"101111111",
  7347=>"111110000",
  7348=>"001101010",
  7349=>"111101111",
  7350=>"000101111",
  7351=>"010001010",
  7352=>"001111001",
  7353=>"010000000",
  7354=>"010101010",
  7355=>"001000011",
  7356=>"110010010",
  7357=>"111011110",
  7358=>"110100110",
  7359=>"110100101",
  7360=>"010000011",
  7361=>"001011001",
  7362=>"110111011",
  7363=>"010011000",
  7364=>"001010100",
  7365=>"000000001",
  7366=>"001101000",
  7367=>"111100111",
  7368=>"111101011",
  7369=>"111111111",
  7370=>"110111110",
  7371=>"001010000",
  7372=>"111011100",
  7373=>"100000001",
  7374=>"000100011",
  7375=>"111000000",
  7376=>"101011001",
  7377=>"000011001",
  7378=>"001000100",
  7379=>"111101101",
  7380=>"000011010",
  7381=>"100110010",
  7382=>"011100010",
  7383=>"000011011",
  7384=>"100000101",
  7385=>"101011100",
  7386=>"011000000",
  7387=>"110010101",
  7388=>"010000110",
  7389=>"101110101",
  7390=>"100101011",
  7391=>"101110111",
  7392=>"010001000",
  7393=>"001111110",
  7394=>"111110011",
  7395=>"100110000",
  7396=>"100011111",
  7397=>"110100000",
  7398=>"111010100",
  7399=>"001100010",
  7400=>"101000110",
  7401=>"100010101",
  7402=>"000111001",
  7403=>"001001001",
  7404=>"111110011",
  7405=>"010110011",
  7406=>"111101111",
  7407=>"000000000",
  7408=>"110101101",
  7409=>"000111100",
  7410=>"001111000",
  7411=>"101010010",
  7412=>"000010010",
  7413=>"010010000",
  7414=>"101100010",
  7415=>"101000101",
  7416=>"010111100",
  7417=>"000101110",
  7418=>"101001100",
  7419=>"000111001",
  7420=>"001100010",
  7421=>"000001101",
  7422=>"100111101",
  7423=>"100010001",
  7424=>"110111110",
  7425=>"011001000",
  7426=>"000000110",
  7427=>"111110000",
  7428=>"000011100",
  7429=>"000011111",
  7430=>"100100001",
  7431=>"100011010",
  7432=>"011101011",
  7433=>"100101010",
  7434=>"000001100",
  7435=>"001000110",
  7436=>"110011110",
  7437=>"111110010",
  7438=>"000001111",
  7439=>"001100010",
  7440=>"011101001",
  7441=>"101100000",
  7442=>"100000101",
  7443=>"111111001",
  7444=>"111110111",
  7445=>"100000001",
  7446=>"100011100",
  7447=>"111011010",
  7448=>"111000001",
  7449=>"101100010",
  7450=>"110001111",
  7451=>"001110110",
  7452=>"101000010",
  7453=>"111010011",
  7454=>"011101100",
  7455=>"100001111",
  7456=>"111000100",
  7457=>"010111110",
  7458=>"000100001",
  7459=>"100010001",
  7460=>"111100100",
  7461=>"110111001",
  7462=>"000000110",
  7463=>"010100100",
  7464=>"000011111",
  7465=>"010000001",
  7466=>"000000100",
  7467=>"111011001",
  7468=>"010100011",
  7469=>"100000111",
  7470=>"100000010",
  7471=>"001111111",
  7472=>"010101110",
  7473=>"011111001",
  7474=>"100100001",
  7475=>"100100111",
  7476=>"110111100",
  7477=>"000101100",
  7478=>"010000100",
  7479=>"110001001",
  7480=>"101000001",
  7481=>"100101110",
  7482=>"010101010",
  7483=>"111111110",
  7484=>"000011000",
  7485=>"001011000",
  7486=>"001101110",
  7487=>"000110000",
  7488=>"101000001",
  7489=>"010101010",
  7490=>"000111010",
  7491=>"001011010",
  7492=>"011011101",
  7493=>"010001011",
  7494=>"110000100",
  7495=>"110100101",
  7496=>"110000000",
  7497=>"010111000",
  7498=>"101011111",
  7499=>"000010000",
  7500=>"111111111",
  7501=>"101101001",
  7502=>"000101101",
  7503=>"111010100",
  7504=>"000111111",
  7505=>"100000111",
  7506=>"110000111",
  7507=>"011011111",
  7508=>"100001001",
  7509=>"111101110",
  7510=>"101000000",
  7511=>"100101001",
  7512=>"101110101",
  7513=>"010111000",
  7514=>"001000001",
  7515=>"001000101",
  7516=>"010110011",
  7517=>"110101110",
  7518=>"110001001",
  7519=>"011001100",
  7520=>"000010110",
  7521=>"001011111",
  7522=>"011011101",
  7523=>"111010001",
  7524=>"011101011",
  7525=>"000011010",
  7526=>"111100110",
  7527=>"110100010",
  7528=>"000100110",
  7529=>"011010101",
  7530=>"101010011",
  7531=>"110111111",
  7532=>"000000000",
  7533=>"111101000",
  7534=>"110000111",
  7535=>"111100011",
  7536=>"110110001",
  7537=>"111100110",
  7538=>"000110110",
  7539=>"111101101",
  7540=>"100011000",
  7541=>"101101001",
  7542=>"010110111",
  7543=>"100000010",
  7544=>"010001001",
  7545=>"011011111",
  7546=>"100110110",
  7547=>"001000111",
  7548=>"010111101",
  7549=>"010000001",
  7550=>"001001010",
  7551=>"100100110",
  7552=>"000000000",
  7553=>"101101010",
  7554=>"011010100",
  7555=>"010100010",
  7556=>"011101110",
  7557=>"101111110",
  7558=>"011101100",
  7559=>"000000101",
  7560=>"001110111",
  7561=>"001111001",
  7562=>"101000001",
  7563=>"110110001",
  7564=>"101011101",
  7565=>"010011011",
  7566=>"010111111",
  7567=>"001010011",
  7568=>"010110011",
  7569=>"110100101",
  7570=>"101101100",
  7571=>"110110111",
  7572=>"111111101",
  7573=>"111001101",
  7574=>"000111001",
  7575=>"100011111",
  7576=>"100010111",
  7577=>"111101110",
  7578=>"111011011",
  7579=>"001000101",
  7580=>"001011111",
  7581=>"000110111",
  7582=>"000001000",
  7583=>"110010000",
  7584=>"111001100",
  7585=>"110100000",
  7586=>"000011001",
  7587=>"101110101",
  7588=>"011110000",
  7589=>"011010000",
  7590=>"111001001",
  7591=>"111111010",
  7592=>"010101111",
  7593=>"001000110",
  7594=>"010111101",
  7595=>"011100111",
  7596=>"100000111",
  7597=>"011000010",
  7598=>"010011001",
  7599=>"001110001",
  7600=>"101100010",
  7601=>"000000101",
  7602=>"101101001",
  7603=>"000000011",
  7604=>"110011110",
  7605=>"111111000",
  7606=>"010000011",
  7607=>"100000001",
  7608=>"101011010",
  7609=>"110001000",
  7610=>"110011111",
  7611=>"001111101",
  7612=>"000010100",
  7613=>"101011010",
  7614=>"101000101",
  7615=>"101011101",
  7616=>"110010010",
  7617=>"111010101",
  7618=>"010110101",
  7619=>"111101101",
  7620=>"100000111",
  7621=>"000001001",
  7622=>"111111111",
  7623=>"100101000",
  7624=>"000101000",
  7625=>"010010000",
  7626=>"101001101",
  7627=>"111111010",
  7628=>"101101000",
  7629=>"101101110",
  7630=>"000010100",
  7631=>"100000100",
  7632=>"101110000",
  7633=>"101010110",
  7634=>"011010010",
  7635=>"111011001",
  7636=>"110111111",
  7637=>"000000101",
  7638=>"011000001",
  7639=>"010101101",
  7640=>"100101001",
  7641=>"101101001",
  7642=>"111110101",
  7643=>"011001001",
  7644=>"110101011",
  7645=>"101011010",
  7646=>"000010111",
  7647=>"000011100",
  7648=>"001001011",
  7649=>"110001101",
  7650=>"110000011",
  7651=>"010001001",
  7652=>"101000100",
  7653=>"010110000",
  7654=>"010011001",
  7655=>"000001111",
  7656=>"110001001",
  7657=>"101000100",
  7658=>"000011100",
  7659=>"011010010",
  7660=>"000110011",
  7661=>"101101011",
  7662=>"011010111",
  7663=>"000001100",
  7664=>"000101110",
  7665=>"100101001",
  7666=>"110000101",
  7667=>"001110011",
  7668=>"111111111",
  7669=>"010100010",
  7670=>"010001000",
  7671=>"101010110",
  7672=>"101111111",
  7673=>"111110111",
  7674=>"000011000",
  7675=>"110101010",
  7676=>"100101001",
  7677=>"111111001",
  7678=>"111011000",
  7679=>"110111111",
  7680=>"010011001",
  7681=>"011101100",
  7682=>"010110111",
  7683=>"010000011",
  7684=>"010011011",
  7685=>"100011000",
  7686=>"010000000",
  7687=>"011010000",
  7688=>"001100101",
  7689=>"110101101",
  7690=>"100011110",
  7691=>"000101000",
  7692=>"100110111",
  7693=>"111100010",
  7694=>"100001110",
  7695=>"110101001",
  7696=>"100101110",
  7697=>"000101110",
  7698=>"111101001",
  7699=>"100010010",
  7700=>"010101111",
  7701=>"110101100",
  7702=>"000010000",
  7703=>"110010110",
  7704=>"001101001",
  7705=>"100110110",
  7706=>"100011111",
  7707=>"000001000",
  7708=>"101111110",
  7709=>"011011011",
  7710=>"000100011",
  7711=>"010110000",
  7712=>"101101011",
  7713=>"000101101",
  7714=>"000010011",
  7715=>"011011000",
  7716=>"101100110",
  7717=>"011010111",
  7718=>"011000111",
  7719=>"100011001",
  7720=>"001110000",
  7721=>"011001100",
  7722=>"011011111",
  7723=>"010101100",
  7724=>"110110101",
  7725=>"100000001",
  7726=>"010110000",
  7727=>"101101111",
  7728=>"111011110",
  7729=>"110110010",
  7730=>"010010010",
  7731=>"110010111",
  7732=>"101100000",
  7733=>"000010111",
  7734=>"010110111",
  7735=>"011101101",
  7736=>"000011010",
  7737=>"010010001",
  7738=>"010011110",
  7739=>"100001011",
  7740=>"001010110",
  7741=>"010000101",
  7742=>"100101000",
  7743=>"000000111",
  7744=>"101000101",
  7745=>"100011011",
  7746=>"000000101",
  7747=>"110111001",
  7748=>"110000000",
  7749=>"010100010",
  7750=>"101001011",
  7751=>"001111001",
  7752=>"111011011",
  7753=>"100110111",
  7754=>"000100010",
  7755=>"100110010",
  7756=>"101111111",
  7757=>"000000000",
  7758=>"110011111",
  7759=>"000011000",
  7760=>"011111100",
  7761=>"011100110",
  7762=>"011111011",
  7763=>"101101010",
  7764=>"101010100",
  7765=>"000111000",
  7766=>"000000010",
  7767=>"100001110",
  7768=>"101011011",
  7769=>"101000010",
  7770=>"111001101",
  7771=>"101111000",
  7772=>"101000001",
  7773=>"011110001",
  7774=>"110110000",
  7775=>"111111110",
  7776=>"011100010",
  7777=>"110010000",
  7778=>"111010111",
  7779=>"010010000",
  7780=>"100110011",
  7781=>"011001000",
  7782=>"000111000",
  7783=>"000110110",
  7784=>"010100111",
  7785=>"000001100",
  7786=>"000111111",
  7787=>"001011111",
  7788=>"001001011",
  7789=>"000110010",
  7790=>"011010101",
  7791=>"010110111",
  7792=>"000011000",
  7793=>"101100100",
  7794=>"000100000",
  7795=>"000101010",
  7796=>"100101100",
  7797=>"011010111",
  7798=>"010100111",
  7799=>"111101101",
  7800=>"100101111",
  7801=>"000110000",
  7802=>"001111111",
  7803=>"001011010",
  7804=>"001110010",
  7805=>"001001000",
  7806=>"011100101",
  7807=>"101101001",
  7808=>"100111001",
  7809=>"100011101",
  7810=>"110100111",
  7811=>"000101010",
  7812=>"010011110",
  7813=>"010010011",
  7814=>"101100101",
  7815=>"000011011",
  7816=>"111010101",
  7817=>"000001010",
  7818=>"110011010",
  7819=>"000101000",
  7820=>"000000110",
  7821=>"010001100",
  7822=>"010000000",
  7823=>"101111100",
  7824=>"010101000",
  7825=>"001101101",
  7826=>"100011110",
  7827=>"100010010",
  7828=>"011011001",
  7829=>"100101100",
  7830=>"010001100",
  7831=>"101001111",
  7832=>"010010001",
  7833=>"110001001",
  7834=>"000000001",
  7835=>"111100101",
  7836=>"000100100",
  7837=>"001000011",
  7838=>"100110001",
  7839=>"100110001",
  7840=>"001111011",
  7841=>"100001111",
  7842=>"001000011",
  7843=>"110101011",
  7844=>"100011011",
  7845=>"000111111",
  7846=>"001011101",
  7847=>"001001000",
  7848=>"111100010",
  7849=>"010100100",
  7850=>"111011101",
  7851=>"000101100",
  7852=>"111011011",
  7853=>"110111100",
  7854=>"101111101",
  7855=>"110110110",
  7856=>"011000000",
  7857=>"000011101",
  7858=>"100110111",
  7859=>"101101101",
  7860=>"010001101",
  7861=>"100100000",
  7862=>"010011101",
  7863=>"000100000",
  7864=>"111111110",
  7865=>"000100111",
  7866=>"000100100",
  7867=>"101101111",
  7868=>"001111100",
  7869=>"011101111",
  7870=>"010011001",
  7871=>"011100111",
  7872=>"010111000",
  7873=>"100101011",
  7874=>"101101101",
  7875=>"010101110",
  7876=>"110111011",
  7877=>"000100011",
  7878=>"010011110",
  7879=>"010100101",
  7880=>"000000000",
  7881=>"011011101",
  7882=>"000111100",
  7883=>"001010010",
  7884=>"100111111",
  7885=>"001100011",
  7886=>"011111111",
  7887=>"110100001",
  7888=>"010000011",
  7889=>"001001111",
  7890=>"100000001",
  7891=>"011111011",
  7892=>"100111111",
  7893=>"110111011",
  7894=>"000111111",
  7895=>"000110000",
  7896=>"000101110",
  7897=>"101110110",
  7898=>"100000110",
  7899=>"000001001",
  7900=>"111010001",
  7901=>"010100101",
  7902=>"001001100",
  7903=>"101000010",
  7904=>"011100000",
  7905=>"000000110",
  7906=>"000000001",
  7907=>"010110011",
  7908=>"010100101",
  7909=>"100011001",
  7910=>"101110000",
  7911=>"101111101",
  7912=>"010100000",
  7913=>"010001100",
  7914=>"100011111",
  7915=>"101001100",
  7916=>"001010001",
  7917=>"110011011",
  7918=>"110100011",
  7919=>"001000000",
  7920=>"101101111",
  7921=>"101000000",
  7922=>"101011000",
  7923=>"110001110",
  7924=>"011100010",
  7925=>"111111111",
  7926=>"011100111",
  7927=>"101101101",
  7928=>"011010101",
  7929=>"001111101",
  7930=>"001111111",
  7931=>"011010101",
  7932=>"010110010",
  7933=>"100111011",
  7934=>"001110010",
  7935=>"101000100",
  7936=>"011100010",
  7937=>"101100001",
  7938=>"111100011",
  7939=>"000011000",
  7940=>"111010101",
  7941=>"000110000",
  7942=>"111000010",
  7943=>"001000001",
  7944=>"101001100",
  7945=>"011001011",
  7946=>"001110011",
  7947=>"000010111",
  7948=>"110011000",
  7949=>"010010000",
  7950=>"010101100",
  7951=>"000110000",
  7952=>"100011001",
  7953=>"100000000",
  7954=>"110011011",
  7955=>"111110111",
  7956=>"100100001",
  7957=>"011010110",
  7958=>"001110101",
  7959=>"101110111",
  7960=>"001101110",
  7961=>"010010010",
  7962=>"110011000",
  7963=>"110011010",
  7964=>"110001101",
  7965=>"111100011",
  7966=>"111001000",
  7967=>"111010100",
  7968=>"111110010",
  7969=>"111000010",
  7970=>"111010110",
  7971=>"100001100",
  7972=>"101011100",
  7973=>"001010001",
  7974=>"000100110",
  7975=>"100000000",
  7976=>"100011001",
  7977=>"001000111",
  7978=>"011011011",
  7979=>"000011100",
  7980=>"000111001",
  7981=>"101101000",
  7982=>"000000000",
  7983=>"111011110",
  7984=>"000111011",
  7985=>"101001011",
  7986=>"010010100",
  7987=>"011111011",
  7988=>"000101101",
  7989=>"100100111",
  7990=>"001001100",
  7991=>"000010001",
  7992=>"101111100",
  7993=>"100100001",
  7994=>"001110111",
  7995=>"000110010",
  7996=>"001000111",
  7997=>"000010101",
  7998=>"010101111",
  7999=>"000001000",
  8000=>"011101100",
  8001=>"001001111",
  8002=>"110001011",
  8003=>"001011011",
  8004=>"110010100",
  8005=>"110010110",
  8006=>"001000010",
  8007=>"101111010",
  8008=>"011111110",
  8009=>"001010001",
  8010=>"101101101",
  8011=>"000100001",
  8012=>"110111101",
  8013=>"101001111",
  8014=>"001110001",
  8015=>"011000000",
  8016=>"001110010",
  8017=>"010101110",
  8018=>"100011100",
  8019=>"010101111",
  8020=>"110011011",
  8021=>"111110001",
  8022=>"000111111",
  8023=>"100000000",
  8024=>"011001111",
  8025=>"011011100",
  8026=>"001110110",
  8027=>"001001000",
  8028=>"100001100",
  8029=>"100100100",
  8030=>"100000101",
  8031=>"000111110",
  8032=>"011000000",
  8033=>"100000001",
  8034=>"011101111",
  8035=>"011111110",
  8036=>"100011111",
  8037=>"000110100",
  8038=>"001010011",
  8039=>"100101001",
  8040=>"111011100",
  8041=>"101001111",
  8042=>"110001111",
  8043=>"010111001",
  8044=>"010011010",
  8045=>"011101011",
  8046=>"101111100",
  8047=>"110010101",
  8048=>"111110110",
  8049=>"011010001",
  8050=>"110110010",
  8051=>"011000101",
  8052=>"000010000",
  8053=>"100110001",
  8054=>"001111000",
  8055=>"011001111",
  8056=>"001101110",
  8057=>"001011001",
  8058=>"100010100",
  8059=>"100010001",
  8060=>"111001000",
  8061=>"110011100",
  8062=>"100111101",
  8063=>"111101010",
  8064=>"111101001",
  8065=>"011111001",
  8066=>"101000011",
  8067=>"010111111",
  8068=>"000000100",
  8069=>"100011010",
  8070=>"101000100",
  8071=>"101110011",
  8072=>"011000110",
  8073=>"111101000",
  8074=>"001001001",
  8075=>"111010001",
  8076=>"011010101",
  8077=>"010110101",
  8078=>"100000110",
  8079=>"010110001",
  8080=>"000111111",
  8081=>"001010101",
  8082=>"110000001",
  8083=>"100110100",
  8084=>"101000011",
  8085=>"100000100",
  8086=>"000101101",
  8087=>"001110001",
  8088=>"101001100",
  8089=>"100111000",
  8090=>"100010000",
  8091=>"110101010",
  8092=>"000011010",
  8093=>"111011000",
  8094=>"111101011",
  8095=>"001000110",
  8096=>"011111011",
  8097=>"000111111",
  8098=>"001001010",
  8099=>"011001010",
  8100=>"000000000",
  8101=>"100111100",
  8102=>"100111011",
  8103=>"001111010",
  8104=>"111111111",
  8105=>"011001110",
  8106=>"000001100",
  8107=>"100010100",
  8108=>"110000111",
  8109=>"101110010",
  8110=>"111011111",
  8111=>"100101010",
  8112=>"111000001",
  8113=>"011100110",
  8114=>"110001000",
  8115=>"001000011",
  8116=>"011100101",
  8117=>"100011000",
  8118=>"100011010",
  8119=>"011001010",
  8120=>"100011101",
  8121=>"101101100",
  8122=>"000100110",
  8123=>"110100000",
  8124=>"110000110",
  8125=>"101001101",
  8126=>"011111111",
  8127=>"011110100",
  8128=>"010110110",
  8129=>"011100010",
  8130=>"011101111",
  8131=>"011111110",
  8132=>"010111001",
  8133=>"111111011",
  8134=>"010011111",
  8135=>"100111101",
  8136=>"000010000",
  8137=>"001100010",
  8138=>"011010001",
  8139=>"000111011",
  8140=>"001010001",
  8141=>"110001100",
  8142=>"110010100",
  8143=>"101100011",
  8144=>"100000001",
  8145=>"011110110",
  8146=>"010010001",
  8147=>"011000110",
  8148=>"000110001",
  8149=>"111011010",
  8150=>"101110101",
  8151=>"101100101",
  8152=>"110000011",
  8153=>"011011100",
  8154=>"001011100",
  8155=>"110101111",
  8156=>"110100010",
  8157=>"011101100",
  8158=>"001110111",
  8159=>"100010001",
  8160=>"011000101",
  8161=>"001101001",
  8162=>"100011100",
  8163=>"011001100",
  8164=>"000110100",
  8165=>"110000110",
  8166=>"001010010",
  8167=>"111100000",
  8168=>"010100001",
  8169=>"010000011",
  8170=>"011100010",
  8171=>"101110010",
  8172=>"100110010",
  8173=>"000011100",
  8174=>"001111011",
  8175=>"101001011",
  8176=>"101010010",
  8177=>"111111010",
  8178=>"000011101",
  8179=>"000011100",
  8180=>"110101011",
  8181=>"000110010",
  8182=>"100011111",
  8183=>"001001001",
  8184=>"010111110",
  8185=>"011001101",
  8186=>"000111001",
  8187=>"110111101",
  8188=>"000000110",
  8189=>"100000011",
  8190=>"000111100",
  8191=>"111001110",
  8192=>"100100001",
  8193=>"000001001",
  8194=>"101010101",
  8195=>"111100101",
  8196=>"011101000",
  8197=>"110010110",
  8198=>"010101100",
  8199=>"101110000",
  8200=>"001010001",
  8201=>"101100000",
  8202=>"001001000",
  8203=>"000100010",
  8204=>"100000000",
  8205=>"100000110",
  8206=>"101011100",
  8207=>"111000110",
  8208=>"000001110",
  8209=>"111110111",
  8210=>"100111111",
  8211=>"011001110",
  8212=>"001110000",
  8213=>"110010011",
  8214=>"111110100",
  8215=>"011000001",
  8216=>"010000010",
  8217=>"100101111",
  8218=>"101001010",
  8219=>"001001110",
  8220=>"001100100",
  8221=>"100000001",
  8222=>"001011100",
  8223=>"110101111",
  8224=>"101100011",
  8225=>"001000110",
  8226=>"000110111",
  8227=>"000011011",
  8228=>"010001011",
  8229=>"100111111",
  8230=>"010110111",
  8231=>"011001100",
  8232=>"001011111",
  8233=>"101011011",
  8234=>"000011110",
  8235=>"111101001",
  8236=>"001010111",
  8237=>"110000000",
  8238=>"100111011",
  8239=>"010001100",
  8240=>"111111011",
  8241=>"100110000",
  8242=>"111111011",
  8243=>"110110101",
  8244=>"101011001",
  8245=>"010100100",
  8246=>"000001010",
  8247=>"110010100",
  8248=>"001010111",
  8249=>"110100101",
  8250=>"011000101",
  8251=>"010000011",
  8252=>"100011000",
  8253=>"100100110",
  8254=>"111011001",
  8255=>"000010001",
  8256=>"000000011",
  8257=>"010100011",
  8258=>"100001000",
  8259=>"111110011",
  8260=>"000000111",
  8261=>"100101111",
  8262=>"110100001",
  8263=>"001001110",
  8264=>"100001110",
  8265=>"011101001",
  8266=>"111001000",
  8267=>"000110100",
  8268=>"000000000",
  8269=>"110101010",
  8270=>"010101111",
  8271=>"011110001",
  8272=>"010110001",
  8273=>"010000010",
  8274=>"010001101",
  8275=>"100111011",
  8276=>"000001000",
  8277=>"100011110",
  8278=>"010111101",
  8279=>"100110110",
  8280=>"100111100",
  8281=>"110111010",
  8282=>"110011000",
  8283=>"000100110",
  8284=>"010010001",
  8285=>"000001111",
  8286=>"111110101",
  8287=>"111010101",
  8288=>"111010100",
  8289=>"101000100",
  8290=>"110110110",
  8291=>"000011000",
  8292=>"101011100",
  8293=>"010010101",
  8294=>"100101111",
  8295=>"100000000",
  8296=>"000100111",
  8297=>"111111010",
  8298=>"110100101",
  8299=>"111001110",
  8300=>"000000100",
  8301=>"101101100",
  8302=>"011011111",
  8303=>"100111010",
  8304=>"111011100",
  8305=>"100110111",
  8306=>"010111010",
  8307=>"100000101",
  8308=>"100010010",
  8309=>"101001100",
  8310=>"000100010",
  8311=>"001101101",
  8312=>"000010001",
  8313=>"110000111",
  8314=>"111010110",
  8315=>"100111111",
  8316=>"011010000",
  8317=>"110100000",
  8318=>"000100111",
  8319=>"111111000",
  8320=>"111011100",
  8321=>"101111000",
  8322=>"000011100",
  8323=>"111001111",
  8324=>"111100010",
  8325=>"000011110",
  8326=>"101100101",
  8327=>"000111111",
  8328=>"011000101",
  8329=>"011111011",
  8330=>"101000100",
  8331=>"000011011",
  8332=>"000100011",
  8333=>"010101110",
  8334=>"000010001",
  8335=>"101001111",
  8336=>"100100100",
  8337=>"010011100",
  8338=>"011001111",
  8339=>"000101011",
  8340=>"001101011",
  8341=>"111110001",
  8342=>"111000100",
  8343=>"001010011",
  8344=>"111000111",
  8345=>"001011111",
  8346=>"101110111",
  8347=>"011110110",
  8348=>"110010001",
  8349=>"110001000",
  8350=>"000000001",
  8351=>"011000110",
  8352=>"110101010",
  8353=>"101010101",
  8354=>"101001111",
  8355=>"101100111",
  8356=>"100001000",
  8357=>"010001010",
  8358=>"001010111",
  8359=>"110100010",
  8360=>"101011100",
  8361=>"001100101",
  8362=>"100010101",
  8363=>"000000100",
  8364=>"100011110",
  8365=>"101101011",
  8366=>"110001101",
  8367=>"000010110",
  8368=>"010111111",
  8369=>"010101000",
  8370=>"010010000",
  8371=>"100111001",
  8372=>"110101001",
  8373=>"100010000",
  8374=>"100101110",
  8375=>"101011011",
  8376=>"001000101",
  8377=>"111100000",
  8378=>"110110100",
  8379=>"011100101",
  8380=>"110001000",
  8381=>"110101000",
  8382=>"010010110",
  8383=>"001101010",
  8384=>"010001100",
  8385=>"000000111",
  8386=>"110111101",
  8387=>"011011101",
  8388=>"110010101",
  8389=>"110010100",
  8390=>"001000110",
  8391=>"010100011",
  8392=>"010001101",
  8393=>"111101000",
  8394=>"000001000",
  8395=>"001101111",
  8396=>"000000100",
  8397=>"111011011",
  8398=>"100000111",
  8399=>"000011011",
  8400=>"011101000",
  8401=>"010011011",
  8402=>"010000110",
  8403=>"001100101",
  8404=>"110011010",
  8405=>"100011110",
  8406=>"000010101",
  8407=>"000000100",
  8408=>"100100011",
  8409=>"001000101",
  8410=>"110110100",
  8411=>"010001000",
  8412=>"001011101",
  8413=>"110101110",
  8414=>"010010010",
  8415=>"001001111",
  8416=>"000000010",
  8417=>"000111001",
  8418=>"011111010",
  8419=>"011111001",
  8420=>"011110111",
  8421=>"110010000",
  8422=>"100100000",
  8423=>"000011111",
  8424=>"100101110",
  8425=>"010111110",
  8426=>"011011110",
  8427=>"101100111",
  8428=>"111011100",
  8429=>"101000110",
  8430=>"010101100",
  8431=>"100111111",
  8432=>"110000101",
  8433=>"110001000",
  8434=>"000001000",
  8435=>"010101111",
  8436=>"100000000",
  8437=>"011011100",
  8438=>"000110101",
  8439=>"000100101",
  8440=>"000101101",
  8441=>"000011100",
  8442=>"101111101",
  8443=>"000010001",
  8444=>"011011001",
  8445=>"101111011",
  8446=>"110101100",
  8447=>"010010110",
  8448=>"110111011",
  8449=>"011011001",
  8450=>"101111010",
  8451=>"010010101",
  8452=>"010111011",
  8453=>"100111010",
  8454=>"101011010",
  8455=>"010011001",
  8456=>"010011000",
  8457=>"010010111",
  8458=>"111111000",
  8459=>"001100001",
  8460=>"110011100",
  8461=>"011001000",
  8462=>"111010101",
  8463=>"111100110",
  8464=>"000010011",
  8465=>"010011110",
  8466=>"101000001",
  8467=>"010000011",
  8468=>"100100011",
  8469=>"100001110",
  8470=>"010111010",
  8471=>"101010010",
  8472=>"010011110",
  8473=>"001001101",
  8474=>"010110100",
  8475=>"101011010",
  8476=>"111001010",
  8477=>"111001110",
  8478=>"100010101",
  8479=>"101100000",
  8480=>"000101011",
  8481=>"011010110",
  8482=>"110111011",
  8483=>"010100111",
  8484=>"100100011",
  8485=>"000001011",
  8486=>"100100100",
  8487=>"000110010",
  8488=>"101000011",
  8489=>"011101101",
  8490=>"010010110",
  8491=>"101111010",
  8492=>"100001010",
  8493=>"110111001",
  8494=>"110000111",
  8495=>"101001010",
  8496=>"011011000",
  8497=>"011111011",
  8498=>"111110010",
  8499=>"000000101",
  8500=>"000100100",
  8501=>"011001111",
  8502=>"010100100",
  8503=>"000011010",
  8504=>"001010010",
  8505=>"011111101",
  8506=>"100110011",
  8507=>"110001110",
  8508=>"111100111",
  8509=>"110000101",
  8510=>"101100001",
  8511=>"110100000",
  8512=>"110101111",
  8513=>"000111111",
  8514=>"101001110",
  8515=>"100011100",
  8516=>"011010010",
  8517=>"100001010",
  8518=>"101100111",
  8519=>"100001111",
  8520=>"011001100",
  8521=>"101111011",
  8522=>"111101110",
  8523=>"111110000",
  8524=>"000011100",
  8525=>"110000100",
  8526=>"001111100",
  8527=>"101001010",
  8528=>"100111011",
  8529=>"011001110",
  8530=>"010101110",
  8531=>"111110001",
  8532=>"011110010",
  8533=>"101110011",
  8534=>"110000110",
  8535=>"001100001",
  8536=>"000101111",
  8537=>"101000101",
  8538=>"101101010",
  8539=>"000100111",
  8540=>"001111001",
  8541=>"001111010",
  8542=>"011001100",
  8543=>"011111001",
  8544=>"100001011",
  8545=>"110110111",
  8546=>"101110000",
  8547=>"111000110",
  8548=>"010111101",
  8549=>"000110001",
  8550=>"100101101",
  8551=>"100001010",
  8552=>"011101011",
  8553=>"001010111",
  8554=>"100100000",
  8555=>"001011011",
  8556=>"100111110",
  8557=>"101000010",
  8558=>"001000000",
  8559=>"100000101",
  8560=>"000100101",
  8561=>"101001111",
  8562=>"010010101",
  8563=>"111100010",
  8564=>"110101010",
  8565=>"001101000",
  8566=>"111110100",
  8567=>"100011110",
  8568=>"011010011",
  8569=>"111011000",
  8570=>"110010100",
  8571=>"111111011",
  8572=>"101011000",
  8573=>"110101001",
  8574=>"111001011",
  8575=>"101101001",
  8576=>"101000101",
  8577=>"011101000",
  8578=>"100101111",
  8579=>"101001001",
  8580=>"110001011",
  8581=>"100100110",
  8582=>"010110101",
  8583=>"011001101",
  8584=>"001001000",
  8585=>"100101000",
  8586=>"101000011",
  8587=>"100010101",
  8588=>"101111110",
  8589=>"110000100",
  8590=>"001000010",
  8591=>"000000100",
  8592=>"101110011",
  8593=>"010100100",
  8594=>"111101111",
  8595=>"001010011",
  8596=>"111011001",
  8597=>"110111110",
  8598=>"100011111",
  8599=>"000010001",
  8600=>"101101000",
  8601=>"111110111",
  8602=>"011101111",
  8603=>"111011000",
  8604=>"110011110",
  8605=>"101100011",
  8606=>"011111001",
  8607=>"010001111",
  8608=>"000000110",
  8609=>"110011101",
  8610=>"111010011",
  8611=>"100000111",
  8612=>"110000010",
  8613=>"000100101",
  8614=>"111101010",
  8615=>"101000101",
  8616=>"101110000",
  8617=>"110011110",
  8618=>"111110111",
  8619=>"111000001",
  8620=>"111101010",
  8621=>"001010101",
  8622=>"011110010",
  8623=>"001111000",
  8624=>"011011011",
  8625=>"110110111",
  8626=>"000011000",
  8627=>"001000010",
  8628=>"100110110",
  8629=>"101100001",
  8630=>"111111111",
  8631=>"110110000",
  8632=>"010010000",
  8633=>"001001101",
  8634=>"011100111",
  8635=>"011101100",
  8636=>"101010110",
  8637=>"100111000",
  8638=>"001101110",
  8639=>"111110110",
  8640=>"111010000",
  8641=>"010000001",
  8642=>"011000100",
  8643=>"000010011",
  8644=>"100100100",
  8645=>"010110101",
  8646=>"111001001",
  8647=>"101011000",
  8648=>"101101000",
  8649=>"010110110",
  8650=>"000011001",
  8651=>"111001010",
  8652=>"110100011",
  8653=>"111101001",
  8654=>"001101011",
  8655=>"011000111",
  8656=>"101110110",
  8657=>"010001110",
  8658=>"001000110",
  8659=>"100001100",
  8660=>"011011101",
  8661=>"101001010",
  8662=>"001110001",
  8663=>"101100110",
  8664=>"010000011",
  8665=>"010000110",
  8666=>"001111000",
  8667=>"110001001",
  8668=>"110000101",
  8669=>"000000010",
  8670=>"101001001",
  8671=>"010100010",
  8672=>"011101011",
  8673=>"111010100",
  8674=>"100011100",
  8675=>"000101000",
  8676=>"111110010",
  8677=>"000001111",
  8678=>"001011011",
  8679=>"011011000",
  8680=>"011110000",
  8681=>"001100111",
  8682=>"001000010",
  8683=>"110100000",
  8684=>"100011001",
  8685=>"011001110",
  8686=>"000000100",
  8687=>"111100001",
  8688=>"110101100",
  8689=>"011110110",
  8690=>"110001000",
  8691=>"000000000",
  8692=>"010101010",
  8693=>"010001110",
  8694=>"110001110",
  8695=>"110000110",
  8696=>"111000011",
  8697=>"011110011",
  8698=>"000010111",
  8699=>"100101101",
  8700=>"010000111",
  8701=>"001010101",
  8702=>"110011111",
  8703=>"010111000",
  8704=>"011000101",
  8705=>"111111010",
  8706=>"111110110",
  8707=>"100100111",
  8708=>"100100111",
  8709=>"010110100",
  8710=>"001001111",
  8711=>"010111111",
  8712=>"100001001",
  8713=>"011010000",
  8714=>"000111101",
  8715=>"000100111",
  8716=>"111001010",
  8717=>"011011100",
  8718=>"100001111",
  8719=>"101101001",
  8720=>"110000111",
  8721=>"111101010",
  8722=>"100101001",
  8723=>"000001000",
  8724=>"101110101",
  8725=>"100100011",
  8726=>"001000010",
  8727=>"011011101",
  8728=>"001111010",
  8729=>"111010101",
  8730=>"101001010",
  8731=>"011011010",
  8732=>"010000000",
  8733=>"000011000",
  8734=>"010111001",
  8735=>"001000101",
  8736=>"000110000",
  8737=>"110000011",
  8738=>"001001110",
  8739=>"011010000",
  8740=>"000000110",
  8741=>"100111111",
  8742=>"011110001",
  8743=>"100011010",
  8744=>"111110101",
  8745=>"011011111",
  8746=>"010010110",
  8747=>"001111001",
  8748=>"001000100",
  8749=>"001101001",
  8750=>"101101011",
  8751=>"000100111",
  8752=>"010010010",
  8753=>"010100101",
  8754=>"111000001",
  8755=>"100000110",
  8756=>"001100101",
  8757=>"001000111",
  8758=>"000000110",
  8759=>"100100101",
  8760=>"000010001",
  8761=>"101100100",
  8762=>"100010011",
  8763=>"110011100",
  8764=>"100110111",
  8765=>"000110100",
  8766=>"101111001",
  8767=>"111001001",
  8768=>"000101111",
  8769=>"001001001",
  8770=>"101000000",
  8771=>"011101000",
  8772=>"101000101",
  8773=>"100001010",
  8774=>"111110111",
  8775=>"011011010",
  8776=>"111100110",
  8777=>"110100100",
  8778=>"011001010",
  8779=>"000010111",
  8780=>"010100101",
  8781=>"010001110",
  8782=>"001101111",
  8783=>"110011101",
  8784=>"000100101",
  8785=>"110101011",
  8786=>"010110101",
  8787=>"011000010",
  8788=>"010010100",
  8789=>"110000111",
  8790=>"110000010",
  8791=>"011001110",
  8792=>"101001010",
  8793=>"101011011",
  8794=>"000100010",
  8795=>"001110101",
  8796=>"110100101",
  8797=>"011001110",
  8798=>"101100100",
  8799=>"000001011",
  8800=>"000000011",
  8801=>"000110111",
  8802=>"111100001",
  8803=>"100101000",
  8804=>"110001011",
  8805=>"111100000",
  8806=>"101101001",
  8807=>"001110011",
  8808=>"100001110",
  8809=>"000001111",
  8810=>"101100000",
  8811=>"100010100",
  8812=>"101101011",
  8813=>"111111000",
  8814=>"110110100",
  8815=>"001111011",
  8816=>"101110000",
  8817=>"000011100",
  8818=>"001111001",
  8819=>"111101001",
  8820=>"011100110",
  8821=>"101010000",
  8822=>"001000011",
  8823=>"000111111",
  8824=>"011101010",
  8825=>"100001100",
  8826=>"001110101",
  8827=>"000000101",
  8828=>"111111111",
  8829=>"001011000",
  8830=>"101010001",
  8831=>"111101100",
  8832=>"010000110",
  8833=>"000110110",
  8834=>"100101100",
  8835=>"011100001",
  8836=>"011001011",
  8837=>"110100011",
  8838=>"010011001",
  8839=>"100101111",
  8840=>"001110111",
  8841=>"001000001",
  8842=>"010011010",
  8843=>"110100110",
  8844=>"001111100",
  8845=>"101110110",
  8846=>"111111101",
  8847=>"010011010",
  8848=>"001000011",
  8849=>"110100101",
  8850=>"000111011",
  8851=>"111001100",
  8852=>"101000111",
  8853=>"000110101",
  8854=>"100101110",
  8855=>"001000010",
  8856=>"110111110",
  8857=>"101101111",
  8858=>"001010001",
  8859=>"010011111",
  8860=>"001000000",
  8861=>"110101110",
  8862=>"011101010",
  8863=>"110001001",
  8864=>"110100011",
  8865=>"000110111",
  8866=>"111001011",
  8867=>"001111110",
  8868=>"001100111",
  8869=>"000101001",
  8870=>"111111101",
  8871=>"000111001",
  8872=>"000000110",
  8873=>"001100110",
  8874=>"001110000",
  8875=>"010001000",
  8876=>"110000000",
  8877=>"110111011",
  8878=>"110001110",
  8879=>"110110110",
  8880=>"011000100",
  8881=>"111001010",
  8882=>"001000101",
  8883=>"110011100",
  8884=>"010001000",
  8885=>"101110010",
  8886=>"100000111",
  8887=>"100110111",
  8888=>"101101000",
  8889=>"010101111",
  8890=>"100111100",
  8891=>"100100110",
  8892=>"100001010",
  8893=>"001000011",
  8894=>"110000101",
  8895=>"000000101",
  8896=>"101000101",
  8897=>"101100111",
  8898=>"010011101",
  8899=>"011010110",
  8900=>"010110001",
  8901=>"101111110",
  8902=>"000010011",
  8903=>"101111111",
  8904=>"010011101",
  8905=>"010011110",
  8906=>"101110110",
  8907=>"111111100",
  8908=>"010101011",
  8909=>"000001000",
  8910=>"110010110",
  8911=>"010000100",
  8912=>"110010100",
  8913=>"001000000",
  8914=>"100111101",
  8915=>"011000111",
  8916=>"111100001",
  8917=>"110000000",
  8918=>"100100101",
  8919=>"110110111",
  8920=>"001010101",
  8921=>"000000010",
  8922=>"111001000",
  8923=>"001010110",
  8924=>"110111101",
  8925=>"111100001",
  8926=>"000011010",
  8927=>"110001111",
  8928=>"010000101",
  8929=>"011010001",
  8930=>"110011000",
  8931=>"110001100",
  8932=>"100000000",
  8933=>"110011011",
  8934=>"010110100",
  8935=>"000000101",
  8936=>"000011110",
  8937=>"110110100",
  8938=>"110000000",
  8939=>"110011000",
  8940=>"000011100",
  8941=>"101111001",
  8942=>"000101111",
  8943=>"101111010",
  8944=>"001111111",
  8945=>"111100111",
  8946=>"100110011",
  8947=>"101101011",
  8948=>"000110010",
  8949=>"101000010",
  8950=>"110100000",
  8951=>"010110010",
  8952=>"001000000",
  8953=>"010100111",
  8954=>"101000001",
  8955=>"110111001",
  8956=>"101101111",
  8957=>"001111010",
  8958=>"101110000",
  8959=>"111001010",
  8960=>"111110101",
  8961=>"000110110",
  8962=>"111000110",
  8963=>"110110001",
  8964=>"001111010",
  8965=>"001001100",
  8966=>"011011111",
  8967=>"100101100",
  8968=>"010100010",
  8969=>"000001100",
  8970=>"111010110",
  8971=>"000101110",
  8972=>"010100000",
  8973=>"000000011",
  8974=>"000110001",
  8975=>"100010010",
  8976=>"000001111",
  8977=>"100010100",
  8978=>"001101100",
  8979=>"011011100",
  8980=>"011011000",
  8981=>"111110010",
  8982=>"101001011",
  8983=>"001010010",
  8984=>"010100001",
  8985=>"001100000",
  8986=>"000001110",
  8987=>"011111011",
  8988=>"010000110",
  8989=>"101011010",
  8990=>"111101111",
  8991=>"010010000",
  8992=>"010111011",
  8993=>"100010000",
  8994=>"101001101",
  8995=>"101011100",
  8996=>"111001111",
  8997=>"110000010",
  8998=>"101000001",
  8999=>"100111101",
  9000=>"111010001",
  9001=>"101001101",
  9002=>"111101101",
  9003=>"011000100",
  9004=>"011110000",
  9005=>"101000010",
  9006=>"000110100",
  9007=>"101101001",
  9008=>"101101011",
  9009=>"010000110",
  9010=>"100011010",
  9011=>"100111010",
  9012=>"011101111",
  9013=>"011110111",
  9014=>"111111101",
  9015=>"110110010",
  9016=>"101111010",
  9017=>"011001111",
  9018=>"110000100",
  9019=>"111010000",
  9020=>"111110110",
  9021=>"001011000",
  9022=>"010010011",
  9023=>"000111000",
  9024=>"010101001",
  9025=>"010011101",
  9026=>"010101010",
  9027=>"000000000",
  9028=>"110111101",
  9029=>"111010011",
  9030=>"101101001",
  9031=>"101000110",
  9032=>"111011000",
  9033=>"100011111",
  9034=>"101010100",
  9035=>"010100001",
  9036=>"101010100",
  9037=>"010000010",
  9038=>"010000000",
  9039=>"001000011",
  9040=>"101111110",
  9041=>"011111001",
  9042=>"001101000",
  9043=>"001000101",
  9044=>"111100110",
  9045=>"110001011",
  9046=>"111101101",
  9047=>"001011111",
  9048=>"110100011",
  9049=>"100010010",
  9050=>"111011011",
  9051=>"111110111",
  9052=>"110100000",
  9053=>"010100010",
  9054=>"011111000",
  9055=>"001000000",
  9056=>"101011101",
  9057=>"000001000",
  9058=>"011001100",
  9059=>"011101000",
  9060=>"110001010",
  9061=>"000101001",
  9062=>"000000101",
  9063=>"000110110",
  9064=>"111000001",
  9065=>"110111100",
  9066=>"000000110",
  9067=>"110110111",
  9068=>"011111000",
  9069=>"101101110",
  9070=>"000001010",
  9071=>"100011000",
  9072=>"000101110",
  9073=>"111110110",
  9074=>"010101111",
  9075=>"011110001",
  9076=>"111111101",
  9077=>"111110100",
  9078=>"110011011",
  9079=>"110010110",
  9080=>"010001000",
  9081=>"111110111",
  9082=>"101111010",
  9083=>"111101111",
  9084=>"011101000",
  9085=>"001000111",
  9086=>"001110110",
  9087=>"001010011",
  9088=>"101001111",
  9089=>"011010101",
  9090=>"000101000",
  9091=>"001101110",
  9092=>"101010011",
  9093=>"001111010",
  9094=>"000100001",
  9095=>"110010101",
  9096=>"000001000",
  9097=>"011011100",
  9098=>"000001110",
  9099=>"011110100",
  9100=>"010110001",
  9101=>"110111011",
  9102=>"110111101",
  9103=>"100011111",
  9104=>"101111111",
  9105=>"010111000",
  9106=>"000111111",
  9107=>"110000110",
  9108=>"101010000",
  9109=>"111011110",
  9110=>"010101110",
  9111=>"011000101",
  9112=>"010010110",
  9113=>"011101110",
  9114=>"011100101",
  9115=>"101110111",
  9116=>"010000011",
  9117=>"010000100",
  9118=>"011101110",
  9119=>"110111000",
  9120=>"011101011",
  9121=>"010111011",
  9122=>"101001011",
  9123=>"011100011",
  9124=>"100100100",
  9125=>"101111011",
  9126=>"011001010",
  9127=>"110010011",
  9128=>"001000110",
  9129=>"101101110",
  9130=>"101111001",
  9131=>"000111101",
  9132=>"101011001",
  9133=>"000010010",
  9134=>"111000101",
  9135=>"011010011",
  9136=>"101101001",
  9137=>"101100111",
  9138=>"101110100",
  9139=>"000000111",
  9140=>"111000000",
  9141=>"110010001",
  9142=>"010100110",
  9143=>"011011001",
  9144=>"000100101",
  9145=>"111101010",
  9146=>"110111110",
  9147=>"001001000",
  9148=>"011110110",
  9149=>"111100110",
  9150=>"001110011",
  9151=>"111111010",
  9152=>"000000000",
  9153=>"110111101",
  9154=>"000001001",
  9155=>"101010111",
  9156=>"111011010",
  9157=>"011111000",
  9158=>"001001101",
  9159=>"010010110",
  9160=>"101111110",
  9161=>"010111011",
  9162=>"010101000",
  9163=>"100111110",
  9164=>"010111011",
  9165=>"111100100",
  9166=>"101011101",
  9167=>"000111101",
  9168=>"100101101",
  9169=>"110010101",
  9170=>"111001000",
  9171=>"011110010",
  9172=>"010110100",
  9173=>"000010110",
  9174=>"001111010",
  9175=>"111111000",
  9176=>"111111100",
  9177=>"000000100",
  9178=>"110111101",
  9179=>"110101010",
  9180=>"110011000",
  9181=>"010001000",
  9182=>"000011111",
  9183=>"011000110",
  9184=>"000100011",
  9185=>"111101000",
  9186=>"001001100",
  9187=>"101011001",
  9188=>"000000111",
  9189=>"100100101",
  9190=>"011011010",
  9191=>"010011100",
  9192=>"000100000",
  9193=>"000100010",
  9194=>"010001001",
  9195=>"001001011",
  9196=>"010111011",
  9197=>"100100000",
  9198=>"101001010",
  9199=>"110100000",
  9200=>"010010111",
  9201=>"011100010",
  9202=>"011010011",
  9203=>"010100111",
  9204=>"010001100",
  9205=>"000010001",
  9206=>"101010101",
  9207=>"000101000",
  9208=>"011111010",
  9209=>"101011101",
  9210=>"010111011",
  9211=>"110110100",
  9212=>"110110101",
  9213=>"001011111",
  9214=>"111100001",
  9215=>"100010000",
  9216=>"111001001",
  9217=>"010111010",
  9218=>"010010011",
  9219=>"100010000",
  9220=>"010111111",
  9221=>"011000000",
  9222=>"011010111",
  9223=>"110111111",
  9224=>"100000000",
  9225=>"111100101",
  9226=>"111101101",
  9227=>"101011000",
  9228=>"001001011",
  9229=>"110001000",
  9230=>"001011111",
  9231=>"011110011",
  9232=>"010001010",
  9233=>"001101001",
  9234=>"110010000",
  9235=>"101001100",
  9236=>"001100000",
  9237=>"001001101",
  9238=>"011100110",
  9239=>"011010011",
  9240=>"000000110",
  9241=>"101001110",
  9242=>"011110000",
  9243=>"011001111",
  9244=>"100110010",
  9245=>"010000110",
  9246=>"001011111",
  9247=>"100011110",
  9248=>"100110010",
  9249=>"111110011",
  9250=>"011000111",
  9251=>"101000001",
  9252=>"100111101",
  9253=>"100010000",
  9254=>"010001000",
  9255=>"010100000",
  9256=>"000101011",
  9257=>"010011111",
  9258=>"011110111",
  9259=>"010010110",
  9260=>"111111000",
  9261=>"111000000",
  9262=>"001001011",
  9263=>"100011011",
  9264=>"111010100",
  9265=>"011000011",
  9266=>"010111111",
  9267=>"111011000",
  9268=>"000011000",
  9269=>"010111001",
  9270=>"000101110",
  9271=>"010111111",
  9272=>"011111000",
  9273=>"011100001",
  9274=>"010101111",
  9275=>"101001001",
  9276=>"100010111",
  9277=>"001010101",
  9278=>"000110101",
  9279=>"000101011",
  9280=>"000100000",
  9281=>"000111111",
  9282=>"001110010",
  9283=>"111100010",
  9284=>"110000001",
  9285=>"011111111",
  9286=>"110010011",
  9287=>"010010011",
  9288=>"111110010",
  9289=>"100000100",
  9290=>"100010000",
  9291=>"000001010",
  9292=>"110010101",
  9293=>"010111010",
  9294=>"100011111",
  9295=>"111111111",
  9296=>"001111100",
  9297=>"010101110",
  9298=>"100101110",
  9299=>"000101100",
  9300=>"010100010",
  9301=>"111000110",
  9302=>"011100001",
  9303=>"111101001",
  9304=>"001111100",
  9305=>"111101101",
  9306=>"001011010",
  9307=>"000001001",
  9308=>"111100111",
  9309=>"010101001",
  9310=>"100110001",
  9311=>"001001101",
  9312=>"000111110",
  9313=>"000111010",
  9314=>"111011011",
  9315=>"101111101",
  9316=>"100110000",
  9317=>"110111111",
  9318=>"110111101",
  9319=>"001010011",
  9320=>"110001001",
  9321=>"011111001",
  9322=>"011100100",
  9323=>"111111101",
  9324=>"100011010",
  9325=>"111000011",
  9326=>"010011001",
  9327=>"001100111",
  9328=>"111100111",
  9329=>"001100110",
  9330=>"100111001",
  9331=>"001010001",
  9332=>"101011101",
  9333=>"100010111",
  9334=>"110100111",
  9335=>"010001110",
  9336=>"101000000",
  9337=>"111111100",
  9338=>"110011110",
  9339=>"000101111",
  9340=>"011100110",
  9341=>"011111100",
  9342=>"010001010",
  9343=>"111001010",
  9344=>"100010101",
  9345=>"100011000",
  9346=>"000001001",
  9347=>"000001101",
  9348=>"110100101",
  9349=>"001010101",
  9350=>"111010100",
  9351=>"101111111",
  9352=>"100001111",
  9353=>"101000000",
  9354=>"011100010",
  9355=>"101000100",
  9356=>"010111101",
  9357=>"000110101",
  9358=>"111010101",
  9359=>"010101110",
  9360=>"010101111",
  9361=>"010010111",
  9362=>"010011001",
  9363=>"111001111",
  9364=>"111110111",
  9365=>"011110010",
  9366=>"111110100",
  9367=>"010111011",
  9368=>"110011010",
  9369=>"010010101",
  9370=>"011101110",
  9371=>"100110001",
  9372=>"101011011",
  9373=>"001011001",
  9374=>"000011011",
  9375=>"011010001",
  9376=>"010100110",
  9377=>"010011010",
  9378=>"010010101",
  9379=>"010110000",
  9380=>"001011101",
  9381=>"010100000",
  9382=>"001000010",
  9383=>"011001001",
  9384=>"110101001",
  9385=>"100010011",
  9386=>"010000010",
  9387=>"000000001",
  9388=>"000101010",
  9389=>"011101010",
  9390=>"001010111",
  9391=>"000101000",
  9392=>"101010011",
  9393=>"110110000",
  9394=>"010110011",
  9395=>"011010111",
  9396=>"111110111",
  9397=>"100110000",
  9398=>"111011011",
  9399=>"110111111",
  9400=>"100010011",
  9401=>"010101010",
  9402=>"000011111",
  9403=>"111010010",
  9404=>"101101110",
  9405=>"000100011",
  9406=>"101010000",
  9407=>"001011000",
  9408=>"100111111",
  9409=>"011001111",
  9410=>"011000011",
  9411=>"010000100",
  9412=>"001000111",
  9413=>"101100110",
  9414=>"001101111",
  9415=>"000111011",
  9416=>"110001010",
  9417=>"100110100",
  9418=>"000010000",
  9419=>"101111011",
  9420=>"101010011",
  9421=>"000110110",
  9422=>"010101010",
  9423=>"100100100",
  9424=>"110001111",
  9425=>"011001101",
  9426=>"100000001",
  9427=>"100011001",
  9428=>"011110100",
  9429=>"011111111",
  9430=>"010011011",
  9431=>"101111001",
  9432=>"010111110",
  9433=>"011111110",
  9434=>"000001000",
  9435=>"111100101",
  9436=>"011110011",
  9437=>"111001101",
  9438=>"100100111",
  9439=>"101110000",
  9440=>"001010110",
  9441=>"111101010",
  9442=>"101001111",
  9443=>"001010111",
  9444=>"011110010",
  9445=>"000001001",
  9446=>"001000011",
  9447=>"010010001",
  9448=>"011111011",
  9449=>"110111111",
  9450=>"111000110",
  9451=>"011000110",
  9452=>"100111110",
  9453=>"010001111",
  9454=>"000000110",
  9455=>"100010100",
  9456=>"101110110",
  9457=>"100010101",
  9458=>"001001011",
  9459=>"000010011",
  9460=>"010101111",
  9461=>"011011101",
  9462=>"110011000",
  9463=>"011101101",
  9464=>"001101111",
  9465=>"011000110",
  9466=>"011110011",
  9467=>"110100101",
  9468=>"011000000",
  9469=>"000001110",
  9470=>"000100001",
  9471=>"111111011",
  9472=>"101011110",
  9473=>"110010010",
  9474=>"010100011",
  9475=>"010101011",
  9476=>"101010000",
  9477=>"111110111",
  9478=>"111110001",
  9479=>"101000100",
  9480=>"011101011",
  9481=>"100000000",
  9482=>"100001110",
  9483=>"111010000",
  9484=>"010001111",
  9485=>"001010011",
  9486=>"010011011",
  9487=>"101101100",
  9488=>"110101100",
  9489=>"010101010",
  9490=>"000100101",
  9491=>"101010000",
  9492=>"101111100",
  9493=>"111001001",
  9494=>"000000000",
  9495=>"111000000",
  9496=>"001111111",
  9497=>"011001000",
  9498=>"111100011",
  9499=>"111101001",
  9500=>"100110010",
  9501=>"011000110",
  9502=>"001001001",
  9503=>"011101011",
  9504=>"000101010",
  9505=>"111111011",
  9506=>"000000100",
  9507=>"100010011",
  9508=>"101010111",
  9509=>"101011100",
  9510=>"000011111",
  9511=>"101011011",
  9512=>"111011111",
  9513=>"110110111",
  9514=>"110110101",
  9515=>"100000001",
  9516=>"101110100",
  9517=>"000000101",
  9518=>"001001101",
  9519=>"100110111",
  9520=>"000010100",
  9521=>"001011100",
  9522=>"111001111",
  9523=>"010001100",
  9524=>"001000101",
  9525=>"001001011",
  9526=>"001111101",
  9527=>"010100111",
  9528=>"001111100",
  9529=>"010011000",
  9530=>"101111011",
  9531=>"100011000",
  9532=>"000001111",
  9533=>"011110001",
  9534=>"011000011",
  9535=>"110010001",
  9536=>"011110100",
  9537=>"000011101",
  9538=>"111101110",
  9539=>"110101000",
  9540=>"111100100",
  9541=>"110001010",
  9542=>"000100110",
  9543=>"111001001",
  9544=>"001000101",
  9545=>"001010100",
  9546=>"101011101",
  9547=>"000100000",
  9548=>"011011101",
  9549=>"010010000",
  9550=>"100101011",
  9551=>"001100000",
  9552=>"001101001",
  9553=>"011110011",
  9554=>"010100100",
  9555=>"010110010",
  9556=>"010101111",
  9557=>"100011111",
  9558=>"000111001",
  9559=>"010101011",
  9560=>"101100011",
  9561=>"110011010",
  9562=>"011100100",
  9563=>"100000000",
  9564=>"010000011",
  9565=>"000100111",
  9566=>"100010000",
  9567=>"010111011",
  9568=>"000001110",
  9569=>"100110100",
  9570=>"000000001",
  9571=>"111101000",
  9572=>"111101011",
  9573=>"111101011",
  9574=>"000010000",
  9575=>"100000000",
  9576=>"000111011",
  9577=>"011100111",
  9578=>"010111010",
  9579=>"000101111",
  9580=>"100000011",
  9581=>"001001000",
  9582=>"000110000",
  9583=>"100010000",
  9584=>"001100001",
  9585=>"011000100",
  9586=>"101111001",
  9587=>"010110111",
  9588=>"100100011",
  9589=>"101111011",
  9590=>"010000010",
  9591=>"101000011",
  9592=>"000110000",
  9593=>"000000010",
  9594=>"011001000",
  9595=>"110001101",
  9596=>"010100111",
  9597=>"010100011",
  9598=>"000011110",
  9599=>"000100010",
  9600=>"000010001",
  9601=>"000101110",
  9602=>"111010001",
  9603=>"010101010",
  9604=>"111000001",
  9605=>"001111010",
  9606=>"100010100",
  9607=>"000111100",
  9608=>"000011111",
  9609=>"000001100",
  9610=>"101001001",
  9611=>"011000010",
  9612=>"011101111",
  9613=>"000000110",
  9614=>"011011011",
  9615=>"111101110",
  9616=>"011110011",
  9617=>"010000011",
  9618=>"000110110",
  9619=>"110111011",
  9620=>"100000100",
  9621=>"101000000",
  9622=>"100011111",
  9623=>"110011111",
  9624=>"010111000",
  9625=>"011001000",
  9626=>"011001100",
  9627=>"001000001",
  9628=>"010011100",
  9629=>"111011111",
  9630=>"100000101",
  9631=>"010010100",
  9632=>"101111111",
  9633=>"011111001",
  9634=>"111110100",
  9635=>"101101101",
  9636=>"011010010",
  9637=>"110101000",
  9638=>"011110010",
  9639=>"010000000",
  9640=>"100101101",
  9641=>"101001011",
  9642=>"000000110",
  9643=>"000011000",
  9644=>"010101111",
  9645=>"010100011",
  9646=>"101101100",
  9647=>"011100101",
  9648=>"010101010",
  9649=>"001001111",
  9650=>"011000011",
  9651=>"111010010",
  9652=>"010010111",
  9653=>"101110001",
  9654=>"110001110",
  9655=>"010111000",
  9656=>"000011110",
  9657=>"010101110",
  9658=>"001010010",
  9659=>"000100100",
  9660=>"111111110",
  9661=>"011100000",
  9662=>"101111111",
  9663=>"100011011",
  9664=>"100010000",
  9665=>"001010010",
  9666=>"000011101",
  9667=>"101110001",
  9668=>"101011101",
  9669=>"001111001",
  9670=>"011111111",
  9671=>"110110010",
  9672=>"010010101",
  9673=>"101101100",
  9674=>"000000011",
  9675=>"110101101",
  9676=>"011110111",
  9677=>"010100100",
  9678=>"100110110",
  9679=>"010010010",
  9680=>"011011011",
  9681=>"001001001",
  9682=>"100000110",
  9683=>"010001100",
  9684=>"001010100",
  9685=>"111001100",
  9686=>"111011011",
  9687=>"111000000",
  9688=>"000111011",
  9689=>"111101100",
  9690=>"000101101",
  9691=>"000000101",
  9692=>"001110111",
  9693=>"011010000",
  9694=>"111000110",
  9695=>"111111011",
  9696=>"000110100",
  9697=>"011101111",
  9698=>"111101111",
  9699=>"011010100",
  9700=>"100000101",
  9701=>"011110111",
  9702=>"010001000",
  9703=>"111110000",
  9704=>"001001001",
  9705=>"000001110",
  9706=>"000101110",
  9707=>"010101100",
  9708=>"000011010",
  9709=>"000011011",
  9710=>"010110010",
  9711=>"001010110",
  9712=>"111100101",
  9713=>"001111110",
  9714=>"100001000",
  9715=>"100010100",
  9716=>"100101111",
  9717=>"111011000",
  9718=>"001000101",
  9719=>"100100001",
  9720=>"010001101",
  9721=>"111010100",
  9722=>"110101101",
  9723=>"101001001",
  9724=>"000111111",
  9725=>"111010111",
  9726=>"001011111",
  9727=>"000000000",
  9728=>"010101001",
  9729=>"001100001",
  9730=>"101110111",
  9731=>"000010000",
  9732=>"011011110",
  9733=>"100111110",
  9734=>"010110000",
  9735=>"000001011",
  9736=>"101101011",
  9737=>"100010010",
  9738=>"010010101",
  9739=>"111110110",
  9740=>"110010111",
  9741=>"000010110",
  9742=>"111111000",
  9743=>"111101001",
  9744=>"000001101",
  9745=>"111011100",
  9746=>"000100010",
  9747=>"011100011",
  9748=>"101101110",
  9749=>"010011111",
  9750=>"011111100",
  9751=>"111011000",
  9752=>"110101011",
  9753=>"001100100",
  9754=>"111101000",
  9755=>"111100000",
  9756=>"001010101",
  9757=>"100000001",
  9758=>"000000000",
  9759=>"011000001",
  9760=>"010010100",
  9761=>"000011100",
  9762=>"000010110",
  9763=>"000100000",
  9764=>"100111110",
  9765=>"000000100",
  9766=>"100101100",
  9767=>"000001000",
  9768=>"000101011",
  9769=>"101100110",
  9770=>"100100000",
  9771=>"110011100",
  9772=>"000111111",
  9773=>"100000101",
  9774=>"000111010",
  9775=>"101011001",
  9776=>"001000011",
  9777=>"110110101",
  9778=>"001000011",
  9779=>"011110111",
  9780=>"101100010",
  9781=>"001010001",
  9782=>"100001100",
  9783=>"110010010",
  9784=>"010101000",
  9785=>"001110010",
  9786=>"100000000",
  9787=>"001101011",
  9788=>"100011100",
  9789=>"100001100",
  9790=>"010100001",
  9791=>"001011000",
  9792=>"001101100",
  9793=>"111010111",
  9794=>"001010100",
  9795=>"110110000",
  9796=>"101110101",
  9797=>"111101001",
  9798=>"001010100",
  9799=>"100000100",
  9800=>"011011111",
  9801=>"110100011",
  9802=>"000001110",
  9803=>"001100000",
  9804=>"101011001",
  9805=>"000010100",
  9806=>"001011010",
  9807=>"101010001",
  9808=>"101100001",
  9809=>"000110100",
  9810=>"001000010",
  9811=>"010010100",
  9812=>"011100111",
  9813=>"010010011",
  9814=>"111111100",
  9815=>"001001011",
  9816=>"011110100",
  9817=>"110001011",
  9818=>"101001011",
  9819=>"000010000",
  9820=>"101000001",
  9821=>"100001010",
  9822=>"000000111",
  9823=>"010101001",
  9824=>"101000001",
  9825=>"000011010",
  9826=>"111110000",
  9827=>"111100101",
  9828=>"011100010",
  9829=>"101010100",
  9830=>"111011110",
  9831=>"100000010",
  9832=>"001001001",
  9833=>"111110010",
  9834=>"001001000",
  9835=>"111110101",
  9836=>"100010011",
  9837=>"010111011",
  9838=>"000111000",
  9839=>"001010100",
  9840=>"101000010",
  9841=>"101110101",
  9842=>"100000010",
  9843=>"101100100",
  9844=>"100101110",
  9845=>"111100010",
  9846=>"101010111",
  9847=>"000010110",
  9848=>"111010001",
  9849=>"110000010",
  9850=>"011011001",
  9851=>"101000100",
  9852=>"000000101",
  9853=>"001110100",
  9854=>"000001000",
  9855=>"000111011",
  9856=>"010011010",
  9857=>"000011000",
  9858=>"001001100",
  9859=>"000000101",
  9860=>"011011101",
  9861=>"111011110",
  9862=>"110000110",
  9863=>"101110000",
  9864=>"110011010",
  9865=>"100000111",
  9866=>"100111111",
  9867=>"010110001",
  9868=>"001110010",
  9869=>"001000110",
  9870=>"111101000",
  9871=>"101101111",
  9872=>"111010110",
  9873=>"000011111",
  9874=>"001010000",
  9875=>"011110011",
  9876=>"111110111",
  9877=>"001011100",
  9878=>"101101001",
  9879=>"110111011",
  9880=>"000010110",
  9881=>"000001010",
  9882=>"100011001",
  9883=>"011001001",
  9884=>"100011011",
  9885=>"011011101",
  9886=>"111101111",
  9887=>"111000011",
  9888=>"111011001",
  9889=>"011100101",
  9890=>"101100011",
  9891=>"011011001",
  9892=>"001010000",
  9893=>"100101101",
  9894=>"100010001",
  9895=>"100001000",
  9896=>"111001000",
  9897=>"111101010",
  9898=>"110111101",
  9899=>"000000000",
  9900=>"010011100",
  9901=>"011001110",
  9902=>"011010011",
  9903=>"110101100",
  9904=>"101000101",
  9905=>"110111111",
  9906=>"110100100",
  9907=>"100010100",
  9908=>"100010111",
  9909=>"101101110",
  9910=>"010010010",
  9911=>"001011110",
  9912=>"001110100",
  9913=>"100111110",
  9914=>"010100001",
  9915=>"001001001",
  9916=>"001000101",
  9917=>"100110000",
  9918=>"010011100",
  9919=>"100010000",
  9920=>"000110011",
  9921=>"101100111",
  9922=>"100100010",
  9923=>"111100000",
  9924=>"000000011",
  9925=>"110001000",
  9926=>"101001010",
  9927=>"000010001",
  9928=>"111010111",
  9929=>"101000001",
  9930=>"101101001",
  9931=>"000000101",
  9932=>"011110010",
  9933=>"010011010",
  9934=>"110011110",
  9935=>"111110011",
  9936=>"011000100",
  9937=>"111000100",
  9938=>"011110100",
  9939=>"011111101",
  9940=>"101111101",
  9941=>"011001010",
  9942=>"111100101",
  9943=>"100000000",
  9944=>"000101010",
  9945=>"010100000",
  9946=>"000001000",
  9947=>"101111110",
  9948=>"101101010",
  9949=>"001001011",
  9950=>"001101011",
  9951=>"010010000",
  9952=>"000010111",
  9953=>"001000000",
  9954=>"000100011",
  9955=>"000101100",
  9956=>"010010111",
  9957=>"011000111",
  9958=>"011101011",
  9959=>"110000000",
  9960=>"000100110",
  9961=>"000010001",
  9962=>"110110110",
  9963=>"111111101",
  9964=>"110000001",
  9965=>"110010000",
  9966=>"101101010",
  9967=>"110101011",
  9968=>"000111101",
  9969=>"010100000",
  9970=>"100001011",
  9971=>"011101010",
  9972=>"010100100",
  9973=>"001001101",
  9974=>"111110010",
  9975=>"010110010",
  9976=>"011111000",
  9977=>"001011101",
  9978=>"000110011",
  9979=>"011000010",
  9980=>"011001000",
  9981=>"111011011",
  9982=>"011110011",
  9983=>"010010110",
  9984=>"101110100",
  9985=>"111101111",
  9986=>"101011000",
  9987=>"100010100",
  9988=>"100011100",
  9989=>"001100110",
  9990=>"001101000",
  9991=>"100110010",
  9992=>"010000010",
  9993=>"011111111",
  9994=>"010100100",
  9995=>"000001000",
  9996=>"111110111",
  9997=>"100111100",
  9998=>"100101011",
  9999=>"000001001",
  10000=>"110000011",
  10001=>"000001101",
  10002=>"001001100",
  10003=>"010001000",
  10004=>"101110100",
  10005=>"110101011",
  10006=>"110100001",
  10007=>"010001000",
  10008=>"000100011",
  10009=>"110010010",
  10010=>"000110100",
  10011=>"101010110",
  10012=>"011001010",
  10013=>"000000101",
  10014=>"101110110",
  10015=>"111010000",
  10016=>"001100101",
  10017=>"011111100",
  10018=>"000000110",
  10019=>"100100111",
  10020=>"011011011",
  10021=>"010111001",
  10022=>"000010001",
  10023=>"111101101",
  10024=>"010000100",
  10025=>"111011101",
  10026=>"011011111",
  10027=>"100010100",
  10028=>"000110001",
  10029=>"010000000",
  10030=>"000011001",
  10031=>"001100001",
  10032=>"100101110",
  10033=>"011011111",
  10034=>"101010000",
  10035=>"111001010",
  10036=>"110111111",
  10037=>"110001011",
  10038=>"000101011",
  10039=>"001110111",
  10040=>"011100011",
  10041=>"101001000",
  10042=>"001110110",
  10043=>"111110011",
  10044=>"111001101",
  10045=>"101000011",
  10046=>"111001110",
  10047=>"101110001",
  10048=>"010001011",
  10049=>"111000000",
  10050=>"111010111",
  10051=>"000010111",
  10052=>"011001101",
  10053=>"100101110",
  10054=>"110110011",
  10055=>"000000101",
  10056=>"001000011",
  10057=>"010010001",
  10058=>"001010101",
  10059=>"110000000",
  10060=>"000010111",
  10061=>"110101000",
  10062=>"110000000",
  10063=>"111111010",
  10064=>"011000000",
  10065=>"010110010",
  10066=>"000000011",
  10067=>"011001000",
  10068=>"100000011",
  10069=>"010011000",
  10070=>"110100010",
  10071=>"100110110",
  10072=>"000000100",
  10073=>"101000011",
  10074=>"001111010",
  10075=>"000001000",
  10076=>"101100001",
  10077=>"000010110",
  10078=>"110100011",
  10079=>"000001101",
  10080=>"011011010",
  10081=>"111001000",
  10082=>"000010100",
  10083=>"101011010",
  10084=>"101111001",
  10085=>"111101101",
  10086=>"111000011",
  10087=>"110100100",
  10088=>"010101010",
  10089=>"010000011",
  10090=>"010101100",
  10091=>"010000111",
  10092=>"100001110",
  10093=>"111011011",
  10094=>"000001110",
  10095=>"101010000",
  10096=>"000101100",
  10097=>"011011000",
  10098=>"011001001",
  10099=>"000110010",
  10100=>"111010010",
  10101=>"100100011",
  10102=>"100001100",
  10103=>"001000111",
  10104=>"111010001",
  10105=>"011100011",
  10106=>"111100110",
  10107=>"101100110",
  10108=>"111001111",
  10109=>"100011010",
  10110=>"000001000",
  10111=>"011111101",
  10112=>"101011111",
  10113=>"100011111",
  10114=>"001101000",
  10115=>"001101101",
  10116=>"001100001",
  10117=>"001011000",
  10118=>"111011111",
  10119=>"101011111",
  10120=>"000000101",
  10121=>"101011100",
  10122=>"101001111",
  10123=>"111101111",
  10124=>"100101011",
  10125=>"010100000",
  10126=>"001000111",
  10127=>"110011001",
  10128=>"110100101",
  10129=>"000010001",
  10130=>"011101010",
  10131=>"010010000",
  10132=>"110111111",
  10133=>"011010011",
  10134=>"101111011",
  10135=>"001000110",
  10136=>"111010000",
  10137=>"000000011",
  10138=>"000100111",
  10139=>"101000110",
  10140=>"100110100",
  10141=>"010001010",
  10142=>"001000001",
  10143=>"100110110",
  10144=>"011111011",
  10145=>"101111100",
  10146=>"011100101",
  10147=>"011100010",
  10148=>"111011101",
  10149=>"100011100",
  10150=>"110100111",
  10151=>"011000110",
  10152=>"110011110",
  10153=>"000101001",
  10154=>"101001010",
  10155=>"111100111",
  10156=>"000110111",
  10157=>"111100010",
  10158=>"100110000",
  10159=>"001100001",
  10160=>"100110101",
  10161=>"001101011",
  10162=>"111111110",
  10163=>"111101011",
  10164=>"111110000",
  10165=>"010100011",
  10166=>"000101010",
  10167=>"000110111",
  10168=>"000100101",
  10169=>"111000100",
  10170=>"110110011",
  10171=>"001000100",
  10172=>"010100011",
  10173=>"001010100",
  10174=>"111110001",
  10175=>"011101111",
  10176=>"110010001",
  10177=>"110100100",
  10178=>"110000110",
  10179=>"101011101",
  10180=>"101110000",
  10181=>"010001001",
  10182=>"101011111",
  10183=>"111101110",
  10184=>"011000110",
  10185=>"100110011",
  10186=>"011000101",
  10187=>"111000111",
  10188=>"000000111",
  10189=>"111110111",
  10190=>"011111000",
  10191=>"101000001",
  10192=>"101110011",
  10193=>"111111100",
  10194=>"110101101",
  10195=>"010100000",
  10196=>"111111111",
  10197=>"011100001",
  10198=>"000000001",
  10199=>"111001010",
  10200=>"000100101",
  10201=>"011110101",
  10202=>"000100100",
  10203=>"010010101",
  10204=>"110110110",
  10205=>"010110101",
  10206=>"101001110",
  10207=>"001000010",
  10208=>"111100011",
  10209=>"110010001",
  10210=>"110111111",
  10211=>"100110000",
  10212=>"110111110",
  10213=>"101011111",
  10214=>"001010111",
  10215=>"101010001",
  10216=>"111001000",
  10217=>"101011001",
  10218=>"010010011",
  10219=>"110010010",
  10220=>"001100010",
  10221=>"111000100",
  10222=>"001111000",
  10223=>"010110000",
  10224=>"111001110",
  10225=>"000000100",
  10226=>"101101010",
  10227=>"101100100",
  10228=>"011010101",
  10229=>"011000001",
  10230=>"011101000",
  10231=>"000010000",
  10232=>"000010001",
  10233=>"000001101",
  10234=>"111111000",
  10235=>"100101000",
  10236=>"000001010",
  10237=>"110111000",
  10238=>"110101010",
  10239=>"011000101",
  10240=>"101111101",
  10241=>"000011111",
  10242=>"001111111",
  10243=>"111000110",
  10244=>"011000111",
  10245=>"101000001",
  10246=>"110010010",
  10247=>"000010100",
  10248=>"110100111",
  10249=>"111001110",
  10250=>"101011010",
  10251=>"010110111",
  10252=>"000100100",
  10253=>"000101000",
  10254=>"000110011",
  10255=>"001010111",
  10256=>"100010101",
  10257=>"001110100",
  10258=>"011000101",
  10259=>"110111110",
  10260=>"001111111",
  10261=>"100101000",
  10262=>"101000111",
  10263=>"000001110",
  10264=>"111101001",
  10265=>"010000110",
  10266=>"001101000",
  10267=>"000001000",
  10268=>"100001100",
  10269=>"101000000",
  10270=>"011010100",
  10271=>"000010100",
  10272=>"001001000",
  10273=>"110111111",
  10274=>"101000010",
  10275=>"001111111",
  10276=>"000011110",
  10277=>"001100101",
  10278=>"111110001",
  10279=>"101111101",
  10280=>"011000000",
  10281=>"010000000",
  10282=>"011010101",
  10283=>"101000011",
  10284=>"101010100",
  10285=>"000100100",
  10286=>"101011000",
  10287=>"101000101",
  10288=>"011111110",
  10289=>"100010000",
  10290=>"000001001",
  10291=>"101011000",
  10292=>"000000010",
  10293=>"000101011",
  10294=>"100111000",
  10295=>"011111100",
  10296=>"101111000",
  10297=>"010011101",
  10298=>"100011100",
  10299=>"100100100",
  10300=>"001110010",
  10301=>"010110001",
  10302=>"100000010",
  10303=>"111000100",
  10304=>"000010110",
  10305=>"000000001",
  10306=>"110011111",
  10307=>"110010000",
  10308=>"110100011",
  10309=>"111010111",
  10310=>"010010010",
  10311=>"101000101",
  10312=>"000110011",
  10313=>"011000011",
  10314=>"000110010",
  10315=>"111111011",
  10316=>"100100000",
  10317=>"101011001",
  10318=>"111100100",
  10319=>"000110011",
  10320=>"011000001",
  10321=>"111111111",
  10322=>"001110110",
  10323=>"011001110",
  10324=>"011111101",
  10325=>"000000001",
  10326=>"000001000",
  10327=>"100110001",
  10328=>"001001100",
  10329=>"110111101",
  10330=>"100000011",
  10331=>"100100111",
  10332=>"101100010",
  10333=>"110011101",
  10334=>"000010111",
  10335=>"010000000",
  10336=>"111111101",
  10337=>"011101100",
  10338=>"101001000",
  10339=>"010010000",
  10340=>"011111110",
  10341=>"000011000",
  10342=>"011011000",
  10343=>"000010100",
  10344=>"111000110",
  10345=>"000101011",
  10346=>"000011010",
  10347=>"111011010",
  10348=>"101100100",
  10349=>"001100010",
  10350=>"010110110",
  10351=>"110100111",
  10352=>"101110111",
  10353=>"011100100",
  10354=>"011000001",
  10355=>"110101000",
  10356=>"111001110",
  10357=>"010001110",
  10358=>"110010110",
  10359=>"101011011",
  10360=>"111010000",
  10361=>"011011110",
  10362=>"100000100",
  10363=>"011001101",
  10364=>"111010100",
  10365=>"001000000",
  10366=>"101101111",
  10367=>"100011011",
  10368=>"100110000",
  10369=>"111101010",
  10370=>"010000011",
  10371=>"011100101",
  10372=>"001010000",
  10373=>"011100100",
  10374=>"110011111",
  10375=>"100111000",
  10376=>"101010100",
  10377=>"010101110",
  10378=>"010001101",
  10379=>"010111010",
  10380=>"010101100",
  10381=>"111001110",
  10382=>"110001011",
  10383=>"100010000",
  10384=>"011011111",
  10385=>"001010101",
  10386=>"010011010",
  10387=>"110110001",
  10388=>"111101111",
  10389=>"000101001",
  10390=>"110010001",
  10391=>"111111000",
  10392=>"000001011",
  10393=>"011100110",
  10394=>"000100101",
  10395=>"110010001",
  10396=>"100010001",
  10397=>"101000100",
  10398=>"011110010",
  10399=>"100111110",
  10400=>"010110111",
  10401=>"101101100",
  10402=>"110111100",
  10403=>"011011111",
  10404=>"001111010",
  10405=>"101000111",
  10406=>"111001111",
  10407=>"011011101",
  10408=>"111101111",
  10409=>"101101101",
  10410=>"101110011",
  10411=>"010111101",
  10412=>"010010010",
  10413=>"110101110",
  10414=>"101100111",
  10415=>"010000011",
  10416=>"111010111",
  10417=>"111000100",
  10418=>"011101100",
  10419=>"101101100",
  10420=>"001101111",
  10421=>"101011011",
  10422=>"100111100",
  10423=>"001000011",
  10424=>"101010000",
  10425=>"000000001",
  10426=>"010001101",
  10427=>"010010000",
  10428=>"001001010",
  10429=>"110011100",
  10430=>"000101100",
  10431=>"010100011",
  10432=>"011110010",
  10433=>"010000101",
  10434=>"001000101",
  10435=>"000000001",
  10436=>"111110000",
  10437=>"000100111",
  10438=>"111101011",
  10439=>"101010010",
  10440=>"010001000",
  10441=>"000101000",
  10442=>"100010100",
  10443=>"101111001",
  10444=>"010000001",
  10445=>"011101101",
  10446=>"111111110",
  10447=>"001001011",
  10448=>"111001111",
  10449=>"100101011",
  10450=>"100010011",
  10451=>"101101101",
  10452=>"000000001",
  10453=>"010110111",
  10454=>"011010000",
  10455=>"111001000",
  10456=>"101000100",
  10457=>"101110000",
  10458=>"000110011",
  10459=>"011010111",
  10460=>"010010001",
  10461=>"110000101",
  10462=>"111001000",
  10463=>"000111101",
  10464=>"101101100",
  10465=>"001110101",
  10466=>"011100110",
  10467=>"101000000",
  10468=>"100100000",
  10469=>"110001010",
  10470=>"101100001",
  10471=>"001100010",
  10472=>"000001101",
  10473=>"100101110",
  10474=>"000111111",
  10475=>"111100000",
  10476=>"000011110",
  10477=>"110110011",
  10478=>"001100101",
  10479=>"001000000",
  10480=>"001001010",
  10481=>"101100000",
  10482=>"010111111",
  10483=>"110001111",
  10484=>"011101000",
  10485=>"100010011",
  10486=>"011010111",
  10487=>"000001111",
  10488=>"101101111",
  10489=>"000101111",
  10490=>"101000010",
  10491=>"010101000",
  10492=>"010100001",
  10493=>"010100111",
  10494=>"001111011",
  10495=>"011001001",
  10496=>"111010111",
  10497=>"011111101",
  10498=>"101101010",
  10499=>"100001011",
  10500=>"110101000",
  10501=>"001110000",
  10502=>"010111100",
  10503=>"101000101",
  10504=>"100110101",
  10505=>"110000111",
  10506=>"011101010",
  10507=>"010110010",
  10508=>"010011111",
  10509=>"000011101",
  10510=>"101111011",
  10511=>"100100101",
  10512=>"000011010",
  10513=>"000011111",
  10514=>"111111101",
  10515=>"101101010",
  10516=>"101000101",
  10517=>"100111000",
  10518=>"110010110",
  10519=>"111011110",
  10520=>"000111111",
  10521=>"111010110",
  10522=>"101100110",
  10523=>"101101001",
  10524=>"000110101",
  10525=>"001000001",
  10526=>"100111010",
  10527=>"000101001",
  10528=>"010010001",
  10529=>"110010110",
  10530=>"100100001",
  10531=>"000011001",
  10532=>"010000011",
  10533=>"111001000",
  10534=>"111011101",
  10535=>"010011011",
  10536=>"100110000",
  10537=>"001010100",
  10538=>"011000000",
  10539=>"010110000",
  10540=>"110100000",
  10541=>"011010100",
  10542=>"010010011",
  10543=>"000110110",
  10544=>"101000100",
  10545=>"100010010",
  10546=>"101010100",
  10547=>"010010011",
  10548=>"010010111",
  10549=>"011111000",
  10550=>"011010110",
  10551=>"010000101",
  10552=>"110000111",
  10553=>"101000000",
  10554=>"110011111",
  10555=>"110001010",
  10556=>"010001010",
  10557=>"100101101",
  10558=>"111110111",
  10559=>"100011000",
  10560=>"100011011",
  10561=>"011001100",
  10562=>"000101001",
  10563=>"010100110",
  10564=>"000111111",
  10565=>"111000101",
  10566=>"001000011",
  10567=>"111001000",
  10568=>"010101110",
  10569=>"000100111",
  10570=>"001001101",
  10571=>"011111110",
  10572=>"101101000",
  10573=>"000001011",
  10574=>"100111001",
  10575=>"000011010",
  10576=>"111001110",
  10577=>"101011100",
  10578=>"111001100",
  10579=>"010111100",
  10580=>"011001001",
  10581=>"110010001",
  10582=>"010011111",
  10583=>"001000011",
  10584=>"011011100",
  10585=>"000110100",
  10586=>"111001110",
  10587=>"000010010",
  10588=>"111110101",
  10589=>"001000010",
  10590=>"000101110",
  10591=>"011010101",
  10592=>"100000011",
  10593=>"000001011",
  10594=>"010111000",
  10595=>"001001010",
  10596=>"010000100",
  10597=>"110110110",
  10598=>"101101001",
  10599=>"000010100",
  10600=>"111001001",
  10601=>"000000111",
  10602=>"111001111",
  10603=>"101000001",
  10604=>"010111111",
  10605=>"110111000",
  10606=>"101000110",
  10607=>"010101011",
  10608=>"100000010",
  10609=>"000011000",
  10610=>"010010010",
  10611=>"011010010",
  10612=>"110010100",
  10613=>"000110111",
  10614=>"101101110",
  10615=>"111010010",
  10616=>"100111010",
  10617=>"001010111",
  10618=>"110100110",
  10619=>"101010111",
  10620=>"000100100",
  10621=>"000111010",
  10622=>"011011011",
  10623=>"110100011",
  10624=>"110010000",
  10625=>"011001010",
  10626=>"100011111",
  10627=>"011100100",
  10628=>"011100000",
  10629=>"100000010",
  10630=>"101111101",
  10631=>"000011100",
  10632=>"000001100",
  10633=>"011010001",
  10634=>"100000011",
  10635=>"011011001",
  10636=>"100101100",
  10637=>"101101111",
  10638=>"100100000",
  10639=>"100100011",
  10640=>"100000011",
  10641=>"001001110",
  10642=>"010011100",
  10643=>"001100100",
  10644=>"010011100",
  10645=>"101000011",
  10646=>"101010000",
  10647=>"000111101",
  10648=>"000010001",
  10649=>"000001100",
  10650=>"111000011",
  10651=>"000010001",
  10652=>"000011111",
  10653=>"011101111",
  10654=>"111111111",
  10655=>"001101010",
  10656=>"100101000",
  10657=>"010110110",
  10658=>"011110001",
  10659=>"010111000",
  10660=>"110110010",
  10661=>"001000000",
  10662=>"111000100",
  10663=>"101001010",
  10664=>"100001110",
  10665=>"000001000",
  10666=>"000010110",
  10667=>"000001101",
  10668=>"000001110",
  10669=>"100110011",
  10670=>"111100010",
  10671=>"111111010",
  10672=>"010011110",
  10673=>"100110010",
  10674=>"011110001",
  10675=>"111001110",
  10676=>"011010000",
  10677=>"111011101",
  10678=>"010100110",
  10679=>"000000000",
  10680=>"010000010",
  10681=>"000010111",
  10682=>"100010110",
  10683=>"111101010",
  10684=>"010000111",
  10685=>"001100011",
  10686=>"101011011",
  10687=>"111011111",
  10688=>"100111000",
  10689=>"111010010",
  10690=>"111110011",
  10691=>"111101111",
  10692=>"101101111",
  10693=>"010001010",
  10694=>"001001110",
  10695=>"101110110",
  10696=>"010011011",
  10697=>"001110000",
  10698=>"111101101",
  10699=>"011110101",
  10700=>"110110110",
  10701=>"010111010",
  10702=>"100011101",
  10703=>"100111001",
  10704=>"110100101",
  10705=>"100100110",
  10706=>"100011111",
  10707=>"000111000",
  10708=>"010001000",
  10709=>"111010001",
  10710=>"100011010",
  10711=>"000110011",
  10712=>"001011000",
  10713=>"010011011",
  10714=>"111001101",
  10715=>"111110100",
  10716=>"110000100",
  10717=>"101000000",
  10718=>"100001111",
  10719=>"000101001",
  10720=>"010111101",
  10721=>"000100010",
  10722=>"010010000",
  10723=>"011100000",
  10724=>"100010011",
  10725=>"010101101",
  10726=>"001001101",
  10727=>"011000000",
  10728=>"111001001",
  10729=>"101000000",
  10730=>"111100100",
  10731=>"000000111",
  10732=>"001001110",
  10733=>"111001011",
  10734=>"011001100",
  10735=>"011000000",
  10736=>"001101101",
  10737=>"011010110",
  10738=>"111010000",
  10739=>"011101111",
  10740=>"010111101",
  10741=>"001100110",
  10742=>"110000001",
  10743=>"010100011",
  10744=>"000111011",
  10745=>"100100010",
  10746=>"010000100",
  10747=>"100011101",
  10748=>"000011111",
  10749=>"101010111",
  10750=>"001111000",
  10751=>"011100001",
  10752=>"110111001",
  10753=>"111010111",
  10754=>"110010100",
  10755=>"111111010",
  10756=>"010010100",
  10757=>"101100000",
  10758=>"001001110",
  10759=>"101111010",
  10760=>"011011101",
  10761=>"000110000",
  10762=>"110000101",
  10763=>"101111010",
  10764=>"111111111",
  10765=>"011011110",
  10766=>"100110001",
  10767=>"010010001",
  10768=>"000100011",
  10769=>"101100001",
  10770=>"001010001",
  10771=>"011111000",
  10772=>"001100001",
  10773=>"111101110",
  10774=>"011000111",
  10775=>"001011001",
  10776=>"110000000",
  10777=>"110010110",
  10778=>"100100100",
  10779=>"011000000",
  10780=>"000110001",
  10781=>"011110011",
  10782=>"100001101",
  10783=>"111100010",
  10784=>"000011011",
  10785=>"010100100",
  10786=>"001000100",
  10787=>"010010000",
  10788=>"001111100",
  10789=>"111001100",
  10790=>"101011011",
  10791=>"101110100",
  10792=>"000100011",
  10793=>"100000001",
  10794=>"100000001",
  10795=>"010101010",
  10796=>"101000000",
  10797=>"000100010",
  10798=>"111111111",
  10799=>"111111111",
  10800=>"100001110",
  10801=>"001111011",
  10802=>"110110101",
  10803=>"010111111",
  10804=>"101001000",
  10805=>"000000100",
  10806=>"010100011",
  10807=>"110001010",
  10808=>"110011001",
  10809=>"000101100",
  10810=>"100101110",
  10811=>"111010010",
  10812=>"001101001",
  10813=>"011011001",
  10814=>"000000001",
  10815=>"111111011",
  10816=>"110111101",
  10817=>"010111101",
  10818=>"011110101",
  10819=>"011010011",
  10820=>"000011000",
  10821=>"101110001",
  10822=>"001101011",
  10823=>"010000000",
  10824=>"100001101",
  10825=>"111111001",
  10826=>"000111111",
  10827=>"011000110",
  10828=>"001110101",
  10829=>"011010001",
  10830=>"010001100",
  10831=>"011001101",
  10832=>"111011111",
  10833=>"100000000",
  10834=>"000000011",
  10835=>"001111010",
  10836=>"011111000",
  10837=>"011001100",
  10838=>"010011110",
  10839=>"100100101",
  10840=>"100101010",
  10841=>"011100100",
  10842=>"000100001",
  10843=>"011001010",
  10844=>"000001110",
  10845=>"000111000",
  10846=>"110011110",
  10847=>"111011010",
  10848=>"100010100",
  10849=>"000001000",
  10850=>"000001001",
  10851=>"000001000",
  10852=>"111100000",
  10853=>"011011001",
  10854=>"001100110",
  10855=>"001101101",
  10856=>"001100110",
  10857=>"001101100",
  10858=>"010000001",
  10859=>"110000000",
  10860=>"110001100",
  10861=>"110101000",
  10862=>"110000101",
  10863=>"110011110",
  10864=>"000010000",
  10865=>"000100010",
  10866=>"100001010",
  10867=>"001010000",
  10868=>"111000100",
  10869=>"010101111",
  10870=>"011100010",
  10871=>"101001001",
  10872=>"100010000",
  10873=>"011101000",
  10874=>"001100110",
  10875=>"010001100",
  10876=>"110010110",
  10877=>"100111000",
  10878=>"100110000",
  10879=>"011000000",
  10880=>"000101011",
  10881=>"000011010",
  10882=>"001001000",
  10883=>"111010100",
  10884=>"000011011",
  10885=>"000110001",
  10886=>"010011100",
  10887=>"011100101",
  10888=>"110010100",
  10889=>"101011000",
  10890=>"001000010",
  10891=>"111100011",
  10892=>"010100001",
  10893=>"010110101",
  10894=>"110110010",
  10895=>"010001000",
  10896=>"001000001",
  10897=>"110001011",
  10898=>"010101100",
  10899=>"111111000",
  10900=>"000010000",
  10901=>"100010010",
  10902=>"101000010",
  10903=>"110001101",
  10904=>"101000000",
  10905=>"000101000",
  10906=>"101100101",
  10907=>"110011111",
  10908=>"001000000",
  10909=>"111100111",
  10910=>"111001010",
  10911=>"110110110",
  10912=>"101000110",
  10913=>"000101110",
  10914=>"011100100",
  10915=>"011110010",
  10916=>"111111011",
  10917=>"100000000",
  10918=>"001101110",
  10919=>"000110010",
  10920=>"111011110",
  10921=>"000110010",
  10922=>"000100000",
  10923=>"001111101",
  10924=>"000100100",
  10925=>"111011010",
  10926=>"100010110",
  10927=>"001100100",
  10928=>"000000101",
  10929=>"010111000",
  10930=>"001110001",
  10931=>"001100000",
  10932=>"001011111",
  10933=>"011001000",
  10934=>"001110110",
  10935=>"101000100",
  10936=>"101001001",
  10937=>"101010010",
  10938=>"001101100",
  10939=>"111111111",
  10940=>"001110101",
  10941=>"001001001",
  10942=>"101011100",
  10943=>"010000000",
  10944=>"011010101",
  10945=>"000001100",
  10946=>"111000101",
  10947=>"110010100",
  10948=>"011111111",
  10949=>"101100001",
  10950=>"000100000",
  10951=>"101001101",
  10952=>"010001000",
  10953=>"101001111",
  10954=>"100010111",
  10955=>"001100000",
  10956=>"101101000",
  10957=>"001101110",
  10958=>"010111010",
  10959=>"100111110",
  10960=>"000000011",
  10961=>"011110100",
  10962=>"101110110",
  10963=>"111001110",
  10964=>"011110001",
  10965=>"101110100",
  10966=>"111110111",
  10967=>"010010010",
  10968=>"000001001",
  10969=>"000000100",
  10970=>"001111011",
  10971=>"011101000",
  10972=>"000011011",
  10973=>"110110011",
  10974=>"011100101",
  10975=>"001000000",
  10976=>"010001010",
  10977=>"101001100",
  10978=>"010111000",
  10979=>"101001000",
  10980=>"011111110",
  10981=>"001010110",
  10982=>"001111101",
  10983=>"001000000",
  10984=>"111110010",
  10985=>"101111101",
  10986=>"000111100",
  10987=>"011100000",
  10988=>"111100011",
  10989=>"100110110",
  10990=>"000110001",
  10991=>"111000101",
  10992=>"001111100",
  10993=>"011010010",
  10994=>"100010010",
  10995=>"011111010",
  10996=>"100010001",
  10997=>"011111010",
  10998=>"110100010",
  10999=>"011111100",
  11000=>"110110011",
  11001=>"110000100",
  11002=>"110010100",
  11003=>"000111011",
  11004=>"101010101",
  11005=>"011110110",
  11006=>"010100100",
  11007=>"101100011",
  11008=>"010111100",
  11009=>"101100010",
  11010=>"010101100",
  11011=>"101100000",
  11012=>"101001100",
  11013=>"000101100",
  11014=>"111111110",
  11015=>"110011011",
  11016=>"011010100",
  11017=>"100000100",
  11018=>"110110101",
  11019=>"000100100",
  11020=>"001111111",
  11021=>"000010111",
  11022=>"101101000",
  11023=>"111011000",
  11024=>"110011111",
  11025=>"100010000",
  11026=>"010010111",
  11027=>"010100110",
  11028=>"101001010",
  11029=>"011001100",
  11030=>"100110101",
  11031=>"100000000",
  11032=>"011100000",
  11033=>"001101010",
  11034=>"011111010",
  11035=>"100100010",
  11036=>"001010110",
  11037=>"111111110",
  11038=>"011100101",
  11039=>"011011001",
  11040=>"000010000",
  11041=>"101101100",
  11042=>"001101011",
  11043=>"011101000",
  11044=>"000011110",
  11045=>"100111101",
  11046=>"101101001",
  11047=>"001110010",
  11048=>"011101010",
  11049=>"010010001",
  11050=>"111011001",
  11051=>"110000011",
  11052=>"110000110",
  11053=>"000110001",
  11054=>"011111010",
  11055=>"111111000",
  11056=>"010010110",
  11057=>"100100010",
  11058=>"100100111",
  11059=>"011101100",
  11060=>"000001111",
  11061=>"011111101",
  11062=>"101110110",
  11063=>"001111111",
  11064=>"111110001",
  11065=>"000000110",
  11066=>"001001100",
  11067=>"111111001",
  11068=>"101001011",
  11069=>"011101010",
  11070=>"000000101",
  11071=>"101001010",
  11072=>"000100011",
  11073=>"001000000",
  11074=>"001100010",
  11075=>"000101000",
  11076=>"110110000",
  11077=>"011110011",
  11078=>"001011011",
  11079=>"110011001",
  11080=>"101010100",
  11081=>"000000110",
  11082=>"110011010",
  11083=>"001111110",
  11084=>"010000001",
  11085=>"111100010",
  11086=>"100000100",
  11087=>"110110000",
  11088=>"110100000",
  11089=>"000100111",
  11090=>"001000010",
  11091=>"101110000",
  11092=>"000011011",
  11093=>"110011101",
  11094=>"011001000",
  11095=>"010001111",
  11096=>"010001111",
  11097=>"111011000",
  11098=>"001000111",
  11099=>"110000111",
  11100=>"001110001",
  11101=>"000001010",
  11102=>"111101011",
  11103=>"010101110",
  11104=>"100110001",
  11105=>"100001111",
  11106=>"011000001",
  11107=>"101100101",
  11108=>"001100000",
  11109=>"000011010",
  11110=>"000010110",
  11111=>"111011000",
  11112=>"111111001",
  11113=>"100011000",
  11114=>"101000110",
  11115=>"000110110",
  11116=>"110010110",
  11117=>"101000000",
  11118=>"110101111",
  11119=>"111100110",
  11120=>"010011010",
  11121=>"001001100",
  11122=>"110101110",
  11123=>"000110001",
  11124=>"001001111",
  11125=>"000011000",
  11126=>"100011000",
  11127=>"010100000",
  11128=>"001011001",
  11129=>"011001000",
  11130=>"101110000",
  11131=>"101111111",
  11132=>"001000100",
  11133=>"101000101",
  11134=>"000010000",
  11135=>"110000100",
  11136=>"101001100",
  11137=>"000100111",
  11138=>"010011000",
  11139=>"001111110",
  11140=>"000000011",
  11141=>"110110100",
  11142=>"100110110",
  11143=>"000101010",
  11144=>"010001101",
  11145=>"110100001",
  11146=>"111101000",
  11147=>"000011010",
  11148=>"000001110",
  11149=>"101111000",
  11150=>"000001010",
  11151=>"001010010",
  11152=>"110111100",
  11153=>"001101011",
  11154=>"000100000",
  11155=>"100001100",
  11156=>"111001111",
  11157=>"010001101",
  11158=>"011111111",
  11159=>"010111011",
  11160=>"011001110",
  11161=>"011100001",
  11162=>"100110111",
  11163=>"001101001",
  11164=>"000000000",
  11165=>"011111000",
  11166=>"000110100",
  11167=>"011001011",
  11168=>"100111100",
  11169=>"111010010",
  11170=>"000010111",
  11171=>"000010011",
  11172=>"000101100",
  11173=>"111110010",
  11174=>"111011010",
  11175=>"100111101",
  11176=>"110010111",
  11177=>"010101000",
  11178=>"010111000",
  11179=>"101111010",
  11180=>"011101010",
  11181=>"111110001",
  11182=>"100000111",
  11183=>"001100110",
  11184=>"000101001",
  11185=>"111000000",
  11186=>"010000101",
  11187=>"011101000",
  11188=>"101000000",
  11189=>"000110011",
  11190=>"110011100",
  11191=>"110000110",
  11192=>"110001010",
  11193=>"010001011",
  11194=>"000111110",
  11195=>"011111001",
  11196=>"111101001",
  11197=>"100100110",
  11198=>"000011011",
  11199=>"101001100",
  11200=>"001101111",
  11201=>"000001001",
  11202=>"000101111",
  11203=>"001110010",
  11204=>"111111101",
  11205=>"001010100",
  11206=>"101000010",
  11207=>"101100110",
  11208=>"111111101",
  11209=>"010000000",
  11210=>"100101101",
  11211=>"111011111",
  11212=>"100010011",
  11213=>"011000000",
  11214=>"110110110",
  11215=>"101111111",
  11216=>"110000001",
  11217=>"000000111",
  11218=>"010001000",
  11219=>"000100111",
  11220=>"011101111",
  11221=>"101111010",
  11222=>"011111100",
  11223=>"001001101",
  11224=>"100100111",
  11225=>"101001111",
  11226=>"001010001",
  11227=>"000111001",
  11228=>"011011111",
  11229=>"101010100",
  11230=>"000110110",
  11231=>"010000100",
  11232=>"100111111",
  11233=>"111011111",
  11234=>"010000110",
  11235=>"000100010",
  11236=>"100000000",
  11237=>"001000011",
  11238=>"110101111",
  11239=>"010111101",
  11240=>"000010111",
  11241=>"000000111",
  11242=>"010100011",
  11243=>"111010101",
  11244=>"101110010",
  11245=>"100000101",
  11246=>"000100110",
  11247=>"000000000",
  11248=>"011100111",
  11249=>"010111011",
  11250=>"011100111",
  11251=>"000010110",
  11252=>"010010011",
  11253=>"011011001",
  11254=>"100001111",
  11255=>"010011001",
  11256=>"000000000",
  11257=>"001111001",
  11258=>"110010110",
  11259=>"100011000",
  11260=>"001101101",
  11261=>"001001110",
  11262=>"011000110",
  11263=>"001001010",
  11264=>"110000000",
  11265=>"011011001",
  11266=>"111100111",
  11267=>"000000110",
  11268=>"001000011",
  11269=>"101101001",
  11270=>"110000111",
  11271=>"111111010",
  11272=>"001000001",
  11273=>"111101000",
  11274=>"110001100",
  11275=>"110100101",
  11276=>"111110110",
  11277=>"111110101",
  11278=>"000011010",
  11279=>"111110001",
  11280=>"010100010",
  11281=>"100110111",
  11282=>"000100011",
  11283=>"101110000",
  11284=>"111111100",
  11285=>"110111011",
  11286=>"001011110",
  11287=>"111000001",
  11288=>"111001010",
  11289=>"100100000",
  11290=>"001111100",
  11291=>"011000001",
  11292=>"101001010",
  11293=>"001010011",
  11294=>"110110011",
  11295=>"010001111",
  11296=>"001000011",
  11297=>"000011000",
  11298=>"100010010",
  11299=>"110100111",
  11300=>"110111000",
  11301=>"001111101",
  11302=>"101101101",
  11303=>"010111111",
  11304=>"010110010",
  11305=>"100110001",
  11306=>"011101111",
  11307=>"100111111",
  11308=>"010010011",
  11309=>"101001011",
  11310=>"111111111",
  11311=>"000000100",
  11312=>"111000000",
  11313=>"100000011",
  11314=>"100011110",
  11315=>"110001011",
  11316=>"010110001",
  11317=>"101001101",
  11318=>"111110101",
  11319=>"100110110",
  11320=>"010010111",
  11321=>"110001011",
  11322=>"010010101",
  11323=>"101010110",
  11324=>"010100111",
  11325=>"111100100",
  11326=>"110100010",
  11327=>"010111000",
  11328=>"001011100",
  11329=>"000000110",
  11330=>"110101110",
  11331=>"000101100",
  11332=>"101110010",
  11333=>"011001011",
  11334=>"011000111",
  11335=>"000011110",
  11336=>"110101110",
  11337=>"100101010",
  11338=>"011001101",
  11339=>"000101100",
  11340=>"100010001",
  11341=>"111000000",
  11342=>"101010000",
  11343=>"001011010",
  11344=>"101110000",
  11345=>"110010010",
  11346=>"000100010",
  11347=>"100000010",
  11348=>"010100110",
  11349=>"011110100",
  11350=>"000000000",
  11351=>"000011100",
  11352=>"011010001",
  11353=>"100101111",
  11354=>"010000000",
  11355=>"011111000",
  11356=>"101111101",
  11357=>"010010001",
  11358=>"111101011",
  11359=>"101000111",
  11360=>"110000101",
  11361=>"000110110",
  11362=>"000101101",
  11363=>"111111101",
  11364=>"110100101",
  11365=>"010000110",
  11366=>"000000011",
  11367=>"010010001",
  11368=>"101000010",
  11369=>"000110010",
  11370=>"000001100",
  11371=>"110000000",
  11372=>"100111100",
  11373=>"010100001",
  11374=>"111000011",
  11375=>"101000111",
  11376=>"011111001",
  11377=>"111011010",
  11378=>"111000111",
  11379=>"000101111",
  11380=>"101111100",
  11381=>"101000010",
  11382=>"011110011",
  11383=>"101000010",
  11384=>"110100100",
  11385=>"001100101",
  11386=>"111001001",
  11387=>"101001101",
  11388=>"100001110",
  11389=>"001000100",
  11390=>"110011111",
  11391=>"101001100",
  11392=>"001000110",
  11393=>"101011000",
  11394=>"010100111",
  11395=>"000100101",
  11396=>"110000010",
  11397=>"100000001",
  11398=>"110011101",
  11399=>"110011011",
  11400=>"010011111",
  11401=>"011101010",
  11402=>"001010011",
  11403=>"011101010",
  11404=>"100010001",
  11405=>"010100000",
  11406=>"011010100",
  11407=>"011110000",
  11408=>"011001111",
  11409=>"010100111",
  11410=>"110100011",
  11411=>"010001001",
  11412=>"011000010",
  11413=>"001011101",
  11414=>"010011011",
  11415=>"010011100",
  11416=>"110111000",
  11417=>"100001001",
  11418=>"010010010",
  11419=>"111101111",
  11420=>"001010100",
  11421=>"001000000",
  11422=>"110100000",
  11423=>"110010000",
  11424=>"110110001",
  11425=>"111001001",
  11426=>"100101111",
  11427=>"011000000",
  11428=>"100001010",
  11429=>"100011011",
  11430=>"000100110",
  11431=>"010100011",
  11432=>"010000010",
  11433=>"100001010",
  11434=>"011101000",
  11435=>"011111010",
  11436=>"010010110",
  11437=>"100011010",
  11438=>"100101100",
  11439=>"101011100",
  11440=>"000110000",
  11441=>"101111010",
  11442=>"110111110",
  11443=>"001011001",
  11444=>"111101101",
  11445=>"001011110",
  11446=>"110000110",
  11447=>"100000101",
  11448=>"111001001",
  11449=>"101100101",
  11450=>"000011101",
  11451=>"111011011",
  11452=>"010111101",
  11453=>"000100000",
  11454=>"100110001",
  11455=>"111111101",
  11456=>"100110101",
  11457=>"101001011",
  11458=>"100011100",
  11459=>"001011100",
  11460=>"110011111",
  11461=>"101111111",
  11462=>"010010100",
  11463=>"011001111",
  11464=>"111001011",
  11465=>"101010110",
  11466=>"101010000",
  11467=>"001011100",
  11468=>"101000101",
  11469=>"000101011",
  11470=>"110100100",
  11471=>"010011000",
  11472=>"111001111",
  11473=>"110000010",
  11474=>"000000110",
  11475=>"110100000",
  11476=>"100011110",
  11477=>"100011101",
  11478=>"010011000",
  11479=>"001101110",
  11480=>"000100101",
  11481=>"001001100",
  11482=>"111101010",
  11483=>"111100111",
  11484=>"010000010",
  11485=>"101010101",
  11486=>"100111111",
  11487=>"011110111",
  11488=>"000010000",
  11489=>"000101001",
  11490=>"111100000",
  11491=>"000000100",
  11492=>"010011111",
  11493=>"111101010",
  11494=>"110110010",
  11495=>"001110100",
  11496=>"100101010",
  11497=>"000100111",
  11498=>"011110001",
  11499=>"100000010",
  11500=>"100100001",
  11501=>"110000011",
  11502=>"000001011",
  11503=>"101010011",
  11504=>"011011000",
  11505=>"101110010",
  11506=>"101101000",
  11507=>"101011010",
  11508=>"000111000",
  11509=>"110100001",
  11510=>"000011000",
  11511=>"000010100",
  11512=>"011010101",
  11513=>"011111000",
  11514=>"111010000",
  11515=>"111001010",
  11516=>"000000110",
  11517=>"010010100",
  11518=>"011100111",
  11519=>"010110001",
  11520=>"010100011",
  11521=>"111011111",
  11522=>"001110100",
  11523=>"000111000",
  11524=>"011000001",
  11525=>"110110101",
  11526=>"101110101",
  11527=>"110001100",
  11528=>"001110100",
  11529=>"000100110",
  11530=>"111110010",
  11531=>"011000000",
  11532=>"100001001",
  11533=>"111111110",
  11534=>"111011101",
  11535=>"001011000",
  11536=>"000100011",
  11537=>"100100100",
  11538=>"000000000",
  11539=>"010001110",
  11540=>"110011010",
  11541=>"100111100",
  11542=>"001001011",
  11543=>"100010110",
  11544=>"101011110",
  11545=>"111111100",
  11546=>"011010101",
  11547=>"001000001",
  11548=>"111000100",
  11549=>"111000010",
  11550=>"011111101",
  11551=>"101100001",
  11552=>"110010101",
  11553=>"000001100",
  11554=>"100011011",
  11555=>"110111111",
  11556=>"110010001",
  11557=>"000010110",
  11558=>"000111001",
  11559=>"111100110",
  11560=>"000001010",
  11561=>"101000100",
  11562=>"010001100",
  11563=>"111110000",
  11564=>"100000110",
  11565=>"001000111",
  11566=>"001000000",
  11567=>"010111110",
  11568=>"111111010",
  11569=>"101001101",
  11570=>"010011000",
  11571=>"101000100",
  11572=>"110000100",
  11573=>"101011000",
  11574=>"001000100",
  11575=>"110010110",
  11576=>"011110101",
  11577=>"111010010",
  11578=>"000000111",
  11579=>"101011000",
  11580=>"001100111",
  11581=>"110111000",
  11582=>"010011000",
  11583=>"000111110",
  11584=>"101000100",
  11585=>"111110111",
  11586=>"101100100",
  11587=>"110100111",
  11588=>"011110101",
  11589=>"101111110",
  11590=>"100001010",
  11591=>"110001010",
  11592=>"011010001",
  11593=>"110001001",
  11594=>"001100111",
  11595=>"010100111",
  11596=>"110111001",
  11597=>"100111001",
  11598=>"000010101",
  11599=>"001111111",
  11600=>"111110101",
  11601=>"000110001",
  11602=>"110110010",
  11603=>"011000011",
  11604=>"001000000",
  11605=>"110111111",
  11606=>"011000011",
  11607=>"110101101",
  11608=>"000101111",
  11609=>"000010000",
  11610=>"011011101",
  11611=>"111000111",
  11612=>"010001011",
  11613=>"110100001",
  11614=>"100000011",
  11615=>"001000000",
  11616=>"010010000",
  11617=>"001011000",
  11618=>"111001000",
  11619=>"011101000",
  11620=>"001110010",
  11621=>"011100000",
  11622=>"001111111",
  11623=>"111101111",
  11624=>"100111001",
  11625=>"010101110",
  11626=>"001010011",
  11627=>"000110101",
  11628=>"100011101",
  11629=>"111111111",
  11630=>"000100110",
  11631=>"001001000",
  11632=>"100011000",
  11633=>"010110110",
  11634=>"010010010",
  11635=>"010110101",
  11636=>"111000000",
  11637=>"101010011",
  11638=>"101000000",
  11639=>"111111110",
  11640=>"001001000",
  11641=>"000000101",
  11642=>"011111100",
  11643=>"100001111",
  11644=>"011110100",
  11645=>"111100011",
  11646=>"110000001",
  11647=>"110001111",
  11648=>"001001001",
  11649=>"100111101",
  11650=>"000111000",
  11651=>"100101110",
  11652=>"010111000",
  11653=>"101101101",
  11654=>"101001010",
  11655=>"001101100",
  11656=>"111001000",
  11657=>"010010000",
  11658=>"000010101",
  11659=>"000111001",
  11660=>"001011010",
  11661=>"111110101",
  11662=>"010010000",
  11663=>"111011110",
  11664=>"110000100",
  11665=>"000000001",
  11666=>"110111010",
  11667=>"010100010",
  11668=>"010111111",
  11669=>"010010001",
  11670=>"100000000",
  11671=>"100111000",
  11672=>"101111010",
  11673=>"000001111",
  11674=>"100111110",
  11675=>"111110110",
  11676=>"010011011",
  11677=>"101100011",
  11678=>"100000011",
  11679=>"100110001",
  11680=>"010111111",
  11681=>"001010100",
  11682=>"101000000",
  11683=>"111000001",
  11684=>"100100010",
  11685=>"010011100",
  11686=>"001010001",
  11687=>"110000101",
  11688=>"100010001",
  11689=>"111010100",
  11690=>"001010011",
  11691=>"101010011",
  11692=>"010001000",
  11693=>"001100111",
  11694=>"000111100",
  11695=>"100111011",
  11696=>"110000001",
  11697=>"011111011",
  11698=>"000101000",
  11699=>"000000011",
  11700=>"011000000",
  11701=>"011110110",
  11702=>"111111010",
  11703=>"001111101",
  11704=>"000111101",
  11705=>"100010110",
  11706=>"110101100",
  11707=>"000001000",
  11708=>"011101101",
  11709=>"001011001",
  11710=>"100100011",
  11711=>"011110001",
  11712=>"001000111",
  11713=>"010000001",
  11714=>"111101110",
  11715=>"101010011",
  11716=>"000011011",
  11717=>"010000110",
  11718=>"000100000",
  11719=>"001100111",
  11720=>"101010011",
  11721=>"000111101",
  11722=>"000011010",
  11723=>"011110111",
  11724=>"100011110",
  11725=>"100111000",
  11726=>"100001100",
  11727=>"011110011",
  11728=>"110011000",
  11729=>"100001001",
  11730=>"001001000",
  11731=>"000000001",
  11732=>"010111011",
  11733=>"001101110",
  11734=>"111011110",
  11735=>"000001010",
  11736=>"101010001",
  11737=>"000001111",
  11738=>"111100001",
  11739=>"101001000",
  11740=>"000111101",
  11741=>"100011011",
  11742=>"001100000",
  11743=>"101000001",
  11744=>"111110100",
  11745=>"111110110",
  11746=>"100000101",
  11747=>"011111110",
  11748=>"000001111",
  11749=>"100000000",
  11750=>"101101000",
  11751=>"010011011",
  11752=>"111111111",
  11753=>"101001110",
  11754=>"100100000",
  11755=>"001011111",
  11756=>"111000000",
  11757=>"000010000",
  11758=>"000010110",
  11759=>"011000100",
  11760=>"000011000",
  11761=>"111100011",
  11762=>"001000010",
  11763=>"000100010",
  11764=>"110001101",
  11765=>"001011110",
  11766=>"001110001",
  11767=>"101100010",
  11768=>"000011010",
  11769=>"010000011",
  11770=>"000011010",
  11771=>"000101001",
  11772=>"000100010",
  11773=>"110100100",
  11774=>"001110100",
  11775=>"001011111",
  11776=>"111000010",
  11777=>"101110111",
  11778=>"111010110",
  11779=>"000000100",
  11780=>"011100010",
  11781=>"111000001",
  11782=>"111100010",
  11783=>"011010000",
  11784=>"110001010",
  11785=>"011110101",
  11786=>"100001110",
  11787=>"010000111",
  11788=>"111111010",
  11789=>"110000111",
  11790=>"010000011",
  11791=>"111100001",
  11792=>"100111101",
  11793=>"001101001",
  11794=>"101100111",
  11795=>"100011011",
  11796=>"000000100",
  11797=>"011101101",
  11798=>"100000100",
  11799=>"011100101",
  11800=>"100001100",
  11801=>"111010110",
  11802=>"011101110",
  11803=>"111111110",
  11804=>"111100000",
  11805=>"000111101",
  11806=>"011011000",
  11807=>"110110000",
  11808=>"110000000",
  11809=>"010000100",
  11810=>"000000001",
  11811=>"100010011",
  11812=>"111111011",
  11813=>"110101011",
  11814=>"101010111",
  11815=>"000110000",
  11816=>"100011000",
  11817=>"011111111",
  11818=>"100001100",
  11819=>"110010010",
  11820=>"101001001",
  11821=>"010101011",
  11822=>"111110011",
  11823=>"111110000",
  11824=>"001100000",
  11825=>"101001010",
  11826=>"111101011",
  11827=>"111011110",
  11828=>"010010011",
  11829=>"111000111",
  11830=>"101011111",
  11831=>"111110101",
  11832=>"011100011",
  11833=>"000010100",
  11834=>"011100010",
  11835=>"100000000",
  11836=>"001110100",
  11837=>"010000001",
  11838=>"110011100",
  11839=>"100000100",
  11840=>"011000001",
  11841=>"111000001",
  11842=>"100011100",
  11843=>"000100000",
  11844=>"111000100",
  11845=>"111110111",
  11846=>"001001110",
  11847=>"010000101",
  11848=>"001110111",
  11849=>"110100111",
  11850=>"110110010",
  11851=>"111011101",
  11852=>"000110000",
  11853=>"100011101",
  11854=>"111000010",
  11855=>"001100100",
  11856=>"111010111",
  11857=>"110011111",
  11858=>"001101110",
  11859=>"101001100",
  11860=>"101111100",
  11861=>"000110001",
  11862=>"101011000",
  11863=>"000110110",
  11864=>"011101100",
  11865=>"001101000",
  11866=>"010000111",
  11867=>"011111000",
  11868=>"100000100",
  11869=>"101000000",
  11870=>"100011000",
  11871=>"010001110",
  11872=>"010110000",
  11873=>"101010101",
  11874=>"111110001",
  11875=>"110110000",
  11876=>"110011101",
  11877=>"111000000",
  11878=>"000000000",
  11879=>"010000100",
  11880=>"001000001",
  11881=>"111010011",
  11882=>"101100101",
  11883=>"000010010",
  11884=>"101010000",
  11885=>"110100000",
  11886=>"011011000",
  11887=>"100000110",
  11888=>"000011100",
  11889=>"110000001",
  11890=>"100001101",
  11891=>"000000101",
  11892=>"110110000",
  11893=>"000001111",
  11894=>"000010111",
  11895=>"110111111",
  11896=>"101010110",
  11897=>"011110010",
  11898=>"011000010",
  11899=>"001101100",
  11900=>"100010111",
  11901=>"011000000",
  11902=>"110110010",
  11903=>"010111011",
  11904=>"010010100",
  11905=>"000110111",
  11906=>"011100101",
  11907=>"001010111",
  11908=>"111100001",
  11909=>"010000101",
  11910=>"011000110",
  11911=>"111001011",
  11912=>"001001111",
  11913=>"100010010",
  11914=>"111100110",
  11915=>"010000000",
  11916=>"000011100",
  11917=>"110000101",
  11918=>"010000011",
  11919=>"011100100",
  11920=>"100110111",
  11921=>"010011010",
  11922=>"101100101",
  11923=>"101111111",
  11924=>"100110110",
  11925=>"110110111",
  11926=>"011100101",
  11927=>"010001100",
  11928=>"100110111",
  11929=>"101000011",
  11930=>"101111101",
  11931=>"000110000",
  11932=>"011110100",
  11933=>"110001011",
  11934=>"100100101",
  11935=>"000100111",
  11936=>"101001011",
  11937=>"010101100",
  11938=>"000010000",
  11939=>"111000000",
  11940=>"111110011",
  11941=>"010000001",
  11942=>"011100101",
  11943=>"101101100",
  11944=>"010110110",
  11945=>"000110000",
  11946=>"000001101",
  11947=>"111110010",
  11948=>"010110000",
  11949=>"001101001",
  11950=>"011001110",
  11951=>"101001000",
  11952=>"001011011",
  11953=>"000110110",
  11954=>"100100100",
  11955=>"011011010",
  11956=>"110010111",
  11957=>"110101010",
  11958=>"001100011",
  11959=>"110010000",
  11960=>"101110010",
  11961=>"010001111",
  11962=>"111111010",
  11963=>"001101001",
  11964=>"101101111",
  11965=>"011000101",
  11966=>"001100100",
  11967=>"111111000",
  11968=>"011100001",
  11969=>"101110010",
  11970=>"001101010",
  11971=>"001011001",
  11972=>"001011000",
  11973=>"010000010",
  11974=>"100000111",
  11975=>"010101000",
  11976=>"111110100",
  11977=>"011111110",
  11978=>"101111001",
  11979=>"101001001",
  11980=>"100011100",
  11981=>"011010110",
  11982=>"110111011",
  11983=>"100101100",
  11984=>"101101111",
  11985=>"100000010",
  11986=>"010010000",
  11987=>"000110011",
  11988=>"100001101",
  11989=>"100011010",
  11990=>"001101010",
  11991=>"010000010",
  11992=>"000001101",
  11993=>"100111111",
  11994=>"111000111",
  11995=>"110011000",
  11996=>"010111011",
  11997=>"000011100",
  11998=>"011111010",
  11999=>"100101000",
  12000=>"001101011",
  12001=>"001001000",
  12002=>"011001000",
  12003=>"110011111",
  12004=>"010011000",
  12005=>"111110101",
  12006=>"000101001",
  12007=>"100110001",
  12008=>"000111011",
  12009=>"100110110",
  12010=>"001101011",
  12011=>"001011101",
  12012=>"010010000",
  12013=>"010110010",
  12014=>"000001100",
  12015=>"110101110",
  12016=>"010101101",
  12017=>"011101101",
  12018=>"100100111",
  12019=>"000100010",
  12020=>"111101111",
  12021=>"011000110",
  12022=>"001101110",
  12023=>"010111110",
  12024=>"101111000",
  12025=>"110111111",
  12026=>"011111101",
  12027=>"110110000",
  12028=>"010000010",
  12029=>"101100011",
  12030=>"001011100",
  12031=>"110100010",
  12032=>"011010011",
  12033=>"000101111",
  12034=>"000010100",
  12035=>"101111101",
  12036=>"100111101",
  12037=>"010000000",
  12038=>"101100100",
  12039=>"110111100",
  12040=>"000110100",
  12041=>"001000100",
  12042=>"110110001",
  12043=>"110100010",
  12044=>"110101101",
  12045=>"111011001",
  12046=>"000000000",
  12047=>"000110110",
  12048=>"001101100",
  12049=>"000011111",
  12050=>"001110101",
  12051=>"000001001",
  12052=>"010001110",
  12053=>"011011011",
  12054=>"100010001",
  12055=>"100100100",
  12056=>"111001110",
  12057=>"000000100",
  12058=>"000110010",
  12059=>"011111100",
  12060=>"101001000",
  12061=>"010010010",
  12062=>"110001100",
  12063=>"111111100",
  12064=>"010110000",
  12065=>"000100100",
  12066=>"100100110",
  12067=>"110110010",
  12068=>"010101101",
  12069=>"100111011",
  12070=>"101110110",
  12071=>"011001010",
  12072=>"000101001",
  12073=>"000010000",
  12074=>"000100110",
  12075=>"111110010",
  12076=>"100101111",
  12077=>"001010110",
  12078=>"101110000",
  12079=>"111111000",
  12080=>"000111011",
  12081=>"100101111",
  12082=>"100010111",
  12083=>"101100010",
  12084=>"001010000",
  12085=>"010011100",
  12086=>"010010010",
  12087=>"100100110",
  12088=>"001111111",
  12089=>"001000010",
  12090=>"110000111",
  12091=>"000001000",
  12092=>"110101011",
  12093=>"110000010",
  12094=>"101001010",
  12095=>"100000011",
  12096=>"011110001",
  12097=>"110001110",
  12098=>"000110110",
  12099=>"010101001",
  12100=>"010001000",
  12101=>"001101101",
  12102=>"001000000",
  12103=>"011000001",
  12104=>"000011000",
  12105=>"010101101",
  12106=>"100000110",
  12107=>"001001100",
  12108=>"010010110",
  12109=>"000000100",
  12110=>"100100111",
  12111=>"000011101",
  12112=>"111101110",
  12113=>"101001100",
  12114=>"110100010",
  12115=>"010110001",
  12116=>"010011110",
  12117=>"100000010",
  12118=>"101100010",
  12119=>"000100001",
  12120=>"001010010",
  12121=>"110100100",
  12122=>"000001101",
  12123=>"110110011",
  12124=>"100110011",
  12125=>"111111000",
  12126=>"010011010",
  12127=>"001000101",
  12128=>"001110110",
  12129=>"111101011",
  12130=>"000111100",
  12131=>"110111110",
  12132=>"010101000",
  12133=>"011101011",
  12134=>"011000101",
  12135=>"011101111",
  12136=>"101000010",
  12137=>"010101100",
  12138=>"011111001",
  12139=>"000010101",
  12140=>"010010110",
  12141=>"001110110",
  12142=>"001110011",
  12143=>"110010100",
  12144=>"011000000",
  12145=>"101101000",
  12146=>"001001111",
  12147=>"100100111",
  12148=>"010100000",
  12149=>"000111111",
  12150=>"100010100",
  12151=>"100001011",
  12152=>"001111011",
  12153=>"000011001",
  12154=>"110010010",
  12155=>"000000100",
  12156=>"111010110",
  12157=>"101010101",
  12158=>"001111010",
  12159=>"111001110",
  12160=>"010100010",
  12161=>"111110111",
  12162=>"011100100",
  12163=>"000011100",
  12164=>"110001101",
  12165=>"110101001",
  12166=>"011100011",
  12167=>"101000000",
  12168=>"101100101",
  12169=>"101011111",
  12170=>"000001111",
  12171=>"110010001",
  12172=>"101010001",
  12173=>"000111011",
  12174=>"110101100",
  12175=>"001011001",
  12176=>"011010011",
  12177=>"011010000",
  12178=>"111000100",
  12179=>"101110111",
  12180=>"000000000",
  12181=>"100010110",
  12182=>"010001101",
  12183=>"100111000",
  12184=>"111101001",
  12185=>"001100110",
  12186=>"101111111",
  12187=>"100110010",
  12188=>"011001110",
  12189=>"101111001",
  12190=>"010100000",
  12191=>"011111111",
  12192=>"001000010",
  12193=>"000100001",
  12194=>"101110100",
  12195=>"110101001",
  12196=>"001001101",
  12197=>"100000000",
  12198=>"011111001",
  12199=>"111100101",
  12200=>"101010111",
  12201=>"011001100",
  12202=>"000001011",
  12203=>"010000010",
  12204=>"101001010",
  12205=>"010001111",
  12206=>"011000100",
  12207=>"000011000",
  12208=>"011110110",
  12209=>"101010001",
  12210=>"011100010",
  12211=>"110101111",
  12212=>"010101010",
  12213=>"111100111",
  12214=>"100010010",
  12215=>"000101010",
  12216=>"101101011",
  12217=>"001011010",
  12218=>"100101000",
  12219=>"100100111",
  12220=>"000010101",
  12221=>"110001101",
  12222=>"111101101",
  12223=>"011001111",
  12224=>"001100111",
  12225=>"000011111",
  12226=>"011111000",
  12227=>"001100100",
  12228=>"010010011",
  12229=>"110011000",
  12230=>"010010111",
  12231=>"001001100",
  12232=>"101100010",
  12233=>"001001111",
  12234=>"010101110",
  12235=>"011010011",
  12236=>"111101000",
  12237=>"001110011",
  12238=>"101100110",
  12239=>"101101000",
  12240=>"010100001",
  12241=>"100010011",
  12242=>"101000010",
  12243=>"000010100",
  12244=>"100111111",
  12245=>"010011011",
  12246=>"110110011",
  12247=>"011111001",
  12248=>"101010111",
  12249=>"110000010",
  12250=>"111000011",
  12251=>"111110011",
  12252=>"100000101",
  12253=>"011010100",
  12254=>"010110111",
  12255=>"101010100",
  12256=>"111111110",
  12257=>"011110001",
  12258=>"001001001",
  12259=>"001100011",
  12260=>"010011110",
  12261=>"011100110",
  12262=>"011011110",
  12263=>"111101100",
  12264=>"000100101",
  12265=>"110001111",
  12266=>"100100010",
  12267=>"111000001",
  12268=>"100011010",
  12269=>"011000010",
  12270=>"110001010",
  12271=>"010010010",
  12272=>"100000000",
  12273=>"010011111",
  12274=>"010100001",
  12275=>"111101010",
  12276=>"011111100",
  12277=>"010000000",
  12278=>"001010001",
  12279=>"000111101",
  12280=>"001111010",
  12281=>"110010101",
  12282=>"000111100",
  12283=>"111101100",
  12284=>"011100100",
  12285=>"000000011",
  12286=>"010010110",
  12287=>"000011000",
  12288=>"010110011",
  12289=>"001100010",
  12290=>"001001110",
  12291=>"101100010",
  12292=>"110000101",
  12293=>"000001010",
  12294=>"110010111",
  12295=>"011000000",
  12296=>"000101000",
  12297=>"100101111",
  12298=>"011110001",
  12299=>"110010110",
  12300=>"011000001",
  12301=>"000110101",
  12302=>"101111100",
  12303=>"001111111",
  12304=>"100101001",
  12305=>"010110110",
  12306=>"111110111",
  12307=>"111111000",
  12308=>"100110101",
  12309=>"001100000",
  12310=>"011111000",
  12311=>"001000101",
  12312=>"110100011",
  12313=>"011010011",
  12314=>"100101001",
  12315=>"100001110",
  12316=>"011011111",
  12317=>"000000011",
  12318=>"100100100",
  12319=>"101101100",
  12320=>"101001111",
  12321=>"100001011",
  12322=>"110000000",
  12323=>"110000101",
  12324=>"000101111",
  12325=>"101000000",
  12326=>"000000100",
  12327=>"000000101",
  12328=>"000001011",
  12329=>"010101111",
  12330=>"011001100",
  12331=>"100110101",
  12332=>"100000011",
  12333=>"010110100",
  12334=>"011010111",
  12335=>"101011100",
  12336=>"010101010",
  12337=>"001111101",
  12338=>"110100110",
  12339=>"101000001",
  12340=>"100011001",
  12341=>"111010011",
  12342=>"100001100",
  12343=>"001101011",
  12344=>"011101011",
  12345=>"110001010",
  12346=>"111001101",
  12347=>"111010001",
  12348=>"001000001",
  12349=>"001000111",
  12350=>"101100001",
  12351=>"110001000",
  12352=>"011010100",
  12353=>"000000010",
  12354=>"101011000",
  12355=>"100010010",
  12356=>"001111100",
  12357=>"011100000",
  12358=>"010011100",
  12359=>"100100011",
  12360=>"010010001",
  12361=>"000110001",
  12362=>"101000010",
  12363=>"100111111",
  12364=>"010100111",
  12365=>"110111111",
  12366=>"101011100",
  12367=>"011110111",
  12368=>"111100100",
  12369=>"010100001",
  12370=>"101001100",
  12371=>"011100001",
  12372=>"110101010",
  12373=>"101001000",
  12374=>"111001011",
  12375=>"001011011",
  12376=>"001000010",
  12377=>"011110010",
  12378=>"100100110",
  12379=>"001001010",
  12380=>"101101010",
  12381=>"010110101",
  12382=>"011001010",
  12383=>"001111000",
  12384=>"011111000",
  12385=>"101001000",
  12386=>"110110101",
  12387=>"000111100",
  12388=>"000110101",
  12389=>"001100100",
  12390=>"110101010",
  12391=>"101010010",
  12392=>"101010000",
  12393=>"101100111",
  12394=>"110011000",
  12395=>"011100110",
  12396=>"010101011",
  12397=>"011101110",
  12398=>"010101110",
  12399=>"100010100",
  12400=>"100000111",
  12401=>"000111011",
  12402=>"000001100",
  12403=>"100011010",
  12404=>"011101100",
  12405=>"110010101",
  12406=>"000110001",
  12407=>"111111111",
  12408=>"010101111",
  12409=>"000010100",
  12410=>"000001101",
  12411=>"010001101",
  12412=>"100111111",
  12413=>"010010111",
  12414=>"111001110",
  12415=>"000010101",
  12416=>"101000010",
  12417=>"100111000",
  12418=>"010001100",
  12419=>"001111100",
  12420=>"001100101",
  12421=>"100011100",
  12422=>"011111110",
  12423=>"010111010",
  12424=>"001000001",
  12425=>"111100010",
  12426=>"100011111",
  12427=>"111100101",
  12428=>"110110100",
  12429=>"000100100",
  12430=>"001010010",
  12431=>"101101100",
  12432=>"000011101",
  12433=>"011010100",
  12434=>"011110111",
  12435=>"011111000",
  12436=>"110010001",
  12437=>"000110101",
  12438=>"110111101",
  12439=>"001111110",
  12440=>"110000110",
  12441=>"100100001",
  12442=>"011101111",
  12443=>"000100111",
  12444=>"011010111",
  12445=>"011100110",
  12446=>"011010000",
  12447=>"000110100",
  12448=>"111000110",
  12449=>"111010001",
  12450=>"010110010",
  12451=>"000010010",
  12452=>"100001111",
  12453=>"111110010",
  12454=>"111111101",
  12455=>"000100110",
  12456=>"010111100",
  12457=>"001010100",
  12458=>"101100011",
  12459=>"100011010",
  12460=>"101001000",
  12461=>"111110101",
  12462=>"100001100",
  12463=>"000110111",
  12464=>"100010001",
  12465=>"011000110",
  12466=>"000110100",
  12467=>"000110100",
  12468=>"000000010",
  12469=>"001010000",
  12470=>"000000110",
  12471=>"010001101",
  12472=>"000011010",
  12473=>"000110111",
  12474=>"011010100",
  12475=>"011111111",
  12476=>"011010101",
  12477=>"011100110",
  12478=>"110011001",
  12479=>"111111100",
  12480=>"100010110",
  12481=>"001000101",
  12482=>"001001001",
  12483=>"011010011",
  12484=>"110000100",
  12485=>"001110111",
  12486=>"001111110",
  12487=>"100101101",
  12488=>"010100111",
  12489=>"100111110",
  12490=>"000001001",
  12491=>"001001001",
  12492=>"011110101",
  12493=>"010111000",
  12494=>"000111100",
  12495=>"010011111",
  12496=>"101111000",
  12497=>"011010000",
  12498=>"100101011",
  12499=>"010110101",
  12500=>"010101010",
  12501=>"111101000",
  12502=>"110111100",
  12503=>"011010001",
  12504=>"010000000",
  12505=>"000001110",
  12506=>"100110011",
  12507=>"010110000",
  12508=>"010001011",
  12509=>"100110000",
  12510=>"010000000",
  12511=>"111111010",
  12512=>"100010000",
  12513=>"011010111",
  12514=>"101101100",
  12515=>"000100100",
  12516=>"001000101",
  12517=>"101011010",
  12518=>"100001011",
  12519=>"111001111",
  12520=>"110100000",
  12521=>"101011011",
  12522=>"001100101",
  12523=>"010110110",
  12524=>"010011110",
  12525=>"000000101",
  12526=>"001011001",
  12527=>"111110000",
  12528=>"111100010",
  12529=>"100010011",
  12530=>"000010000",
  12531=>"100100100",
  12532=>"101010101",
  12533=>"111111111",
  12534=>"000001101",
  12535=>"000000100",
  12536=>"010000111",
  12537=>"101000010",
  12538=>"101111111",
  12539=>"000011100",
  12540=>"110100001",
  12541=>"000100110",
  12542=>"001000110",
  12543=>"110001010",
  12544=>"100011110",
  12545=>"001010111",
  12546=>"001010110",
  12547=>"100111011",
  12548=>"001011111",
  12549=>"000110110",
  12550=>"100010110",
  12551=>"111100001",
  12552=>"000101000",
  12553=>"010111110",
  12554=>"000011010",
  12555=>"100000101",
  12556=>"001110100",
  12557=>"001001001",
  12558=>"101001101",
  12559=>"101110001",
  12560=>"111100111",
  12561=>"101110000",
  12562=>"111111101",
  12563=>"110111100",
  12564=>"101111000",
  12565=>"011000000",
  12566=>"001100111",
  12567=>"100110101",
  12568=>"000111000",
  12569=>"100001001",
  12570=>"010010000",
  12571=>"010101010",
  12572=>"100101000",
  12573=>"100000110",
  12574=>"000000000",
  12575=>"000101011",
  12576=>"000101111",
  12577=>"111111111",
  12578=>"000100001",
  12579=>"100111100",
  12580=>"101000110",
  12581=>"011011111",
  12582=>"010010101",
  12583=>"101111100",
  12584=>"010001111",
  12585=>"000001011",
  12586=>"011100101",
  12587=>"110111010",
  12588=>"111001011",
  12589=>"011100101",
  12590=>"111000000",
  12591=>"111101011",
  12592=>"001011101",
  12593=>"111101000",
  12594=>"100101110",
  12595=>"101000001",
  12596=>"101101010",
  12597=>"000010110",
  12598=>"110101110",
  12599=>"101011000",
  12600=>"000110010",
  12601=>"010100101",
  12602=>"111010000",
  12603=>"100010001",
  12604=>"001110000",
  12605=>"101111000",
  12606=>"100000101",
  12607=>"110100101",
  12608=>"110111110",
  12609=>"111101001",
  12610=>"010001100",
  12611=>"110110001",
  12612=>"101010100",
  12613=>"110010000",
  12614=>"011011100",
  12615=>"100101110",
  12616=>"101011100",
  12617=>"011011100",
  12618=>"100101010",
  12619=>"010010011",
  12620=>"110101001",
  12621=>"100110010",
  12622=>"000000101",
  12623=>"111110000",
  12624=>"100111110",
  12625=>"000000101",
  12626=>"001001100",
  12627=>"000100010",
  12628=>"000000000",
  12629=>"011000001",
  12630=>"111001011",
  12631=>"100001000",
  12632=>"010110010",
  12633=>"000110000",
  12634=>"000100000",
  12635=>"100011001",
  12636=>"110111011",
  12637=>"011111111",
  12638=>"010111110",
  12639=>"111001000",
  12640=>"001110000",
  12641=>"110101110",
  12642=>"001011010",
  12643=>"101101011",
  12644=>"101011011",
  12645=>"000111000",
  12646=>"000011010",
  12647=>"010110010",
  12648=>"101100010",
  12649=>"100001010",
  12650=>"011011010",
  12651=>"010010011",
  12652=>"000001100",
  12653=>"111011001",
  12654=>"100010000",
  12655=>"001010101",
  12656=>"000011001",
  12657=>"001011111",
  12658=>"001011011",
  12659=>"101110100",
  12660=>"110010101",
  12661=>"111010101",
  12662=>"101001101",
  12663=>"001010010",
  12664=>"011010010",
  12665=>"011110110",
  12666=>"111010011",
  12667=>"101000101",
  12668=>"101010100",
  12669=>"101101111",
  12670=>"111111010",
  12671=>"101101001",
  12672=>"100100101",
  12673=>"010010100",
  12674=>"101110000",
  12675=>"111110110",
  12676=>"010100001",
  12677=>"100111100",
  12678=>"101001011",
  12679=>"010111100",
  12680=>"010010101",
  12681=>"010010010",
  12682=>"000001000",
  12683=>"001000101",
  12684=>"010110001",
  12685=>"111101000",
  12686=>"110000100",
  12687=>"001000000",
  12688=>"001010101",
  12689=>"100011011",
  12690=>"110010000",
  12691=>"100111111",
  12692=>"100101100",
  12693=>"010011111",
  12694=>"111000001",
  12695=>"110111000",
  12696=>"000110101",
  12697=>"110000001",
  12698=>"111011001",
  12699=>"000000111",
  12700=>"111001111",
  12701=>"100000001",
  12702=>"001111110",
  12703=>"001000001",
  12704=>"101100110",
  12705=>"010111110",
  12706=>"000001010",
  12707=>"111101010",
  12708=>"110010010",
  12709=>"000000001",
  12710=>"110011100",
  12711=>"110111011",
  12712=>"000011010",
  12713=>"000101000",
  12714=>"001011010",
  12715=>"010101010",
  12716=>"110110110",
  12717=>"111111101",
  12718=>"000100001",
  12719=>"100011100",
  12720=>"100011111",
  12721=>"111111110",
  12722=>"010110000",
  12723=>"110011111",
  12724=>"110000111",
  12725=>"111111010",
  12726=>"111110001",
  12727=>"111010110",
  12728=>"100101001",
  12729=>"011100010",
  12730=>"011101010",
  12731=>"011100011",
  12732=>"100101011",
  12733=>"100001110",
  12734=>"111100101",
  12735=>"001101110",
  12736=>"100010001",
  12737=>"001011011",
  12738=>"000010110",
  12739=>"110110011",
  12740=>"000000110",
  12741=>"011000001",
  12742=>"110101100",
  12743=>"100110001",
  12744=>"010100010",
  12745=>"010001000",
  12746=>"100001001",
  12747=>"001110001",
  12748=>"010111100",
  12749=>"001111110",
  12750=>"000000101",
  12751=>"010110000",
  12752=>"010101011",
  12753=>"000001000",
  12754=>"001000010",
  12755=>"110010101",
  12756=>"100001110",
  12757=>"010101000",
  12758=>"001010000",
  12759=>"000111010",
  12760=>"001010100",
  12761=>"110100110",
  12762=>"010001100",
  12763=>"100100011",
  12764=>"100011001",
  12765=>"011100111",
  12766=>"000111111",
  12767=>"010111011",
  12768=>"010100010",
  12769=>"111000111",
  12770=>"000000001",
  12771=>"110110001",
  12772=>"010101101",
  12773=>"111101000",
  12774=>"001000000",
  12775=>"101010001",
  12776=>"010110100",
  12777=>"100101100",
  12778=>"010000100",
  12779=>"010000001",
  12780=>"110100101",
  12781=>"110001011",
  12782=>"001011100",
  12783=>"000011011",
  12784=>"010100100",
  12785=>"111010100",
  12786=>"110101001",
  12787=>"000001001",
  12788=>"000011011",
  12789=>"000100001",
  12790=>"111010111",
  12791=>"011111000",
  12792=>"110101011",
  12793=>"101111000",
  12794=>"010010110",
  12795=>"110111000",
  12796=>"111010000",
  12797=>"010000100",
  12798=>"111101000",
  12799=>"001000001",
  12800=>"010011101",
  12801=>"101111110",
  12802=>"010111011",
  12803=>"100100101",
  12804=>"010010010",
  12805=>"001000110",
  12806=>"000000010",
  12807=>"000010100",
  12808=>"000011100",
  12809=>"010010001",
  12810=>"100111001",
  12811=>"100101000",
  12812=>"000000010",
  12813=>"110001100",
  12814=>"001001001",
  12815=>"010010001",
  12816=>"010100111",
  12817=>"001110100",
  12818=>"100001111",
  12819=>"001100001",
  12820=>"110001101",
  12821=>"001010011",
  12822=>"011111010",
  12823=>"110010111",
  12824=>"110110011",
  12825=>"001000110",
  12826=>"001011100",
  12827=>"101110110",
  12828=>"111101000",
  12829=>"101010000",
  12830=>"100001110",
  12831=>"001000011",
  12832=>"100000101",
  12833=>"000000100",
  12834=>"011100110",
  12835=>"000100100",
  12836=>"111111111",
  12837=>"011101100",
  12838=>"111010001",
  12839=>"100001010",
  12840=>"010100110",
  12841=>"100101100",
  12842=>"111010110",
  12843=>"010110110",
  12844=>"010010011",
  12845=>"000101100",
  12846=>"100100000",
  12847=>"010100111",
  12848=>"101000000",
  12849=>"001111010",
  12850=>"110100000",
  12851=>"011001010",
  12852=>"000001000",
  12853=>"100110010",
  12854=>"010000011",
  12855=>"110000101",
  12856=>"010000000",
  12857=>"101101110",
  12858=>"111111011",
  12859=>"100100100",
  12860=>"110111101",
  12861=>"010001000",
  12862=>"001111001",
  12863=>"100100001",
  12864=>"110101010",
  12865=>"100001101",
  12866=>"000001101",
  12867=>"111111100",
  12868=>"001100000",
  12869=>"010101010",
  12870=>"100101001",
  12871=>"010000000",
  12872=>"010110101",
  12873=>"111110001",
  12874=>"011110101",
  12875=>"101010101",
  12876=>"111110001",
  12877=>"100001110",
  12878=>"001110111",
  12879=>"101001010",
  12880=>"101110100",
  12881=>"011101001",
  12882=>"111000000",
  12883=>"110001110",
  12884=>"010010011",
  12885=>"001111101",
  12886=>"101000000",
  12887=>"100001011",
  12888=>"111101111",
  12889=>"001001100",
  12890=>"100000001",
  12891=>"001000110",
  12892=>"100111011",
  12893=>"001010011",
  12894=>"100100010",
  12895=>"110001011",
  12896=>"010100100",
  12897=>"011111000",
  12898=>"011100100",
  12899=>"010010010",
  12900=>"111011111",
  12901=>"001100101",
  12902=>"000111011",
  12903=>"000011111",
  12904=>"101001010",
  12905=>"011010011",
  12906=>"011100101",
  12907=>"100101001",
  12908=>"001101111",
  12909=>"010011110",
  12910=>"001101010",
  12911=>"000111001",
  12912=>"000010001",
  12913=>"010001100",
  12914=>"101110001",
  12915=>"011100010",
  12916=>"000000110",
  12917=>"110100111",
  12918=>"110000000",
  12919=>"001111010",
  12920=>"011011000",
  12921=>"111111001",
  12922=>"001110001",
  12923=>"001110110",
  12924=>"001000010",
  12925=>"100100000",
  12926=>"111000011",
  12927=>"101100010",
  12928=>"110010001",
  12929=>"111100110",
  12930=>"110110100",
  12931=>"110111011",
  12932=>"001110010",
  12933=>"100001001",
  12934=>"110011011",
  12935=>"010101010",
  12936=>"100001011",
  12937=>"010100101",
  12938=>"110100010",
  12939=>"101000011",
  12940=>"100100000",
  12941=>"000101011",
  12942=>"011000000",
  12943=>"000011101",
  12944=>"100111101",
  12945=>"001000101",
  12946=>"010101100",
  12947=>"000011100",
  12948=>"010001100",
  12949=>"011110100",
  12950=>"111111011",
  12951=>"001011110",
  12952=>"111100011",
  12953=>"011110000",
  12954=>"000101111",
  12955=>"110100110",
  12956=>"110010100",
  12957=>"001110001",
  12958=>"111010100",
  12959=>"111100010",
  12960=>"000111111",
  12961=>"111111000",
  12962=>"010100011",
  12963=>"110011001",
  12964=>"000010111",
  12965=>"100011100",
  12966=>"010111010",
  12967=>"100010010",
  12968=>"111111110",
  12969=>"001101100",
  12970=>"100011001",
  12971=>"011010001",
  12972=>"110101000",
  12973=>"000100000",
  12974=>"010110101",
  12975=>"101101000",
  12976=>"011000110",
  12977=>"001110010",
  12978=>"000101101",
  12979=>"101011011",
  12980=>"000011010",
  12981=>"011101000",
  12982=>"110111000",
  12983=>"101001111",
  12984=>"100100100",
  12985=>"100110110",
  12986=>"000000001",
  12987=>"001111010",
  12988=>"000100110",
  12989=>"001011011",
  12990=>"110111011",
  12991=>"110101111",
  12992=>"111001100",
  12993=>"010011010",
  12994=>"000111110",
  12995=>"100100000",
  12996=>"101010011",
  12997=>"001101111",
  12998=>"110100011",
  12999=>"010110001",
  13000=>"100110000",
  13001=>"000011001",
  13002=>"011001011",
  13003=>"111000111",
  13004=>"100110111",
  13005=>"001010000",
  13006=>"101011111",
  13007=>"011100010",
  13008=>"010010100",
  13009=>"001011010",
  13010=>"110111110",
  13011=>"110001011",
  13012=>"001100111",
  13013=>"011110110",
  13014=>"001101001",
  13015=>"001111100",
  13016=>"100110011",
  13017=>"110100101",
  13018=>"101010101",
  13019=>"110001000",
  13020=>"001011110",
  13021=>"000000101",
  13022=>"000001000",
  13023=>"011111001",
  13024=>"001000010",
  13025=>"001001000",
  13026=>"010101011",
  13027=>"000000101",
  13028=>"110011110",
  13029=>"111101011",
  13030=>"101101101",
  13031=>"000001001",
  13032=>"000110010",
  13033=>"110110000",
  13034=>"001110010",
  13035=>"000100010",
  13036=>"101010000",
  13037=>"010011010",
  13038=>"000101101",
  13039=>"001101001",
  13040=>"100010101",
  13041=>"101000011",
  13042=>"111110000",
  13043=>"010101111",
  13044=>"101101100",
  13045=>"001000010",
  13046=>"001000011",
  13047=>"011110110",
  13048=>"010111000",
  13049=>"101001110",
  13050=>"010000111",
  13051=>"000010101",
  13052=>"111111110",
  13053=>"000110011",
  13054=>"010110011",
  13055=>"010000111",
  13056=>"111100011",
  13057=>"110100011",
  13058=>"001010111",
  13059=>"010000110",
  13060=>"110110100",
  13061=>"000110011",
  13062=>"101111001",
  13063=>"000010001",
  13064=>"100101100",
  13065=>"010000110",
  13066=>"011111101",
  13067=>"111000100",
  13068=>"000001000",
  13069=>"110000110",
  13070=>"000110010",
  13071=>"101111011",
  13072=>"001001100",
  13073=>"111101011",
  13074=>"000111100",
  13075=>"110111001",
  13076=>"011011000",
  13077=>"011100001",
  13078=>"001010001",
  13079=>"111001010",
  13080=>"010011010",
  13081=>"001101100",
  13082=>"011010010",
  13083=>"101011111",
  13084=>"101111001",
  13085=>"001000111",
  13086=>"001000111",
  13087=>"100011000",
  13088=>"011010101",
  13089=>"000000111",
  13090=>"001111011",
  13091=>"111011101",
  13092=>"011101100",
  13093=>"100101010",
  13094=>"111011011",
  13095=>"111011011",
  13096=>"111100110",
  13097=>"000100011",
  13098=>"001101111",
  13099=>"010001001",
  13100=>"000101100",
  13101=>"100101001",
  13102=>"011100100",
  13103=>"101111100",
  13104=>"110000100",
  13105=>"010010101",
  13106=>"100001010",
  13107=>"110100011",
  13108=>"101110010",
  13109=>"010101011",
  13110=>"110101000",
  13111=>"001110111",
  13112=>"011010010",
  13113=>"110011000",
  13114=>"011110110",
  13115=>"101100000",
  13116=>"010110001",
  13117=>"100001010",
  13118=>"001010001",
  13119=>"110111010",
  13120=>"110010000",
  13121=>"111011001",
  13122=>"000111011",
  13123=>"110000100",
  13124=>"111011011",
  13125=>"001110101",
  13126=>"100000101",
  13127=>"000001101",
  13128=>"101001000",
  13129=>"011010110",
  13130=>"011011011",
  13131=>"000100010",
  13132=>"100010100",
  13133=>"100001110",
  13134=>"110111100",
  13135=>"010010010",
  13136=>"100110111",
  13137=>"011111000",
  13138=>"100000111",
  13139=>"100110110",
  13140=>"110011111",
  13141=>"011010100",
  13142=>"110000110",
  13143=>"111010000",
  13144=>"010110100",
  13145=>"100011101",
  13146=>"000000001",
  13147=>"100011101",
  13148=>"110110110",
  13149=>"100001111",
  13150=>"000010001",
  13151=>"000001000",
  13152=>"010000111",
  13153=>"010010010",
  13154=>"010001100",
  13155=>"100100011",
  13156=>"000011011",
  13157=>"100110000",
  13158=>"110100001",
  13159=>"010110010",
  13160=>"101011110",
  13161=>"011010111",
  13162=>"000010100",
  13163=>"010010010",
  13164=>"011111000",
  13165=>"111000111",
  13166=>"110011000",
  13167=>"001100010",
  13168=>"100111100",
  13169=>"110111011",
  13170=>"001000011",
  13171=>"001111111",
  13172=>"101001000",
  13173=>"100100001",
  13174=>"001100011",
  13175=>"101000000",
  13176=>"100001111",
  13177=>"000001001",
  13178=>"001001110",
  13179=>"010010111",
  13180=>"010001000",
  13181=>"011000100",
  13182=>"101101110",
  13183=>"000010000",
  13184=>"011101001",
  13185=>"110011101",
  13186=>"000111101",
  13187=>"001011001",
  13188=>"011010110",
  13189=>"010100010",
  13190=>"010111111",
  13191=>"011011101",
  13192=>"110111011",
  13193=>"111111111",
  13194=>"101011011",
  13195=>"011110100",
  13196=>"100010011",
  13197=>"100000000",
  13198=>"010111001",
  13199=>"101110000",
  13200=>"001000010",
  13201=>"101100111",
  13202=>"100000000",
  13203=>"010001000",
  13204=>"001100010",
  13205=>"110001110",
  13206=>"110100010",
  13207=>"110101111",
  13208=>"101010101",
  13209=>"001101001",
  13210=>"001110110",
  13211=>"111010101",
  13212=>"011101101",
  13213=>"000100010",
  13214=>"000111101",
  13215=>"100100101",
  13216=>"011011010",
  13217=>"011100100",
  13218=>"010110001",
  13219=>"100001011",
  13220=>"100000011",
  13221=>"000110111",
  13222=>"010010011",
  13223=>"010011000",
  13224=>"101110001",
  13225=>"000000110",
  13226=>"001101101",
  13227=>"110110111",
  13228=>"111100000",
  13229=>"000100111",
  13230=>"101101000",
  13231=>"101101110",
  13232=>"101011011",
  13233=>"100010111",
  13234=>"000100110",
  13235=>"110100001",
  13236=>"110000110",
  13237=>"110100111",
  13238=>"110001001",
  13239=>"000010101",
  13240=>"010110100",
  13241=>"000010100",
  13242=>"110011001",
  13243=>"011101010",
  13244=>"011111101",
  13245=>"010001111",
  13246=>"111001101",
  13247=>"100010111",
  13248=>"100110101",
  13249=>"000111110",
  13250=>"010101001",
  13251=>"100001110",
  13252=>"110000010",
  13253=>"011011110",
  13254=>"101010000",
  13255=>"010101001",
  13256=>"001100100",
  13257=>"001111001",
  13258=>"011011011",
  13259=>"010000111",
  13260=>"010011000",
  13261=>"000001111",
  13262=>"000000011",
  13263=>"100010111",
  13264=>"010001011",
  13265=>"000011110",
  13266=>"101010101",
  13267=>"111111111",
  13268=>"111011111",
  13269=>"011100010",
  13270=>"000001111",
  13271=>"010011100",
  13272=>"010000111",
  13273=>"000001101",
  13274=>"001010010",
  13275=>"000110011",
  13276=>"011111010",
  13277=>"110100001",
  13278=>"011011111",
  13279=>"011000100",
  13280=>"000111011",
  13281=>"101110001",
  13282=>"001110111",
  13283=>"101111101",
  13284=>"001010101",
  13285=>"010010101",
  13286=>"011111011",
  13287=>"010101101",
  13288=>"000001000",
  13289=>"111100010",
  13290=>"001000001",
  13291=>"001100100",
  13292=>"111111001",
  13293=>"110001000",
  13294=>"101001000",
  13295=>"001111111",
  13296=>"000001101",
  13297=>"010101010",
  13298=>"000101000",
  13299=>"010101101",
  13300=>"110101110",
  13301=>"010010111",
  13302=>"000101000",
  13303=>"101010110",
  13304=>"000111101",
  13305=>"010100111",
  13306=>"110100010",
  13307=>"111000000",
  13308=>"000100000",
  13309=>"010000001",
  13310=>"010110111",
  13311=>"101101000",
  13312=>"010011000",
  13313=>"101011010",
  13314=>"000101001",
  13315=>"000000110",
  13316=>"010101111",
  13317=>"010101000",
  13318=>"010000000",
  13319=>"111111110",
  13320=>"001001010",
  13321=>"010000000",
  13322=>"000011100",
  13323=>"001010011",
  13324=>"000011011",
  13325=>"111000001",
  13326=>"110000101",
  13327=>"111011101",
  13328=>"101011010",
  13329=>"000000000",
  13330=>"101101111",
  13331=>"010100010",
  13332=>"010000111",
  13333=>"101010010",
  13334=>"111100101",
  13335=>"110010001",
  13336=>"101001000",
  13337=>"010000000",
  13338=>"110010111",
  13339=>"011111011",
  13340=>"101111101",
  13341=>"101011100",
  13342=>"110110011",
  13343=>"111011000",
  13344=>"110111010",
  13345=>"000000100",
  13346=>"001110001",
  13347=>"110011011",
  13348=>"000000110",
  13349=>"110100000",
  13350=>"110111110",
  13351=>"100000111",
  13352=>"101000010",
  13353=>"000000011",
  13354=>"111110111",
  13355=>"010000111",
  13356=>"100001011",
  13357=>"111001010",
  13358=>"010111110",
  13359=>"111011110",
  13360=>"110111111",
  13361=>"001000111",
  13362=>"011100011",
  13363=>"100111100",
  13364=>"000000000",
  13365=>"010000010",
  13366=>"011110001",
  13367=>"100011011",
  13368=>"001001111",
  13369=>"110110110",
  13370=>"100101101",
  13371=>"000100000",
  13372=>"001111011",
  13373=>"100100010",
  13374=>"100000111",
  13375=>"110000001",
  13376=>"111001011",
  13377=>"001010100",
  13378=>"000111100",
  13379=>"011000100",
  13380=>"000010100",
  13381=>"010110000",
  13382=>"000010110",
  13383=>"111010000",
  13384=>"000011101",
  13385=>"110011010",
  13386=>"010111001",
  13387=>"000000011",
  13388=>"000001000",
  13389=>"000000111",
  13390=>"111111100",
  13391=>"001010010",
  13392=>"000101111",
  13393=>"111111000",
  13394=>"010001001",
  13395=>"000001111",
  13396=>"000101110",
  13397=>"000000110",
  13398=>"110011100",
  13399=>"010011110",
  13400=>"101000011",
  13401=>"110110000",
  13402=>"000010100",
  13403=>"001010001",
  13404=>"111001110",
  13405=>"000100011",
  13406=>"001010010",
  13407=>"100011101",
  13408=>"111100110",
  13409=>"001001000",
  13410=>"000011101",
  13411=>"011000010",
  13412=>"011111101",
  13413=>"100011101",
  13414=>"101011111",
  13415=>"011101001",
  13416=>"111100010",
  13417=>"101101001",
  13418=>"100110111",
  13419=>"111010111",
  13420=>"010000101",
  13421=>"100101100",
  13422=>"111001101",
  13423=>"000110011",
  13424=>"111000010",
  13425=>"001100101",
  13426=>"011000110",
  13427=>"000010011",
  13428=>"000010100",
  13429=>"100100010",
  13430=>"110100000",
  13431=>"001111010",
  13432=>"011011010",
  13433=>"100110110",
  13434=>"000010000",
  13435=>"110011110",
  13436=>"101111010",
  13437=>"001000010",
  13438=>"001010010",
  13439=>"011101011",
  13440=>"101000010",
  13441=>"010100010",
  13442=>"011000111",
  13443=>"110111011",
  13444=>"111101101",
  13445=>"000010011",
  13446=>"000000011",
  13447=>"101111010",
  13448=>"110111000",
  13449=>"001000101",
  13450=>"100101110",
  13451=>"101110010",
  13452=>"100111101",
  13453=>"010111001",
  13454=>"101011010",
  13455=>"011110010",
  13456=>"110101111",
  13457=>"100100010",
  13458=>"110000111",
  13459=>"110100100",
  13460=>"110000101",
  13461=>"000000000",
  13462=>"001111110",
  13463=>"110110100",
  13464=>"010110000",
  13465=>"011100110",
  13466=>"001001110",
  13467=>"110000111",
  13468=>"100011100",
  13469=>"111101100",
  13470=>"101011011",
  13471=>"011001010",
  13472=>"100010100",
  13473=>"111110111",
  13474=>"001010111",
  13475=>"101100001",
  13476=>"110010100",
  13477=>"100100110",
  13478=>"000010100",
  13479=>"010000000",
  13480=>"111001000",
  13481=>"111000000",
  13482=>"001000101",
  13483=>"011111010",
  13484=>"101011011",
  13485=>"001011011",
  13486=>"110111101",
  13487=>"100000000",
  13488=>"010000010",
  13489=>"110101100",
  13490=>"110111110",
  13491=>"101000010",
  13492=>"011110100",
  13493=>"000000111",
  13494=>"110001001",
  13495=>"000110100",
  13496=>"101001100",
  13497=>"100010101",
  13498=>"000011110",
  13499=>"001000100",
  13500=>"101000011",
  13501=>"110111101",
  13502=>"010101111",
  13503=>"110001011",
  13504=>"011010101",
  13505=>"010001010",
  13506=>"011110111",
  13507=>"110001010",
  13508=>"010000010",
  13509=>"110010111",
  13510=>"111000101",
  13511=>"000110010",
  13512=>"111011111",
  13513=>"000001010",
  13514=>"101000110",
  13515=>"101001101",
  13516=>"111110101",
  13517=>"100001111",
  13518=>"001001001",
  13519=>"100111000",
  13520=>"001100010",
  13521=>"000101111",
  13522=>"001101011",
  13523=>"110011000",
  13524=>"011111111",
  13525=>"010000000",
  13526=>"101111101",
  13527=>"101111000",
  13528=>"101111001",
  13529=>"101101111",
  13530=>"110011100",
  13531=>"110101101",
  13532=>"110000001",
  13533=>"000100010",
  13534=>"111100011",
  13535=>"101110100",
  13536=>"011111010",
  13537=>"111101011",
  13538=>"110010000",
  13539=>"101101001",
  13540=>"110011111",
  13541=>"100110101",
  13542=>"000010001",
  13543=>"010110111",
  13544=>"010001010",
  13545=>"001010001",
  13546=>"000000111",
  13547=>"101110011",
  13548=>"000000100",
  13549=>"110111001",
  13550=>"011010100",
  13551=>"000000101",
  13552=>"001111110",
  13553=>"110101010",
  13554=>"100110100",
  13555=>"101001011",
  13556=>"110001010",
  13557=>"000010101",
  13558=>"110000101",
  13559=>"000100101",
  13560=>"111111111",
  13561=>"111100110",
  13562=>"100011111",
  13563=>"010101000",
  13564=>"010011101",
  13565=>"111010000",
  13566=>"000100010",
  13567=>"111111111",
  13568=>"111100110",
  13569=>"101101101",
  13570=>"111000011",
  13571=>"101001010",
  13572=>"010010101",
  13573=>"101111001",
  13574=>"001011011",
  13575=>"111010001",
  13576=>"000010000",
  13577=>"100000110",
  13578=>"110011111",
  13579=>"111110011",
  13580=>"011001110",
  13581=>"111001010",
  13582=>"101001010",
  13583=>"010101110",
  13584=>"101100101",
  13585=>"100110110",
  13586=>"001111111",
  13587=>"111001111",
  13588=>"011011111",
  13589=>"110101111",
  13590=>"000001001",
  13591=>"101001110",
  13592=>"101001001",
  13593=>"011100000",
  13594=>"011010010",
  13595=>"111100011",
  13596=>"001011001",
  13597=>"111110101",
  13598=>"100111111",
  13599=>"000000010",
  13600=>"010000110",
  13601=>"101001100",
  13602=>"111101010",
  13603=>"000011010",
  13604=>"111000111",
  13605=>"100000100",
  13606=>"110010010",
  13607=>"000010001",
  13608=>"100000101",
  13609=>"000111111",
  13610=>"101101111",
  13611=>"011100010",
  13612=>"000010000",
  13613=>"111010100",
  13614=>"010011111",
  13615=>"010001100",
  13616=>"011101100",
  13617=>"111100000",
  13618=>"100010100",
  13619=>"011100110",
  13620=>"001110111",
  13621=>"011110101",
  13622=>"111001111",
  13623=>"111101001",
  13624=>"101011010",
  13625=>"010010110",
  13626=>"000010110",
  13627=>"101110000",
  13628=>"111010011",
  13629=>"001111101",
  13630=>"100000110",
  13631=>"100000101",
  13632=>"000010101",
  13633=>"000000101",
  13634=>"000000001",
  13635=>"111100000",
  13636=>"001010010",
  13637=>"011101101",
  13638=>"011101001",
  13639=>"100100000",
  13640=>"001111000",
  13641=>"111101110",
  13642=>"000010001",
  13643=>"111110001",
  13644=>"011011001",
  13645=>"111101101",
  13646=>"111001011",
  13647=>"011111111",
  13648=>"010011110",
  13649=>"110011010",
  13650=>"111000010",
  13651=>"001111001",
  13652=>"110000101",
  13653=>"111111111",
  13654=>"000010010",
  13655=>"000110001",
  13656=>"000010111",
  13657=>"101011110",
  13658=>"110010110",
  13659=>"111001101",
  13660=>"000101100",
  13661=>"100010000",
  13662=>"111101101",
  13663=>"000110011",
  13664=>"101101111",
  13665=>"101010010",
  13666=>"101110101",
  13667=>"000011011",
  13668=>"100100100",
  13669=>"000100000",
  13670=>"101011100",
  13671=>"101101101",
  13672=>"110001110",
  13673=>"100110000",
  13674=>"010001011",
  13675=>"101101101",
  13676=>"111101101",
  13677=>"111101000",
  13678=>"101100110",
  13679=>"110101011",
  13680=>"100110000",
  13681=>"010101000",
  13682=>"100001101",
  13683=>"001001111",
  13684=>"100111010",
  13685=>"000110100",
  13686=>"110100110",
  13687=>"000110111",
  13688=>"101101011",
  13689=>"011100111",
  13690=>"111010011",
  13691=>"011001110",
  13692=>"101010101",
  13693=>"011111111",
  13694=>"000001001",
  13695=>"110111100",
  13696=>"000000110",
  13697=>"011100100",
  13698=>"111001100",
  13699=>"111101001",
  13700=>"011000011",
  13701=>"111001111",
  13702=>"010101111",
  13703=>"110011010",
  13704=>"110110111",
  13705=>"110111111",
  13706=>"001011000",
  13707=>"000010010",
  13708=>"110001111",
  13709=>"110111001",
  13710=>"100111101",
  13711=>"010001111",
  13712=>"000000011",
  13713=>"001010000",
  13714=>"001110101",
  13715=>"011000110",
  13716=>"011001010",
  13717=>"000011100",
  13718=>"001011101",
  13719=>"010000011",
  13720=>"111000001",
  13721=>"000010010",
  13722=>"111111001",
  13723=>"000001000",
  13724=>"111011000",
  13725=>"011111010",
  13726=>"111001110",
  13727=>"101110000",
  13728=>"010001011",
  13729=>"010010000",
  13730=>"101001111",
  13731=>"101001011",
  13732=>"101001110",
  13733=>"011111111",
  13734=>"111101000",
  13735=>"000000111",
  13736=>"010100110",
  13737=>"001001100",
  13738=>"110111110",
  13739=>"010110110",
  13740=>"100111111",
  13741=>"000000101",
  13742=>"101100100",
  13743=>"111000011",
  13744=>"100101000",
  13745=>"010111101",
  13746=>"010011001",
  13747=>"001001111",
  13748=>"111100011",
  13749=>"101001010",
  13750=>"100110000",
  13751=>"010100100",
  13752=>"000110101",
  13753=>"011110101",
  13754=>"010000110",
  13755=>"011010000",
  13756=>"111010111",
  13757=>"000011011",
  13758=>"001110110",
  13759=>"111011111",
  13760=>"110010001",
  13761=>"010011110",
  13762=>"110011111",
  13763=>"000110111",
  13764=>"000000000",
  13765=>"000100001",
  13766=>"111000010",
  13767=>"100010010",
  13768=>"100010010",
  13769=>"110010001",
  13770=>"010111100",
  13771=>"110000001",
  13772=>"111100010",
  13773=>"110110110",
  13774=>"110001011",
  13775=>"101011101",
  13776=>"111100010",
  13777=>"111110110",
  13778=>"000000001",
  13779=>"110111010",
  13780=>"000111011",
  13781=>"110000001",
  13782=>"110101111",
  13783=>"010100010",
  13784=>"101110110",
  13785=>"100101111",
  13786=>"110000001",
  13787=>"001000111",
  13788=>"101001011",
  13789=>"011010110",
  13790=>"001101111",
  13791=>"111110111",
  13792=>"111010010",
  13793=>"001001101",
  13794=>"100101000",
  13795=>"010010100",
  13796=>"001110011",
  13797=>"000101001",
  13798=>"110111100",
  13799=>"000001000",
  13800=>"000111001",
  13801=>"100101111",
  13802=>"010111000",
  13803=>"110111010",
  13804=>"010011010",
  13805=>"011000100",
  13806=>"111100011",
  13807=>"000110000",
  13808=>"011101111",
  13809=>"000001101",
  13810=>"101011101",
  13811=>"011011100",
  13812=>"011010011",
  13813=>"010001111",
  13814=>"111101010",
  13815=>"011001100",
  13816=>"000110010",
  13817=>"011010100",
  13818=>"001111101",
  13819=>"101010101",
  13820=>"111000001",
  13821=>"100111101",
  13822=>"001011000",
  13823=>"011011100",
  13824=>"101100011",
  13825=>"010111100",
  13826=>"101000111",
  13827=>"100011011",
  13828=>"011110010",
  13829=>"100000100",
  13830=>"000010000",
  13831=>"000111001",
  13832=>"000100111",
  13833=>"010010000",
  13834=>"100101101",
  13835=>"110101000",
  13836=>"101101100",
  13837=>"001111110",
  13838=>"100000001",
  13839=>"001001010",
  13840=>"100010001",
  13841=>"000011100",
  13842=>"100101111",
  13843=>"101110110",
  13844=>"000110010",
  13845=>"010111100",
  13846=>"111101001",
  13847=>"001101101",
  13848=>"001111100",
  13849=>"010010001",
  13850=>"000100001",
  13851=>"001110101",
  13852=>"101011100",
  13853=>"010111111",
  13854=>"001010110",
  13855=>"100101000",
  13856=>"111010100",
  13857=>"110110011",
  13858=>"000111101",
  13859=>"101100001",
  13860=>"110001001",
  13861=>"100011100",
  13862=>"000111001",
  13863=>"010010111",
  13864=>"001111000",
  13865=>"001101010",
  13866=>"101000001",
  13867=>"101010000",
  13868=>"111010101",
  13869=>"101001101",
  13870=>"000100100",
  13871=>"100100011",
  13872=>"100000111",
  13873=>"000000000",
  13874=>"010111010",
  13875=>"101010001",
  13876=>"110010000",
  13877=>"010100100",
  13878=>"010100100",
  13879=>"100001011",
  13880=>"101011001",
  13881=>"100110100",
  13882=>"011010000",
  13883=>"011111111",
  13884=>"101111011",
  13885=>"010111111",
  13886=>"101101000",
  13887=>"100000110",
  13888=>"111000100",
  13889=>"101101010",
  13890=>"010111110",
  13891=>"010110000",
  13892=>"101011101",
  13893=>"001001100",
  13894=>"100000010",
  13895=>"010111010",
  13896=>"101100011",
  13897=>"000100000",
  13898=>"011110101",
  13899=>"111011100",
  13900=>"110111101",
  13901=>"101010100",
  13902=>"001010111",
  13903=>"110111101",
  13904=>"010101000",
  13905=>"000001000",
  13906=>"110101101",
  13907=>"110000011",
  13908=>"011010000",
  13909=>"000001001",
  13910=>"001111101",
  13911=>"011110011",
  13912=>"110011111",
  13913=>"001011001",
  13914=>"001110001",
  13915=>"001011000",
  13916=>"100111100",
  13917=>"111011011",
  13918=>"101011001",
  13919=>"100000101",
  13920=>"100011101",
  13921=>"100010001",
  13922=>"001101100",
  13923=>"010010110",
  13924=>"000101000",
  13925=>"101010010",
  13926=>"011010011",
  13927=>"001110011",
  13928=>"110001111",
  13929=>"101001100",
  13930=>"111111100",
  13931=>"000000000",
  13932=>"111010011",
  13933=>"101100101",
  13934=>"110100111",
  13935=>"111011101",
  13936=>"100001111",
  13937=>"001110111",
  13938=>"010110110",
  13939=>"110011010",
  13940=>"111110101",
  13941=>"101101010",
  13942=>"111101000",
  13943=>"111000111",
  13944=>"000000110",
  13945=>"000101100",
  13946=>"000011000",
  13947=>"100001001",
  13948=>"001101000",
  13949=>"000001010",
  13950=>"101111001",
  13951=>"100010011",
  13952=>"011111000",
  13953=>"110000101",
  13954=>"001010110",
  13955=>"011001011",
  13956=>"111001000",
  13957=>"000000010",
  13958=>"001011011",
  13959=>"011110100",
  13960=>"101010101",
  13961=>"000101110",
  13962=>"101000001",
  13963=>"001110100",
  13964=>"001111111",
  13965=>"001011100",
  13966=>"000111000",
  13967=>"100010100",
  13968=>"111001101",
  13969=>"100000000",
  13970=>"011110101",
  13971=>"011011101",
  13972=>"111010001",
  13973=>"111011011",
  13974=>"011111111",
  13975=>"101111101",
  13976=>"001100100",
  13977=>"001010000",
  13978=>"000101111",
  13979=>"001001000",
  13980=>"111100011",
  13981=>"110111110",
  13982=>"001100011",
  13983=>"011100001",
  13984=>"010010101",
  13985=>"111101011",
  13986=>"000100010",
  13987=>"001000001",
  13988=>"111001101",
  13989=>"011111000",
  13990=>"011101010",
  13991=>"111100000",
  13992=>"001100100",
  13993=>"010001000",
  13994=>"000010100",
  13995=>"001010010",
  13996=>"101101111",
  13997=>"110100010",
  13998=>"000100011",
  13999=>"000000100",
  14000=>"110110000",
  14001=>"111000001",
  14002=>"111001101",
  14003=>"100010100",
  14004=>"001001000",
  14005=>"111100000",
  14006=>"101011111",
  14007=>"010111101",
  14008=>"001100011",
  14009=>"010100000",
  14010=>"111100011",
  14011=>"101010100",
  14012=>"001000110",
  14013=>"010110000",
  14014=>"110001000",
  14015=>"101010110",
  14016=>"000010111",
  14017=>"001110100",
  14018=>"111111010",
  14019=>"011110001",
  14020=>"001001111",
  14021=>"110000000",
  14022=>"010011010",
  14023=>"011001110",
  14024=>"101111100",
  14025=>"100001010",
  14026=>"010100100",
  14027=>"000011011",
  14028=>"011010111",
  14029=>"001111101",
  14030=>"111000111",
  14031=>"001000101",
  14032=>"100111000",
  14033=>"111111100",
  14034=>"111101001",
  14035=>"010101000",
  14036=>"011111001",
  14037=>"010000000",
  14038=>"000110001",
  14039=>"010100011",
  14040=>"000000000",
  14041=>"110110110",
  14042=>"111111111",
  14043=>"010010000",
  14044=>"110001101",
  14045=>"010001111",
  14046=>"111001001",
  14047=>"110001000",
  14048=>"111010011",
  14049=>"011001101",
  14050=>"010111110",
  14051=>"110010001",
  14052=>"111101000",
  14053=>"100100111",
  14054=>"111000010",
  14055=>"110001111",
  14056=>"010011010",
  14057=>"111110111",
  14058=>"010001011",
  14059=>"011001011",
  14060=>"011010010",
  14061=>"110010011",
  14062=>"001000111",
  14063=>"110001110",
  14064=>"111011010",
  14065=>"001110110",
  14066=>"111011111",
  14067=>"010110111",
  14068=>"001001010",
  14069=>"001000010",
  14070=>"000101010",
  14071=>"100010011",
  14072=>"011010000",
  14073=>"110110111",
  14074=>"001110001",
  14075=>"100000010",
  14076=>"001110011",
  14077=>"011101000",
  14078=>"000111000",
  14079=>"011100000",
  14080=>"001001001",
  14081=>"111011111",
  14082=>"111101101",
  14083=>"101000001",
  14084=>"101010001",
  14085=>"000000011",
  14086=>"001010001",
  14087=>"111110001",
  14088=>"111011101",
  14089=>"110111000",
  14090=>"001110110",
  14091=>"100111111",
  14092=>"001100000",
  14093=>"111010111",
  14094=>"000001100",
  14095=>"110000001",
  14096=>"101100101",
  14097=>"000000111",
  14098=>"101111101",
  14099=>"001110101",
  14100=>"111100111",
  14101=>"000001001",
  14102=>"000111100",
  14103=>"110110100",
  14104=>"100011011",
  14105=>"001001100",
  14106=>"011111010",
  14107=>"111011010",
  14108=>"100001010",
  14109=>"010101011",
  14110=>"000111010",
  14111=>"010100011",
  14112=>"101100010",
  14113=>"110100100",
  14114=>"010011000",
  14115=>"100100001",
  14116=>"100011100",
  14117=>"010111000",
  14118=>"011111011",
  14119=>"110010111",
  14120=>"111110001",
  14121=>"010100100",
  14122=>"001100100",
  14123=>"011100001",
  14124=>"100101001",
  14125=>"111010100",
  14126=>"000010001",
  14127=>"000011011",
  14128=>"011001010",
  14129=>"001111001",
  14130=>"111110001",
  14131=>"011010010",
  14132=>"111011110",
  14133=>"100001101",
  14134=>"100111101",
  14135=>"011110001",
  14136=>"000001100",
  14137=>"100001000",
  14138=>"001011111",
  14139=>"100100101",
  14140=>"110011100",
  14141=>"111010011",
  14142=>"101101010",
  14143=>"110110111",
  14144=>"101001000",
  14145=>"010001100",
  14146=>"110100101",
  14147=>"101100110",
  14148=>"001010001",
  14149=>"111000000",
  14150=>"001001111",
  14151=>"000001100",
  14152=>"000100101",
  14153=>"011101000",
  14154=>"101100010",
  14155=>"001111100",
  14156=>"001101111",
  14157=>"111100110",
  14158=>"101000100",
  14159=>"101101100",
  14160=>"010111001",
  14161=>"101001100",
  14162=>"001111000",
  14163=>"000000010",
  14164=>"111111110",
  14165=>"111111000",
  14166=>"111010110",
  14167=>"101101100",
  14168=>"010110001",
  14169=>"000000001",
  14170=>"001101100",
  14171=>"010010100",
  14172=>"010010001",
  14173=>"101100011",
  14174=>"001101111",
  14175=>"100100011",
  14176=>"100111101",
  14177=>"110011101",
  14178=>"010111111",
  14179=>"110100100",
  14180=>"000010111",
  14181=>"000010110",
  14182=>"101001110",
  14183=>"011001111",
  14184=>"100100111",
  14185=>"010011111",
  14186=>"101110011",
  14187=>"110001110",
  14188=>"110011010",
  14189=>"011100001",
  14190=>"101100100",
  14191=>"111111100",
  14192=>"111010111",
  14193=>"000100110",
  14194=>"111101101",
  14195=>"001001000",
  14196=>"110101101",
  14197=>"111100111",
  14198=>"110000000",
  14199=>"100000100",
  14200=>"001010111",
  14201=>"111001111",
  14202=>"110011000",
  14203=>"111001111",
  14204=>"100101000",
  14205=>"111111111",
  14206=>"011011011",
  14207=>"101101111",
  14208=>"100001010",
  14209=>"011110000",
  14210=>"001011111",
  14211=>"111111100",
  14212=>"101000110",
  14213=>"010111111",
  14214=>"101001110",
  14215=>"100101110",
  14216=>"110001000",
  14217=>"010011101",
  14218=>"011110001",
  14219=>"001010011",
  14220=>"100100001",
  14221=>"111111011",
  14222=>"100110010",
  14223=>"100010111",
  14224=>"010111100",
  14225=>"110001000",
  14226=>"000010010",
  14227=>"101110010",
  14228=>"100000111",
  14229=>"100110000",
  14230=>"111111000",
  14231=>"111111001",
  14232=>"110111110",
  14233=>"000001010",
  14234=>"110011010",
  14235=>"010010001",
  14236=>"000100100",
  14237=>"111011111",
  14238=>"000011101",
  14239=>"101110010",
  14240=>"001001011",
  14241=>"101100100",
  14242=>"101110001",
  14243=>"000101110",
  14244=>"001110010",
  14245=>"101001010",
  14246=>"001001100",
  14247=>"010101101",
  14248=>"000001100",
  14249=>"110111010",
  14250=>"010100110",
  14251=>"100001100",
  14252=>"101101110",
  14253=>"010111101",
  14254=>"001010100",
  14255=>"111100100",
  14256=>"001101010",
  14257=>"111111001",
  14258=>"100100000",
  14259=>"010100011",
  14260=>"111010000",
  14261=>"111100110",
  14262=>"100000110",
  14263=>"001001111",
  14264=>"010111100",
  14265=>"100100011",
  14266=>"001001001",
  14267=>"000110100",
  14268=>"101010111",
  14269=>"000111000",
  14270=>"111010111",
  14271=>"110001011",
  14272=>"011101000",
  14273=>"110101101",
  14274=>"100100001",
  14275=>"001110011",
  14276=>"110010011",
  14277=>"010111101",
  14278=>"111110000",
  14279=>"001001101",
  14280=>"010111110",
  14281=>"001010101",
  14282=>"011010001",
  14283=>"111111011",
  14284=>"000101000",
  14285=>"111100100",
  14286=>"001100111",
  14287=>"011110000",
  14288=>"110111110",
  14289=>"000111001",
  14290=>"011011110",
  14291=>"111100101",
  14292=>"101100001",
  14293=>"001111111",
  14294=>"010100110",
  14295=>"101111000",
  14296=>"010111110",
  14297=>"001000100",
  14298=>"111001011",
  14299=>"110001010",
  14300=>"111101100",
  14301=>"011000111",
  14302=>"010010110",
  14303=>"010011011",
  14304=>"101011110",
  14305=>"111110001",
  14306=>"011111100",
  14307=>"001000101",
  14308=>"011111000",
  14309=>"000010010",
  14310=>"111110110",
  14311=>"011001100",
  14312=>"111100010",
  14313=>"101011001",
  14314=>"000110010",
  14315=>"011101010",
  14316=>"101100011",
  14317=>"010110000",
  14318=>"011101111",
  14319=>"101001001",
  14320=>"000011000",
  14321=>"011111101",
  14322=>"010101010",
  14323=>"000111010",
  14324=>"011100000",
  14325=>"100000000",
  14326=>"110110100",
  14327=>"110111111",
  14328=>"111010110",
  14329=>"111101110",
  14330=>"110000100",
  14331=>"101110100",
  14332=>"110011011",
  14333=>"101001011",
  14334=>"001110011",
  14335=>"100001010",
  14336=>"110111001",
  14337=>"100011000",
  14338=>"010001001",
  14339=>"101001000",
  14340=>"000001000",
  14341=>"011110110",
  14342=>"010011111",
  14343=>"011110111",
  14344=>"110011100",
  14345=>"001100110",
  14346=>"011001010",
  14347=>"110001001",
  14348=>"110100100",
  14349=>"001101011",
  14350=>"001111010",
  14351=>"110000110",
  14352=>"101110101",
  14353=>"101001101",
  14354=>"100100101",
  14355=>"111010011",
  14356=>"111101100",
  14357=>"100000110",
  14358=>"111101111",
  14359=>"100100000",
  14360=>"111100010",
  14361=>"111101111",
  14362=>"001001011",
  14363=>"001111010",
  14364=>"111100101",
  14365=>"011000101",
  14366=>"111011000",
  14367=>"100110111",
  14368=>"011011001",
  14369=>"000010101",
  14370=>"000000101",
  14371=>"111010100",
  14372=>"000011110",
  14373=>"101100000",
  14374=>"000010100",
  14375=>"110000011",
  14376=>"101001001",
  14377=>"000100011",
  14378=>"010110111",
  14379=>"000011100",
  14380=>"110011110",
  14381=>"111000110",
  14382=>"111101011",
  14383=>"010001110",
  14384=>"010111110",
  14385=>"110110000",
  14386=>"000111110",
  14387=>"010111100",
  14388=>"111011001",
  14389=>"010101011",
  14390=>"000010000",
  14391=>"001100100",
  14392=>"011011001",
  14393=>"110000111",
  14394=>"001110000",
  14395=>"101010101",
  14396=>"010001110",
  14397=>"011111000",
  14398=>"001101100",
  14399=>"101111001",
  14400=>"000001101",
  14401=>"111001001",
  14402=>"110111010",
  14403=>"111101000",
  14404=>"000100110",
  14405=>"000100001",
  14406=>"101101010",
  14407=>"001001110",
  14408=>"100111010",
  14409=>"110001101",
  14410=>"001110110",
  14411=>"111100000",
  14412=>"101010001",
  14413=>"001010001",
  14414=>"001010001",
  14415=>"111100111",
  14416=>"000100101",
  14417=>"000000101",
  14418=>"010111011",
  14419=>"000000000",
  14420=>"001000001",
  14421=>"000000111",
  14422=>"000100011",
  14423=>"011001000",
  14424=>"111111011",
  14425=>"011001000",
  14426=>"100001000",
  14427=>"011010111",
  14428=>"000011010",
  14429=>"101011001",
  14430=>"010001001",
  14431=>"000110100",
  14432=>"101101001",
  14433=>"110111101",
  14434=>"100011101",
  14435=>"011010101",
  14436=>"111111100",
  14437=>"001010011",
  14438=>"001111111",
  14439=>"001101000",
  14440=>"101001111",
  14441=>"000101100",
  14442=>"011100110",
  14443=>"101101000",
  14444=>"001101000",
  14445=>"010000000",
  14446=>"101110100",
  14447=>"111110111",
  14448=>"111111000",
  14449=>"000110110",
  14450=>"110111111",
  14451=>"110111001",
  14452=>"011110101",
  14453=>"111110011",
  14454=>"001010111",
  14455=>"011100001",
  14456=>"110111010",
  14457=>"001000100",
  14458=>"111011001",
  14459=>"011001001",
  14460=>"001000111",
  14461=>"111101100",
  14462=>"111111010",
  14463=>"000101011",
  14464=>"000000010",
  14465=>"111111011",
  14466=>"010010111",
  14467=>"110101001",
  14468=>"001010000",
  14469=>"100011000",
  14470=>"111010001",
  14471=>"001111101",
  14472=>"100001111",
  14473=>"001010001",
  14474=>"110010110",
  14475=>"111101010",
  14476=>"000101001",
  14477=>"111100100",
  14478=>"000001111",
  14479=>"100101000",
  14480=>"010100010",
  14481=>"111010001",
  14482=>"111111000",
  14483=>"010000111",
  14484=>"101000101",
  14485=>"000110001",
  14486=>"010010000",
  14487=>"001110000",
  14488=>"000001000",
  14489=>"110000011",
  14490=>"010010000",
  14491=>"110111010",
  14492=>"000110000",
  14493=>"000010101",
  14494=>"100011111",
  14495=>"001001100",
  14496=>"101000101",
  14497=>"110101101",
  14498=>"111001000",
  14499=>"110010110",
  14500=>"101111001",
  14501=>"100010100",
  14502=>"001001100",
  14503=>"100000000",
  14504=>"111111111",
  14505=>"001101011",
  14506=>"100101011",
  14507=>"110101100",
  14508=>"011101110",
  14509=>"010010111",
  14510=>"010101110",
  14511=>"000010101",
  14512=>"110000001",
  14513=>"110111101",
  14514=>"101000101",
  14515=>"000110010",
  14516=>"111000011",
  14517=>"001011101",
  14518=>"110111110",
  14519=>"110110011",
  14520=>"000000000",
  14521=>"110110000",
  14522=>"011110010",
  14523=>"110001010",
  14524=>"111010110",
  14525=>"010000001",
  14526=>"101111000",
  14527=>"111001111",
  14528=>"111000111",
  14529=>"101100010",
  14530=>"011010110",
  14531=>"110110111",
  14532=>"001101101",
  14533=>"010010011",
  14534=>"111010101",
  14535=>"011100000",
  14536=>"011010100",
  14537=>"010001101",
  14538=>"011111111",
  14539=>"101001001",
  14540=>"111011010",
  14541=>"010101111",
  14542=>"001000110",
  14543=>"110011000",
  14544=>"110010100",
  14545=>"000101110",
  14546=>"111000111",
  14547=>"110011010",
  14548=>"100110000",
  14549=>"110001110",
  14550=>"001110100",
  14551=>"010100101",
  14552=>"001100000",
  14553=>"100000110",
  14554=>"011100100",
  14555=>"100101000",
  14556=>"100010000",
  14557=>"110000101",
  14558=>"100011110",
  14559=>"000110110",
  14560=>"000101100",
  14561=>"111101011",
  14562=>"000000100",
  14563=>"111000000",
  14564=>"001000111",
  14565=>"000010101",
  14566=>"110111110",
  14567=>"111101101",
  14568=>"101000100",
  14569=>"011010000",
  14570=>"100010110",
  14571=>"001001010",
  14572=>"101001000",
  14573=>"010110100",
  14574=>"101010100",
  14575=>"011110111",
  14576=>"001111100",
  14577=>"100001101",
  14578=>"001111000",
  14579=>"110111101",
  14580=>"011110000",
  14581=>"111001000",
  14582=>"110001110",
  14583=>"010100110",
  14584=>"110000100",
  14585=>"111100111",
  14586=>"001111101",
  14587=>"110011010",
  14588=>"111100101",
  14589=>"011001110",
  14590=>"000100001",
  14591=>"111001110",
  14592=>"010000000",
  14593=>"011101111",
  14594=>"011110111",
  14595=>"010011111",
  14596=>"010000110",
  14597=>"000000001",
  14598=>"111011000",
  14599=>"101011001",
  14600=>"111011100",
  14601=>"101110010",
  14602=>"111011111",
  14603=>"100100000",
  14604=>"000111000",
  14605=>"110111010",
  14606=>"001101000",
  14607=>"111111001",
  14608=>"111100100",
  14609=>"101110100",
  14610=>"111100111",
  14611=>"010101101",
  14612=>"001010111",
  14613=>"100010100",
  14614=>"000111110",
  14615=>"100000100",
  14616=>"100010001",
  14617=>"000101001",
  14618=>"100011001",
  14619=>"110010100",
  14620=>"011000010",
  14621=>"011111000",
  14622=>"111110000",
  14623=>"111001101",
  14624=>"110001100",
  14625=>"001001011",
  14626=>"101110011",
  14627=>"111011010",
  14628=>"110011101",
  14629=>"001011100",
  14630=>"000100101",
  14631=>"000001111",
  14632=>"001110111",
  14633=>"110111001",
  14634=>"001010000",
  14635=>"111010110",
  14636=>"100111111",
  14637=>"011100000",
  14638=>"100001010",
  14639=>"111111101",
  14640=>"011101100",
  14641=>"111111111",
  14642=>"110101110",
  14643=>"000010110",
  14644=>"101000001",
  14645=>"011001101",
  14646=>"001010110",
  14647=>"111110010",
  14648=>"111011000",
  14649=>"111101001",
  14650=>"111100101",
  14651=>"010101101",
  14652=>"111101111",
  14653=>"000011110",
  14654=>"111110100",
  14655=>"101010000",
  14656=>"001111011",
  14657=>"011011101",
  14658=>"101110000",
  14659=>"110111000",
  14660=>"000001010",
  14661=>"111001001",
  14662=>"011000101",
  14663=>"110100101",
  14664=>"100010100",
  14665=>"000110000",
  14666=>"101011011",
  14667=>"110000000",
  14668=>"000111100",
  14669=>"111011111",
  14670=>"000010000",
  14671=>"010110001",
  14672=>"110010101",
  14673=>"011000101",
  14674=>"100001011",
  14675=>"111101110",
  14676=>"001010111",
  14677=>"110101011",
  14678=>"000110000",
  14679=>"101101001",
  14680=>"000000000",
  14681=>"100000101",
  14682=>"000000010",
  14683=>"011100110",
  14684=>"111111101",
  14685=>"011010101",
  14686=>"111010111",
  14687=>"100011100",
  14688=>"000100010",
  14689=>"101010110",
  14690=>"000000000",
  14691=>"000011010",
  14692=>"001000101",
  14693=>"011000111",
  14694=>"100101101",
  14695=>"001011011",
  14696=>"010011100",
  14697=>"011001001",
  14698=>"011100001",
  14699=>"111101000",
  14700=>"001001010",
  14701=>"110110010",
  14702=>"111100100",
  14703=>"011100101",
  14704=>"000100011",
  14705=>"000011100",
  14706=>"110000010",
  14707=>"001110000",
  14708=>"000110010",
  14709=>"101011111",
  14710=>"000101001",
  14711=>"011100101",
  14712=>"101100011",
  14713=>"001111100",
  14714=>"100111100",
  14715=>"110110111",
  14716=>"100001010",
  14717=>"000011111",
  14718=>"000001101",
  14719=>"110111100",
  14720=>"111110111",
  14721=>"000011000",
  14722=>"010110101",
  14723=>"100011101",
  14724=>"101100011",
  14725=>"111101010",
  14726=>"011101110",
  14727=>"100100010",
  14728=>"001001001",
  14729=>"111111001",
  14730=>"100111001",
  14731=>"100110000",
  14732=>"001010111",
  14733=>"010110110",
  14734=>"001010011",
  14735=>"011110111",
  14736=>"011001010",
  14737=>"000010011",
  14738=>"001011100",
  14739=>"010110010",
  14740=>"100011011",
  14741=>"000001110",
  14742=>"001100000",
  14743=>"001110111",
  14744=>"010100001",
  14745=>"101111100",
  14746=>"010000011",
  14747=>"010010010",
  14748=>"111001100",
  14749=>"101101101",
  14750=>"000111011",
  14751=>"010100101",
  14752=>"010000000",
  14753=>"111011100",
  14754=>"011001101",
  14755=>"011100110",
  14756=>"000001111",
  14757=>"110001101",
  14758=>"101001101",
  14759=>"001100111",
  14760=>"111010111",
  14761=>"001001010",
  14762=>"000111110",
  14763=>"111111010",
  14764=>"111110101",
  14765=>"110010110",
  14766=>"000010011",
  14767=>"111110001",
  14768=>"001100001",
  14769=>"110110000",
  14770=>"100110011",
  14771=>"010101101",
  14772=>"001010100",
  14773=>"000001100",
  14774=>"101001101",
  14775=>"000101010",
  14776=>"101000010",
  14777=>"111001100",
  14778=>"101111010",
  14779=>"011100001",
  14780=>"111101010",
  14781=>"011001010",
  14782=>"000001011",
  14783=>"001100100",
  14784=>"001000001",
  14785=>"110111001",
  14786=>"001011110",
  14787=>"110101111",
  14788=>"010101001",
  14789=>"000001000",
  14790=>"001100001",
  14791=>"110111100",
  14792=>"110101011",
  14793=>"101001000",
  14794=>"101100111",
  14795=>"100110101",
  14796=>"001000010",
  14797=>"110011101",
  14798=>"100001011",
  14799=>"000110110",
  14800=>"110010101",
  14801=>"011011110",
  14802=>"011001011",
  14803=>"111011010",
  14804=>"100001101",
  14805=>"110001100",
  14806=>"111111101",
  14807=>"111111100",
  14808=>"111010111",
  14809=>"000001010",
  14810=>"111100010",
  14811=>"110110101",
  14812=>"111000001",
  14813=>"111101000",
  14814=>"001001001",
  14815=>"011010000",
  14816=>"001010111",
  14817=>"111100001",
  14818=>"010101000",
  14819=>"111000100",
  14820=>"010100110",
  14821=>"101001101",
  14822=>"110000100",
  14823=>"101000101",
  14824=>"110000011",
  14825=>"100101100",
  14826=>"110101000",
  14827=>"100001100",
  14828=>"010001011",
  14829=>"000011110",
  14830=>"001001110",
  14831=>"010110000",
  14832=>"111110000",
  14833=>"110000111",
  14834=>"101110010",
  14835=>"010110001",
  14836=>"001101101",
  14837=>"001000001",
  14838=>"010100011",
  14839=>"001010010",
  14840=>"111000000",
  14841=>"001011101",
  14842=>"000101001",
  14843=>"111100110",
  14844=>"010101100",
  14845=>"010111010",
  14846=>"101110010",
  14847=>"010011010",
  14848=>"000110011",
  14849=>"111010100",
  14850=>"101011011",
  14851=>"000011000",
  14852=>"011000000",
  14853=>"000001001",
  14854=>"111011011",
  14855=>"101110001",
  14856=>"000000001",
  14857=>"110001001",
  14858=>"000101101",
  14859=>"111111110",
  14860=>"000010010",
  14861=>"000110001",
  14862=>"100100111",
  14863=>"011001111",
  14864=>"111111110",
  14865=>"011101010",
  14866=>"000100000",
  14867=>"011101001",
  14868=>"000001010",
  14869=>"110001111",
  14870=>"100110011",
  14871=>"011010000",
  14872=>"000110000",
  14873=>"100100111",
  14874=>"110101000",
  14875=>"011101001",
  14876=>"010111111",
  14877=>"010000011",
  14878=>"111001010",
  14879=>"010001110",
  14880=>"100101010",
  14881=>"011011001",
  14882=>"100100011",
  14883=>"100001010",
  14884=>"101111111",
  14885=>"011111000",
  14886=>"110100111",
  14887=>"100101100",
  14888=>"100001001",
  14889=>"111011001",
  14890=>"100010100",
  14891=>"100100000",
  14892=>"001100101",
  14893=>"011001101",
  14894=>"100001111",
  14895=>"111010111",
  14896=>"101100010",
  14897=>"011101111",
  14898=>"100101001",
  14899=>"000011111",
  14900=>"100000001",
  14901=>"001011111",
  14902=>"110110000",
  14903=>"011110101",
  14904=>"111000100",
  14905=>"111110101",
  14906=>"000011001",
  14907=>"010111100",
  14908=>"000011010",
  14909=>"011010001",
  14910=>"111010100",
  14911=>"001101111",
  14912=>"000110000",
  14913=>"110111110",
  14914=>"111011100",
  14915=>"011000101",
  14916=>"100100001",
  14917=>"101000100",
  14918=>"100100110",
  14919=>"100100100",
  14920=>"011000111",
  14921=>"001001101",
  14922=>"111000101",
  14923=>"110100001",
  14924=>"000101101",
  14925=>"110111010",
  14926=>"010110100",
  14927=>"001011011",
  14928=>"001001011",
  14929=>"010110011",
  14930=>"010100000",
  14931=>"110001001",
  14932=>"111010100",
  14933=>"100111101",
  14934=>"000011001",
  14935=>"010011111",
  14936=>"111010011",
  14937=>"101110100",
  14938=>"111101100",
  14939=>"010111010",
  14940=>"110100100",
  14941=>"110100010",
  14942=>"111010011",
  14943=>"100000111",
  14944=>"001101000",
  14945=>"000110010",
  14946=>"110011101",
  14947=>"101100111",
  14948=>"100111110",
  14949=>"000111101",
  14950=>"010010110",
  14951=>"000110010",
  14952=>"101001010",
  14953=>"010000000",
  14954=>"010111011",
  14955=>"010110000",
  14956=>"111010111",
  14957=>"111101011",
  14958=>"110010001",
  14959=>"110010100",
  14960=>"000101001",
  14961=>"111101101",
  14962=>"011000000",
  14963=>"111000011",
  14964=>"010001111",
  14965=>"110011100",
  14966=>"101111011",
  14967=>"101100100",
  14968=>"010010010",
  14969=>"010100010",
  14970=>"000010111",
  14971=>"001011100",
  14972=>"011011101",
  14973=>"011001100",
  14974=>"010110100",
  14975=>"011111100",
  14976=>"011111101",
  14977=>"011001011",
  14978=>"110011100",
  14979=>"110110110",
  14980=>"000010010",
  14981=>"011100101",
  14982=>"110001101",
  14983=>"010001100",
  14984=>"010110011",
  14985=>"000001001",
  14986=>"011111000",
  14987=>"111101011",
  14988=>"010000001",
  14989=>"000101110",
  14990=>"111111101",
  14991=>"010100111",
  14992=>"011011010",
  14993=>"111000100",
  14994=>"010110101",
  14995=>"010111111",
  14996=>"000000001",
  14997=>"110101011",
  14998=>"011110010",
  14999=>"100101000",
  15000=>"101111111",
  15001=>"010100000",
  15002=>"001000111",
  15003=>"001001111",
  15004=>"000010111",
  15005=>"000110000",
  15006=>"101011111",
  15007=>"101110000",
  15008=>"100011011",
  15009=>"101010111",
  15010=>"001000110",
  15011=>"010001000",
  15012=>"010001000",
  15013=>"000101101",
  15014=>"100000110",
  15015=>"101111000",
  15016=>"001001101",
  15017=>"000100001",
  15018=>"010000000",
  15019=>"110110001",
  15020=>"011010111",
  15021=>"100101111",
  15022=>"010111111",
  15023=>"010011011",
  15024=>"101011011",
  15025=>"101110100",
  15026=>"100101110",
  15027=>"110110000",
  15028=>"111111010",
  15029=>"111011010",
  15030=>"101001111",
  15031=>"111010100",
  15032=>"111001100",
  15033=>"110111101",
  15034=>"000100001",
  15035=>"000011001",
  15036=>"000110101",
  15037=>"001010101",
  15038=>"111101101",
  15039=>"000000111",
  15040=>"111110100",
  15041=>"111011001",
  15042=>"010100000",
  15043=>"011111001",
  15044=>"111111010",
  15045=>"100100100",
  15046=>"000100011",
  15047=>"001011000",
  15048=>"011001101",
  15049=>"010000000",
  15050=>"110110010",
  15051=>"110100111",
  15052=>"010010011",
  15053=>"101010001",
  15054=>"111110000",
  15055=>"000010101",
  15056=>"111010111",
  15057=>"100011110",
  15058=>"111101100",
  15059=>"100100011",
  15060=>"101011101",
  15061=>"011111001",
  15062=>"001001110",
  15063=>"001101111",
  15064=>"101001001",
  15065=>"110101011",
  15066=>"000010001",
  15067=>"101110001",
  15068=>"001101101",
  15069=>"100111110",
  15070=>"001011111",
  15071=>"001110100",
  15072=>"110001110",
  15073=>"010000000",
  15074=>"111100001",
  15075=>"001111001",
  15076=>"111000000",
  15077=>"011110100",
  15078=>"111111010",
  15079=>"100100100",
  15080=>"101101011",
  15081=>"011100110",
  15082=>"011010010",
  15083=>"101100000",
  15084=>"111100010",
  15085=>"100101111",
  15086=>"001101101",
  15087=>"110000100",
  15088=>"110011100",
  15089=>"000010111",
  15090=>"001001010",
  15091=>"000100000",
  15092=>"110001011",
  15093=>"111011000",
  15094=>"011001011",
  15095=>"001001001",
  15096=>"101001111",
  15097=>"101101101",
  15098=>"011011101",
  15099=>"100101111",
  15100=>"100000011",
  15101=>"110000100",
  15102=>"100010101",
  15103=>"000111011",
  15104=>"111100110",
  15105=>"001011001",
  15106=>"110100111",
  15107=>"001000001",
  15108=>"000101001",
  15109=>"010011001",
  15110=>"001000111",
  15111=>"011111001",
  15112=>"110100101",
  15113=>"101111010",
  15114=>"110111001",
  15115=>"000000010",
  15116=>"111000010",
  15117=>"000001110",
  15118=>"001010010",
  15119=>"000010010",
  15120=>"100101101",
  15121=>"001000001",
  15122=>"011110000",
  15123=>"010000010",
  15124=>"011011100",
  15125=>"011110001",
  15126=>"100111111",
  15127=>"001001100",
  15128=>"001011010",
  15129=>"010011010",
  15130=>"010110001",
  15131=>"010101001",
  15132=>"100000001",
  15133=>"011100100",
  15134=>"000110011",
  15135=>"001101001",
  15136=>"000000101",
  15137=>"010111111",
  15138=>"111001011",
  15139=>"110101100",
  15140=>"000001100",
  15141=>"111111101",
  15142=>"111111110",
  15143=>"011001111",
  15144=>"001000000",
  15145=>"000011011",
  15146=>"100011010",
  15147=>"001111000",
  15148=>"011011101",
  15149=>"000000100",
  15150=>"010001010",
  15151=>"100100001",
  15152=>"011101101",
  15153=>"010001011",
  15154=>"011010001",
  15155=>"001001001",
  15156=>"011001000",
  15157=>"011111111",
  15158=>"100110011",
  15159=>"000100100",
  15160=>"011011010",
  15161=>"001101110",
  15162=>"100000010",
  15163=>"011101010",
  15164=>"111110010",
  15165=>"001110110",
  15166=>"100011101",
  15167=>"000110110",
  15168=>"101100101",
  15169=>"111010011",
  15170=>"011000100",
  15171=>"111011111",
  15172=>"001000100",
  15173=>"010101100",
  15174=>"110011110",
  15175=>"111010100",
  15176=>"011101101",
  15177=>"111111011",
  15178=>"101001001",
  15179=>"001001101",
  15180=>"011101100",
  15181=>"100101011",
  15182=>"010110001",
  15183=>"011100001",
  15184=>"100000010",
  15185=>"100101101",
  15186=>"000000100",
  15187=>"000000101",
  15188=>"110010011",
  15189=>"001110111",
  15190=>"001100000",
  15191=>"111111001",
  15192=>"101000011",
  15193=>"011110110",
  15194=>"111001001",
  15195=>"111000011",
  15196=>"000010001",
  15197=>"001111101",
  15198=>"100101111",
  15199=>"000111001",
  15200=>"000010110",
  15201=>"100110110",
  15202=>"111000111",
  15203=>"111000101",
  15204=>"100000010",
  15205=>"000110101",
  15206=>"110110010",
  15207=>"111000000",
  15208=>"111100000",
  15209=>"110100001",
  15210=>"011110001",
  15211=>"001111111",
  15212=>"011000101",
  15213=>"101101001",
  15214=>"000001111",
  15215=>"010010101",
  15216=>"011101100",
  15217=>"011100000",
  15218=>"000011011",
  15219=>"101011101",
  15220=>"100011110",
  15221=>"011011011",
  15222=>"010111000",
  15223=>"000101000",
  15224=>"001000110",
  15225=>"010101111",
  15226=>"111110010",
  15227=>"011110001",
  15228=>"100000000",
  15229=>"001000111",
  15230=>"000000010",
  15231=>"000011111",
  15232=>"000110010",
  15233=>"010010101",
  15234=>"101101100",
  15235=>"111000011",
  15236=>"111000000",
  15237=>"110010101",
  15238=>"110000110",
  15239=>"111101001",
  15240=>"001000111",
  15241=>"001101100",
  15242=>"100001111",
  15243=>"010101011",
  15244=>"000001001",
  15245=>"110011101",
  15246=>"011101011",
  15247=>"111001110",
  15248=>"110000110",
  15249=>"000000001",
  15250=>"000011111",
  15251=>"110001010",
  15252=>"101001101",
  15253=>"110001110",
  15254=>"000000101",
  15255=>"010010010",
  15256=>"110110110",
  15257=>"011100010",
  15258=>"101001010",
  15259=>"010010101",
  15260=>"000100010",
  15261=>"110010001",
  15262=>"100001000",
  15263=>"111011101",
  15264=>"011111100",
  15265=>"100001000",
  15266=>"101001000",
  15267=>"010010100",
  15268=>"110111000",
  15269=>"001010110",
  15270=>"101001110",
  15271=>"011001101",
  15272=>"001011001",
  15273=>"000110000",
  15274=>"001100101",
  15275=>"001100010",
  15276=>"011101001",
  15277=>"111111100",
  15278=>"110011000",
  15279=>"111101101",
  15280=>"100011000",
  15281=>"011010001",
  15282=>"010001000",
  15283=>"000100000",
  15284=>"111011111",
  15285=>"001100011",
  15286=>"011010000",
  15287=>"111100110",
  15288=>"011110111",
  15289=>"010011010",
  15290=>"000011010",
  15291=>"011011010",
  15292=>"010011001",
  15293=>"101001011",
  15294=>"001000110",
  15295=>"100011110",
  15296=>"011100111",
  15297=>"001101110",
  15298=>"101100101",
  15299=>"110010011",
  15300=>"101001001",
  15301=>"110000000",
  15302=>"001111100",
  15303=>"010100000",
  15304=>"011000111",
  15305=>"011111001",
  15306=>"000001011",
  15307=>"100011100",
  15308=>"110001111",
  15309=>"111010110",
  15310=>"111111110",
  15311=>"100001010",
  15312=>"111000111",
  15313=>"011100100",
  15314=>"000011011",
  15315=>"000011000",
  15316=>"101100000",
  15317=>"101110001",
  15318=>"111101011",
  15319=>"001001111",
  15320=>"110111100",
  15321=>"101100111",
  15322=>"100001001",
  15323=>"001000001",
  15324=>"010010101",
  15325=>"010101011",
  15326=>"111111100",
  15327=>"001101010",
  15328=>"111101110",
  15329=>"101101011",
  15330=>"011110010",
  15331=>"110001111",
  15332=>"011000000",
  15333=>"110011100",
  15334=>"111010111",
  15335=>"111100111",
  15336=>"011101100",
  15337=>"010011000",
  15338=>"010111001",
  15339=>"110000011",
  15340=>"111011011",
  15341=>"000000011",
  15342=>"011001001",
  15343=>"101101000",
  15344=>"010010000",
  15345=>"010010100",
  15346=>"001001010",
  15347=>"100100101",
  15348=>"110111111",
  15349=>"011100000",
  15350=>"100100111",
  15351=>"000111011",
  15352=>"111110110",
  15353=>"000011101",
  15354=>"101101101",
  15355=>"100100001",
  15356=>"010010101",
  15357=>"100101010",
  15358=>"111000100",
  15359=>"111111011",
  15360=>"101101001",
  15361=>"101010101",
  15362=>"010110000",
  15363=>"111010110",
  15364=>"110111011",
  15365=>"111111100",
  15366=>"010000000",
  15367=>"010001110",
  15368=>"001011010",
  15369=>"101100001",
  15370=>"010111101",
  15371=>"101110000",
  15372=>"011001100",
  15373=>"011010000",
  15374=>"001101101",
  15375=>"000001100",
  15376=>"001010110",
  15377=>"001110000",
  15378=>"001001001",
  15379=>"010000110",
  15380=>"101010100",
  15381=>"001011011",
  15382=>"111101000",
  15383=>"010010011",
  15384=>"111010101",
  15385=>"010011000",
  15386=>"001011111",
  15387=>"101001101",
  15388=>"101010010",
  15389=>"101001111",
  15390=>"000011101",
  15391=>"000100010",
  15392=>"111000011",
  15393=>"000010110",
  15394=>"010010000",
  15395=>"010001000",
  15396=>"001100100",
  15397=>"110001111",
  15398=>"100101110",
  15399=>"110011011",
  15400=>"000000000",
  15401=>"010111101",
  15402=>"100111001",
  15403=>"100110111",
  15404=>"101001010",
  15405=>"110100010",
  15406=>"010100110",
  15407=>"101011001",
  15408=>"101011101",
  15409=>"011010111",
  15410=>"000011010",
  15411=>"111111001",
  15412=>"000001010",
  15413=>"111010000",
  15414=>"011111011",
  15415=>"111100111",
  15416=>"001000000",
  15417=>"000001000",
  15418=>"000100010",
  15419=>"110111111",
  15420=>"010000010",
  15421=>"100001111",
  15422=>"001000011",
  15423=>"101101101",
  15424=>"101001110",
  15425=>"000010110",
  15426=>"001011101",
  15427=>"011000011",
  15428=>"001010000",
  15429=>"000011010",
  15430=>"011100110",
  15431=>"011010000",
  15432=>"010001100",
  15433=>"011110111",
  15434=>"000010000",
  15435=>"111111101",
  15436=>"011100000",
  15437=>"111010101",
  15438=>"001101101",
  15439=>"111001001",
  15440=>"100101100",
  15441=>"111110100",
  15442=>"011100011",
  15443=>"011110100",
  15444=>"000110000",
  15445=>"111010101",
  15446=>"010110011",
  15447=>"010010110",
  15448=>"100111000",
  15449=>"001101101",
  15450=>"001110000",
  15451=>"001001111",
  15452=>"111111100",
  15453=>"000001101",
  15454=>"100100010",
  15455=>"000101101",
  15456=>"101000111",
  15457=>"001001010",
  15458=>"000110111",
  15459=>"010001111",
  15460=>"001110010",
  15461=>"110101110",
  15462=>"010001000",
  15463=>"101111100",
  15464=>"100111010",
  15465=>"101001001",
  15466=>"110010110",
  15467=>"101111110",
  15468=>"000100111",
  15469=>"011010011",
  15470=>"110110000",
  15471=>"111101000",
  15472=>"111101000",
  15473=>"110110000",
  15474=>"010100101",
  15475=>"011111000",
  15476=>"000000001",
  15477=>"101111110",
  15478=>"000010101",
  15479=>"110101010",
  15480=>"110010000",
  15481=>"101100010",
  15482=>"000000111",
  15483=>"000011011",
  15484=>"111110111",
  15485=>"011100010",
  15486=>"000100100",
  15487=>"101001000",
  15488=>"101000011",
  15489=>"110110010",
  15490=>"010110011",
  15491=>"100111111",
  15492=>"010101001",
  15493=>"001100111",
  15494=>"101110110",
  15495=>"010001111",
  15496=>"010001111",
  15497=>"000001001",
  15498=>"001010010",
  15499=>"100110110",
  15500=>"011101110",
  15501=>"110111110",
  15502=>"011010101",
  15503=>"111001111",
  15504=>"011011111",
  15505=>"010100000",
  15506=>"100100010",
  15507=>"010001100",
  15508=>"000001011",
  15509=>"110100011",
  15510=>"000100000",
  15511=>"110101101",
  15512=>"000000100",
  15513=>"000100001",
  15514=>"011001010",
  15515=>"100000010",
  15516=>"000110011",
  15517=>"111011011",
  15518=>"101110010",
  15519=>"011100001",
  15520=>"100110100",
  15521=>"001000101",
  15522=>"001010101",
  15523=>"001100010",
  15524=>"110111101",
  15525=>"101100001",
  15526=>"101101100",
  15527=>"010001101",
  15528=>"011011001",
  15529=>"110100110",
  15530=>"001110000",
  15531=>"000110110",
  15532=>"101101000",
  15533=>"111110001",
  15534=>"011111011",
  15535=>"011101001",
  15536=>"000011110",
  15537=>"111101111",
  15538=>"010111000",
  15539=>"100101100",
  15540=>"101100011",
  15541=>"111010011",
  15542=>"100010000",
  15543=>"011111011",
  15544=>"001010000",
  15545=>"101100101",
  15546=>"000011111",
  15547=>"011011001",
  15548=>"011011001",
  15549=>"010010100",
  15550=>"100110010",
  15551=>"010101010",
  15552=>"011000010",
  15553=>"110111000",
  15554=>"011111001",
  15555=>"110110011",
  15556=>"001010111",
  15557=>"010001010",
  15558=>"011001110",
  15559=>"101101011",
  15560=>"010100110",
  15561=>"100011111",
  15562=>"001101010",
  15563=>"110011111",
  15564=>"011101001",
  15565=>"000111101",
  15566=>"111101111",
  15567=>"100101000",
  15568=>"011111111",
  15569=>"100111111",
  15570=>"110000010",
  15571=>"000000101",
  15572=>"100101100",
  15573=>"001000100",
  15574=>"010010111",
  15575=>"111111000",
  15576=>"110000101",
  15577=>"000001000",
  15578=>"110011111",
  15579=>"101101100",
  15580=>"011011101",
  15581=>"001110100",
  15582=>"010111100",
  15583=>"100110000",
  15584=>"010000110",
  15585=>"111101110",
  15586=>"010101001",
  15587=>"110110000",
  15588=>"011110100",
  15589=>"000001110",
  15590=>"010000010",
  15591=>"000110010",
  15592=>"000000011",
  15593=>"011110000",
  15594=>"011110101",
  15595=>"010100010",
  15596=>"101110101",
  15597=>"000101011",
  15598=>"111000101",
  15599=>"000100000",
  15600=>"110010011",
  15601=>"000011101",
  15602=>"110001101",
  15603=>"110110100",
  15604=>"011100011",
  15605=>"101111110",
  15606=>"100111000",
  15607=>"011011000",
  15608=>"001111101",
  15609=>"000110100",
  15610=>"110011000",
  15611=>"000101001",
  15612=>"001100101",
  15613=>"000101101",
  15614=>"011110101",
  15615=>"010010011",
  15616=>"001110000",
  15617=>"101001001",
  15618=>"101101110",
  15619=>"111110111",
  15620=>"110010101",
  15621=>"101111010",
  15622=>"001000011",
  15623=>"001100001",
  15624=>"101011100",
  15625=>"011110001",
  15626=>"101110100",
  15627=>"010000001",
  15628=>"100110110",
  15629=>"000110111",
  15630=>"010101001",
  15631=>"101110111",
  15632=>"101100000",
  15633=>"100111000",
  15634=>"100101111",
  15635=>"100101100",
  15636=>"001001011",
  15637=>"110111111",
  15638=>"100011011",
  15639=>"000011101",
  15640=>"110001010",
  15641=>"011110011",
  15642=>"100101111",
  15643=>"011100110",
  15644=>"100001011",
  15645=>"000011000",
  15646=>"001100111",
  15647=>"100000111",
  15648=>"011101011",
  15649=>"000010010",
  15650=>"100100000",
  15651=>"000100100",
  15652=>"110101111",
  15653=>"100010000",
  15654=>"111111111",
  15655=>"011100101",
  15656=>"110010010",
  15657=>"101010010",
  15658=>"001001000",
  15659=>"100101001",
  15660=>"110000110",
  15661=>"001000001",
  15662=>"001000110",
  15663=>"101001110",
  15664=>"111110100",
  15665=>"101000010",
  15666=>"111011111",
  15667=>"001000000",
  15668=>"000001001",
  15669=>"010110011",
  15670=>"110101001",
  15671=>"000010101",
  15672=>"101111011",
  15673=>"101001111",
  15674=>"000011100",
  15675=>"001100110",
  15676=>"000000001",
  15677=>"111001011",
  15678=>"011100010",
  15679=>"011100110",
  15680=>"111100010",
  15681=>"000100110",
  15682=>"111000111",
  15683=>"110011100",
  15684=>"110011110",
  15685=>"111001000",
  15686=>"101001000",
  15687=>"111111001",
  15688=>"100111110",
  15689=>"101100011",
  15690=>"101011011",
  15691=>"110000101",
  15692=>"101011111",
  15693=>"010010000",
  15694=>"011100111",
  15695=>"011001101",
  15696=>"100100110",
  15697=>"001110101",
  15698=>"100000000",
  15699=>"111111111",
  15700=>"000011100",
  15701=>"000101100",
  15702=>"100101110",
  15703=>"010111001",
  15704=>"101110000",
  15705=>"110101010",
  15706=>"011001011",
  15707=>"001010110",
  15708=>"011011110",
  15709=>"001111101",
  15710=>"011101100",
  15711=>"100000000",
  15712=>"001000010",
  15713=>"000010100",
  15714=>"010111000",
  15715=>"001000011",
  15716=>"001100101",
  15717=>"101111111",
  15718=>"111111000",
  15719=>"100100011",
  15720=>"110010101",
  15721=>"110000000",
  15722=>"110011001",
  15723=>"101110010",
  15724=>"010011011",
  15725=>"101000000",
  15726=>"011011100",
  15727=>"010010000",
  15728=>"111101101",
  15729=>"011010100",
  15730=>"011111001",
  15731=>"101110001",
  15732=>"101001011",
  15733=>"111101001",
  15734=>"001000011",
  15735=>"000100111",
  15736=>"010011011",
  15737=>"101010110",
  15738=>"011100000",
  15739=>"001110110",
  15740=>"010010011",
  15741=>"011111111",
  15742=>"110100011",
  15743=>"011001000",
  15744=>"100111001",
  15745=>"111100000",
  15746=>"100011001",
  15747=>"010111101",
  15748=>"101101100",
  15749=>"010001100",
  15750=>"111011100",
  15751=>"010011010",
  15752=>"110100011",
  15753=>"001111100",
  15754=>"011001100",
  15755=>"110011010",
  15756=>"011010001",
  15757=>"010110001",
  15758=>"011001001",
  15759=>"010011000",
  15760=>"001011010",
  15761=>"000110110",
  15762=>"000010101",
  15763=>"101000001",
  15764=>"011000011",
  15765=>"010100010",
  15766=>"010001001",
  15767=>"000000000",
  15768=>"000101100",
  15769=>"011110011",
  15770=>"001010100",
  15771=>"101001111",
  15772=>"011000000",
  15773=>"101011101",
  15774=>"000100001",
  15775=>"100010001",
  15776=>"100100000",
  15777=>"001111101",
  15778=>"010111000",
  15779=>"000010100",
  15780=>"011001000",
  15781=>"001001100",
  15782=>"011010111",
  15783=>"110011001",
  15784=>"000100111",
  15785=>"010100100",
  15786=>"001010111",
  15787=>"001010011",
  15788=>"101111001",
  15789=>"001111001",
  15790=>"011000001",
  15791=>"110000101",
  15792=>"000110111",
  15793=>"100100000",
  15794=>"011000000",
  15795=>"111011101",
  15796=>"101111010",
  15797=>"011100000",
  15798=>"100011000",
  15799=>"000110010",
  15800=>"010101010",
  15801=>"111001110",
  15802=>"111110101",
  15803=>"101110110",
  15804=>"111011110",
  15805=>"100111101",
  15806=>"100111011",
  15807=>"111101000",
  15808=>"101010001",
  15809=>"000100100",
  15810=>"010101000",
  15811=>"010000000",
  15812=>"001000001",
  15813=>"100011000",
  15814=>"110011010",
  15815=>"111100101",
  15816=>"100011100",
  15817=>"000100011",
  15818=>"111001101",
  15819=>"111000100",
  15820=>"010010110",
  15821=>"011110010",
  15822=>"010101110",
  15823=>"100000001",
  15824=>"101100101",
  15825=>"001010110",
  15826=>"100101000",
  15827=>"110100010",
  15828=>"010101111",
  15829=>"110011011",
  15830=>"100011001",
  15831=>"101100000",
  15832=>"011100011",
  15833=>"101001100",
  15834=>"000011111",
  15835=>"010100101",
  15836=>"100111011",
  15837=>"101000011",
  15838=>"001000001",
  15839=>"010101011",
  15840=>"000000001",
  15841=>"000001000",
  15842=>"101011111",
  15843=>"111111100",
  15844=>"010000001",
  15845=>"110011101",
  15846=>"011011101",
  15847=>"110100100",
  15848=>"111000000",
  15849=>"000010111",
  15850=>"111000101",
  15851=>"000100010",
  15852=>"101110011",
  15853=>"000011001",
  15854=>"000111011",
  15855=>"011111110",
  15856=>"110101101",
  15857=>"011100110",
  15858=>"011011110",
  15859=>"000101011",
  15860=>"010001111",
  15861=>"000010111",
  15862=>"110001001",
  15863=>"101110111",
  15864=>"011010010",
  15865=>"110111011",
  15866=>"011010000",
  15867=>"110101010",
  15868=>"111011000",
  15869=>"101111110",
  15870=>"011010001",
  15871=>"010001010",
  15872=>"110000100",
  15873=>"010110111",
  15874=>"000110011",
  15875=>"010011010",
  15876=>"111000111",
  15877=>"101111000",
  15878=>"000101111",
  15879=>"100000100",
  15880=>"110010101",
  15881=>"101000000",
  15882=>"000100100",
  15883=>"111111111",
  15884=>"011011010",
  15885=>"011101100",
  15886=>"000110001",
  15887=>"101100100",
  15888=>"010110010",
  15889=>"001000111",
  15890=>"001111000",
  15891=>"101010010",
  15892=>"011100011",
  15893=>"111111010",
  15894=>"011000001",
  15895=>"111100010",
  15896=>"100111110",
  15897=>"010111000",
  15898=>"111100000",
  15899=>"010100011",
  15900=>"110010100",
  15901=>"110111001",
  15902=>"000010011",
  15903=>"111100101",
  15904=>"000010011",
  15905=>"010100000",
  15906=>"111000101",
  15907=>"010101001",
  15908=>"000010010",
  15909=>"111011011",
  15910=>"110010111",
  15911=>"000000101",
  15912=>"100000011",
  15913=>"111000110",
  15914=>"000010000",
  15915=>"111110111",
  15916=>"010111001",
  15917=>"100001001",
  15918=>"010101111",
  15919=>"101101110",
  15920=>"000000101",
  15921=>"110101111",
  15922=>"110000110",
  15923=>"010001000",
  15924=>"101010000",
  15925=>"100101110",
  15926=>"110011011",
  15927=>"001010111",
  15928=>"101001010",
  15929=>"001010011",
  15930=>"101000011",
  15931=>"011010110",
  15932=>"101101101",
  15933=>"100100111",
  15934=>"111000000",
  15935=>"011110000",
  15936=>"011110000",
  15937=>"010000010",
  15938=>"111011000",
  15939=>"000101000",
  15940=>"111110001",
  15941=>"001110000",
  15942=>"110101000",
  15943=>"011100011",
  15944=>"100110100",
  15945=>"110100100",
  15946=>"101010101",
  15947=>"111101100",
  15948=>"111100000",
  15949=>"001111010",
  15950=>"101100111",
  15951=>"011111101",
  15952=>"000010111",
  15953=>"001111110",
  15954=>"111001000",
  15955=>"000011001",
  15956=>"110100110",
  15957=>"110001100",
  15958=>"100111010",
  15959=>"010101011",
  15960=>"111100111",
  15961=>"101011011",
  15962=>"011001100",
  15963=>"000010100",
  15964=>"111011001",
  15965=>"010100011",
  15966=>"000011101",
  15967=>"010000000",
  15968=>"111111000",
  15969=>"001111110",
  15970=>"000100011",
  15971=>"001100111",
  15972=>"011000000",
  15973=>"000111011",
  15974=>"011101101",
  15975=>"011101111",
  15976=>"111101110",
  15977=>"001001101",
  15978=>"110111010",
  15979=>"111010001",
  15980=>"101111111",
  15981=>"001011000",
  15982=>"011000110",
  15983=>"100110111",
  15984=>"000000001",
  15985=>"000111110",
  15986=>"010000100",
  15987=>"111101100",
  15988=>"000010011",
  15989=>"011111101",
  15990=>"110011101",
  15991=>"100110100",
  15992=>"110111001",
  15993=>"111111110",
  15994=>"111101101",
  15995=>"001111100",
  15996=>"001000110",
  15997=>"010110001",
  15998=>"100110100",
  15999=>"110001111",
  16000=>"001111000",
  16001=>"011101000",
  16002=>"011101110",
  16003=>"001000011",
  16004=>"100111101",
  16005=>"100101000",
  16006=>"111000110",
  16007=>"110110011",
  16008=>"111011100",
  16009=>"000100001",
  16010=>"101000101",
  16011=>"001000101",
  16012=>"110000101",
  16013=>"010010111",
  16014=>"000111111",
  16015=>"110100110",
  16016=>"011100101",
  16017=>"001101001",
  16018=>"110010010",
  16019=>"110010110",
  16020=>"011111000",
  16021=>"011111010",
  16022=>"011101000",
  16023=>"011111110",
  16024=>"111110011",
  16025=>"011000010",
  16026=>"110000110",
  16027=>"010101001",
  16028=>"101111001",
  16029=>"011110010",
  16030=>"111110100",
  16031=>"110100000",
  16032=>"110100111",
  16033=>"010101101",
  16034=>"100001110",
  16035=>"000010001",
  16036=>"100011000",
  16037=>"101011101",
  16038=>"001001101",
  16039=>"110011010",
  16040=>"001011111",
  16041=>"111100011",
  16042=>"010100001",
  16043=>"000100010",
  16044=>"100110001",
  16045=>"010110010",
  16046=>"111111100",
  16047=>"001110110",
  16048=>"101001100",
  16049=>"010000100",
  16050=>"101001011",
  16051=>"000111101",
  16052=>"000101101",
  16053=>"000101011",
  16054=>"011000011",
  16055=>"000000010",
  16056=>"011010001",
  16057=>"110101001",
  16058=>"010111010",
  16059=>"001001011",
  16060=>"011011111",
  16061=>"010011110",
  16062=>"010000000",
  16063=>"011111010",
  16064=>"001011011",
  16065=>"111001011",
  16066=>"000101110",
  16067=>"000101000",
  16068=>"101100000",
  16069=>"101101100",
  16070=>"011101001",
  16071=>"010101011",
  16072=>"010010010",
  16073=>"000010110",
  16074=>"100100110",
  16075=>"110011101",
  16076=>"000101101",
  16077=>"000101111",
  16078=>"100110110",
  16079=>"110101111",
  16080=>"010011101",
  16081=>"010101111",
  16082=>"000000010",
  16083=>"111001110",
  16084=>"101010101",
  16085=>"010100000",
  16086=>"110111000",
  16087=>"001010100",
  16088=>"011101111",
  16089=>"001111100",
  16090=>"110010000",
  16091=>"011100100",
  16092=>"010001110",
  16093=>"111110111",
  16094=>"111001111",
  16095=>"101001001",
  16096=>"011011110",
  16097=>"101101001",
  16098=>"001100100",
  16099=>"010010001",
  16100=>"001010011",
  16101=>"110100010",
  16102=>"011111001",
  16103=>"000001111",
  16104=>"010010000",
  16105=>"000110001",
  16106=>"101010010",
  16107=>"010100001",
  16108=>"010001110",
  16109=>"111111100",
  16110=>"010111110",
  16111=>"100110100",
  16112=>"011011001",
  16113=>"000111101",
  16114=>"000000110",
  16115=>"110000010",
  16116=>"011110001",
  16117=>"100010110",
  16118=>"100101000",
  16119=>"111111111",
  16120=>"010010010",
  16121=>"110100101",
  16122=>"110000111",
  16123=>"111011100",
  16124=>"110101110",
  16125=>"111111110",
  16126=>"100100110",
  16127=>"001000110",
  16128=>"110111111",
  16129=>"100010011",
  16130=>"001101011",
  16131=>"100100100",
  16132=>"111001000",
  16133=>"100100000",
  16134=>"000001101",
  16135=>"101100001",
  16136=>"111010111",
  16137=>"001000011",
  16138=>"110001101",
  16139=>"010010001",
  16140=>"110100010",
  16141=>"101110101",
  16142=>"100000110",
  16143=>"100100010",
  16144=>"111111111",
  16145=>"100101111",
  16146=>"101100100",
  16147=>"100000111",
  16148=>"000100001",
  16149=>"100000011",
  16150=>"010110101",
  16151=>"110010111",
  16152=>"001101111",
  16153=>"111000001",
  16154=>"001000011",
  16155=>"111111100",
  16156=>"111101101",
  16157=>"010100111",
  16158=>"011010001",
  16159=>"001001111",
  16160=>"100011001",
  16161=>"101111110",
  16162=>"100101101",
  16163=>"000011000",
  16164=>"000001000",
  16165=>"111111111",
  16166=>"110001100",
  16167=>"110000111",
  16168=>"101011100",
  16169=>"010100000",
  16170=>"101010101",
  16171=>"010011110",
  16172=>"110110010",
  16173=>"000011101",
  16174=>"011101000",
  16175=>"000011100",
  16176=>"100000100",
  16177=>"010100100",
  16178=>"010010000",
  16179=>"111110110",
  16180=>"100110111",
  16181=>"101001100",
  16182=>"011101000",
  16183=>"010100000",
  16184=>"001100100",
  16185=>"001111110",
  16186=>"000111110",
  16187=>"010010010",
  16188=>"001111001",
  16189=>"111110101",
  16190=>"000001111",
  16191=>"010101111",
  16192=>"100101111",
  16193=>"000100001",
  16194=>"000110000",
  16195=>"111110100",
  16196=>"001000000",
  16197=>"000011110",
  16198=>"111010011",
  16199=>"011110001",
  16200=>"101111001",
  16201=>"010011110",
  16202=>"111111111",
  16203=>"111010001",
  16204=>"111011000",
  16205=>"000101111",
  16206=>"110110101",
  16207=>"110101000",
  16208=>"011111101",
  16209=>"000000111",
  16210=>"111000010",
  16211=>"001110000",
  16212=>"111001000",
  16213=>"100011011",
  16214=>"001100101",
  16215=>"010101011",
  16216=>"000010010",
  16217=>"101111110",
  16218=>"000001010",
  16219=>"011011010",
  16220=>"101001100",
  16221=>"011010010",
  16222=>"010111001",
  16223=>"111111110",
  16224=>"010011011",
  16225=>"001111100",
  16226=>"110000101",
  16227=>"111010001",
  16228=>"000110101",
  16229=>"000111100",
  16230=>"100110110",
  16231=>"000101100",
  16232=>"111001011",
  16233=>"101001011",
  16234=>"111111010",
  16235=>"010111011",
  16236=>"010110111",
  16237=>"011110000",
  16238=>"111111100",
  16239=>"000110110",
  16240=>"000100000",
  16241=>"110001101",
  16242=>"001110000",
  16243=>"001101101",
  16244=>"010011111",
  16245=>"111111111",
  16246=>"110100011",
  16247=>"010101011",
  16248=>"111110001",
  16249=>"001101011",
  16250=>"000100000",
  16251=>"000101000",
  16252=>"110011001",
  16253=>"111011110",
  16254=>"000101111",
  16255=>"000110100",
  16256=>"111001011",
  16257=>"100111011",
  16258=>"000110100",
  16259=>"000011000",
  16260=>"100100000",
  16261=>"100011110",
  16262=>"001100010",
  16263=>"110111111",
  16264=>"110100000",
  16265=>"000000011",
  16266=>"000000110",
  16267=>"011000101",
  16268=>"010110001",
  16269=>"111011001",
  16270=>"111101011",
  16271=>"000111111",
  16272=>"010101001",
  16273=>"011001100",
  16274=>"111011000",
  16275=>"000001001",
  16276=>"110001000",
  16277=>"110100100",
  16278=>"101110111",
  16279=>"011011001",
  16280=>"010000000",
  16281=>"000101010",
  16282=>"001110100",
  16283=>"000011010",
  16284=>"001001101",
  16285=>"000011001",
  16286=>"111100101",
  16287=>"011001110",
  16288=>"010011010",
  16289=>"110101000",
  16290=>"010000010",
  16291=>"101000000",
  16292=>"001000001",
  16293=>"001011000",
  16294=>"111111111",
  16295=>"001101011",
  16296=>"110110100",
  16297=>"000100000",
  16298=>"000011100",
  16299=>"001000010",
  16300=>"111000101",
  16301=>"111100111",
  16302=>"101010100",
  16303=>"010111010",
  16304=>"100010001",
  16305=>"000011101",
  16306=>"101011000",
  16307=>"011110000",
  16308=>"101110100",
  16309=>"000110100",
  16310=>"011001010",
  16311=>"001011011",
  16312=>"101111011",
  16313=>"000101111",
  16314=>"011101010",
  16315=>"011111101",
  16316=>"100100111",
  16317=>"010010000",
  16318=>"011111010",
  16319=>"011100010",
  16320=>"000010010",
  16321=>"110111101",
  16322=>"111010110",
  16323=>"001000000",
  16324=>"010001100",
  16325=>"001010100",
  16326=>"101100110",
  16327=>"001100110",
  16328=>"111001001",
  16329=>"011001000",
  16330=>"001111011",
  16331=>"001100001",
  16332=>"001111100",
  16333=>"001110011",
  16334=>"111101011",
  16335=>"100001101",
  16336=>"111000100",
  16337=>"111001111",
  16338=>"011100100",
  16339=>"001101000",
  16340=>"111110101",
  16341=>"010000010",
  16342=>"001110110",
  16343=>"010010111",
  16344=>"100001010",
  16345=>"011100000",
  16346=>"110000100",
  16347=>"111111110",
  16348=>"100101000",
  16349=>"100011011",
  16350=>"100010111",
  16351=>"000010010",
  16352=>"000001001",
  16353=>"011000011",
  16354=>"111011111",
  16355=>"110101101",
  16356=>"010000001",
  16357=>"000010011",
  16358=>"011100110",
  16359=>"010100110",
  16360=>"110010110",
  16361=>"001110001",
  16362=>"010000101",
  16363=>"010011001",
  16364=>"111010010",
  16365=>"010000011",
  16366=>"000001001",
  16367=>"100101001",
  16368=>"010000000",
  16369=>"111100000",
  16370=>"010011101",
  16371=>"000110001",
  16372=>"000100111",
  16373=>"100111000",
  16374=>"100110010",
  16375=>"010001111",
  16376=>"100011100",
  16377=>"111000000",
  16378=>"001011011",
  16379=>"101111001",
  16380=>"100111010",
  16381=>"101010111",
  16382=>"111011010",
  16383=>"111111100",
  16384=>"110011001",
  16385=>"111001010",
  16386=>"111011101",
  16387=>"101111000",
  16388=>"101110000",
  16389=>"100101100",
  16390=>"001111111",
  16391=>"110111000",
  16392=>"111010001",
  16393=>"001111010",
  16394=>"010001011",
  16395=>"100000111",
  16396=>"101000111",
  16397=>"100001001",
  16398=>"011110111",
  16399=>"100001111",
  16400=>"101101111",
  16401=>"111010001",
  16402=>"001001011",
  16403=>"100111001",
  16404=>"011100111",
  16405=>"000010011",
  16406=>"101011010",
  16407=>"100100000",
  16408=>"001101000",
  16409=>"101011101",
  16410=>"000000000",
  16411=>"100010111",
  16412=>"010001011",
  16413=>"001110010",
  16414=>"110101000",
  16415=>"111010101",
  16416=>"000011010",
  16417=>"010011010",
  16418=>"000011111",
  16419=>"001110001",
  16420=>"001001110",
  16421=>"000100100",
  16422=>"101100101",
  16423=>"101100010",
  16424=>"100000010",
  16425=>"011111001",
  16426=>"111000001",
  16427=>"000011000",
  16428=>"001111010",
  16429=>"101110001",
  16430=>"111100100",
  16431=>"100110100",
  16432=>"111000111",
  16433=>"101111011",
  16434=>"100101001",
  16435=>"101111110",
  16436=>"111111111",
  16437=>"000011011",
  16438=>"110100100",
  16439=>"110110000",
  16440=>"000011010",
  16441=>"101100000",
  16442=>"101101110",
  16443=>"101000001",
  16444=>"110011111",
  16445=>"010100010",
  16446=>"000101010",
  16447=>"101101001",
  16448=>"001100000",
  16449=>"010111000",
  16450=>"111011000",
  16451=>"000010111",
  16452=>"100000000",
  16453=>"011011011",
  16454=>"011010000",
  16455=>"001010110",
  16456=>"000101001",
  16457=>"000010010",
  16458=>"011000001",
  16459=>"001101000",
  16460=>"110110000",
  16461=>"100110100",
  16462=>"110100010",
  16463=>"001010111",
  16464=>"101010100",
  16465=>"110010111",
  16466=>"110110000",
  16467=>"000010001",
  16468=>"000010111",
  16469=>"000010110",
  16470=>"011101101",
  16471=>"101001111",
  16472=>"111101010",
  16473=>"011111001",
  16474=>"101011000",
  16475=>"000100110",
  16476=>"010111000",
  16477=>"100001011",
  16478=>"100000100",
  16479=>"110001010",
  16480=>"100001111",
  16481=>"110110101",
  16482=>"010100010",
  16483=>"110010011",
  16484=>"011100110",
  16485=>"010111100",
  16486=>"000101111",
  16487=>"100000011",
  16488=>"111110101",
  16489=>"101010000",
  16490=>"111110010",
  16491=>"100011100",
  16492=>"011100111",
  16493=>"111001010",
  16494=>"000010101",
  16495=>"100011000",
  16496=>"011010011",
  16497=>"011101111",
  16498=>"000000111",
  16499=>"011101000",
  16500=>"010010100",
  16501=>"000000000",
  16502=>"101000110",
  16503=>"000110110",
  16504=>"011010101",
  16505=>"110100011",
  16506=>"100110010",
  16507=>"001110010",
  16508=>"000000000",
  16509=>"011100000",
  16510=>"110101000",
  16511=>"110111000",
  16512=>"000110110",
  16513=>"011010010",
  16514=>"000101010",
  16515=>"000010110",
  16516=>"001101000",
  16517=>"011000010",
  16518=>"000100000",
  16519=>"001001011",
  16520=>"010110100",
  16521=>"110100010",
  16522=>"101110000",
  16523=>"010111111",
  16524=>"111001101",
  16525=>"111001111",
  16526=>"000111111",
  16527=>"011001100",
  16528=>"111110110",
  16529=>"110010001",
  16530=>"010111010",
  16531=>"011001110",
  16532=>"111000010",
  16533=>"100001101",
  16534=>"111111000",
  16535=>"010010010",
  16536=>"000110000",
  16537=>"110100000",
  16538=>"010010010",
  16539=>"010000001",
  16540=>"100001110",
  16541=>"000000100",
  16542=>"111000001",
  16543=>"011001011",
  16544=>"000010001",
  16545=>"111110101",
  16546=>"001111110",
  16547=>"011010111",
  16548=>"000110110",
  16549=>"000100111",
  16550=>"010010010",
  16551=>"101001000",
  16552=>"010010110",
  16553=>"000101010",
  16554=>"010001011",
  16555=>"001111101",
  16556=>"000101100",
  16557=>"101011110",
  16558=>"011000011",
  16559=>"110111000",
  16560=>"100111010",
  16561=>"101111110",
  16562=>"111110000",
  16563=>"001001111",
  16564=>"000101111",
  16565=>"001101100",
  16566=>"001011011",
  16567=>"111000100",
  16568=>"110000001",
  16569=>"111010011",
  16570=>"101001111",
  16571=>"011001010",
  16572=>"110101111",
  16573=>"011000111",
  16574=>"111010001",
  16575=>"000001010",
  16576=>"001100111",
  16577=>"011101110",
  16578=>"001000001",
  16579=>"010000011",
  16580=>"111111111",
  16581=>"001111101",
  16582=>"010110100",
  16583=>"100111111",
  16584=>"001000111",
  16585=>"010011110",
  16586=>"111101011",
  16587=>"100100100",
  16588=>"100101110",
  16589=>"110111111",
  16590=>"001101000",
  16591=>"010010001",
  16592=>"001010011",
  16593=>"010100011",
  16594=>"111101000",
  16595=>"101100101",
  16596=>"000000010",
  16597=>"010010011",
  16598=>"110000000",
  16599=>"011111011",
  16600=>"101011010",
  16601=>"001100100",
  16602=>"010111011",
  16603=>"010001100",
  16604=>"010110010",
  16605=>"111110011",
  16606=>"100010000",
  16607=>"101111000",
  16608=>"010111000",
  16609=>"110110111",
  16610=>"100010010",
  16611=>"111111101",
  16612=>"101000010",
  16613=>"010000000",
  16614=>"100100011",
  16615=>"101000000",
  16616=>"110111100",
  16617=>"001110010",
  16618=>"100111101",
  16619=>"100101011",
  16620=>"111011111",
  16621=>"110000101",
  16622=>"110111111",
  16623=>"010100010",
  16624=>"101001000",
  16625=>"110010001",
  16626=>"110101010",
  16627=>"010001011",
  16628=>"101011011",
  16629=>"111001111",
  16630=>"100000011",
  16631=>"110010011",
  16632=>"101010000",
  16633=>"110100011",
  16634=>"010000111",
  16635=>"101101111",
  16636=>"111011100",
  16637=>"001010101",
  16638=>"101000011",
  16639=>"011101100",
  16640=>"000101011",
  16641=>"111010000",
  16642=>"010110111",
  16643=>"000011100",
  16644=>"110000101",
  16645=>"010011010",
  16646=>"110001011",
  16647=>"101011001",
  16648=>"101101111",
  16649=>"001101111",
  16650=>"010111101",
  16651=>"011000000",
  16652=>"010100011",
  16653=>"101111101",
  16654=>"111100000",
  16655=>"011101011",
  16656=>"111010101",
  16657=>"101011101",
  16658=>"110011001",
  16659=>"101110000",
  16660=>"000010010",
  16661=>"001101110",
  16662=>"110111000",
  16663=>"111001000",
  16664=>"010011010",
  16665=>"111100011",
  16666=>"100111011",
  16667=>"000100110",
  16668=>"111110111",
  16669=>"110110100",
  16670=>"000011100",
  16671=>"000011011",
  16672=>"000100011",
  16673=>"100100111",
  16674=>"111111101",
  16675=>"100011111",
  16676=>"100111100",
  16677=>"001011011",
  16678=>"001100010",
  16679=>"000100010",
  16680=>"100111111",
  16681=>"001001010",
  16682=>"111110100",
  16683=>"111100110",
  16684=>"100110010",
  16685=>"010000100",
  16686=>"000001011",
  16687=>"100101110",
  16688=>"100000001",
  16689=>"011001010",
  16690=>"111100101",
  16691=>"010011101",
  16692=>"110111110",
  16693=>"100101110",
  16694=>"010100000",
  16695=>"110110111",
  16696=>"101101101",
  16697=>"011100100",
  16698=>"001001111",
  16699=>"010111111",
  16700=>"111011000",
  16701=>"000111011",
  16702=>"111010110",
  16703=>"010011000",
  16704=>"000011100",
  16705=>"000100110",
  16706=>"101100100",
  16707=>"011000101",
  16708=>"000000101",
  16709=>"111110110",
  16710=>"001010001",
  16711=>"000000011",
  16712=>"110000011",
  16713=>"010111101",
  16714=>"001010001",
  16715=>"100101010",
  16716=>"010101010",
  16717=>"010111111",
  16718=>"101000000",
  16719=>"100110101",
  16720=>"011101100",
  16721=>"010111010",
  16722=>"000000110",
  16723=>"111111110",
  16724=>"000101001",
  16725=>"001010010",
  16726=>"101000111",
  16727=>"011000101",
  16728=>"111011101",
  16729=>"101001000",
  16730=>"010001101",
  16731=>"100111011",
  16732=>"010111011",
  16733=>"000001010",
  16734=>"101001101",
  16735=>"110110111",
  16736=>"111011000",
  16737=>"001011000",
  16738=>"000010001",
  16739=>"001000110",
  16740=>"000101101",
  16741=>"100100110",
  16742=>"101100001",
  16743=>"101110001",
  16744=>"011110101",
  16745=>"000000010",
  16746=>"111100101",
  16747=>"101000000",
  16748=>"001111110",
  16749=>"000110001",
  16750=>"111000001",
  16751=>"110011101",
  16752=>"101100111",
  16753=>"011000110",
  16754=>"011010011",
  16755=>"010000100",
  16756=>"000011111",
  16757=>"111010111",
  16758=>"000101100",
  16759=>"000001010",
  16760=>"111110010",
  16761=>"011110101",
  16762=>"100110111",
  16763=>"011110011",
  16764=>"111110111",
  16765=>"001000011",
  16766=>"110100011",
  16767=>"101001101",
  16768=>"000111101",
  16769=>"111100011",
  16770=>"010001011",
  16771=>"010110001",
  16772=>"000000110",
  16773=>"010101000",
  16774=>"100101101",
  16775=>"010010010",
  16776=>"111000011",
  16777=>"000110111",
  16778=>"011010000",
  16779=>"110000110",
  16780=>"010010001",
  16781=>"001011101",
  16782=>"001010011",
  16783=>"111000000",
  16784=>"011001101",
  16785=>"000100010",
  16786=>"010001000",
  16787=>"110010110",
  16788=>"010010101",
  16789=>"101011010",
  16790=>"000000101",
  16791=>"101011101",
  16792=>"011010101",
  16793=>"101100000",
  16794=>"000010010",
  16795=>"100000100",
  16796=>"100110001",
  16797=>"010100100",
  16798=>"011000110",
  16799=>"101010111",
  16800=>"001100000",
  16801=>"101000000",
  16802=>"111110011",
  16803=>"111111100",
  16804=>"100110001",
  16805=>"001111101",
  16806=>"111100000",
  16807=>"101100001",
  16808=>"010001010",
  16809=>"111111001",
  16810=>"000111110",
  16811=>"110100100",
  16812=>"100101110",
  16813=>"001011011",
  16814=>"111100110",
  16815=>"110000000",
  16816=>"101001100",
  16817=>"111100110",
  16818=>"000010001",
  16819=>"111011111",
  16820=>"010000110",
  16821=>"010011100",
  16822=>"011111010",
  16823=>"011011110",
  16824=>"110110101",
  16825=>"000101100",
  16826=>"000011010",
  16827=>"100100011",
  16828=>"000010010",
  16829=>"100110011",
  16830=>"111010011",
  16831=>"110011111",
  16832=>"010001010",
  16833=>"010010011",
  16834=>"100011111",
  16835=>"010000101",
  16836=>"010000010",
  16837=>"010100011",
  16838=>"011100011",
  16839=>"010000100",
  16840=>"101111100",
  16841=>"110111110",
  16842=>"011000000",
  16843=>"000111001",
  16844=>"010110101",
  16845=>"111100101",
  16846=>"000010101",
  16847=>"110010100",
  16848=>"100110110",
  16849=>"110111100",
  16850=>"011100100",
  16851=>"101111111",
  16852=>"101100010",
  16853=>"100010101",
  16854=>"001101011",
  16855=>"101010010",
  16856=>"010011110",
  16857=>"111001010",
  16858=>"011011111",
  16859=>"111001010",
  16860=>"100100110",
  16861=>"111101001",
  16862=>"001101001",
  16863=>"111100000",
  16864=>"010010000",
  16865=>"001011100",
  16866=>"011010100",
  16867=>"000111111",
  16868=>"110001110",
  16869=>"111111101",
  16870=>"000100011",
  16871=>"101111000",
  16872=>"111010010",
  16873=>"111001101",
  16874=>"100000010",
  16875=>"111111100",
  16876=>"001111010",
  16877=>"010111010",
  16878=>"110000001",
  16879=>"001100110",
  16880=>"001000100",
  16881=>"100000110",
  16882=>"111001000",
  16883=>"110110101",
  16884=>"101010111",
  16885=>"111000001",
  16886=>"010001000",
  16887=>"110101000",
  16888=>"101001101",
  16889=>"110111101",
  16890=>"010110000",
  16891=>"010100000",
  16892=>"101101011",
  16893=>"011000000",
  16894=>"110111110",
  16895=>"000101001",
  16896=>"001101111",
  16897=>"000001010",
  16898=>"011010001",
  16899=>"001100010",
  16900=>"011011000",
  16901=>"101001111",
  16902=>"011001001",
  16903=>"011100101",
  16904=>"000000001",
  16905=>"100011110",
  16906=>"110100010",
  16907=>"010001010",
  16908=>"101001001",
  16909=>"010010111",
  16910=>"101100011",
  16911=>"111111011",
  16912=>"010100001",
  16913=>"101011100",
  16914=>"011011100",
  16915=>"111111111",
  16916=>"110101000",
  16917=>"001010011",
  16918=>"110101111",
  16919=>"010010100",
  16920=>"101110101",
  16921=>"001000000",
  16922=>"010101011",
  16923=>"011100100",
  16924=>"100100011",
  16925=>"111100001",
  16926=>"001111011",
  16927=>"100101001",
  16928=>"010100101",
  16929=>"001100111",
  16930=>"000001010",
  16931=>"100101000",
  16932=>"110100001",
  16933=>"011010000",
  16934=>"110000111",
  16935=>"010010100",
  16936=>"010101011",
  16937=>"111110100",
  16938=>"110111101",
  16939=>"011111111",
  16940=>"101111000",
  16941=>"101101111",
  16942=>"101111111",
  16943=>"010001110",
  16944=>"001010110",
  16945=>"110111100",
  16946=>"000001001",
  16947=>"011100110",
  16948=>"010001101",
  16949=>"110101001",
  16950=>"110111010",
  16951=>"111111110",
  16952=>"111010110",
  16953=>"110110101",
  16954=>"111100110",
  16955=>"000111001",
  16956=>"011011100",
  16957=>"100110111",
  16958=>"000111001",
  16959=>"011011101",
  16960=>"001011111",
  16961=>"000011111",
  16962=>"010001001",
  16963=>"111001011",
  16964=>"111011101",
  16965=>"010000000",
  16966=>"001100110",
  16967=>"110111010",
  16968=>"000110010",
  16969=>"011001010",
  16970=>"100000001",
  16971=>"010011110",
  16972=>"010000000",
  16973=>"001000111",
  16974=>"110011101",
  16975=>"111011000",
  16976=>"001000010",
  16977=>"000101111",
  16978=>"101111011",
  16979=>"100001101",
  16980=>"001010110",
  16981=>"001000110",
  16982=>"101010000",
  16983=>"011110001",
  16984=>"100111110",
  16985=>"110111100",
  16986=>"111010111",
  16987=>"100111010",
  16988=>"111001010",
  16989=>"101000000",
  16990=>"101001111",
  16991=>"011010100",
  16992=>"000101011",
  16993=>"010010000",
  16994=>"010100000",
  16995=>"110001001",
  16996=>"100110010",
  16997=>"010101011",
  16998=>"000000000",
  16999=>"101101011",
  17000=>"000000000",
  17001=>"000001000",
  17002=>"000111001",
  17003=>"001001010",
  17004=>"001100001",
  17005=>"110111010",
  17006=>"110101000",
  17007=>"001101010",
  17008=>"010110110",
  17009=>"011011101",
  17010=>"010010100",
  17011=>"110101011",
  17012=>"110110111",
  17013=>"001000000",
  17014=>"101011011",
  17015=>"001110011",
  17016=>"011101100",
  17017=>"101101001",
  17018=>"100011110",
  17019=>"101110010",
  17020=>"110101001",
  17021=>"101010101",
  17022=>"000100010",
  17023=>"111000101",
  17024=>"110110100",
  17025=>"101001001",
  17026=>"001000101",
  17027=>"111111001",
  17028=>"111011111",
  17029=>"011011000",
  17030=>"000100111",
  17031=>"000000001",
  17032=>"000111011",
  17033=>"110010011",
  17034=>"111111010",
  17035=>"010110000",
  17036=>"100101100",
  17037=>"010111011",
  17038=>"000110100",
  17039=>"111110101",
  17040=>"100010101",
  17041=>"010101010",
  17042=>"110001010",
  17043=>"111010101",
  17044=>"001011111",
  17045=>"100010100",
  17046=>"000111110",
  17047=>"100011011",
  17048=>"100000110",
  17049=>"100011001",
  17050=>"101010100",
  17051=>"101010100",
  17052=>"110111010",
  17053=>"100010000",
  17054=>"010000101",
  17055=>"001111110",
  17056=>"100010010",
  17057=>"010100001",
  17058=>"100101011",
  17059=>"011110011",
  17060=>"011001111",
  17061=>"010010001",
  17062=>"101011010",
  17063=>"111011011",
  17064=>"111111110",
  17065=>"111000000",
  17066=>"111000100",
  17067=>"001100011",
  17068=>"010101011",
  17069=>"011011011",
  17070=>"111110110",
  17071=>"111001001",
  17072=>"001110010",
  17073=>"010101111",
  17074=>"110100100",
  17075=>"011001110",
  17076=>"100100010",
  17077=>"111111010",
  17078=>"000110100",
  17079=>"011101100",
  17080=>"001101111",
  17081=>"110111110",
  17082=>"100010011",
  17083=>"101001001",
  17084=>"011001111",
  17085=>"000010010",
  17086=>"111010100",
  17087=>"100010011",
  17088=>"011111011",
  17089=>"101111111",
  17090=>"000010000",
  17091=>"000001100",
  17092=>"100010110",
  17093=>"001110000",
  17094=>"100111100",
  17095=>"111100010",
  17096=>"101110101",
  17097=>"001010010",
  17098=>"010100010",
  17099=>"100110001",
  17100=>"100100110",
  17101=>"000011111",
  17102=>"111111010",
  17103=>"011000000",
  17104=>"110010000",
  17105=>"100011111",
  17106=>"000101111",
  17107=>"101000100",
  17108=>"001101011",
  17109=>"101001010",
  17110=>"010111101",
  17111=>"010101000",
  17112=>"101110100",
  17113=>"110111111",
  17114=>"101010101",
  17115=>"110111011",
  17116=>"001000000",
  17117=>"101010111",
  17118=>"011101010",
  17119=>"010100110",
  17120=>"001001000",
  17121=>"000101101",
  17122=>"011110101",
  17123=>"000000110",
  17124=>"010101101",
  17125=>"001011100",
  17126=>"000100011",
  17127=>"000010100",
  17128=>"000101110",
  17129=>"000101111",
  17130=>"000011011",
  17131=>"110011111",
  17132=>"000001001",
  17133=>"101000010",
  17134=>"100111011",
  17135=>"111111111",
  17136=>"010011100",
  17137=>"101001110",
  17138=>"101011100",
  17139=>"111100000",
  17140=>"100100010",
  17141=>"010111100",
  17142=>"110110101",
  17143=>"000000011",
  17144=>"101110001",
  17145=>"101111010",
  17146=>"101000000",
  17147=>"110101010",
  17148=>"100011010",
  17149=>"110100111",
  17150=>"100001001",
  17151=>"101010000",
  17152=>"101001010",
  17153=>"001000001",
  17154=>"011011001",
  17155=>"000010010",
  17156=>"000010010",
  17157=>"001111011",
  17158=>"000000010",
  17159=>"101000100",
  17160=>"110111010",
  17161=>"111101000",
  17162=>"001001001",
  17163=>"000111010",
  17164=>"001011001",
  17165=>"010111101",
  17166=>"101111111",
  17167=>"010111100",
  17168=>"111101111",
  17169=>"001100011",
  17170=>"010101001",
  17171=>"100010100",
  17172=>"000100000",
  17173=>"000010001",
  17174=>"001101100",
  17175=>"111010011",
  17176=>"000001100",
  17177=>"111010011",
  17178=>"000111111",
  17179=>"101010100",
  17180=>"011100010",
  17181=>"001101000",
  17182=>"011111111",
  17183=>"001100101",
  17184=>"110010011",
  17185=>"100110111",
  17186=>"111100101",
  17187=>"110101011",
  17188=>"101111110",
  17189=>"101110111",
  17190=>"000100010",
  17191=>"100110100",
  17192=>"101100000",
  17193=>"111001101",
  17194=>"101101011",
  17195=>"110101111",
  17196=>"010011010",
  17197=>"110100000",
  17198=>"000111010",
  17199=>"100101110",
  17200=>"111110101",
  17201=>"010000000",
  17202=>"011000000",
  17203=>"011000001",
  17204=>"000110110",
  17205=>"100001111",
  17206=>"001100001",
  17207=>"000011100",
  17208=>"111011010",
  17209=>"011111111",
  17210=>"100111010",
  17211=>"111101110",
  17212=>"010010101",
  17213=>"111010010",
  17214=>"110001100",
  17215=>"110110001",
  17216=>"011011111",
  17217=>"000101100",
  17218=>"001000010",
  17219=>"000100101",
  17220=>"001101000",
  17221=>"111110011",
  17222=>"111111111",
  17223=>"010110000",
  17224=>"010010001",
  17225=>"100010000",
  17226=>"101100100",
  17227=>"101000110",
  17228=>"000011010",
  17229=>"101100110",
  17230=>"010001010",
  17231=>"110000101",
  17232=>"011100101",
  17233=>"011000010",
  17234=>"000111011",
  17235=>"110000101",
  17236=>"111011000",
  17237=>"010100111",
  17238=>"101110101",
  17239=>"001111100",
  17240=>"001111100",
  17241=>"011100100",
  17242=>"111011011",
  17243=>"011000011",
  17244=>"110110010",
  17245=>"001001101",
  17246=>"111010001",
  17247=>"010000110",
  17248=>"111000110",
  17249=>"101101110",
  17250=>"011100111",
  17251=>"100110110",
  17252=>"110011101",
  17253=>"000000110",
  17254=>"001100100",
  17255=>"110010111",
  17256=>"100100010",
  17257=>"011111100",
  17258=>"100101111",
  17259=>"110111010",
  17260=>"110101110",
  17261=>"111110111",
  17262=>"010110000",
  17263=>"101001011",
  17264=>"101001011",
  17265=>"110011000",
  17266=>"011010011",
  17267=>"110111000",
  17268=>"011100000",
  17269=>"110110111",
  17270=>"001101000",
  17271=>"010001010",
  17272=>"100101111",
  17273=>"100000001",
  17274=>"100000110",
  17275=>"100110010",
  17276=>"001111100",
  17277=>"000001110",
  17278=>"100100100",
  17279=>"101001101",
  17280=>"100011011",
  17281=>"011000111",
  17282=>"111101010",
  17283=>"011010011",
  17284=>"001000110",
  17285=>"100010001",
  17286=>"001111010",
  17287=>"001101100",
  17288=>"101000100",
  17289=>"101100011",
  17290=>"101111110",
  17291=>"001011001",
  17292=>"010011100",
  17293=>"110010001",
  17294=>"011101100",
  17295=>"101100100",
  17296=>"101111010",
  17297=>"010011101",
  17298=>"100010111",
  17299=>"100100010",
  17300=>"111011111",
  17301=>"101000000",
  17302=>"110011110",
  17303=>"101111110",
  17304=>"011000000",
  17305=>"000100000",
  17306=>"011011011",
  17307=>"111001011",
  17308=>"000011101",
  17309=>"110110110",
  17310=>"101001000",
  17311=>"111100011",
  17312=>"010001101",
  17313=>"111111101",
  17314=>"111000001",
  17315=>"011001001",
  17316=>"010101001",
  17317=>"111000011",
  17318=>"110000000",
  17319=>"100000110",
  17320=>"101010101",
  17321=>"010000100",
  17322=>"000000111",
  17323=>"101011101",
  17324=>"000110001",
  17325=>"001001000",
  17326=>"101100000",
  17327=>"000000000",
  17328=>"101000000",
  17329=>"010110101",
  17330=>"001001100",
  17331=>"000001010",
  17332=>"101011010",
  17333=>"101000111",
  17334=>"110110000",
  17335=>"001010101",
  17336=>"010111110",
  17337=>"110101000",
  17338=>"111110000",
  17339=>"101000110",
  17340=>"010111100",
  17341=>"001110111",
  17342=>"100011000",
  17343=>"011000001",
  17344=>"000011110",
  17345=>"000100001",
  17346=>"111110100",
  17347=>"011010001",
  17348=>"110000011",
  17349=>"100010011",
  17350=>"110011000",
  17351=>"010100010",
  17352=>"000000010",
  17353=>"000011101",
  17354=>"001100101",
  17355=>"001001100",
  17356=>"111000011",
  17357=>"001100100",
  17358=>"011110000",
  17359=>"101000001",
  17360=>"001010101",
  17361=>"111001011",
  17362=>"000000000",
  17363=>"000011100",
  17364=>"011111101",
  17365=>"000101110",
  17366=>"000010111",
  17367=>"010110101",
  17368=>"011101000",
  17369=>"011111000",
  17370=>"111001010",
  17371=>"000010001",
  17372=>"001011101",
  17373=>"110110000",
  17374=>"010001111",
  17375=>"010110011",
  17376=>"010111001",
  17377=>"011010101",
  17378=>"110001011",
  17379=>"000000101",
  17380=>"000000100",
  17381=>"010100100",
  17382=>"000000011",
  17383=>"000000101",
  17384=>"111100010",
  17385=>"010101110",
  17386=>"000011011",
  17387=>"110000100",
  17388=>"001100111",
  17389=>"111111010",
  17390=>"100110101",
  17391=>"111111101",
  17392=>"101110111",
  17393=>"111111111",
  17394=>"000111110",
  17395=>"000100010",
  17396=>"111001010",
  17397=>"011011111",
  17398=>"111111110",
  17399=>"001011011",
  17400=>"000001010",
  17401=>"010001010",
  17402=>"110000010",
  17403=>"100010110",
  17404=>"010001111",
  17405=>"011101101",
  17406=>"111101101",
  17407=>"110000001",
  17408=>"010111111",
  17409=>"100111000",
  17410=>"100101011",
  17411=>"110111111",
  17412=>"110100110",
  17413=>"111110010",
  17414=>"111111111",
  17415=>"100001010",
  17416=>"111010110",
  17417=>"111001101",
  17418=>"010000011",
  17419=>"011111010",
  17420=>"100001100",
  17421=>"101010111",
  17422=>"101110000",
  17423=>"111011010",
  17424=>"011101011",
  17425=>"100101011",
  17426=>"110111010",
  17427=>"000111001",
  17428=>"101100010",
  17429=>"111101100",
  17430=>"100001110",
  17431=>"010111101",
  17432=>"100100101",
  17433=>"100011000",
  17434=>"010011111",
  17435=>"010101001",
  17436=>"001110111",
  17437=>"000100110",
  17438=>"110111110",
  17439=>"110110111",
  17440=>"111101010",
  17441=>"001110101",
  17442=>"011001100",
  17443=>"100100001",
  17444=>"000011001",
  17445=>"001010000",
  17446=>"101101010",
  17447=>"100101010",
  17448=>"110101000",
  17449=>"001001111",
  17450=>"101101110",
  17451=>"111111011",
  17452=>"101000001",
  17453=>"010101111",
  17454=>"111010100",
  17455=>"001101111",
  17456=>"111011111",
  17457=>"001000001",
  17458=>"100100101",
  17459=>"010011001",
  17460=>"100011000",
  17461=>"000001010",
  17462=>"110000110",
  17463=>"011011000",
  17464=>"000011111",
  17465=>"111100011",
  17466=>"000110011",
  17467=>"100000111",
  17468=>"001010111",
  17469=>"011000010",
  17470=>"011000011",
  17471=>"101111011",
  17472=>"111100000",
  17473=>"100111111",
  17474=>"001111000",
  17475=>"010000110",
  17476=>"110001000",
  17477=>"110111110",
  17478=>"011100011",
  17479=>"000110110",
  17480=>"001100010",
  17481=>"000111000",
  17482=>"000100010",
  17483=>"010101111",
  17484=>"111000101",
  17485=>"110111010",
  17486=>"100011111",
  17487=>"001001010",
  17488=>"000001011",
  17489=>"000001100",
  17490=>"100110011",
  17491=>"010001010",
  17492=>"000100110",
  17493=>"111001010",
  17494=>"000000011",
  17495=>"010010001",
  17496=>"101000100",
  17497=>"100110111",
  17498=>"100010001",
  17499=>"000001101",
  17500=>"101100100",
  17501=>"111110111",
  17502=>"011000001",
  17503=>"001111111",
  17504=>"000010001",
  17505=>"001000010",
  17506=>"010011010",
  17507=>"000101010",
  17508=>"111110001",
  17509=>"100100101",
  17510=>"011100001",
  17511=>"011100010",
  17512=>"100001101",
  17513=>"110011010",
  17514=>"100000111",
  17515=>"000011001",
  17516=>"111000110",
  17517=>"000101100",
  17518=>"110010100",
  17519=>"010001110",
  17520=>"110111011",
  17521=>"100111000",
  17522=>"011001100",
  17523=>"110100000",
  17524=>"101100100",
  17525=>"100100110",
  17526=>"000000101",
  17527=>"001101000",
  17528=>"110110011",
  17529=>"010010010",
  17530=>"101001110",
  17531=>"110110001",
  17532=>"010011101",
  17533=>"010101001",
  17534=>"101011010",
  17535=>"011000000",
  17536=>"010000100",
  17537=>"001001101",
  17538=>"111110010",
  17539=>"000111010",
  17540=>"111110111",
  17541=>"001011111",
  17542=>"111101111",
  17543=>"100001100",
  17544=>"000011001",
  17545=>"100001111",
  17546=>"111011111",
  17547=>"100000100",
  17548=>"011000010",
  17549=>"010111101",
  17550=>"001000001",
  17551=>"111000101",
  17552=>"111010010",
  17553=>"000111011",
  17554=>"111011000",
  17555=>"010010000",
  17556=>"100111000",
  17557=>"111101101",
  17558=>"001011000",
  17559=>"111001010",
  17560=>"100000110",
  17561=>"110001011",
  17562=>"101010110",
  17563=>"100001001",
  17564=>"011111011",
  17565=>"000111100",
  17566=>"100011111",
  17567=>"001000000",
  17568=>"100010111",
  17569=>"100010000",
  17570=>"000100010",
  17571=>"101110001",
  17572=>"010010000",
  17573=>"000000000",
  17574=>"100100000",
  17575=>"001010010",
  17576=>"000011110",
  17577=>"010101100",
  17578=>"000011010",
  17579=>"010000101",
  17580=>"011110011",
  17581=>"001011111",
  17582=>"000110100",
  17583=>"011011111",
  17584=>"100001110",
  17585=>"000010001",
  17586=>"111110010",
  17587=>"011100011",
  17588=>"110101100",
  17589=>"010100110",
  17590=>"010101000",
  17591=>"001000101",
  17592=>"000101100",
  17593=>"011001011",
  17594=>"010000101",
  17595=>"011101110",
  17596=>"110100110",
  17597=>"000001110",
  17598=>"101110011",
  17599=>"011000100",
  17600=>"011101110",
  17601=>"110111001",
  17602=>"111001110",
  17603=>"110010000",
  17604=>"001001100",
  17605=>"101001101",
  17606=>"011110001",
  17607=>"000100001",
  17608=>"000011001",
  17609=>"111011111",
  17610=>"111111100",
  17611=>"011011001",
  17612=>"111000000",
  17613=>"101000110",
  17614=>"110100100",
  17615=>"000101101",
  17616=>"111101101",
  17617=>"001111111",
  17618=>"101110010",
  17619=>"100100011",
  17620=>"101110001",
  17621=>"111001001",
  17622=>"100001001",
  17623=>"111110101",
  17624=>"100001110",
  17625=>"101100001",
  17626=>"111111101",
  17627=>"101010001",
  17628=>"100010000",
  17629=>"011111101",
  17630=>"010000011",
  17631=>"001101001",
  17632=>"100001000",
  17633=>"001101100",
  17634=>"100011001",
  17635=>"010111100",
  17636=>"111111111",
  17637=>"010000001",
  17638=>"000100000",
  17639=>"100101011",
  17640=>"001000011",
  17641=>"111110011",
  17642=>"001010110",
  17643=>"101101001",
  17644=>"110110100",
  17645=>"000110100",
  17646=>"111110101",
  17647=>"010000100",
  17648=>"010000111",
  17649=>"111101100",
  17650=>"101010101",
  17651=>"000000110",
  17652=>"110101000",
  17653=>"011010101",
  17654=>"010000011",
  17655=>"100001010",
  17656=>"000000001",
  17657=>"011011001",
  17658=>"111001101",
  17659=>"111111011",
  17660=>"100011011",
  17661=>"101110100",
  17662=>"011000111",
  17663=>"011000111",
  17664=>"011011101",
  17665=>"111001000",
  17666=>"100110111",
  17667=>"000011100",
  17668=>"011011101",
  17669=>"111100011",
  17670=>"000101011",
  17671=>"011111010",
  17672=>"111010010",
  17673=>"010100011",
  17674=>"000001010",
  17675=>"101000111",
  17676=>"101011011",
  17677=>"011101001",
  17678=>"111100101",
  17679=>"011111100",
  17680=>"001111111",
  17681=>"010000100",
  17682=>"001111001",
  17683=>"001001000",
  17684=>"111000001",
  17685=>"000101100",
  17686=>"011101110",
  17687=>"111111110",
  17688=>"000101000",
  17689=>"111100011",
  17690=>"000110011",
  17691=>"011010001",
  17692=>"011111101",
  17693=>"011100010",
  17694=>"101000101",
  17695=>"010000111",
  17696=>"011001100",
  17697=>"001010000",
  17698=>"111111110",
  17699=>"100011000",
  17700=>"010101101",
  17701=>"101001011",
  17702=>"000001011",
  17703=>"011111101",
  17704=>"000011101",
  17705=>"110011010",
  17706=>"000111101",
  17707=>"100110000",
  17708=>"111110001",
  17709=>"011010111",
  17710=>"000000000",
  17711=>"110000101",
  17712=>"000110100",
  17713=>"110111011",
  17714=>"110111010",
  17715=>"110011110",
  17716=>"000100101",
  17717=>"100010011",
  17718=>"011000100",
  17719=>"111000111",
  17720=>"001100000",
  17721=>"011010101",
  17722=>"101011110",
  17723=>"001100101",
  17724=>"100100100",
  17725=>"001101101",
  17726=>"010011011",
  17727=>"100010111",
  17728=>"000110000",
  17729=>"000000000",
  17730=>"000000000",
  17731=>"100011000",
  17732=>"101011000",
  17733=>"100001000",
  17734=>"100101000",
  17735=>"111001100",
  17736=>"111010110",
  17737=>"101110010",
  17738=>"100010110",
  17739=>"010100100",
  17740=>"001111011",
  17741=>"011101001",
  17742=>"101110111",
  17743=>"111111001",
  17744=>"010101110",
  17745=>"111010100",
  17746=>"001101011",
  17747=>"101000000",
  17748=>"110001111",
  17749=>"010011010",
  17750=>"110010000",
  17751=>"110100001",
  17752=>"000100010",
  17753=>"011001010",
  17754=>"110000101",
  17755=>"001110011",
  17756=>"110100101",
  17757=>"010000110",
  17758=>"111110000",
  17759=>"111111101",
  17760=>"110011110",
  17761=>"111010001",
  17762=>"111001010",
  17763=>"000101000",
  17764=>"110011111",
  17765=>"001100111",
  17766=>"000100101",
  17767=>"001001101",
  17768=>"111001010",
  17769=>"110010001",
  17770=>"001010000",
  17771=>"000000100",
  17772=>"000000000",
  17773=>"110010000",
  17774=>"001110110",
  17775=>"100010000",
  17776=>"100010001",
  17777=>"100111100",
  17778=>"011110010",
  17779=>"011011111",
  17780=>"111110010",
  17781=>"110100011",
  17782=>"101101011",
  17783=>"101101100",
  17784=>"100100010",
  17785=>"000000101",
  17786=>"110001111",
  17787=>"101100000",
  17788=>"111010100",
  17789=>"001100110",
  17790=>"010001001",
  17791=>"010101001",
  17792=>"111111000",
  17793=>"111101001",
  17794=>"110101111",
  17795=>"100010001",
  17796=>"101000000",
  17797=>"111100000",
  17798=>"101111110",
  17799=>"111111001",
  17800=>"001000101",
  17801=>"001001010",
  17802=>"110010000",
  17803=>"000010011",
  17804=>"111010101",
  17805=>"101000111",
  17806=>"011001110",
  17807=>"000100010",
  17808=>"010101010",
  17809=>"001101011",
  17810=>"010111111",
  17811=>"001001011",
  17812=>"101010001",
  17813=>"011000000",
  17814=>"001000100",
  17815=>"111010001",
  17816=>"010010100",
  17817=>"010100100",
  17818=>"101010100",
  17819=>"000110110",
  17820=>"110001100",
  17821=>"000100000",
  17822=>"100101010",
  17823=>"010000110",
  17824=>"100101011",
  17825=>"000110000",
  17826=>"110011100",
  17827=>"010110001",
  17828=>"001111000",
  17829=>"000000111",
  17830=>"001111110",
  17831=>"001100011",
  17832=>"011110111",
  17833=>"001110111",
  17834=>"000100000",
  17835=>"111011000",
  17836=>"001010011",
  17837=>"010011110",
  17838=>"000010011",
  17839=>"001100110",
  17840=>"101111111",
  17841=>"010010101",
  17842=>"111111000",
  17843=>"000011000",
  17844=>"111101100",
  17845=>"011010100",
  17846=>"101011010",
  17847=>"101001111",
  17848=>"001111010",
  17849=>"111111110",
  17850=>"101101101",
  17851=>"011100101",
  17852=>"111101001",
  17853=>"101000000",
  17854=>"101111001",
  17855=>"101111011",
  17856=>"110110011",
  17857=>"001101011",
  17858=>"100110000",
  17859=>"111110010",
  17860=>"000100010",
  17861=>"110010100",
  17862=>"101100100",
  17863=>"010110110",
  17864=>"110010111",
  17865=>"001001000",
  17866=>"111000111",
  17867=>"011111101",
  17868=>"011110101",
  17869=>"000100100",
  17870=>"101111010",
  17871=>"111110100",
  17872=>"001010000",
  17873=>"010111000",
  17874=>"010011000",
  17875=>"111001110",
  17876=>"111100000",
  17877=>"010000000",
  17878=>"100110011",
  17879=>"111100001",
  17880=>"101110010",
  17881=>"010000000",
  17882=>"110101011",
  17883=>"101111011",
  17884=>"100111010",
  17885=>"000110110",
  17886=>"010010000",
  17887=>"100000101",
  17888=>"101111101",
  17889=>"110010001",
  17890=>"101100001",
  17891=>"000011110",
  17892=>"100000110",
  17893=>"110111110",
  17894=>"010000000",
  17895=>"101010111",
  17896=>"011011100",
  17897=>"000111011",
  17898=>"101100101",
  17899=>"100000111",
  17900=>"011101000",
  17901=>"100110000",
  17902=>"111110011",
  17903=>"000110111",
  17904=>"111010001",
  17905=>"100110101",
  17906=>"100011111",
  17907=>"110010010",
  17908=>"001011011",
  17909=>"001000001",
  17910=>"111010110",
  17911=>"111101111",
  17912=>"010110110",
  17913=>"111111001",
  17914=>"110010110",
  17915=>"101001000",
  17916=>"111011110",
  17917=>"001001001",
  17918=>"000001000",
  17919=>"110000010",
  17920=>"101011010",
  17921=>"000101011",
  17922=>"001001100",
  17923=>"101000100",
  17924=>"110110101",
  17925=>"011111101",
  17926=>"011110100",
  17927=>"011100101",
  17928=>"010100000",
  17929=>"000110110",
  17930=>"000011000",
  17931=>"000000100",
  17932=>"011011101",
  17933=>"010001010",
  17934=>"001000110",
  17935=>"010010001",
  17936=>"011100001",
  17937=>"101001000",
  17938=>"011111001",
  17939=>"011111111",
  17940=>"110111010",
  17941=>"100001001",
  17942=>"100101011",
  17943=>"000000111",
  17944=>"001110100",
  17945=>"100000001",
  17946=>"011101011",
  17947=>"000000100",
  17948=>"101001111",
  17949=>"100000110",
  17950=>"001101110",
  17951=>"101001110",
  17952=>"000010000",
  17953=>"010100101",
  17954=>"110100011",
  17955=>"000111111",
  17956=>"001111001",
  17957=>"011010100",
  17958=>"010100110",
  17959=>"110010001",
  17960=>"100010001",
  17961=>"010110100",
  17962=>"000011000",
  17963=>"101101101",
  17964=>"010101111",
  17965=>"011110100",
  17966=>"110011100",
  17967=>"101101111",
  17968=>"010010000",
  17969=>"000010101",
  17970=>"000100111",
  17971=>"010000100",
  17972=>"111111001",
  17973=>"001011101",
  17974=>"111100100",
  17975=>"011100010",
  17976=>"111000101",
  17977=>"110001110",
  17978=>"011100010",
  17979=>"101011011",
  17980=>"110001000",
  17981=>"000010000",
  17982=>"110001110",
  17983=>"110001001",
  17984=>"000110101",
  17985=>"000111110",
  17986=>"110011010",
  17987=>"100101110",
  17988=>"011111000",
  17989=>"100010011",
  17990=>"101001111",
  17991=>"000100001",
  17992=>"100000101",
  17993=>"101001001",
  17994=>"110101010",
  17995=>"010011011",
  17996=>"100000111",
  17997=>"010011001",
  17998=>"011011100",
  17999=>"000011101",
  18000=>"011101000",
  18001=>"111100101",
  18002=>"000111101",
  18003=>"101111000",
  18004=>"101001111",
  18005=>"010010001",
  18006=>"101111001",
  18007=>"010001011",
  18008=>"111010011",
  18009=>"110110100",
  18010=>"111000111",
  18011=>"010101101",
  18012=>"100100010",
  18013=>"101110100",
  18014=>"100010101",
  18015=>"101000100",
  18016=>"001010110",
  18017=>"000101000",
  18018=>"001011110",
  18019=>"010011001",
  18020=>"110101101",
  18021=>"000101000",
  18022=>"000001111",
  18023=>"000110101",
  18024=>"101000101",
  18025=>"000011100",
  18026=>"010110000",
  18027=>"111001000",
  18028=>"100001000",
  18029=>"010000000",
  18030=>"100100110",
  18031=>"000000111",
  18032=>"000110110",
  18033=>"100101101",
  18034=>"110110000",
  18035=>"011000010",
  18036=>"011100100",
  18037=>"010001001",
  18038=>"101111111",
  18039=>"001010010",
  18040=>"111101000",
  18041=>"010000010",
  18042=>"110110001",
  18043=>"100010010",
  18044=>"100000000",
  18045=>"110101001",
  18046=>"001011001",
  18047=>"100010110",
  18048=>"001000100",
  18049=>"001101111",
  18050=>"101001101",
  18051=>"011010110",
  18052=>"000010011",
  18053=>"100111011",
  18054=>"000111110",
  18055=>"110010000",
  18056=>"101100011",
  18057=>"011100100",
  18058=>"110011011",
  18059=>"101010110",
  18060=>"101001000",
  18061=>"100110111",
  18062=>"101001001",
  18063=>"010111011",
  18064=>"000000100",
  18065=>"100111001",
  18066=>"001011001",
  18067=>"110101101",
  18068=>"011101000",
  18069=>"101011011",
  18070=>"100001111",
  18071=>"010010111",
  18072=>"011110000",
  18073=>"000010011",
  18074=>"000010111",
  18075=>"001010010",
  18076=>"100110010",
  18077=>"001000111",
  18078=>"111111011",
  18079=>"100111010",
  18080=>"111101110",
  18081=>"101111000",
  18082=>"101100000",
  18083=>"001111110",
  18084=>"011111000",
  18085=>"111101101",
  18086=>"010010010",
  18087=>"000011011",
  18088=>"111010111",
  18089=>"001000010",
  18090=>"100001000",
  18091=>"011100100",
  18092=>"101010111",
  18093=>"000000001",
  18094=>"100010001",
  18095=>"100100101",
  18096=>"101001100",
  18097=>"010111110",
  18098=>"000010010",
  18099=>"001011100",
  18100=>"101110000",
  18101=>"000110011",
  18102=>"011101001",
  18103=>"100110011",
  18104=>"100000011",
  18105=>"010000110",
  18106=>"111111011",
  18107=>"000001001",
  18108=>"000010000",
  18109=>"000100010",
  18110=>"010000111",
  18111=>"010101100",
  18112=>"110101111",
  18113=>"100010011",
  18114=>"100000100",
  18115=>"110010100",
  18116=>"110111110",
  18117=>"111001110",
  18118=>"110110001",
  18119=>"011101100",
  18120=>"000000111",
  18121=>"110111001",
  18122=>"001011001",
  18123=>"111101101",
  18124=>"101111110",
  18125=>"001010101",
  18126=>"101001011",
  18127=>"100100110",
  18128=>"100110110",
  18129=>"110101011",
  18130=>"000110111",
  18131=>"010001000",
  18132=>"100001010",
  18133=>"110100111",
  18134=>"111000111",
  18135=>"011111111",
  18136=>"010110001",
  18137=>"001110111",
  18138=>"111011100",
  18139=>"110000101",
  18140=>"101011101",
  18141=>"100111100",
  18142=>"001111100",
  18143=>"100100000",
  18144=>"001100010",
  18145=>"000111100",
  18146=>"000000110",
  18147=>"101101011",
  18148=>"101001101",
  18149=>"011000100",
  18150=>"000000110",
  18151=>"100010001",
  18152=>"101101011",
  18153=>"100101001",
  18154=>"001111001",
  18155=>"101001010",
  18156=>"111001101",
  18157=>"101011001",
  18158=>"001111101",
  18159=>"100100111",
  18160=>"011100111",
  18161=>"100011100",
  18162=>"001001111",
  18163=>"100000001",
  18164=>"011000011",
  18165=>"100000100",
  18166=>"000001110",
  18167=>"010000000",
  18168=>"000010011",
  18169=>"110110110",
  18170=>"110101111",
  18171=>"000011111",
  18172=>"000001011",
  18173=>"111001011",
  18174=>"011010000",
  18175=>"100000101",
  18176=>"110100010",
  18177=>"111111101",
  18178=>"100100111",
  18179=>"001100011",
  18180=>"010000010",
  18181=>"010101110",
  18182=>"011110110",
  18183=>"011000111",
  18184=>"101000000",
  18185=>"000000011",
  18186=>"000110011",
  18187=>"100010110",
  18188=>"001110111",
  18189=>"110101010",
  18190=>"000010000",
  18191=>"100000001",
  18192=>"011111001",
  18193=>"011001000",
  18194=>"101000000",
  18195=>"110110010",
  18196=>"001001111",
  18197=>"101100100",
  18198=>"101010110",
  18199=>"000000000",
  18200=>"111100000",
  18201=>"110010110",
  18202=>"101010010",
  18203=>"001010001",
  18204=>"010010011",
  18205=>"100001000",
  18206=>"001101011",
  18207=>"110010111",
  18208=>"100011101",
  18209=>"000100111",
  18210=>"000001110",
  18211=>"100010101",
  18212=>"000110101",
  18213=>"011000110",
  18214=>"001010100",
  18215=>"101111110",
  18216=>"001100010",
  18217=>"100000010",
  18218=>"011011100",
  18219=>"101101100",
  18220=>"110000000",
  18221=>"100110010",
  18222=>"111001100",
  18223=>"010011010",
  18224=>"001110011",
  18225=>"010110111",
  18226=>"111111111",
  18227=>"110011101",
  18228=>"110010101",
  18229=>"011100111",
  18230=>"010111111",
  18231=>"000001010",
  18232=>"111011011",
  18233=>"001100000",
  18234=>"100011110",
  18235=>"101011111",
  18236=>"101000000",
  18237=>"000100101",
  18238=>"000011010",
  18239=>"110000110",
  18240=>"111011111",
  18241=>"100011000",
  18242=>"010110100",
  18243=>"010110011",
  18244=>"000011100",
  18245=>"001101111",
  18246=>"010010000",
  18247=>"011011010",
  18248=>"111110100",
  18249=>"000101111",
  18250=>"100111111",
  18251=>"011100101",
  18252=>"110001000",
  18253=>"111111110",
  18254=>"101110101",
  18255=>"101100001",
  18256=>"111001100",
  18257=>"101010011",
  18258=>"100101001",
  18259=>"100101100",
  18260=>"100100110",
  18261=>"011110011",
  18262=>"110111110",
  18263=>"001110110",
  18264=>"111011001",
  18265=>"110111001",
  18266=>"000111011",
  18267=>"001100101",
  18268=>"000011000",
  18269=>"100101001",
  18270=>"100110011",
  18271=>"000111010",
  18272=>"011110100",
  18273=>"110011000",
  18274=>"000010000",
  18275=>"101111101",
  18276=>"111001100",
  18277=>"100001000",
  18278=>"001101100",
  18279=>"010110101",
  18280=>"000011101",
  18281=>"000001011",
  18282=>"101001110",
  18283=>"101100110",
  18284=>"100111101",
  18285=>"000000101",
  18286=>"010111100",
  18287=>"010011100",
  18288=>"001111010",
  18289=>"100010110",
  18290=>"110011010",
  18291=>"101001101",
  18292=>"100111000",
  18293=>"111011010",
  18294=>"011011111",
  18295=>"111000100",
  18296=>"000100001",
  18297=>"011010110",
  18298=>"111011010",
  18299=>"000011111",
  18300=>"010111000",
  18301=>"111111100",
  18302=>"000001110",
  18303=>"100010001",
  18304=>"010010011",
  18305=>"010101111",
  18306=>"000111000",
  18307=>"010100000",
  18308=>"010110000",
  18309=>"110101101",
  18310=>"001001101",
  18311=>"000111011",
  18312=>"011101111",
  18313=>"011110111",
  18314=>"000011110",
  18315=>"100001000",
  18316=>"010001010",
  18317=>"100011101",
  18318=>"000100110",
  18319=>"111110111",
  18320=>"100001000",
  18321=>"010100010",
  18322=>"100000010",
  18323=>"110011000",
  18324=>"110000111",
  18325=>"100011110",
  18326=>"100001001",
  18327=>"011010111",
  18328=>"010100000",
  18329=>"011000000",
  18330=>"011100011",
  18331=>"011100101",
  18332=>"000110010",
  18333=>"101101000",
  18334=>"110110101",
  18335=>"001100111",
  18336=>"101011010",
  18337=>"101011100",
  18338=>"111011110",
  18339=>"000000110",
  18340=>"101000101",
  18341=>"010011111",
  18342=>"110111110",
  18343=>"011000011",
  18344=>"100010001",
  18345=>"101010100",
  18346=>"110110111",
  18347=>"100111100",
  18348=>"000010100",
  18349=>"011110100",
  18350=>"100010110",
  18351=>"010111011",
  18352=>"111111101",
  18353=>"011010010",
  18354=>"111111111",
  18355=>"010001100",
  18356=>"000000101",
  18357=>"101011000",
  18358=>"011101000",
  18359=>"101001111",
  18360=>"101110110",
  18361=>"110010001",
  18362=>"100000101",
  18363=>"110010000",
  18364=>"010010011",
  18365=>"000011001",
  18366=>"101011110",
  18367=>"001011001",
  18368=>"100010110",
  18369=>"100110001",
  18370=>"101001111",
  18371=>"001100000",
  18372=>"000110000",
  18373=>"111111010",
  18374=>"011000100",
  18375=>"111101111",
  18376=>"110011100",
  18377=>"010100001",
  18378=>"100101011",
  18379=>"100100101",
  18380=>"010101011",
  18381=>"100010000",
  18382=>"110111101",
  18383=>"011011110",
  18384=>"010000010",
  18385=>"000110001",
  18386=>"101011010",
  18387=>"101101111",
  18388=>"011001001",
  18389=>"100010000",
  18390=>"100111011",
  18391=>"110110111",
  18392=>"000101000",
  18393=>"100101100",
  18394=>"010001111",
  18395=>"111101101",
  18396=>"100111011",
  18397=>"010110011",
  18398=>"010100010",
  18399=>"000001000",
  18400=>"100001101",
  18401=>"010010000",
  18402=>"100111111",
  18403=>"011110101",
  18404=>"000001100",
  18405=>"111000001",
  18406=>"101010101",
  18407=>"011000000",
  18408=>"011101100",
  18409=>"000001100",
  18410=>"100101101",
  18411=>"111011010",
  18412=>"011010110",
  18413=>"000000011",
  18414=>"010101101",
  18415=>"111101110",
  18416=>"101000100",
  18417=>"010011100",
  18418=>"101111010",
  18419=>"111100110",
  18420=>"101010001",
  18421=>"010101000",
  18422=>"110111100",
  18423=>"111000111",
  18424=>"110101011",
  18425=>"010100111",
  18426=>"100100101",
  18427=>"100110111",
  18428=>"000000110",
  18429=>"100101010",
  18430=>"011101110",
  18431=>"110000000",
  18432=>"011110100",
  18433=>"110110011",
  18434=>"111000100",
  18435=>"010000010",
  18436=>"111100001",
  18437=>"111010111",
  18438=>"000001000",
  18439=>"100101010",
  18440=>"101010001",
  18441=>"001000010",
  18442=>"001011011",
  18443=>"001111101",
  18444=>"100110011",
  18445=>"101101101",
  18446=>"010000101",
  18447=>"010101000",
  18448=>"010110100",
  18449=>"101000101",
  18450=>"101110011",
  18451=>"101001010",
  18452=>"111111111",
  18453=>"111111001",
  18454=>"000010010",
  18455=>"100000111",
  18456=>"000110001",
  18457=>"101010011",
  18458=>"011100010",
  18459=>"011101111",
  18460=>"001110111",
  18461=>"101100100",
  18462=>"111010110",
  18463=>"100100000",
  18464=>"101000101",
  18465=>"110110110",
  18466=>"011111100",
  18467=>"011001010",
  18468=>"010001100",
  18469=>"111010110",
  18470=>"000100010",
  18471=>"000001010",
  18472=>"100100100",
  18473=>"010011000",
  18474=>"101011010",
  18475=>"011010001",
  18476=>"010000000",
  18477=>"110001110",
  18478=>"000100101",
  18479=>"111101100",
  18480=>"111000101",
  18481=>"111111011",
  18482=>"000000010",
  18483=>"011011110",
  18484=>"111100011",
  18485=>"000000000",
  18486=>"110011010",
  18487=>"110101000",
  18488=>"101110100",
  18489=>"110011001",
  18490=>"001010010",
  18491=>"001011000",
  18492=>"010111101",
  18493=>"110011111",
  18494=>"000000000",
  18495=>"110010111",
  18496=>"001000011",
  18497=>"001010101",
  18498=>"110000010",
  18499=>"001001011",
  18500=>"110000010",
  18501=>"011100001",
  18502=>"010001011",
  18503=>"101110001",
  18504=>"101110000",
  18505=>"111000000",
  18506=>"101100000",
  18507=>"110001000",
  18508=>"011001101",
  18509=>"000111100",
  18510=>"111011110",
  18511=>"010101111",
  18512=>"000011000",
  18513=>"111011010",
  18514=>"000010010",
  18515=>"011010010",
  18516=>"010110110",
  18517=>"001100010",
  18518=>"001111010",
  18519=>"011101000",
  18520=>"110000001",
  18521=>"111011100",
  18522=>"000000011",
  18523=>"111101110",
  18524=>"000000101",
  18525=>"000100000",
  18526=>"010011000",
  18527=>"000001011",
  18528=>"000010000",
  18529=>"010001001",
  18530=>"010000011",
  18531=>"010111011",
  18532=>"010001101",
  18533=>"111111100",
  18534=>"100001101",
  18535=>"000010001",
  18536=>"010000110",
  18537=>"100001010",
  18538=>"010101011",
  18539=>"100010111",
  18540=>"111100000",
  18541=>"010010101",
  18542=>"111000000",
  18543=>"000000001",
  18544=>"010111001",
  18545=>"000001111",
  18546=>"010000110",
  18547=>"110011010",
  18548=>"010101101",
  18549=>"000001010",
  18550=>"101110000",
  18551=>"000101010",
  18552=>"110000001",
  18553=>"000001001",
  18554=>"111010101",
  18555=>"101000100",
  18556=>"111100010",
  18557=>"111110110",
  18558=>"100011101",
  18559=>"110111000",
  18560=>"111011000",
  18561=>"100111001",
  18562=>"011001001",
  18563=>"010010000",
  18564=>"010000000",
  18565=>"010110010",
  18566=>"000011110",
  18567=>"111010111",
  18568=>"110101111",
  18569=>"101110001",
  18570=>"110000111",
  18571=>"111000000",
  18572=>"000100100",
  18573=>"111010101",
  18574=>"101101010",
  18575=>"110100100",
  18576=>"011100010",
  18577=>"100000101",
  18578=>"111100110",
  18579=>"011001110",
  18580=>"101110001",
  18581=>"111000101",
  18582=>"001100010",
  18583=>"110101101",
  18584=>"011101110",
  18585=>"000110101",
  18586=>"111010100",
  18587=>"011011101",
  18588=>"000101000",
  18589=>"011110011",
  18590=>"101111010",
  18591=>"011001101",
  18592=>"101100001",
  18593=>"111100101",
  18594=>"101100111",
  18595=>"001110111",
  18596=>"001011111",
  18597=>"011000111",
  18598=>"001011011",
  18599=>"000111011",
  18600=>"010111101",
  18601=>"000100011",
  18602=>"010011100",
  18603=>"110011111",
  18604=>"010010110",
  18605=>"100101001",
  18606=>"100010100",
  18607=>"111001101",
  18608=>"011010001",
  18609=>"010010000",
  18610=>"010000010",
  18611=>"000100001",
  18612=>"011010001",
  18613=>"101111101",
  18614=>"110011101",
  18615=>"100111011",
  18616=>"001111111",
  18617=>"101010111",
  18618=>"100001111",
  18619=>"011101011",
  18620=>"011011111",
  18621=>"011000110",
  18622=>"001101011",
  18623=>"001110111",
  18624=>"010111111",
  18625=>"101101101",
  18626=>"001110011",
  18627=>"011110111",
  18628=>"111101010",
  18629=>"110101000",
  18630=>"000010100",
  18631=>"100101011",
  18632=>"001100010",
  18633=>"111000111",
  18634=>"000101100",
  18635=>"000010110",
  18636=>"011001101",
  18637=>"000101010",
  18638=>"010001010",
  18639=>"011111111",
  18640=>"010010111",
  18641=>"001101101",
  18642=>"010101111",
  18643=>"000000100",
  18644=>"010101011",
  18645=>"110000110",
  18646=>"110000111",
  18647=>"001111110",
  18648=>"001100010",
  18649=>"011111111",
  18650=>"110111100",
  18651=>"111110011",
  18652=>"101000101",
  18653=>"000010001",
  18654=>"101100010",
  18655=>"011100010",
  18656=>"111011110",
  18657=>"100110010",
  18658=>"110110110",
  18659=>"001010100",
  18660=>"101001011",
  18661=>"101010000",
  18662=>"001100001",
  18663=>"111100000",
  18664=>"010011010",
  18665=>"100110101",
  18666=>"110000000",
  18667=>"000001111",
  18668=>"010000100",
  18669=>"000100100",
  18670=>"000010011",
  18671=>"111000111",
  18672=>"101100000",
  18673=>"110111011",
  18674=>"010110000",
  18675=>"011010110",
  18676=>"011110101",
  18677=>"001111111",
  18678=>"111001010",
  18679=>"000100000",
  18680=>"011010111",
  18681=>"101000101",
  18682=>"010000010",
  18683=>"010000100",
  18684=>"010000101",
  18685=>"100110110",
  18686=>"000011110",
  18687=>"010001000",
  18688=>"111110000",
  18689=>"000110101",
  18690=>"111101101",
  18691=>"000101100",
  18692=>"101011101",
  18693=>"101010000",
  18694=>"000100000",
  18695=>"111010110",
  18696=>"100101011",
  18697=>"010101101",
  18698=>"011111010",
  18699=>"010010001",
  18700=>"001100001",
  18701=>"001111110",
  18702=>"110101100",
  18703=>"000101100",
  18704=>"000001000",
  18705=>"100011011",
  18706=>"111001010",
  18707=>"110101100",
  18708=>"011011011",
  18709=>"011011001",
  18710=>"011001101",
  18711=>"100110111",
  18712=>"011010110",
  18713=>"010010100",
  18714=>"001011000",
  18715=>"100001101",
  18716=>"000000110",
  18717=>"111011101",
  18718=>"110100111",
  18719=>"101000110",
  18720=>"010001101",
  18721=>"101011101",
  18722=>"100011000",
  18723=>"000101010",
  18724=>"111101111",
  18725=>"001100001",
  18726=>"110110011",
  18727=>"111000101",
  18728=>"111010010",
  18729=>"001100000",
  18730=>"001010011",
  18731=>"110100000",
  18732=>"111110010",
  18733=>"110000100",
  18734=>"010011010",
  18735=>"001011011",
  18736=>"101101001",
  18737=>"000101111",
  18738=>"100010000",
  18739=>"101101000",
  18740=>"100100101",
  18741=>"100010110",
  18742=>"000111011",
  18743=>"011010101",
  18744=>"011011001",
  18745=>"001001001",
  18746=>"000110101",
  18747=>"101101111",
  18748=>"011111111",
  18749=>"101001001",
  18750=>"100010001",
  18751=>"111011010",
  18752=>"010100001",
  18753=>"010110110",
  18754=>"011110001",
  18755=>"001010100",
  18756=>"001101000",
  18757=>"001011100",
  18758=>"110000010",
  18759=>"111011110",
  18760=>"010001000",
  18761=>"101110111",
  18762=>"101110101",
  18763=>"011101011",
  18764=>"010000010",
  18765=>"111010110",
  18766=>"100110100",
  18767=>"000011010",
  18768=>"000110101",
  18769=>"010010110",
  18770=>"111101101",
  18771=>"000111001",
  18772=>"010001011",
  18773=>"001000110",
  18774=>"111000101",
  18775=>"001011011",
  18776=>"001000011",
  18777=>"101010011",
  18778=>"011111101",
  18779=>"011010111",
  18780=>"000111110",
  18781=>"011110011",
  18782=>"010111000",
  18783=>"010100101",
  18784=>"111011101",
  18785=>"111110101",
  18786=>"111111001",
  18787=>"001111101",
  18788=>"010000101",
  18789=>"110001001",
  18790=>"100111100",
  18791=>"000011010",
  18792=>"000010101",
  18793=>"000011001",
  18794=>"111000000",
  18795=>"010110100",
  18796=>"011110001",
  18797=>"100001111",
  18798=>"100010000",
  18799=>"100000001",
  18800=>"001100101",
  18801=>"110110100",
  18802=>"001000111",
  18803=>"100111101",
  18804=>"000100101",
  18805=>"011100111",
  18806=>"011111000",
  18807=>"111100111",
  18808=>"011110110",
  18809=>"011111110",
  18810=>"011101101",
  18811=>"101000101",
  18812=>"011000001",
  18813=>"111010001",
  18814=>"011100110",
  18815=>"100100010",
  18816=>"101110001",
  18817=>"000000001",
  18818=>"011110001",
  18819=>"011110000",
  18820=>"000010101",
  18821=>"100010101",
  18822=>"100111011",
  18823=>"101010000",
  18824=>"010111010",
  18825=>"011111101",
  18826=>"110000111",
  18827=>"100001000",
  18828=>"001111100",
  18829=>"101011011",
  18830=>"100111111",
  18831=>"100100111",
  18832=>"110010110",
  18833=>"000001100",
  18834=>"100110111",
  18835=>"000011010",
  18836=>"110101111",
  18837=>"000110101",
  18838=>"000101000",
  18839=>"000000010",
  18840=>"011010010",
  18841=>"001011101",
  18842=>"010111000",
  18843=>"011000000",
  18844=>"000011111",
  18845=>"000110111",
  18846=>"110001110",
  18847=>"010110100",
  18848=>"111010100",
  18849=>"000011010",
  18850=>"011110101",
  18851=>"001001000",
  18852=>"010100101",
  18853=>"100100011",
  18854=>"110110101",
  18855=>"001011011",
  18856=>"101001100",
  18857=>"001001011",
  18858=>"100111001",
  18859=>"001110111",
  18860=>"000001100",
  18861=>"111110001",
  18862=>"011011000",
  18863=>"010111000",
  18864=>"001011000",
  18865=>"000000101",
  18866=>"110000100",
  18867=>"000100011",
  18868=>"010100100",
  18869=>"000111000",
  18870=>"010001010",
  18871=>"101101111",
  18872=>"010110110",
  18873=>"110111001",
  18874=>"110111100",
  18875=>"001011101",
  18876=>"100110110",
  18877=>"111110011",
  18878=>"110010001",
  18879=>"111100001",
  18880=>"001011111",
  18881=>"001100100",
  18882=>"000101110",
  18883=>"110100000",
  18884=>"100000000",
  18885=>"101100100",
  18886=>"110110000",
  18887=>"000111011",
  18888=>"011111000",
  18889=>"100010011",
  18890=>"010101010",
  18891=>"110100111",
  18892=>"001110101",
  18893=>"111011111",
  18894=>"000100100",
  18895=>"010100010",
  18896=>"110101011",
  18897=>"000001100",
  18898=>"100001011",
  18899=>"011010100",
  18900=>"110100111",
  18901=>"100000101",
  18902=>"111100010",
  18903=>"010111011",
  18904=>"010001001",
  18905=>"000100010",
  18906=>"110101001",
  18907=>"001111000",
  18908=>"000011111",
  18909=>"100010110",
  18910=>"010011010",
  18911=>"100001110",
  18912=>"111101111",
  18913=>"010010000",
  18914=>"000001110",
  18915=>"110001101",
  18916=>"001100000",
  18917=>"000101100",
  18918=>"011000011",
  18919=>"100110001",
  18920=>"110000000",
  18921=>"001001111",
  18922=>"000100001",
  18923=>"110011010",
  18924=>"101010111",
  18925=>"111011010",
  18926=>"000010000",
  18927=>"011010001",
  18928=>"011110010",
  18929=>"110000100",
  18930=>"110110101",
  18931=>"101111000",
  18932=>"000100101",
  18933=>"011011100",
  18934=>"111010001",
  18935=>"110000111",
  18936=>"010001000",
  18937=>"110001010",
  18938=>"001001001",
  18939=>"111010110",
  18940=>"001110101",
  18941=>"101011001",
  18942=>"111111011",
  18943=>"000110100",
  18944=>"111001111",
  18945=>"100000011",
  18946=>"001110011",
  18947=>"000101010",
  18948=>"010000011",
  18949=>"101111010",
  18950=>"101010100",
  18951=>"010011000",
  18952=>"101110000",
  18953=>"011001000",
  18954=>"011101101",
  18955=>"110101000",
  18956=>"000100110",
  18957=>"011111001",
  18958=>"000001000",
  18959=>"100011111",
  18960=>"010101011",
  18961=>"000101101",
  18962=>"101101100",
  18963=>"011101010",
  18964=>"000111000",
  18965=>"000011111",
  18966=>"000111110",
  18967=>"111110011",
  18968=>"110011110",
  18969=>"010011010",
  18970=>"001000001",
  18971=>"100000100",
  18972=>"110111101",
  18973=>"000010000",
  18974=>"001011101",
  18975=>"011011100",
  18976=>"011110101",
  18977=>"000100010",
  18978=>"001010000",
  18979=>"111100010",
  18980=>"010001000",
  18981=>"010100101",
  18982=>"000100000",
  18983=>"110110101",
  18984=>"111110011",
  18985=>"001010001",
  18986=>"001100110",
  18987=>"111001101",
  18988=>"000111110",
  18989=>"000110101",
  18990=>"001000001",
  18991=>"101000100",
  18992=>"100101000",
  18993=>"111011000",
  18994=>"101000011",
  18995=>"110100011",
  18996=>"111110110",
  18997=>"101111011",
  18998=>"010010100",
  18999=>"000110111",
  19000=>"111101010",
  19001=>"110100011",
  19002=>"001110110",
  19003=>"010011111",
  19004=>"001100100",
  19005=>"100001100",
  19006=>"101011111",
  19007=>"000010110",
  19008=>"001000111",
  19009=>"001000001",
  19010=>"110000000",
  19011=>"111000001",
  19012=>"010111101",
  19013=>"010100110",
  19014=>"000000010",
  19015=>"101111111",
  19016=>"001000111",
  19017=>"111010001",
  19018=>"011111110",
  19019=>"011111100",
  19020=>"000001001",
  19021=>"010000011",
  19022=>"100001010",
  19023=>"011010000",
  19024=>"000011001",
  19025=>"001101001",
  19026=>"111011010",
  19027=>"001011111",
  19028=>"000010111",
  19029=>"011001000",
  19030=>"110011100",
  19031=>"110001110",
  19032=>"000101110",
  19033=>"111111111",
  19034=>"011111000",
  19035=>"011110111",
  19036=>"100000011",
  19037=>"000010111",
  19038=>"111110101",
  19039=>"000100001",
  19040=>"001110010",
  19041=>"011000111",
  19042=>"010110111",
  19043=>"111100001",
  19044=>"111111011",
  19045=>"111110100",
  19046=>"001101111",
  19047=>"101100110",
  19048=>"001100110",
  19049=>"011001001",
  19050=>"111110000",
  19051=>"010001001",
  19052=>"101001101",
  19053=>"100101000",
  19054=>"011010101",
  19055=>"000110110",
  19056=>"011110000",
  19057=>"011010100",
  19058=>"100000110",
  19059=>"100000111",
  19060=>"101000110",
  19061=>"011011001",
  19062=>"111010111",
  19063=>"111010011",
  19064=>"011111000",
  19065=>"011111110",
  19066=>"100011000",
  19067=>"001010000",
  19068=>"111010111",
  19069=>"101101101",
  19070=>"001010001",
  19071=>"000101001",
  19072=>"111011100",
  19073=>"111001011",
  19074=>"010000000",
  19075=>"000001111",
  19076=>"110100000",
  19077=>"000011010",
  19078=>"100101010",
  19079=>"111110110",
  19080=>"011000000",
  19081=>"000010001",
  19082=>"010010011",
  19083=>"100001011",
  19084=>"011110101",
  19085=>"110000101",
  19086=>"110001000",
  19087=>"000011000",
  19088=>"001011011",
  19089=>"001011001",
  19090=>"010001001",
  19091=>"100010110",
  19092=>"001101111",
  19093=>"000001101",
  19094=>"110011110",
  19095=>"000001000",
  19096=>"000100100",
  19097=>"111100111",
  19098=>"011110011",
  19099=>"101001000",
  19100=>"001111000",
  19101=>"011000010",
  19102=>"010110010",
  19103=>"011101011",
  19104=>"111101111",
  19105=>"011110110",
  19106=>"111001111",
  19107=>"000110000",
  19108=>"001100110",
  19109=>"100010111",
  19110=>"100111000",
  19111=>"011000000",
  19112=>"000000100",
  19113=>"001100011",
  19114=>"110000100",
  19115=>"110101100",
  19116=>"000001001",
  19117=>"000000000",
  19118=>"001001010",
  19119=>"000110111",
  19120=>"001000100",
  19121=>"101010010",
  19122=>"110101101",
  19123=>"110000001",
  19124=>"001100111",
  19125=>"101010100",
  19126=>"101111000",
  19127=>"101011010",
  19128=>"101001011",
  19129=>"110000010",
  19130=>"100101111",
  19131=>"011000011",
  19132=>"000100000",
  19133=>"001000011",
  19134=>"001101110",
  19135=>"110010101",
  19136=>"110101110",
  19137=>"010110111",
  19138=>"000010011",
  19139=>"111000111",
  19140=>"010011101",
  19141=>"100000100",
  19142=>"111100011",
  19143=>"100010011",
  19144=>"001000000",
  19145=>"101111101",
  19146=>"010111010",
  19147=>"011010110",
  19148=>"100011011",
  19149=>"100110101",
  19150=>"001110011",
  19151=>"001101011",
  19152=>"000011100",
  19153=>"000101111",
  19154=>"101010001",
  19155=>"000111001",
  19156=>"101000101",
  19157=>"010011111",
  19158=>"010110011",
  19159=>"010111011",
  19160=>"110010100",
  19161=>"100100110",
  19162=>"101100101",
  19163=>"101001001",
  19164=>"100100010",
  19165=>"010010001",
  19166=>"100111001",
  19167=>"010011000",
  19168=>"011101010",
  19169=>"101010100",
  19170=>"010110000",
  19171=>"101101011",
  19172=>"000110100",
  19173=>"110110011",
  19174=>"011010000",
  19175=>"100010100",
  19176=>"000010110",
  19177=>"110101101",
  19178=>"100010101",
  19179=>"010010100",
  19180=>"101101100",
  19181=>"111111101",
  19182=>"110111001",
  19183=>"111111111",
  19184=>"101101010",
  19185=>"000100001",
  19186=>"101010011",
  19187=>"000001000",
  19188=>"100001000",
  19189=>"110101011",
  19190=>"110100011",
  19191=>"111011010",
  19192=>"100111000",
  19193=>"111101101",
  19194=>"100101000",
  19195=>"000010110",
  19196=>"110011100",
  19197=>"000000010",
  19198=>"010111100",
  19199=>"110110011",
  19200=>"010000000",
  19201=>"110111011",
  19202=>"101011111",
  19203=>"111110110",
  19204=>"010000100",
  19205=>"000011110",
  19206=>"101010101",
  19207=>"100000110",
  19208=>"100110000",
  19209=>"000111001",
  19210=>"010110111",
  19211=>"100001100",
  19212=>"011111100",
  19213=>"011010010",
  19214=>"001100001",
  19215=>"110011101",
  19216=>"000011011",
  19217=>"010001110",
  19218=>"011000011",
  19219=>"100010100",
  19220=>"111111101",
  19221=>"111110110",
  19222=>"111110001",
  19223=>"110111010",
  19224=>"010100000",
  19225=>"111001101",
  19226=>"111101110",
  19227=>"000011100",
  19228=>"010010010",
  19229=>"011110111",
  19230=>"000000100",
  19231=>"100101001",
  19232=>"111111000",
  19233=>"001001100",
  19234=>"111110101",
  19235=>"001011010",
  19236=>"111111110",
  19237=>"000110100",
  19238=>"111001011",
  19239=>"110010110",
  19240=>"001101111",
  19241=>"111011111",
  19242=>"001010000",
  19243=>"111100110",
  19244=>"010011010",
  19245=>"101101011",
  19246=>"101001101",
  19247=>"111101100",
  19248=>"001100111",
  19249=>"101001001",
  19250=>"110111111",
  19251=>"000000010",
  19252=>"000011101",
  19253=>"001001000",
  19254=>"011010000",
  19255=>"100001100",
  19256=>"010001100",
  19257=>"010101101",
  19258=>"111101110",
  19259=>"010000100",
  19260=>"100100000",
  19261=>"000101010",
  19262=>"001001111",
  19263=>"101100100",
  19264=>"101000100",
  19265=>"000110110",
  19266=>"001100110",
  19267=>"001010011",
  19268=>"001010011",
  19269=>"101110111",
  19270=>"100011000",
  19271=>"000110100",
  19272=>"011100101",
  19273=>"110010101",
  19274=>"100100101",
  19275=>"001001100",
  19276=>"010100000",
  19277=>"010000001",
  19278=>"000001010",
  19279=>"110110010",
  19280=>"111101001",
  19281=>"000010111",
  19282=>"000110011",
  19283=>"000110010",
  19284=>"110100110",
  19285=>"010100000",
  19286=>"100010111",
  19287=>"000110110",
  19288=>"011111111",
  19289=>"000010011",
  19290=>"111101001",
  19291=>"000100101",
  19292=>"001001010",
  19293=>"100011001",
  19294=>"101111111",
  19295=>"001110011",
  19296=>"100111100",
  19297=>"100100010",
  19298=>"010111110",
  19299=>"110111111",
  19300=>"101100100",
  19301=>"110010011",
  19302=>"100010110",
  19303=>"011110111",
  19304=>"101010110",
  19305=>"111110010",
  19306=>"100101100",
  19307=>"011111101",
  19308=>"010110010",
  19309=>"101010011",
  19310=>"110011100",
  19311=>"101101001",
  19312=>"010000000",
  19313=>"110111110",
  19314=>"101011010",
  19315=>"010001110",
  19316=>"000000001",
  19317=>"001100001",
  19318=>"011100011",
  19319=>"001010100",
  19320=>"011111001",
  19321=>"000001100",
  19322=>"001000010",
  19323=>"010111111",
  19324=>"000000001",
  19325=>"000011010",
  19326=>"101111111",
  19327=>"101001100",
  19328=>"101111110",
  19329=>"010011000",
  19330=>"100110011",
  19331=>"000101010",
  19332=>"100001010",
  19333=>"101100011",
  19334=>"111110010",
  19335=>"110101010",
  19336=>"110100100",
  19337=>"010010001",
  19338=>"000000100",
  19339=>"001100100",
  19340=>"000111111",
  19341=>"010010111",
  19342=>"111010000",
  19343=>"001011100",
  19344=>"000011001",
  19345=>"100001011",
  19346=>"010110101",
  19347=>"111100000",
  19348=>"000110001",
  19349=>"110010110",
  19350=>"100001000",
  19351=>"110111010",
  19352=>"101000110",
  19353=>"101000001",
  19354=>"000110111",
  19355=>"011101000",
  19356=>"101011111",
  19357=>"101110000",
  19358=>"101010100",
  19359=>"110111101",
  19360=>"000000000",
  19361=>"000111000",
  19362=>"100011111",
  19363=>"000001100",
  19364=>"001010000",
  19365=>"000110100",
  19366=>"111111111",
  19367=>"001000100",
  19368=>"000010010",
  19369=>"111111000",
  19370=>"111001001",
  19371=>"001001111",
  19372=>"010000111",
  19373=>"101101111",
  19374=>"100010011",
  19375=>"110000101",
  19376=>"000001011",
  19377=>"110101100",
  19378=>"000100011",
  19379=>"001101001",
  19380=>"011011001",
  19381=>"001100100",
  19382=>"001001010",
  19383=>"101101100",
  19384=>"011101111",
  19385=>"110110000",
  19386=>"100001111",
  19387=>"010110010",
  19388=>"001010000",
  19389=>"010100100",
  19390=>"001110010",
  19391=>"001000001",
  19392=>"000100011",
  19393=>"110010110",
  19394=>"011111101",
  19395=>"100011110",
  19396=>"011111110",
  19397=>"011000000",
  19398=>"111101010",
  19399=>"101100111",
  19400=>"000000010",
  19401=>"011011111",
  19402=>"111111001",
  19403=>"010000110",
  19404=>"010111101",
  19405=>"000010001",
  19406=>"100011110",
  19407=>"011101110",
  19408=>"111100110",
  19409=>"011010010",
  19410=>"110011101",
  19411=>"001100101",
  19412=>"100000000",
  19413=>"110101101",
  19414=>"101110101",
  19415=>"001001100",
  19416=>"111011111",
  19417=>"010010100",
  19418=>"011101101",
  19419=>"101111001",
  19420=>"111011000",
  19421=>"100100010",
  19422=>"100000010",
  19423=>"011001111",
  19424=>"011001110",
  19425=>"011110001",
  19426=>"111011111",
  19427=>"110010010",
  19428=>"000011001",
  19429=>"111000000",
  19430=>"010011010",
  19431=>"100110111",
  19432=>"000001001",
  19433=>"000100101",
  19434=>"010101100",
  19435=>"010010101",
  19436=>"000010100",
  19437=>"001011111",
  19438=>"111111010",
  19439=>"101111111",
  19440=>"000111110",
  19441=>"001100110",
  19442=>"000111010",
  19443=>"011110111",
  19444=>"011010010",
  19445=>"110110111",
  19446=>"111101110",
  19447=>"110100010",
  19448=>"010111101",
  19449=>"100110110",
  19450=>"101011101",
  19451=>"101010000",
  19452=>"110011000",
  19453=>"101100111",
  19454=>"100110010",
  19455=>"110010000",
  19456=>"011111110",
  19457=>"111100111",
  19458=>"000100001",
  19459=>"110110101",
  19460=>"000011000",
  19461=>"011000110",
  19462=>"010101111",
  19463=>"111011001",
  19464=>"110100100",
  19465=>"111011001",
  19466=>"110011001",
  19467=>"001100000",
  19468=>"011011011",
  19469=>"000100011",
  19470=>"110010110",
  19471=>"010100110",
  19472=>"000101011",
  19473=>"100111111",
  19474=>"110010111",
  19475=>"011001110",
  19476=>"001110101",
  19477=>"111010010",
  19478=>"001101111",
  19479=>"101100101",
  19480=>"110110001",
  19481=>"101001000",
  19482=>"100100111",
  19483=>"111111101",
  19484=>"111101001",
  19485=>"001100100",
  19486=>"010100101",
  19487=>"000001110",
  19488=>"100101001",
  19489=>"110111010",
  19490=>"011001110",
  19491=>"001100111",
  19492=>"111011000",
  19493=>"000101010",
  19494=>"101101001",
  19495=>"110000110",
  19496=>"001110111",
  19497=>"111001110",
  19498=>"110100110",
  19499=>"000111001",
  19500=>"001010101",
  19501=>"000011110",
  19502=>"101000100",
  19503=>"111111001",
  19504=>"111101010",
  19505=>"001010011",
  19506=>"101110110",
  19507=>"100001100",
  19508=>"001101000",
  19509=>"110100010",
  19510=>"111110111",
  19511=>"000110011",
  19512=>"101000110",
  19513=>"010101000",
  19514=>"111101110",
  19515=>"000000000",
  19516=>"010000001",
  19517=>"011000011",
  19518=>"111001011",
  19519=>"000011000",
  19520=>"110011101",
  19521=>"001100010",
  19522=>"111111010",
  19523=>"100011111",
  19524=>"110111011",
  19525=>"111111101",
  19526=>"100101011",
  19527=>"001010001",
  19528=>"110000101",
  19529=>"001110100",
  19530=>"011000101",
  19531=>"110111000",
  19532=>"000100010",
  19533=>"111000000",
  19534=>"111010100",
  19535=>"111111110",
  19536=>"000000100",
  19537=>"111100111",
  19538=>"100111001",
  19539=>"010101101",
  19540=>"110001111",
  19541=>"000001110",
  19542=>"001001011",
  19543=>"111011001",
  19544=>"011000100",
  19545=>"000110011",
  19546=>"001100111",
  19547=>"001001010",
  19548=>"000011010",
  19549=>"100000010",
  19550=>"100110111",
  19551=>"110100001",
  19552=>"101011111",
  19553=>"111001001",
  19554=>"101010100",
  19555=>"111110001",
  19556=>"001100111",
  19557=>"000010100",
  19558=>"000100011",
  19559=>"001010011",
  19560=>"101100011",
  19561=>"000000101",
  19562=>"001111100",
  19563=>"011010001",
  19564=>"010011000",
  19565=>"100000100",
  19566=>"111000011",
  19567=>"010101001",
  19568=>"110100111",
  19569=>"111101010",
  19570=>"111111111",
  19571=>"111110001",
  19572=>"100110111",
  19573=>"000111101",
  19574=>"000100101",
  19575=>"000101111",
  19576=>"100011000",
  19577=>"011101100",
  19578=>"110010100",
  19579=>"100010100",
  19580=>"000111001",
  19581=>"011010000",
  19582=>"101001000",
  19583=>"011000111",
  19584=>"011111101",
  19585=>"111110101",
  19586=>"010010010",
  19587=>"001101101",
  19588=>"011101000",
  19589=>"111101111",
  19590=>"111110110",
  19591=>"111010010",
  19592=>"100100101",
  19593=>"100111011",
  19594=>"011100000",
  19595=>"001110010",
  19596=>"011001001",
  19597=>"000111101",
  19598=>"100011100",
  19599=>"000011110",
  19600=>"101001100",
  19601=>"110111011",
  19602=>"110011000",
  19603=>"010100001",
  19604=>"000010111",
  19605=>"111000010",
  19606=>"000110101",
  19607=>"110010110",
  19608=>"110110101",
  19609=>"010111100",
  19610=>"000011001",
  19611=>"011100101",
  19612=>"011011000",
  19613=>"000001010",
  19614=>"010101010",
  19615=>"100100100",
  19616=>"010001100",
  19617=>"011001011",
  19618=>"101000110",
  19619=>"101111001",
  19620=>"111110001",
  19621=>"100101110",
  19622=>"111000100",
  19623=>"000111111",
  19624=>"011110000",
  19625=>"011111010",
  19626=>"111100111",
  19627=>"111001010",
  19628=>"001101110",
  19629=>"000001001",
  19630=>"011011111",
  19631=>"001111110",
  19632=>"000110011",
  19633=>"000000111",
  19634=>"101011110",
  19635=>"111101010",
  19636=>"010010011",
  19637=>"111010110",
  19638=>"110000001",
  19639=>"011000101",
  19640=>"110100001",
  19641=>"011001110",
  19642=>"011010100",
  19643=>"011000101",
  19644=>"000011011",
  19645=>"110100100",
  19646=>"110110000",
  19647=>"011101111",
  19648=>"110001100",
  19649=>"010010100",
  19650=>"100010110",
  19651=>"110000001",
  19652=>"100100110",
  19653=>"101011001",
  19654=>"100010110",
  19655=>"001011100",
  19656=>"111111011",
  19657=>"100010101",
  19658=>"111001101",
  19659=>"111111100",
  19660=>"001001001",
  19661=>"001011101",
  19662=>"110011101",
  19663=>"010001101",
  19664=>"110010000",
  19665=>"101110101",
  19666=>"010001101",
  19667=>"100001000",
  19668=>"111001011",
  19669=>"111101100",
  19670=>"011000010",
  19671=>"001110001",
  19672=>"001100110",
  19673=>"000110101",
  19674=>"100100100",
  19675=>"110101000",
  19676=>"111000100",
  19677=>"010111011",
  19678=>"001010110",
  19679=>"001110000",
  19680=>"010100011",
  19681=>"111100110",
  19682=>"101001111",
  19683=>"001111111",
  19684=>"001101001",
  19685=>"110100111",
  19686=>"111011001",
  19687=>"100001001",
  19688=>"101010011",
  19689=>"100010111",
  19690=>"110011101",
  19691=>"100110100",
  19692=>"011101110",
  19693=>"110101101",
  19694=>"000001101",
  19695=>"011010111",
  19696=>"100010000",
  19697=>"110111000",
  19698=>"010110001",
  19699=>"101011101",
  19700=>"111010000",
  19701=>"111111111",
  19702=>"110101011",
  19703=>"011100001",
  19704=>"100100010",
  19705=>"110110000",
  19706=>"110000010",
  19707=>"001001110",
  19708=>"100111011",
  19709=>"010101111",
  19710=>"000001110",
  19711=>"100100000",
  19712=>"101110101",
  19713=>"001001010",
  19714=>"001000000",
  19715=>"000000010",
  19716=>"101011000",
  19717=>"001100010",
  19718=>"010100010",
  19719=>"111010110",
  19720=>"000111000",
  19721=>"011101101",
  19722=>"001011000",
  19723=>"111100011",
  19724=>"000011101",
  19725=>"001100011",
  19726=>"000011010",
  19727=>"000000000",
  19728=>"100110111",
  19729=>"100001101",
  19730=>"000100011",
  19731=>"100111011",
  19732=>"000010100",
  19733=>"011101010",
  19734=>"100110010",
  19735=>"101001000",
  19736=>"111110111",
  19737=>"010110010",
  19738=>"111110010",
  19739=>"100010111",
  19740=>"001111110",
  19741=>"011111001",
  19742=>"000000010",
  19743=>"010010001",
  19744=>"100111101",
  19745=>"000000110",
  19746=>"001011001",
  19747=>"100101001",
  19748=>"001111110",
  19749=>"001010001",
  19750=>"011110000",
  19751=>"110011100",
  19752=>"000101100",
  19753=>"111110001",
  19754=>"010001110",
  19755=>"001110001",
  19756=>"110001101",
  19757=>"110101110",
  19758=>"000111010",
  19759=>"111011010",
  19760=>"100001000",
  19761=>"011000010",
  19762=>"011110001",
  19763=>"000100011",
  19764=>"001011011",
  19765=>"011010000",
  19766=>"100001111",
  19767=>"011111001",
  19768=>"000111100",
  19769=>"100111011",
  19770=>"111111011",
  19771=>"001000001",
  19772=>"110111010",
  19773=>"100110110",
  19774=>"011100101",
  19775=>"101101001",
  19776=>"101101001",
  19777=>"010000010",
  19778=>"111100000",
  19779=>"000101100",
  19780=>"001100110",
  19781=>"010011010",
  19782=>"001110000",
  19783=>"010000101",
  19784=>"000000010",
  19785=>"011010101",
  19786=>"001011010",
  19787=>"110110010",
  19788=>"001001010",
  19789=>"011110111",
  19790=>"101100001",
  19791=>"001100100",
  19792=>"011100110",
  19793=>"100101001",
  19794=>"101110011",
  19795=>"001010111",
  19796=>"000000000",
  19797=>"111111101",
  19798=>"100001101",
  19799=>"111011100",
  19800=>"100001000",
  19801=>"100111000",
  19802=>"100111001",
  19803=>"011010101",
  19804=>"000100110",
  19805=>"111110100",
  19806=>"110110111",
  19807=>"010010011",
  19808=>"110000110",
  19809=>"111000011",
  19810=>"011000010",
  19811=>"101010111",
  19812=>"000101000",
  19813=>"111001101",
  19814=>"001001011",
  19815=>"100011110",
  19816=>"111101001",
  19817=>"101100001",
  19818=>"010111010",
  19819=>"001011001",
  19820=>"010010000",
  19821=>"011011010",
  19822=>"011110100",
  19823=>"000110110",
  19824=>"011000010",
  19825=>"111110100",
  19826=>"110011110",
  19827=>"010010100",
  19828=>"101001111",
  19829=>"001001001",
  19830=>"010001101",
  19831=>"111010110",
  19832=>"111000010",
  19833=>"111000111",
  19834=>"001000100",
  19835=>"000010000",
  19836=>"001001111",
  19837=>"111101111",
  19838=>"100000000",
  19839=>"001001010",
  19840=>"111100010",
  19841=>"000101001",
  19842=>"000111000",
  19843=>"100000100",
  19844=>"001101001",
  19845=>"000000000",
  19846=>"010110111",
  19847=>"111011010",
  19848=>"000001000",
  19849=>"110101111",
  19850=>"011101011",
  19851=>"100100010",
  19852=>"011101111",
  19853=>"010110101",
  19854=>"000100101",
  19855=>"010011011",
  19856=>"101111100",
  19857=>"000010001",
  19858=>"001001010",
  19859=>"111110101",
  19860=>"000110111",
  19861=>"101011011",
  19862=>"111001000",
  19863=>"010111100",
  19864=>"001111100",
  19865=>"010011010",
  19866=>"110111110",
  19867=>"110110010",
  19868=>"100111100",
  19869=>"001010000",
  19870=>"100011011",
  19871=>"101011111",
  19872=>"001001011",
  19873=>"100011110",
  19874=>"010111010",
  19875=>"110111101",
  19876=>"100001111",
  19877=>"010000101",
  19878=>"000011011",
  19879=>"000111001",
  19880=>"110010010",
  19881=>"000111011",
  19882=>"000100001",
  19883=>"000010000",
  19884=>"110111010",
  19885=>"010010111",
  19886=>"110110100",
  19887=>"100011000",
  19888=>"011101101",
  19889=>"011000000",
  19890=>"111101010",
  19891=>"101011000",
  19892=>"010110000",
  19893=>"100111011",
  19894=>"110011000",
  19895=>"011010000",
  19896=>"110101000",
  19897=>"100101000",
  19898=>"000000001",
  19899=>"100111010",
  19900=>"101000000",
  19901=>"111010011",
  19902=>"001111001",
  19903=>"111001101",
  19904=>"110010111",
  19905=>"010000101",
  19906=>"101111110",
  19907=>"100001100",
  19908=>"101001001",
  19909=>"110110100",
  19910=>"111100011",
  19911=>"100010100",
  19912=>"110110101",
  19913=>"001011110",
  19914=>"011010001",
  19915=>"110111011",
  19916=>"000001001",
  19917=>"100010011",
  19918=>"101011011",
  19919=>"000110001",
  19920=>"000000111",
  19921=>"111111000",
  19922=>"101111010",
  19923=>"111101110",
  19924=>"100100111",
  19925=>"101100101",
  19926=>"000000011",
  19927=>"100101111",
  19928=>"100011010",
  19929=>"100001100",
  19930=>"001001101",
  19931=>"111000000",
  19932=>"001010101",
  19933=>"101110010",
  19934=>"100000010",
  19935=>"010110101",
  19936=>"100010011",
  19937=>"001000110",
  19938=>"000001101",
  19939=>"101001001",
  19940=>"100100111",
  19941=>"111011000",
  19942=>"011101110",
  19943=>"110110101",
  19944=>"000000100",
  19945=>"000100101",
  19946=>"110001101",
  19947=>"000000100",
  19948=>"000001110",
  19949=>"110010101",
  19950=>"111001000",
  19951=>"100010101",
  19952=>"010111001",
  19953=>"001111101",
  19954=>"110001110",
  19955=>"100011001",
  19956=>"001011011",
  19957=>"110111101",
  19958=>"010010100",
  19959=>"001010111",
  19960=>"110111100",
  19961=>"101000110",
  19962=>"100111000",
  19963=>"001101000",
  19964=>"110101010",
  19965=>"111000111",
  19966=>"000111011",
  19967=>"111111110",
  19968=>"110110101",
  19969=>"110111100",
  19970=>"100110110",
  19971=>"011011111",
  19972=>"111011010",
  19973=>"011010100",
  19974=>"111010000",
  19975=>"111111111",
  19976=>"001110011",
  19977=>"010101001",
  19978=>"000000001",
  19979=>"111111000",
  19980=>"111111111",
  19981=>"111000101",
  19982=>"011000010",
  19983=>"101100100",
  19984=>"011111101",
  19985=>"000001110",
  19986=>"000100101",
  19987=>"100011100",
  19988=>"101001100",
  19989=>"001011110",
  19990=>"011011010",
  19991=>"010100111",
  19992=>"111111101",
  19993=>"010000001",
  19994=>"011011110",
  19995=>"101100010",
  19996=>"000010000",
  19997=>"101001101",
  19998=>"010011001",
  19999=>"111100101",
  20000=>"010100000",
  20001=>"111100110",
  20002=>"110110000",
  20003=>"001000111",
  20004=>"100000010",
  20005=>"111111111",
  20006=>"101111010",
  20007=>"000000101",
  20008=>"110000101",
  20009=>"110010111",
  20010=>"010111111",
  20011=>"010001110",
  20012=>"110001100",
  20013=>"000110001",
  20014=>"001010010",
  20015=>"000011000",
  20016=>"011011110",
  20017=>"101111111",
  20018=>"110011011",
  20019=>"000000110",
  20020=>"001000000",
  20021=>"001111100",
  20022=>"011010111",
  20023=>"010001010",
  20024=>"010110110",
  20025=>"111110011",
  20026=>"001011101",
  20027=>"011001111",
  20028=>"010111010",
  20029=>"100000011",
  20030=>"100111100",
  20031=>"011100110",
  20032=>"101111001",
  20033=>"010000101",
  20034=>"111111111",
  20035=>"111100001",
  20036=>"100011100",
  20037=>"010110100",
  20038=>"001000000",
  20039=>"001000111",
  20040=>"000000011",
  20041=>"010010000",
  20042=>"111111001",
  20043=>"011010010",
  20044=>"010000110",
  20045=>"001111111",
  20046=>"111100111",
  20047=>"111101111",
  20048=>"000111101",
  20049=>"110011000",
  20050=>"011001101",
  20051=>"011100101",
  20052=>"001001010",
  20053=>"110100000",
  20054=>"000001100",
  20055=>"101000000",
  20056=>"010001000",
  20057=>"111110111",
  20058=>"110000111",
  20059=>"100001011",
  20060=>"001010010",
  20061=>"110010010",
  20062=>"000001000",
  20063=>"110110111",
  20064=>"011100010",
  20065=>"001110001",
  20066=>"001101100",
  20067=>"111101010",
  20068=>"110100111",
  20069=>"000010000",
  20070=>"110010010",
  20071=>"000000101",
  20072=>"010101100",
  20073=>"111111011",
  20074=>"000100011",
  20075=>"011111001",
  20076=>"100000111",
  20077=>"101101001",
  20078=>"100010001",
  20079=>"001010101",
  20080=>"001001100",
  20081=>"010001011",
  20082=>"010010110",
  20083=>"100110001",
  20084=>"100011010",
  20085=>"101100111",
  20086=>"100001011",
  20087=>"101100101",
  20088=>"101101110",
  20089=>"011101111",
  20090=>"111011001",
  20091=>"001000101",
  20092=>"111100001",
  20093=>"000110010",
  20094=>"000001011",
  20095=>"110001011",
  20096=>"000001101",
  20097=>"011001100",
  20098=>"011000010",
  20099=>"010000100",
  20100=>"011001001",
  20101=>"111000011",
  20102=>"001100110",
  20103=>"011111011",
  20104=>"110011000",
  20105=>"100100101",
  20106=>"100000110",
  20107=>"100010000",
  20108=>"100101110",
  20109=>"100000100",
  20110=>"100010000",
  20111=>"110010010",
  20112=>"001001010",
  20113=>"101101001",
  20114=>"100101101",
  20115=>"110010101",
  20116=>"111110010",
  20117=>"001111101",
  20118=>"110011101",
  20119=>"111010000",
  20120=>"110110001",
  20121=>"000001001",
  20122=>"011111101",
  20123=>"111000000",
  20124=>"011000000",
  20125=>"000110111",
  20126=>"000001100",
  20127=>"011010111",
  20128=>"011011110",
  20129=>"111101100",
  20130=>"001100111",
  20131=>"010110100",
  20132=>"010001101",
  20133=>"010000110",
  20134=>"111010000",
  20135=>"000000101",
  20136=>"111001000",
  20137=>"001000110",
  20138=>"011101010",
  20139=>"101011010",
  20140=>"100111101",
  20141=>"011010110",
  20142=>"101110011",
  20143=>"001000110",
  20144=>"111110010",
  20145=>"011100111",
  20146=>"001001011",
  20147=>"011000000",
  20148=>"011101101",
  20149=>"011000100",
  20150=>"100011000",
  20151=>"101110100",
  20152=>"011000000",
  20153=>"101111000",
  20154=>"110011011",
  20155=>"001100000",
  20156=>"111001111",
  20157=>"000010101",
  20158=>"110011001",
  20159=>"000000110",
  20160=>"100110100",
  20161=>"100010100",
  20162=>"100000100",
  20163=>"000001010",
  20164=>"110110100",
  20165=>"001111000",
  20166=>"000100110",
  20167=>"010001110",
  20168=>"011101010",
  20169=>"001010011",
  20170=>"110110100",
  20171=>"010110001",
  20172=>"000001000",
  20173=>"101110011",
  20174=>"001100010",
  20175=>"100000010",
  20176=>"001000010",
  20177=>"011000110",
  20178=>"000010010",
  20179=>"110110001",
  20180=>"100110010",
  20181=>"000110010",
  20182=>"000101010",
  20183=>"100011101",
  20184=>"111001010",
  20185=>"111100101",
  20186=>"111101110",
  20187=>"001100110",
  20188=>"000000000",
  20189=>"101010101",
  20190=>"010100001",
  20191=>"001101110",
  20192=>"110001100",
  20193=>"110110001",
  20194=>"000010001",
  20195=>"110011110",
  20196=>"000101010",
  20197=>"011000011",
  20198=>"010010010",
  20199=>"110000010",
  20200=>"000110010",
  20201=>"100110111",
  20202=>"101011011",
  20203=>"101001010",
  20204=>"000110000",
  20205=>"101110001",
  20206=>"110100000",
  20207=>"110000111",
  20208=>"000010000",
  20209=>"000101110",
  20210=>"011110100",
  20211=>"110110001",
  20212=>"000010101",
  20213=>"000010000",
  20214=>"011111110",
  20215=>"011011000",
  20216=>"000011100",
  20217=>"100010100",
  20218=>"011010110",
  20219=>"101010110",
  20220=>"100011100",
  20221=>"000010011",
  20222=>"101011100",
  20223=>"111100011",
  20224=>"110110001",
  20225=>"001101101",
  20226=>"111011000",
  20227=>"000010010",
  20228=>"110011111",
  20229=>"110001000",
  20230=>"110010110",
  20231=>"101110000",
  20232=>"101110101",
  20233=>"100101111",
  20234=>"000010010",
  20235=>"100100000",
  20236=>"010101011",
  20237=>"111011101",
  20238=>"010001101",
  20239=>"100001100",
  20240=>"000011001",
  20241=>"010011100",
  20242=>"011001011",
  20243=>"001101101",
  20244=>"011011011",
  20245=>"101010111",
  20246=>"000100111",
  20247=>"011000000",
  20248=>"001100011",
  20249=>"110001100",
  20250=>"110001011",
  20251=>"110110110",
  20252=>"001111010",
  20253=>"010111110",
  20254=>"101011011",
  20255=>"100010011",
  20256=>"011000111",
  20257=>"111101111",
  20258=>"101100101",
  20259=>"010111011",
  20260=>"010001101",
  20261=>"111011101",
  20262=>"100000101",
  20263=>"111101001",
  20264=>"111001111",
  20265=>"010101001",
  20266=>"000100100",
  20267=>"100000010",
  20268=>"101001100",
  20269=>"000000000",
  20270=>"101110100",
  20271=>"001000001",
  20272=>"110001001",
  20273=>"010000111",
  20274=>"110010100",
  20275=>"001101101",
  20276=>"110011111",
  20277=>"111101111",
  20278=>"011110000",
  20279=>"111111111",
  20280=>"011000011",
  20281=>"101010011",
  20282=>"000111111",
  20283=>"100111011",
  20284=>"111110111",
  20285=>"010101011",
  20286=>"010111000",
  20287=>"011000111",
  20288=>"011110011",
  20289=>"000110000",
  20290=>"110010100",
  20291=>"100001111",
  20292=>"000101110",
  20293=>"101100000",
  20294=>"010111011",
  20295=>"111101001",
  20296=>"111001001",
  20297=>"110101001",
  20298=>"000110000",
  20299=>"111010011",
  20300=>"110001101",
  20301=>"111010110",
  20302=>"010110011",
  20303=>"001111101",
  20304=>"110101100",
  20305=>"101100011",
  20306=>"111001101",
  20307=>"001010011",
  20308=>"000110110",
  20309=>"011111110",
  20310=>"100011011",
  20311=>"010000010",
  20312=>"000100100",
  20313=>"101110001",
  20314=>"100010101",
  20315=>"011101110",
  20316=>"111001010",
  20317=>"101011101",
  20318=>"101000110",
  20319=>"110101000",
  20320=>"101010100",
  20321=>"111011001",
  20322=>"001011110",
  20323=>"010011011",
  20324=>"011101011",
  20325=>"001010011",
  20326=>"000110101",
  20327=>"111001010",
  20328=>"101011001",
  20329=>"111000111",
  20330=>"010000110",
  20331=>"111011000",
  20332=>"000110001",
  20333=>"000001100",
  20334=>"101011101",
  20335=>"111110110",
  20336=>"000100011",
  20337=>"001000011",
  20338=>"110101011",
  20339=>"010010101",
  20340=>"100001000",
  20341=>"111010000",
  20342=>"000001010",
  20343=>"101001111",
  20344=>"001010000",
  20345=>"110111100",
  20346=>"011100010",
  20347=>"101110001",
  20348=>"101010010",
  20349=>"010001110",
  20350=>"001111111",
  20351=>"111101100",
  20352=>"010011000",
  20353=>"001010111",
  20354=>"101010111",
  20355=>"000101101",
  20356=>"110011011",
  20357=>"010000010",
  20358=>"000010000",
  20359=>"011101010",
  20360=>"100110111",
  20361=>"010100101",
  20362=>"000001000",
  20363=>"101100111",
  20364=>"100010110",
  20365=>"101101011",
  20366=>"001100010",
  20367=>"111110000",
  20368=>"111010111",
  20369=>"010101110",
  20370=>"101101111",
  20371=>"101111011",
  20372=>"100000000",
  20373=>"110111100",
  20374=>"000000100",
  20375=>"100001000",
  20376=>"010101000",
  20377=>"101101111",
  20378=>"011100101",
  20379=>"011000111",
  20380=>"011010011",
  20381=>"110110100",
  20382=>"000101110",
  20383=>"000111101",
  20384=>"000000110",
  20385=>"100010001",
  20386=>"001000000",
  20387=>"010001111",
  20388=>"111000111",
  20389=>"001101110",
  20390=>"110000000",
  20391=>"000110010",
  20392=>"000100100",
  20393=>"101110011",
  20394=>"000100000",
  20395=>"010111110",
  20396=>"111001001",
  20397=>"111111110",
  20398=>"000011001",
  20399=>"001000101",
  20400=>"000100000",
  20401=>"111100110",
  20402=>"101111011",
  20403=>"110001010",
  20404=>"110110111",
  20405=>"100100010",
  20406=>"001011101",
  20407=>"001100100",
  20408=>"011110111",
  20409=>"010000010",
  20410=>"100111010",
  20411=>"110110111",
  20412=>"100000110",
  20413=>"110110000",
  20414=>"110101000",
  20415=>"010110001",
  20416=>"000110101",
  20417=>"000001000",
  20418=>"000110101",
  20419=>"000110001",
  20420=>"000000110",
  20421=>"101111000",
  20422=>"011000011",
  20423=>"100010011",
  20424=>"110001100",
  20425=>"000110010",
  20426=>"000010001",
  20427=>"111000101",
  20428=>"100011110",
  20429=>"110101100",
  20430=>"000011101",
  20431=>"010001010",
  20432=>"010101100",
  20433=>"100001001",
  20434=>"101100011",
  20435=>"110000001",
  20436=>"111010111",
  20437=>"000111010",
  20438=>"011011000",
  20439=>"111111111",
  20440=>"010111000",
  20441=>"110000000",
  20442=>"110011000",
  20443=>"010011010",
  20444=>"001011101",
  20445=>"000010001",
  20446=>"000010110",
  20447=>"000100110",
  20448=>"010101111",
  20449=>"110011101",
  20450=>"011101100",
  20451=>"010100100",
  20452=>"111100011",
  20453=>"110111000",
  20454=>"101010010",
  20455=>"010100000",
  20456=>"001000011",
  20457=>"010010111",
  20458=>"101011101",
  20459=>"110010110",
  20460=>"010010001",
  20461=>"101001001",
  20462=>"111110111",
  20463=>"000110100",
  20464=>"010111011",
  20465=>"111110101",
  20466=>"100100011",
  20467=>"010010011",
  20468=>"001110000",
  20469=>"000101111",
  20470=>"111011101",
  20471=>"110011100",
  20472=>"001010100",
  20473=>"000100010",
  20474=>"000001111",
  20475=>"100010000",
  20476=>"000011100",
  20477=>"101100010",
  20478=>"001110011",
  20479=>"110100000",
  20480=>"100001100",
  20481=>"000001001",
  20482=>"111101111",
  20483=>"010010111",
  20484=>"010001110",
  20485=>"101010110",
  20486=>"001101111",
  20487=>"001000010",
  20488=>"001100001",
  20489=>"000011000",
  20490=>"011101000",
  20491=>"100101100",
  20492=>"101110011",
  20493=>"010000100",
  20494=>"100001011",
  20495=>"111110110",
  20496=>"111101111",
  20497=>"101100000",
  20498=>"100101000",
  20499=>"110110110",
  20500=>"111001001",
  20501=>"000111111",
  20502=>"111111001",
  20503=>"011000011",
  20504=>"010101111",
  20505=>"011110111",
  20506=>"011100011",
  20507=>"010100010",
  20508=>"000001101",
  20509=>"111011011",
  20510=>"110111010",
  20511=>"111000101",
  20512=>"001001101",
  20513=>"001111011",
  20514=>"100011000",
  20515=>"010111000",
  20516=>"110011010",
  20517=>"010110100",
  20518=>"100100010",
  20519=>"100101011",
  20520=>"000100010",
  20521=>"000110011",
  20522=>"111111110",
  20523=>"100000100",
  20524=>"000010110",
  20525=>"000011111",
  20526=>"100110011",
  20527=>"001111101",
  20528=>"001110110",
  20529=>"111001101",
  20530=>"101000001",
  20531=>"110101111",
  20532=>"000001010",
  20533=>"110001010",
  20534=>"010011101",
  20535=>"001110001",
  20536=>"000001100",
  20537=>"000000011",
  20538=>"000010110",
  20539=>"101100101",
  20540=>"111001001",
  20541=>"010011011",
  20542=>"100000111",
  20543=>"111001011",
  20544=>"100001101",
  20545=>"010010000",
  20546=>"010110001",
  20547=>"000000101",
  20548=>"000001101",
  20549=>"100001011",
  20550=>"101011101",
  20551=>"110000111",
  20552=>"100111011",
  20553=>"000101011",
  20554=>"001011100",
  20555=>"111001011",
  20556=>"110001100",
  20557=>"110000000",
  20558=>"010010110",
  20559=>"010100000",
  20560=>"110000010",
  20561=>"010110010",
  20562=>"011100101",
  20563=>"101001110",
  20564=>"111000000",
  20565=>"000100000",
  20566=>"101001011",
  20567=>"000101100",
  20568=>"000001100",
  20569=>"110011101",
  20570=>"100000000",
  20571=>"010000100",
  20572=>"101101101",
  20573=>"100000110",
  20574=>"011000000",
  20575=>"001110111",
  20576=>"011111011",
  20577=>"100110110",
  20578=>"110001000",
  20579=>"101011011",
  20580=>"111100001",
  20581=>"011000110",
  20582=>"101110010",
  20583=>"111011001",
  20584=>"010011110",
  20585=>"001111001",
  20586=>"100101111",
  20587=>"111110100",
  20588=>"011101111",
  20589=>"011100101",
  20590=>"100001110",
  20591=>"011001111",
  20592=>"100000101",
  20593=>"000111101",
  20594=>"001101111",
  20595=>"010101011",
  20596=>"000010000",
  20597=>"110101100",
  20598=>"011011001",
  20599=>"010111010",
  20600=>"000111011",
  20601=>"101110100",
  20602=>"011110010",
  20603=>"110100100",
  20604=>"101000000",
  20605=>"000100111",
  20606=>"101011000",
  20607=>"100111011",
  20608=>"101111111",
  20609=>"000101110",
  20610=>"011101110",
  20611=>"010000100",
  20612=>"001000101",
  20613=>"011000010",
  20614=>"110001100",
  20615=>"010000000",
  20616=>"010100110",
  20617=>"010111110",
  20618=>"100010011",
  20619=>"000101000",
  20620=>"000000101",
  20621=>"111001101",
  20622=>"000110111",
  20623=>"000110001",
  20624=>"011100010",
  20625=>"011110101",
  20626=>"001110101",
  20627=>"010001010",
  20628=>"101011100",
  20629=>"101101001",
  20630=>"101100110",
  20631=>"101001100",
  20632=>"010010001",
  20633=>"101000000",
  20634=>"101011101",
  20635=>"111111000",
  20636=>"001001001",
  20637=>"100101001",
  20638=>"001111111",
  20639=>"111100110",
  20640=>"110111101",
  20641=>"110111110",
  20642=>"000000001",
  20643=>"010110001",
  20644=>"100011110",
  20645=>"001011111",
  20646=>"001011101",
  20647=>"111101111",
  20648=>"101100111",
  20649=>"001101010",
  20650=>"001101011",
  20651=>"010000001",
  20652=>"011100101",
  20653=>"010001111",
  20654=>"011001101",
  20655=>"011111011",
  20656=>"001000101",
  20657=>"011000000",
  20658=>"101000000",
  20659=>"100101011",
  20660=>"011101111",
  20661=>"110011001",
  20662=>"101111101",
  20663=>"000111001",
  20664=>"000010111",
  20665=>"001010111",
  20666=>"110011010",
  20667=>"000010110",
  20668=>"110010011",
  20669=>"110010111",
  20670=>"001110010",
  20671=>"000101100",
  20672=>"110100001",
  20673=>"001000011",
  20674=>"101101000",
  20675=>"011011010",
  20676=>"000100010",
  20677=>"001010011",
  20678=>"111111111",
  20679=>"000111010",
  20680=>"001011001",
  20681=>"010010110",
  20682=>"101010110",
  20683=>"001000011",
  20684=>"000111010",
  20685=>"011100111",
  20686=>"111001110",
  20687=>"010100101",
  20688=>"101111011",
  20689=>"101100000",
  20690=>"001001000",
  20691=>"000001000",
  20692=>"011001101",
  20693=>"011010000",
  20694=>"001011101",
  20695=>"110111111",
  20696=>"011011000",
  20697=>"001100010",
  20698=>"100000000",
  20699=>"011001100",
  20700=>"100011100",
  20701=>"110100010",
  20702=>"101110100",
  20703=>"101111010",
  20704=>"100001000",
  20705=>"001101001",
  20706=>"011001100",
  20707=>"100000001",
  20708=>"000011001",
  20709=>"101011100",
  20710=>"010011101",
  20711=>"010010000",
  20712=>"101001001",
  20713=>"011001010",
  20714=>"011110010",
  20715=>"010101000",
  20716=>"010110011",
  20717=>"100001101",
  20718=>"010001011",
  20719=>"001010100",
  20720=>"110010011",
  20721=>"011110100",
  20722=>"100001100",
  20723=>"111011110",
  20724=>"110111000",
  20725=>"010011011",
  20726=>"100000110",
  20727=>"001100110",
  20728=>"101101100",
  20729=>"000001111",
  20730=>"001000110",
  20731=>"011001011",
  20732=>"011100101",
  20733=>"010011111",
  20734=>"110010101",
  20735=>"111000111",
  20736=>"001111111",
  20737=>"001000110",
  20738=>"001011111",
  20739=>"000111110",
  20740=>"100011011",
  20741=>"010100000",
  20742=>"001110000",
  20743=>"111000011",
  20744=>"111100010",
  20745=>"101101100",
  20746=>"111100101",
  20747=>"010001001",
  20748=>"111101000",
  20749=>"011110111",
  20750=>"101000111",
  20751=>"010001000",
  20752=>"001111001",
  20753=>"010110100",
  20754=>"011001010",
  20755=>"000110000",
  20756=>"001110001",
  20757=>"000001110",
  20758=>"010001010",
  20759=>"000101010",
  20760=>"011001010",
  20761=>"001010111",
  20762=>"100110000",
  20763=>"100000100",
  20764=>"000110101",
  20765=>"011101111",
  20766=>"000110111",
  20767=>"110001000",
  20768=>"010010111",
  20769=>"111011101",
  20770=>"110110011",
  20771=>"100010101",
  20772=>"001101101",
  20773=>"011110010",
  20774=>"110000010",
  20775=>"011000100",
  20776=>"111011111",
  20777=>"000111011",
  20778=>"110010000",
  20779=>"010101111",
  20780=>"001011010",
  20781=>"001100000",
  20782=>"010000101",
  20783=>"100011011",
  20784=>"100101100",
  20785=>"001111101",
  20786=>"110110011",
  20787=>"111111111",
  20788=>"000011111",
  20789=>"100100111",
  20790=>"110110011",
  20791=>"000011010",
  20792=>"111001101",
  20793=>"010010001",
  20794=>"101011110",
  20795=>"100000111",
  20796=>"110111010",
  20797=>"001011100",
  20798=>"111000010",
  20799=>"111111001",
  20800=>"100011110",
  20801=>"010000011",
  20802=>"001110001",
  20803=>"101101101",
  20804=>"111000101",
  20805=>"111101010",
  20806=>"011010100",
  20807=>"101111011",
  20808=>"110000010",
  20809=>"101010110",
  20810=>"010000010",
  20811=>"000011110",
  20812=>"110010010",
  20813=>"011101001",
  20814=>"101000111",
  20815=>"101100111",
  20816=>"111001011",
  20817=>"111010001",
  20818=>"011001100",
  20819=>"111100100",
  20820=>"100010001",
  20821=>"111111011",
  20822=>"101001111",
  20823=>"000101111",
  20824=>"100111100",
  20825=>"001000000",
  20826=>"000011110",
  20827=>"000000001",
  20828=>"110001101",
  20829=>"010010110",
  20830=>"001110111",
  20831=>"101111101",
  20832=>"001001100",
  20833=>"011001100",
  20834=>"111100110",
  20835=>"110000010",
  20836=>"101110010",
  20837=>"010101101",
  20838=>"101110100",
  20839=>"011111111",
  20840=>"100010000",
  20841=>"000011110",
  20842=>"110111101",
  20843=>"000110110",
  20844=>"111011111",
  20845=>"111000010",
  20846=>"010111101",
  20847=>"001000001",
  20848=>"111110001",
  20849=>"000101001",
  20850=>"010100110",
  20851=>"111110001",
  20852=>"111110101",
  20853=>"111101101",
  20854=>"111110101",
  20855=>"000001010",
  20856=>"011110001",
  20857=>"011110001",
  20858=>"111000011",
  20859=>"110100011",
  20860=>"011101000",
  20861=>"100010001",
  20862=>"000100001",
  20863=>"010010101",
  20864=>"111000111",
  20865=>"100101011",
  20866=>"111100000",
  20867=>"001110110",
  20868=>"100100111",
  20869=>"000111001",
  20870=>"110110011",
  20871=>"000111111",
  20872=>"111111111",
  20873=>"110101101",
  20874=>"110100010",
  20875=>"111110011",
  20876=>"000100111",
  20877=>"000101101",
  20878=>"001010111",
  20879=>"111111000",
  20880=>"001010011",
  20881=>"111111001",
  20882=>"111010000",
  20883=>"111100101",
  20884=>"100001111",
  20885=>"100011111",
  20886=>"100111101",
  20887=>"110100110",
  20888=>"000000010",
  20889=>"001000110",
  20890=>"111100111",
  20891=>"100011010",
  20892=>"010011011",
  20893=>"101001011",
  20894=>"100101101",
  20895=>"100110101",
  20896=>"001000001",
  20897=>"110010001",
  20898=>"000110110",
  20899=>"111010001",
  20900=>"101011011",
  20901=>"110100100",
  20902=>"000101010",
  20903=>"000111111",
  20904=>"000000010",
  20905=>"110010001",
  20906=>"111011011",
  20907=>"111111111",
  20908=>"101011101",
  20909=>"100001000",
  20910=>"010110001",
  20911=>"111011101",
  20912=>"111111111",
  20913=>"000100101",
  20914=>"000100000",
  20915=>"001011000",
  20916=>"000111011",
  20917=>"011010110",
  20918=>"101011000",
  20919=>"111100010",
  20920=>"000111111",
  20921=>"110000110",
  20922=>"100101110",
  20923=>"101011111",
  20924=>"001100000",
  20925=>"000000100",
  20926=>"110010100",
  20927=>"111000001",
  20928=>"000010111",
  20929=>"101010010",
  20930=>"111101111",
  20931=>"110110100",
  20932=>"011011111",
  20933=>"010100011",
  20934=>"101100110",
  20935=>"010000111",
  20936=>"111001011",
  20937=>"101011001",
  20938=>"111111101",
  20939=>"000100011",
  20940=>"101110001",
  20941=>"100111101",
  20942=>"100000000",
  20943=>"100100101",
  20944=>"101101100",
  20945=>"111101100",
  20946=>"010001000",
  20947=>"100001111",
  20948=>"100001100",
  20949=>"100101100",
  20950=>"111101111",
  20951=>"000000000",
  20952=>"001011111",
  20953=>"110100111",
  20954=>"001110010",
  20955=>"001101011",
  20956=>"000000010",
  20957=>"101000000",
  20958=>"000100101",
  20959=>"110011101",
  20960=>"111011110",
  20961=>"000010001",
  20962=>"000011001",
  20963=>"110001110",
  20964=>"111100001",
  20965=>"011000000",
  20966=>"101011100",
  20967=>"010001001",
  20968=>"000110110",
  20969=>"110100010",
  20970=>"100000000",
  20971=>"000000001",
  20972=>"000010010",
  20973=>"000010101",
  20974=>"110110000",
  20975=>"010000111",
  20976=>"010110100",
  20977=>"000010011",
  20978=>"010000111",
  20979=>"000101111",
  20980=>"110010011",
  20981=>"011011000",
  20982=>"010011010",
  20983=>"000100100",
  20984=>"111100111",
  20985=>"011001111",
  20986=>"010111111",
  20987=>"010001101",
  20988=>"110110010",
  20989=>"000111100",
  20990=>"001100111",
  20991=>"101000110",
  20992=>"101000011",
  20993=>"110010010",
  20994=>"111000011",
  20995=>"100111110",
  20996=>"110001010",
  20997=>"101010001",
  20998=>"110000000",
  20999=>"011001010",
  21000=>"010000011",
  21001=>"101110100",
  21002=>"011010001",
  21003=>"011110001",
  21004=>"011010001",
  21005=>"110111011",
  21006=>"000011011",
  21007=>"010000100",
  21008=>"101111001",
  21009=>"111101110",
  21010=>"111101011",
  21011=>"101100001",
  21012=>"011100011",
  21013=>"100000001",
  21014=>"101110001",
  21015=>"100101100",
  21016=>"101010101",
  21017=>"001110101",
  21018=>"010110000",
  21019=>"100111101",
  21020=>"011010001",
  21021=>"101000000",
  21022=>"010110000",
  21023=>"001010001",
  21024=>"010111001",
  21025=>"100111101",
  21026=>"000000001",
  21027=>"111100100",
  21028=>"001001010",
  21029=>"010000010",
  21030=>"111101010",
  21031=>"110011110",
  21032=>"011001010",
  21033=>"010000110",
  21034=>"101110010",
  21035=>"001010001",
  21036=>"101010011",
  21037=>"111101101",
  21038=>"001010011",
  21039=>"110010110",
  21040=>"011101111",
  21041=>"010010001",
  21042=>"000011001",
  21043=>"000101000",
  21044=>"010101101",
  21045=>"001010000",
  21046=>"010000011",
  21047=>"001000000",
  21048=>"001000011",
  21049=>"101110010",
  21050=>"101000110",
  21051=>"000010011",
  21052=>"001011001",
  21053=>"101111110",
  21054=>"110010100",
  21055=>"000000001",
  21056=>"010100101",
  21057=>"101100110",
  21058=>"000100111",
  21059=>"000100100",
  21060=>"010100101",
  21061=>"010000011",
  21062=>"110010101",
  21063=>"100000000",
  21064=>"101001101",
  21065=>"011000110",
  21066=>"111101110",
  21067=>"001111000",
  21068=>"010000001",
  21069=>"000001000",
  21070=>"001100011",
  21071=>"010010100",
  21072=>"000011000",
  21073=>"111110101",
  21074=>"110000111",
  21075=>"001010100",
  21076=>"111001111",
  21077=>"001010010",
  21078=>"011110111",
  21079=>"010011001",
  21080=>"101000010",
  21081=>"011010011",
  21082=>"011011111",
  21083=>"111011011",
  21084=>"111100010",
  21085=>"001001100",
  21086=>"100010101",
  21087=>"001101010",
  21088=>"010000001",
  21089=>"101010000",
  21090=>"100110111",
  21091=>"001011011",
  21092=>"100111100",
  21093=>"111010001",
  21094=>"111101100",
  21095=>"001001011",
  21096=>"100000000",
  21097=>"011000111",
  21098=>"111101101",
  21099=>"000001011",
  21100=>"001110111",
  21101=>"011011011",
  21102=>"100110101",
  21103=>"011010100",
  21104=>"101100010",
  21105=>"101111001",
  21106=>"011100010",
  21107=>"011011001",
  21108=>"010110000",
  21109=>"010110111",
  21110=>"111110011",
  21111=>"111110101",
  21112=>"110111110",
  21113=>"001110000",
  21114=>"010110101",
  21115=>"100111100",
  21116=>"010000111",
  21117=>"001010000",
  21118=>"000011011",
  21119=>"001011101",
  21120=>"101101011",
  21121=>"011101101",
  21122=>"111110001",
  21123=>"011100000",
  21124=>"100010001",
  21125=>"101111000",
  21126=>"011011010",
  21127=>"010000100",
  21128=>"000100000",
  21129=>"101001010",
  21130=>"111000101",
  21131=>"011001110",
  21132=>"110001001",
  21133=>"011000011",
  21134=>"101011111",
  21135=>"110101001",
  21136=>"111111100",
  21137=>"100001000",
  21138=>"101000101",
  21139=>"111001111",
  21140=>"010001101",
  21141=>"110101101",
  21142=>"101110110",
  21143=>"100100110",
  21144=>"110111111",
  21145=>"000100001",
  21146=>"100100011",
  21147=>"111001000",
  21148=>"010101111",
  21149=>"110100000",
  21150=>"010001001",
  21151=>"111111001",
  21152=>"111111111",
  21153=>"011111101",
  21154=>"000111110",
  21155=>"111110001",
  21156=>"100101011",
  21157=>"101101111",
  21158=>"111111010",
  21159=>"111101101",
  21160=>"000111010",
  21161=>"111001111",
  21162=>"000110101",
  21163=>"010001000",
  21164=>"000111101",
  21165=>"101101000",
  21166=>"001111011",
  21167=>"000001100",
  21168=>"111000001",
  21169=>"011110010",
  21170=>"010010001",
  21171=>"111001001",
  21172=>"010011011",
  21173=>"001110111",
  21174=>"001101110",
  21175=>"110111000",
  21176=>"101000011",
  21177=>"011101111",
  21178=>"000001001",
  21179=>"001111100",
  21180=>"000010110",
  21181=>"001001000",
  21182=>"100011100",
  21183=>"111000001",
  21184=>"011101001",
  21185=>"010000000",
  21186=>"100101001",
  21187=>"110011110",
  21188=>"000100000",
  21189=>"101100101",
  21190=>"111011100",
  21191=>"100100100",
  21192=>"110001000",
  21193=>"000000000",
  21194=>"100111101",
  21195=>"100110001",
  21196=>"000011100",
  21197=>"000100010",
  21198=>"111111011",
  21199=>"010001001",
  21200=>"000011010",
  21201=>"101101100",
  21202=>"000011111",
  21203=>"101011011",
  21204=>"000011011",
  21205=>"001111000",
  21206=>"000010111",
  21207=>"001100010",
  21208=>"001100101",
  21209=>"011101101",
  21210=>"000011001",
  21211=>"011011010",
  21212=>"100001001",
  21213=>"011011010",
  21214=>"010000110",
  21215=>"110111000",
  21216=>"110100001",
  21217=>"110110000",
  21218=>"100010010",
  21219=>"110111110",
  21220=>"110111001",
  21221=>"011010111",
  21222=>"110010101",
  21223=>"111110111",
  21224=>"110010000",
  21225=>"010000111",
  21226=>"100110001",
  21227=>"001010000",
  21228=>"100111011",
  21229=>"000000001",
  21230=>"100111001",
  21231=>"000010111",
  21232=>"001110001",
  21233=>"011000010",
  21234=>"011101001",
  21235=>"110011010",
  21236=>"010001100",
  21237=>"011011101",
  21238=>"000010100",
  21239=>"111111111",
  21240=>"101111100",
  21241=>"011100110",
  21242=>"111100011",
  21243=>"111010000",
  21244=>"100110001",
  21245=>"110000100",
  21246=>"111100001",
  21247=>"110010001",
  21248=>"111011010",
  21249=>"011110001",
  21250=>"110010111",
  21251=>"100010011",
  21252=>"001110011",
  21253=>"000100111",
  21254=>"110111000",
  21255=>"100111000",
  21256=>"100111001",
  21257=>"010010101",
  21258=>"011100000",
  21259=>"110111101",
  21260=>"001011110",
  21261=>"111101100",
  21262=>"001000110",
  21263=>"001010111",
  21264=>"001011011",
  21265=>"110010100",
  21266=>"010111010",
  21267=>"111011011",
  21268=>"011010001",
  21269=>"110011011",
  21270=>"111001100",
  21271=>"111111110",
  21272=>"101100111",
  21273=>"111011011",
  21274=>"100000001",
  21275=>"111001000",
  21276=>"100101111",
  21277=>"110101010",
  21278=>"000000101",
  21279=>"011001001",
  21280=>"011101000",
  21281=>"101000000",
  21282=>"011001101",
  21283=>"101111111",
  21284=>"101110101",
  21285=>"010111101",
  21286=>"000010100",
  21287=>"111001001",
  21288=>"111001110",
  21289=>"100100000",
  21290=>"000101010",
  21291=>"100100010",
  21292=>"010111000",
  21293=>"001000100",
  21294=>"110001000",
  21295=>"111010001",
  21296=>"010101010",
  21297=>"010010101",
  21298=>"011010011",
  21299=>"110001110",
  21300=>"011011010",
  21301=>"101011000",
  21302=>"010001000",
  21303=>"010011011",
  21304=>"110000100",
  21305=>"001100100",
  21306=>"100100110",
  21307=>"100000000",
  21308=>"001111101",
  21309=>"001010111",
  21310=>"010011001",
  21311=>"110010001",
  21312=>"111010101",
  21313=>"010010000",
  21314=>"100110000",
  21315=>"000011010",
  21316=>"010010100",
  21317=>"000001000",
  21318=>"011011110",
  21319=>"000101001",
  21320=>"000101110",
  21321=>"010101010",
  21322=>"100010011",
  21323=>"011001010",
  21324=>"110100010",
  21325=>"110010110",
  21326=>"111101100",
  21327=>"010001000",
  21328=>"111001011",
  21329=>"000000010",
  21330=>"001000011",
  21331=>"001001101",
  21332=>"001010111",
  21333=>"111001110",
  21334=>"010001001",
  21335=>"101111100",
  21336=>"110110001",
  21337=>"000000001",
  21338=>"011010010",
  21339=>"000001111",
  21340=>"011101011",
  21341=>"010110100",
  21342=>"011011000",
  21343=>"001001101",
  21344=>"100100000",
  21345=>"001101111",
  21346=>"111100101",
  21347=>"101010111",
  21348=>"001110111",
  21349=>"010101101",
  21350=>"000110100",
  21351=>"111000111",
  21352=>"111110010",
  21353=>"110111100",
  21354=>"110110110",
  21355=>"101100100",
  21356=>"001000111",
  21357=>"110011011",
  21358=>"111100101",
  21359=>"000001011",
  21360=>"001001000",
  21361=>"010101000",
  21362=>"111101110",
  21363=>"111110110",
  21364=>"001101111",
  21365=>"101101101",
  21366=>"000001001",
  21367=>"101011001",
  21368=>"001111110",
  21369=>"101110100",
  21370=>"101011110",
  21371=>"111011001",
  21372=>"100001100",
  21373=>"111011111",
  21374=>"110001110",
  21375=>"110110010",
  21376=>"110011011",
  21377=>"000100000",
  21378=>"001100010",
  21379=>"010110011",
  21380=>"101110011",
  21381=>"010000101",
  21382=>"011011111",
  21383=>"111010001",
  21384=>"110000010",
  21385=>"101001111",
  21386=>"001111100",
  21387=>"100000100",
  21388=>"101000111",
  21389=>"100111011",
  21390=>"101000110",
  21391=>"110111011",
  21392=>"000101010",
  21393=>"101000101",
  21394=>"011010010",
  21395=>"100000001",
  21396=>"011011011",
  21397=>"011001100",
  21398=>"100000111",
  21399=>"000001110",
  21400=>"110011011",
  21401=>"100000001",
  21402=>"101000111",
  21403=>"101111100",
  21404=>"100001001",
  21405=>"000010101",
  21406=>"110110001",
  21407=>"001000101",
  21408=>"110100111",
  21409=>"000101111",
  21410=>"001000000",
  21411=>"001100011",
  21412=>"001110110",
  21413=>"111010001",
  21414=>"000001111",
  21415=>"011010000",
  21416=>"010111011",
  21417=>"111111111",
  21418=>"110101010",
  21419=>"110011000",
  21420=>"000010110",
  21421=>"110101100",
  21422=>"111010010",
  21423=>"001011001",
  21424=>"100101101",
  21425=>"100011101",
  21426=>"000101010",
  21427=>"001101110",
  21428=>"111111010",
  21429=>"110101101",
  21430=>"100111011",
  21431=>"011101000",
  21432=>"100100010",
  21433=>"100001101",
  21434=>"000010110",
  21435=>"010100100",
  21436=>"001000111",
  21437=>"000010110",
  21438=>"111111001",
  21439=>"000000111",
  21440=>"001100001",
  21441=>"001000001",
  21442=>"100110001",
  21443=>"010111011",
  21444=>"000110001",
  21445=>"011001000",
  21446=>"111011101",
  21447=>"010011110",
  21448=>"010000000",
  21449=>"011101000",
  21450=>"111100011",
  21451=>"101101111",
  21452=>"101000011",
  21453=>"100000110",
  21454=>"011110010",
  21455=>"100010101",
  21456=>"000101000",
  21457=>"010110111",
  21458=>"110110010",
  21459=>"010001010",
  21460=>"001000010",
  21461=>"001010000",
  21462=>"111100110",
  21463=>"110000100",
  21464=>"010000100",
  21465=>"000011100",
  21466=>"101100110",
  21467=>"101011111",
  21468=>"010001001",
  21469=>"000000101",
  21470=>"100101100",
  21471=>"011101111",
  21472=>"100001110",
  21473=>"110101101",
  21474=>"010011010",
  21475=>"110100011",
  21476=>"100000010",
  21477=>"010000000",
  21478=>"111100000",
  21479=>"101101001",
  21480=>"011110011",
  21481=>"000000111",
  21482=>"001001001",
  21483=>"110100001",
  21484=>"101100000",
  21485=>"000100010",
  21486=>"100010100",
  21487=>"111111001",
  21488=>"000011000",
  21489=>"001001111",
  21490=>"111000010",
  21491=>"110110000",
  21492=>"111101100",
  21493=>"000011010",
  21494=>"110101100",
  21495=>"011001001",
  21496=>"100011000",
  21497=>"100001110",
  21498=>"011100010",
  21499=>"011110001",
  21500=>"110000111",
  21501=>"100100110",
  21502=>"100011111",
  21503=>"100101100",
  21504=>"010100011",
  21505=>"110111001",
  21506=>"100010110",
  21507=>"101110000",
  21508=>"000111010",
  21509=>"111110101",
  21510=>"010111011",
  21511=>"111110000",
  21512=>"111001000",
  21513=>"001001100",
  21514=>"000101101",
  21515=>"100001010",
  21516=>"111110001",
  21517=>"111101000",
  21518=>"111110111",
  21519=>"100111101",
  21520=>"001100011",
  21521=>"011110001",
  21522=>"101011011",
  21523=>"010011111",
  21524=>"010000110",
  21525=>"100111110",
  21526=>"100100101",
  21527=>"000000111",
  21528=>"000001010",
  21529=>"110010010",
  21530=>"111101111",
  21531=>"000100000",
  21532=>"010010101",
  21533=>"111000100",
  21534=>"101011010",
  21535=>"011110000",
  21536=>"111100011",
  21537=>"110100111",
  21538=>"010100101",
  21539=>"100010011",
  21540=>"101110001",
  21541=>"000001000",
  21542=>"010011010",
  21543=>"101011110",
  21544=>"010000000",
  21545=>"000011111",
  21546=>"001011011",
  21547=>"011110100",
  21548=>"001100011",
  21549=>"000110101",
  21550=>"101000000",
  21551=>"101011100",
  21552=>"110111111",
  21553=>"101011000",
  21554=>"101110111",
  21555=>"000101000",
  21556=>"100000111",
  21557=>"000110110",
  21558=>"101000001",
  21559=>"000111101",
  21560=>"000000000",
  21561=>"110101010",
  21562=>"000110000",
  21563=>"101001000",
  21564=>"101000010",
  21565=>"000101000",
  21566=>"101101000",
  21567=>"110011111",
  21568=>"101011100",
  21569=>"000111001",
  21570=>"100101000",
  21571=>"011011101",
  21572=>"101111010",
  21573=>"100110100",
  21574=>"100010110",
  21575=>"101011000",
  21576=>"001101111",
  21577=>"011000101",
  21578=>"001011101",
  21579=>"010111000",
  21580=>"101000001",
  21581=>"101100000",
  21582=>"011100111",
  21583=>"001001011",
  21584=>"000110010",
  21585=>"011011011",
  21586=>"000111101",
  21587=>"111111111",
  21588=>"111110000",
  21589=>"000001100",
  21590=>"011110000",
  21591=>"100100000",
  21592=>"111000101",
  21593=>"111011110",
  21594=>"001001010",
  21595=>"111101101",
  21596=>"001010010",
  21597=>"110110000",
  21598=>"011111001",
  21599=>"110110100",
  21600=>"001000101",
  21601=>"001000011",
  21602=>"100100111",
  21603=>"011001010",
  21604=>"000010111",
  21605=>"101111110",
  21606=>"101111111",
  21607=>"010000101",
  21608=>"111111000",
  21609=>"100101000",
  21610=>"110111111",
  21611=>"001101001",
  21612=>"100010011",
  21613=>"001110111",
  21614=>"111111000",
  21615=>"010101010",
  21616=>"010000000",
  21617=>"000000111",
  21618=>"001100101",
  21619=>"001011011",
  21620=>"010001110",
  21621=>"001110101",
  21622=>"111110000",
  21623=>"001100010",
  21624=>"010011010",
  21625=>"001101110",
  21626=>"000000100",
  21627=>"001111001",
  21628=>"000111111",
  21629=>"101001001",
  21630=>"001000000",
  21631=>"100011010",
  21632=>"001101100",
  21633=>"001000101",
  21634=>"001000010",
  21635=>"101000000",
  21636=>"100001001",
  21637=>"000101111",
  21638=>"111111111",
  21639=>"101111101",
  21640=>"000000100",
  21641=>"011001000",
  21642=>"110000000",
  21643=>"101101110",
  21644=>"110000101",
  21645=>"110101110",
  21646=>"111011100",
  21647=>"100111101",
  21648=>"000001110",
  21649=>"101110000",
  21650=>"110101101",
  21651=>"111110101",
  21652=>"101111001",
  21653=>"111011101",
  21654=>"010010001",
  21655=>"000110100",
  21656=>"011110100",
  21657=>"111100110",
  21658=>"110110100",
  21659=>"011001100",
  21660=>"111010001",
  21661=>"011010110",
  21662=>"000000101",
  21663=>"101000100",
  21664=>"001111101",
  21665=>"000001111",
  21666=>"010100110",
  21667=>"101001001",
  21668=>"101000111",
  21669=>"100110111",
  21670=>"000001010",
  21671=>"111010100",
  21672=>"000111000",
  21673=>"001011010",
  21674=>"010010010",
  21675=>"011101100",
  21676=>"101111001",
  21677=>"111111001",
  21678=>"000110011",
  21679=>"001000110",
  21680=>"100011101",
  21681=>"000011111",
  21682=>"101000010",
  21683=>"010111100",
  21684=>"110001101",
  21685=>"000011100",
  21686=>"011111110",
  21687=>"000000110",
  21688=>"001011001",
  21689=>"011011011",
  21690=>"100001010",
  21691=>"111100101",
  21692=>"011111001",
  21693=>"101001000",
  21694=>"011001111",
  21695=>"100100110",
  21696=>"000101111",
  21697=>"110111100",
  21698=>"001100011",
  21699=>"101100100",
  21700=>"111111100",
  21701=>"111101111",
  21702=>"111111110",
  21703=>"110110000",
  21704=>"101011110",
  21705=>"000010100",
  21706=>"001110111",
  21707=>"001011101",
  21708=>"110001000",
  21709=>"011111011",
  21710=>"000101011",
  21711=>"001100001",
  21712=>"010011011",
  21713=>"010110001",
  21714=>"010100000",
  21715=>"001001010",
  21716=>"011101010",
  21717=>"111111101",
  21718=>"010000101",
  21719=>"001100000",
  21720=>"100001010",
  21721=>"001111011",
  21722=>"110111101",
  21723=>"110011101",
  21724=>"001101000",
  21725=>"000111110",
  21726=>"001001110",
  21727=>"000101000",
  21728=>"101111001",
  21729=>"000001010",
  21730=>"001011100",
  21731=>"000001110",
  21732=>"101001100",
  21733=>"100101111",
  21734=>"001011101",
  21735=>"010100011",
  21736=>"101010111",
  21737=>"001100111",
  21738=>"001011111",
  21739=>"001001111",
  21740=>"000010101",
  21741=>"110100001",
  21742=>"101101000",
  21743=>"000100001",
  21744=>"100000010",
  21745=>"110111010",
  21746=>"100101010",
  21747=>"101100100",
  21748=>"111011111",
  21749=>"000010010",
  21750=>"111110001",
  21751=>"011111111",
  21752=>"000111101",
  21753=>"100000011",
  21754=>"001110110",
  21755=>"111110110",
  21756=>"100000010",
  21757=>"011100000",
  21758=>"100000110",
  21759=>"001000100",
  21760=>"110011010",
  21761=>"000011111",
  21762=>"110001101",
  21763=>"001100100",
  21764=>"001011101",
  21765=>"010110010",
  21766=>"111010000",
  21767=>"111010001",
  21768=>"100011101",
  21769=>"011101010",
  21770=>"011100010",
  21771=>"001011000",
  21772=>"001100111",
  21773=>"000111000",
  21774=>"000110101",
  21775=>"010000000",
  21776=>"011010111",
  21777=>"100111110",
  21778=>"101111011",
  21779=>"110001001",
  21780=>"000001110",
  21781=>"010000000",
  21782=>"000001110",
  21783=>"101110001",
  21784=>"110011100",
  21785=>"000011010",
  21786=>"001010101",
  21787=>"000100001",
  21788=>"110010000",
  21789=>"111010000",
  21790=>"001001001",
  21791=>"100000100",
  21792=>"111110111",
  21793=>"100010100",
  21794=>"101101010",
  21795=>"100111010",
  21796=>"001001010",
  21797=>"000101011",
  21798=>"010000000",
  21799=>"000000001",
  21800=>"100011101",
  21801=>"101001001",
  21802=>"001000110",
  21803=>"001100001",
  21804=>"111001100",
  21805=>"000001000",
  21806=>"001100010",
  21807=>"101010001",
  21808=>"010001011",
  21809=>"010000001",
  21810=>"000101010",
  21811=>"110111111",
  21812=>"000100010",
  21813=>"011000110",
  21814=>"101010000",
  21815=>"110001101",
  21816=>"100100001",
  21817=>"010111111",
  21818=>"101001011",
  21819=>"101000000",
  21820=>"111101111",
  21821=>"111111000",
  21822=>"000100110",
  21823=>"000111001",
  21824=>"001111111",
  21825=>"111101011",
  21826=>"011111101",
  21827=>"111011101",
  21828=>"100110010",
  21829=>"011111111",
  21830=>"101010000",
  21831=>"101111110",
  21832=>"111011110",
  21833=>"011100011",
  21834=>"000010000",
  21835=>"010111111",
  21836=>"110000010",
  21837=>"111111100",
  21838=>"000111101",
  21839=>"110011110",
  21840=>"100011101",
  21841=>"000101000",
  21842=>"100011100",
  21843=>"110111101",
  21844=>"111011110",
  21845=>"010010100",
  21846=>"110010011",
  21847=>"011101000",
  21848=>"111010001",
  21849=>"101011101",
  21850=>"110110100",
  21851=>"011011011",
  21852=>"000010000",
  21853=>"110111011",
  21854=>"000011010",
  21855=>"100110110",
  21856=>"110110011",
  21857=>"110110110",
  21858=>"100100111",
  21859=>"001111011",
  21860=>"010101000",
  21861=>"000100100",
  21862=>"100010111",
  21863=>"011110011",
  21864=>"110010101",
  21865=>"100010011",
  21866=>"111110010",
  21867=>"111011010",
  21868=>"101000011",
  21869=>"000011101",
  21870=>"101111111",
  21871=>"100001010",
  21872=>"000011100",
  21873=>"100110010",
  21874=>"111000110",
  21875=>"110100110",
  21876=>"000000110",
  21877=>"010011011",
  21878=>"000110111",
  21879=>"011011101",
  21880=>"111111000",
  21881=>"101000101",
  21882=>"001100110",
  21883=>"110001111",
  21884=>"111110001",
  21885=>"001001010",
  21886=>"010011111",
  21887=>"010110110",
  21888=>"000000010",
  21889=>"000001011",
  21890=>"110111011",
  21891=>"000010110",
  21892=>"010110101",
  21893=>"111011101",
  21894=>"000001010",
  21895=>"011011011",
  21896=>"000001100",
  21897=>"101001000",
  21898=>"110111101",
  21899=>"001000001",
  21900=>"000110011",
  21901=>"000110101",
  21902=>"010000011",
  21903=>"001010111",
  21904=>"011101010",
  21905=>"001101011",
  21906=>"111100000",
  21907=>"111011110",
  21908=>"111110011",
  21909=>"110110110",
  21910=>"100110010",
  21911=>"111001010",
  21912=>"000011000",
  21913=>"000111011",
  21914=>"000000010",
  21915=>"100000011",
  21916=>"100010100",
  21917=>"010101111",
  21918=>"110010011",
  21919=>"010000000",
  21920=>"110011001",
  21921=>"110100101",
  21922=>"000010111",
  21923=>"101001010",
  21924=>"011110001",
  21925=>"001000111",
  21926=>"001000000",
  21927=>"111111010",
  21928=>"100110111",
  21929=>"000110100",
  21930=>"000001110",
  21931=>"010000011",
  21932=>"010010110",
  21933=>"000101001",
  21934=>"000010111",
  21935=>"000011011",
  21936=>"000110101",
  21937=>"111101011",
  21938=>"010100110",
  21939=>"111010101",
  21940=>"000010000",
  21941=>"111011110",
  21942=>"101101111",
  21943=>"010100000",
  21944=>"111100111",
  21945=>"011000100",
  21946=>"100101001",
  21947=>"100111010",
  21948=>"101111010",
  21949=>"001111111",
  21950=>"000011011",
  21951=>"100111110",
  21952=>"111010110",
  21953=>"001010111",
  21954=>"010111000",
  21955=>"101101001",
  21956=>"010100111",
  21957=>"100001110",
  21958=>"101110111",
  21959=>"001101001",
  21960=>"001111111",
  21961=>"101101111",
  21962=>"011110010",
  21963=>"001001101",
  21964=>"110001001",
  21965=>"000001111",
  21966=>"100010101",
  21967=>"011101111",
  21968=>"110000101",
  21969=>"001010100",
  21970=>"100000001",
  21971=>"110100100",
  21972=>"011101001",
  21973=>"111111011",
  21974=>"000010101",
  21975=>"101011111",
  21976=>"100001110",
  21977=>"100000110",
  21978=>"001101001",
  21979=>"101111011",
  21980=>"111011001",
  21981=>"111110000",
  21982=>"011110011",
  21983=>"111110111",
  21984=>"101011000",
  21985=>"001100000",
  21986=>"011010111",
  21987=>"111111110",
  21988=>"010001010",
  21989=>"000010011",
  21990=>"000001110",
  21991=>"010011001",
  21992=>"101001101",
  21993=>"111011110",
  21994=>"000101000",
  21995=>"110111100",
  21996=>"010001011",
  21997=>"001001000",
  21998=>"000100000",
  21999=>"110001001",
  22000=>"010111000",
  22001=>"001111110",
  22002=>"100100100",
  22003=>"111110000",
  22004=>"101101001",
  22005=>"111000000",
  22006=>"001110001",
  22007=>"000101011",
  22008=>"101100101",
  22009=>"011110010",
  22010=>"010001110",
  22011=>"010100010",
  22012=>"000011001",
  22013=>"000001100",
  22014=>"001110111",
  22015=>"011000001",
  22016=>"001100111",
  22017=>"100000000",
  22018=>"111111001",
  22019=>"010001010",
  22020=>"010101101",
  22021=>"001001001",
  22022=>"000011000",
  22023=>"001011000",
  22024=>"010111100",
  22025=>"111011001",
  22026=>"001110111",
  22027=>"000000001",
  22028=>"010000000",
  22029=>"100101010",
  22030=>"010000110",
  22031=>"111101010",
  22032=>"100101001",
  22033=>"010100010",
  22034=>"101101000",
  22035=>"000010110",
  22036=>"000000000",
  22037=>"111000101",
  22038=>"111111101",
  22039=>"111001101",
  22040=>"110001001",
  22041=>"001101111",
  22042=>"111111011",
  22043=>"100001100",
  22044=>"000001101",
  22045=>"011100010",
  22046=>"110101101",
  22047=>"110101011",
  22048=>"100101011",
  22049=>"101100110",
  22050=>"000000010",
  22051=>"010010010",
  22052=>"010111001",
  22053=>"100001110",
  22054=>"001111110",
  22055=>"001101100",
  22056=>"010101000",
  22057=>"000000011",
  22058=>"111110110",
  22059=>"110001110",
  22060=>"101100110",
  22061=>"010010000",
  22062=>"001110011",
  22063=>"100011010",
  22064=>"010100100",
  22065=>"000010110",
  22066=>"010110010",
  22067=>"010101111",
  22068=>"100101000",
  22069=>"100011000",
  22070=>"101110010",
  22071=>"011110011",
  22072=>"110011010",
  22073=>"010101010",
  22074=>"010110011",
  22075=>"000000110",
  22076=>"000000111",
  22077=>"010101110",
  22078=>"111111010",
  22079=>"110010010",
  22080=>"111011001",
  22081=>"000110111",
  22082=>"001100000",
  22083=>"110111110",
  22084=>"001001011",
  22085=>"100001000",
  22086=>"100100000",
  22087=>"110001101",
  22088=>"000000111",
  22089=>"000110111",
  22090=>"110110110",
  22091=>"010110000",
  22092=>"111011111",
  22093=>"110110100",
  22094=>"111000000",
  22095=>"100100001",
  22096=>"111011111",
  22097=>"001001001",
  22098=>"001110010",
  22099=>"001001111",
  22100=>"110100001",
  22101=>"010110101",
  22102=>"010101001",
  22103=>"100100110",
  22104=>"000101100",
  22105=>"001001001",
  22106=>"010010000",
  22107=>"000111010",
  22108=>"110011011",
  22109=>"000000011",
  22110=>"110111011",
  22111=>"111000110",
  22112=>"010011101",
  22113=>"010010001",
  22114=>"010000101",
  22115=>"101011010",
  22116=>"110011111",
  22117=>"110101000",
  22118=>"011011000",
  22119=>"100101111",
  22120=>"100000110",
  22121=>"110100010",
  22122=>"101111001",
  22123=>"101011001",
  22124=>"000101111",
  22125=>"101011111",
  22126=>"011110001",
  22127=>"001000101",
  22128=>"001010010",
  22129=>"001101110",
  22130=>"110100001",
  22131=>"101110110",
  22132=>"001011001",
  22133=>"100011000",
  22134=>"110010110",
  22135=>"001000010",
  22136=>"011011011",
  22137=>"001001100",
  22138=>"001001000",
  22139=>"001000000",
  22140=>"001010001",
  22141=>"110100100",
  22142=>"101111101",
  22143=>"000011011",
  22144=>"110111000",
  22145=>"110111000",
  22146=>"000000110",
  22147=>"110000011",
  22148=>"000010101",
  22149=>"001111000",
  22150=>"111110000",
  22151=>"011111001",
  22152=>"011111111",
  22153=>"010100000",
  22154=>"000001001",
  22155=>"001111100",
  22156=>"011100010",
  22157=>"001101010",
  22158=>"010001010",
  22159=>"100001000",
  22160=>"110000100",
  22161=>"100110010",
  22162=>"111010011",
  22163=>"011011011",
  22164=>"000111100",
  22165=>"110111110",
  22166=>"100000101",
  22167=>"011100111",
  22168=>"110000001",
  22169=>"101011101",
  22170=>"101000011",
  22171=>"111000101",
  22172=>"000010100",
  22173=>"001101111",
  22174=>"101111110",
  22175=>"001000110",
  22176=>"000001010",
  22177=>"110110111",
  22178=>"101110000",
  22179=>"111110101",
  22180=>"111100100",
  22181=>"111110000",
  22182=>"000010000",
  22183=>"000011010",
  22184=>"000001011",
  22185=>"000001110",
  22186=>"101100010",
  22187=>"011000001",
  22188=>"011001010",
  22189=>"101010111",
  22190=>"000001101",
  22191=>"010100000",
  22192=>"000001001",
  22193=>"010110001",
  22194=>"011010010",
  22195=>"111110000",
  22196=>"100111101",
  22197=>"011111011",
  22198=>"111000010",
  22199=>"000011001",
  22200=>"000100111",
  22201=>"111010100",
  22202=>"000100010",
  22203=>"111111011",
  22204=>"010100110",
  22205=>"111110111",
  22206=>"010110001",
  22207=>"101100001",
  22208=>"111010100",
  22209=>"101001110",
  22210=>"111111000",
  22211=>"100100100",
  22212=>"101001101",
  22213=>"101111001",
  22214=>"110101001",
  22215=>"000001000",
  22216=>"101011010",
  22217=>"111110111",
  22218=>"011110111",
  22219=>"001100110",
  22220=>"111001010",
  22221=>"101110100",
  22222=>"111000010",
  22223=>"110000011",
  22224=>"110100000",
  22225=>"010010000",
  22226=>"001110000",
  22227=>"001001000",
  22228=>"110000110",
  22229=>"110111001",
  22230=>"010001001",
  22231=>"000000111",
  22232=>"000011101",
  22233=>"110001001",
  22234=>"101110111",
  22235=>"011111000",
  22236=>"111101101",
  22237=>"110011000",
  22238=>"110001100",
  22239=>"101111100",
  22240=>"101111001",
  22241=>"000010010",
  22242=>"100011010",
  22243=>"100101000",
  22244=>"110110100",
  22245=>"101000001",
  22246=>"010010010",
  22247=>"101110010",
  22248=>"101101111",
  22249=>"111000101",
  22250=>"011001100",
  22251=>"010101110",
  22252=>"001011111",
  22253=>"111110001",
  22254=>"111000010",
  22255=>"000110011",
  22256=>"000000000",
  22257=>"100101101",
  22258=>"111010011",
  22259=>"011111111",
  22260=>"011110100",
  22261=>"111110001",
  22262=>"111101101",
  22263=>"100111110",
  22264=>"101011100",
  22265=>"111100100",
  22266=>"010001001",
  22267=>"010011100",
  22268=>"110101000",
  22269=>"010101000",
  22270=>"110110010",
  22271=>"110101000",
  22272=>"011001011",
  22273=>"000111010",
  22274=>"010010000",
  22275=>"111010100",
  22276=>"000100000",
  22277=>"101111111",
  22278=>"001111011",
  22279=>"000110111",
  22280=>"111101111",
  22281=>"010110111",
  22282=>"010101100",
  22283=>"001111001",
  22284=>"011111101",
  22285=>"110111111",
  22286=>"110010000",
  22287=>"111011111",
  22288=>"000011001",
  22289=>"101110000",
  22290=>"101111111",
  22291=>"110101101",
  22292=>"001000001",
  22293=>"000110111",
  22294=>"011110100",
  22295=>"110011000",
  22296=>"000011000",
  22297=>"010000111",
  22298=>"111011110",
  22299=>"100001110",
  22300=>"110100001",
  22301=>"010111100",
  22302=>"000010100",
  22303=>"011111001",
  22304=>"010010110",
  22305=>"110110100",
  22306=>"100011010",
  22307=>"101111110",
  22308=>"111111000",
  22309=>"001001010",
  22310=>"010110101",
  22311=>"101000111",
  22312=>"101001100",
  22313=>"101100001",
  22314=>"010110110",
  22315=>"110100011",
  22316=>"100000111",
  22317=>"011001000",
  22318=>"111100110",
  22319=>"011110000",
  22320=>"010000000",
  22321=>"111010101",
  22322=>"001011110",
  22323=>"010000101",
  22324=>"110011010",
  22325=>"111001100",
  22326=>"000001110",
  22327=>"000100001",
  22328=>"011101001",
  22329=>"011110110",
  22330=>"100111001",
  22331=>"001011001",
  22332=>"100001011",
  22333=>"000010010",
  22334=>"100100111",
  22335=>"011011010",
  22336=>"000111111",
  22337=>"000000111",
  22338=>"011101100",
  22339=>"000100100",
  22340=>"000100010",
  22341=>"110100010",
  22342=>"100011010",
  22343=>"000011010",
  22344=>"010110000",
  22345=>"010000100",
  22346=>"110111010",
  22347=>"111001000",
  22348=>"000001010",
  22349=>"101011110",
  22350=>"100001100",
  22351=>"001110100",
  22352=>"110011011",
  22353=>"100000000",
  22354=>"011100110",
  22355=>"000100010",
  22356=>"110010110",
  22357=>"010011111",
  22358=>"010000010",
  22359=>"010010001",
  22360=>"101011111",
  22361=>"001111011",
  22362=>"000100010",
  22363=>"000010101",
  22364=>"000111010",
  22365=>"110101101",
  22366=>"101110010",
  22367=>"000001011",
  22368=>"101010011",
  22369=>"101100001",
  22370=>"101111011",
  22371=>"010111011",
  22372=>"100101011",
  22373=>"111000101",
  22374=>"000101001",
  22375=>"111111100",
  22376=>"010001000",
  22377=>"010100111",
  22378=>"110010000",
  22379=>"010000110",
  22380=>"111111110",
  22381=>"110011110",
  22382=>"111010001",
  22383=>"010100010",
  22384=>"000111100",
  22385=>"101110000",
  22386=>"101011101",
  22387=>"000111000",
  22388=>"111111111",
  22389=>"000110001",
  22390=>"010100011",
  22391=>"100001000",
  22392=>"010000011",
  22393=>"001001101",
  22394=>"111111101",
  22395=>"000110111",
  22396=>"010101011",
  22397=>"000011100",
  22398=>"001011000",
  22399=>"010100011",
  22400=>"101111110",
  22401=>"111101101",
  22402=>"001110111",
  22403=>"111001111",
  22404=>"000010110",
  22405=>"101110010",
  22406=>"111101010",
  22407=>"100100011",
  22408=>"100001111",
  22409=>"001010001",
  22410=>"110101110",
  22411=>"001110001",
  22412=>"011011000",
  22413=>"101001100",
  22414=>"100110010",
  22415=>"110101101",
  22416=>"010111100",
  22417=>"010100101",
  22418=>"000000011",
  22419=>"011010001",
  22420=>"000111100",
  22421=>"001001100",
  22422=>"100000100",
  22423=>"001010001",
  22424=>"001010110",
  22425=>"100100001",
  22426=>"101100001",
  22427=>"110010001",
  22428=>"011010000",
  22429=>"011001100",
  22430=>"011100001",
  22431=>"001011001",
  22432=>"001010000",
  22433=>"111101010",
  22434=>"011100111",
  22435=>"111110110",
  22436=>"000100110",
  22437=>"100001110",
  22438=>"101111010",
  22439=>"100111111",
  22440=>"001001000",
  22441=>"001100011",
  22442=>"001110111",
  22443=>"111010110",
  22444=>"000111101",
  22445=>"111111110",
  22446=>"110011010",
  22447=>"110101000",
  22448=>"111110011",
  22449=>"101000000",
  22450=>"010101011",
  22451=>"111011111",
  22452=>"110110000",
  22453=>"111100110",
  22454=>"110110110",
  22455=>"001100011",
  22456=>"111101011",
  22457=>"110010001",
  22458=>"000011001",
  22459=>"111101101",
  22460=>"101001000",
  22461=>"111001000",
  22462=>"011011000",
  22463=>"010101101",
  22464=>"010011111",
  22465=>"000001011",
  22466=>"101101111",
  22467=>"010010000",
  22468=>"010101011",
  22469=>"011111101",
  22470=>"101010100",
  22471=>"101001101",
  22472=>"001000101",
  22473=>"110000000",
  22474=>"100001110",
  22475=>"101001000",
  22476=>"000011001",
  22477=>"001001101",
  22478=>"111111101",
  22479=>"100110110",
  22480=>"100111000",
  22481=>"000011001",
  22482=>"001111111",
  22483=>"101101010",
  22484=>"100101101",
  22485=>"110010010",
  22486=>"011110010",
  22487=>"010100100",
  22488=>"111111011",
  22489=>"000100001",
  22490=>"100110111",
  22491=>"001101000",
  22492=>"000110101",
  22493=>"111100000",
  22494=>"001101000",
  22495=>"000100111",
  22496=>"000001001",
  22497=>"111101000",
  22498=>"010011001",
  22499=>"100011110",
  22500=>"000111000",
  22501=>"110011001",
  22502=>"101101111",
  22503=>"000101000",
  22504=>"001011011",
  22505=>"001101110",
  22506=>"101011100",
  22507=>"000100100",
  22508=>"011001110",
  22509=>"110101011",
  22510=>"011000111",
  22511=>"000001001",
  22512=>"001011110",
  22513=>"110010000",
  22514=>"110101110",
  22515=>"110100100",
  22516=>"001110100",
  22517=>"001001111",
  22518=>"001001111",
  22519=>"101000100",
  22520=>"000001001",
  22521=>"110101001",
  22522=>"100001000",
  22523=>"000000110",
  22524=>"010100001",
  22525=>"000111000",
  22526=>"101101011",
  22527=>"010101111",
  22528=>"001101001",
  22529=>"100000101",
  22530=>"000010010",
  22531=>"000100011",
  22532=>"000001000",
  22533=>"010001001",
  22534=>"111001010",
  22535=>"100000100",
  22536=>"111110001",
  22537=>"010000100",
  22538=>"000000000",
  22539=>"101010111",
  22540=>"111000000",
  22541=>"101110000",
  22542=>"001101100",
  22543=>"000010100",
  22544=>"111001101",
  22545=>"010010001",
  22546=>"000101111",
  22547=>"000100101",
  22548=>"000011111",
  22549=>"000101011",
  22550=>"101100001",
  22551=>"000000100",
  22552=>"100000101",
  22553=>"001000000",
  22554=>"100011100",
  22555=>"111111110",
  22556=>"111110000",
  22557=>"110111100",
  22558=>"111000101",
  22559=>"101110110",
  22560=>"010100111",
  22561=>"011110011",
  22562=>"000001100",
  22563=>"110101001",
  22564=>"010000011",
  22565=>"110001100",
  22566=>"010111110",
  22567=>"000000110",
  22568=>"100101011",
  22569=>"000010001",
  22570=>"011001110",
  22571=>"100001111",
  22572=>"010011010",
  22573=>"000001110",
  22574=>"101101011",
  22575=>"101010010",
  22576=>"100100111",
  22577=>"100110010",
  22578=>"110010100",
  22579=>"000010001",
  22580=>"100111011",
  22581=>"010110101",
  22582=>"011111101",
  22583=>"000111011",
  22584=>"100001101",
  22585=>"111001111",
  22586=>"100011101",
  22587=>"100000000",
  22588=>"000010011",
  22589=>"110011100",
  22590=>"101110110",
  22591=>"101011111",
  22592=>"010000000",
  22593=>"000001110",
  22594=>"100000110",
  22595=>"100011110",
  22596=>"000110001",
  22597=>"011001110",
  22598=>"010110110",
  22599=>"010100100",
  22600=>"010010010",
  22601=>"010111100",
  22602=>"000111101",
  22603=>"000101101",
  22604=>"110000000",
  22605=>"010100111",
  22606=>"011010100",
  22607=>"001001001",
  22608=>"111101110",
  22609=>"000001011",
  22610=>"010100100",
  22611=>"001001011",
  22612=>"000011000",
  22613=>"101110111",
  22614=>"101011100",
  22615=>"001001000",
  22616=>"110111101",
  22617=>"010110010",
  22618=>"000001001",
  22619=>"000000001",
  22620=>"000100101",
  22621=>"100110001",
  22622=>"110101000",
  22623=>"010010001",
  22624=>"101000100",
  22625=>"001100100",
  22626=>"100111001",
  22627=>"110001001",
  22628=>"111110101",
  22629=>"101011111",
  22630=>"011000101",
  22631=>"000011011",
  22632=>"011000010",
  22633=>"101010001",
  22634=>"111100000",
  22635=>"010101100",
  22636=>"101111001",
  22637=>"110010001",
  22638=>"100000000",
  22639=>"111101000",
  22640=>"111010101",
  22641=>"111010111",
  22642=>"100011011",
  22643=>"101010000",
  22644=>"011111101",
  22645=>"001001001",
  22646=>"010100110",
  22647=>"000100101",
  22648=>"000010110",
  22649=>"101010101",
  22650=>"010100011",
  22651=>"110100101",
  22652=>"001010111",
  22653=>"100110010",
  22654=>"100011111",
  22655=>"100100110",
  22656=>"001100111",
  22657=>"110001010",
  22658=>"100101000",
  22659=>"101100101",
  22660=>"111110001",
  22661=>"101000101",
  22662=>"000111111",
  22663=>"001101111",
  22664=>"010011101",
  22665=>"010100010",
  22666=>"011010110",
  22667=>"000100101",
  22668=>"000000011",
  22669=>"101110111",
  22670=>"111111111",
  22671=>"110010110",
  22672=>"100101001",
  22673=>"010011011",
  22674=>"100011101",
  22675=>"111011110",
  22676=>"110001110",
  22677=>"010011001",
  22678=>"011101001",
  22679=>"010000110",
  22680=>"110101000",
  22681=>"000101000",
  22682=>"010010101",
  22683=>"110001000",
  22684=>"100011000",
  22685=>"100110000",
  22686=>"010010010",
  22687=>"001100101",
  22688=>"111100010",
  22689=>"011101011",
  22690=>"010101011",
  22691=>"010000100",
  22692=>"100111000",
  22693=>"100111011",
  22694=>"101100101",
  22695=>"101000011",
  22696=>"010011100",
  22697=>"001001110",
  22698=>"001000110",
  22699=>"011111100",
  22700=>"011101100",
  22701=>"101110111",
  22702=>"011110010",
  22703=>"110000111",
  22704=>"101010111",
  22705=>"011100010",
  22706=>"111010100",
  22707=>"100001001",
  22708=>"000000101",
  22709=>"110100011",
  22710=>"100100100",
  22711=>"000110011",
  22712=>"011000011",
  22713=>"101001001",
  22714=>"010110000",
  22715=>"110000011",
  22716=>"010001101",
  22717=>"010000001",
  22718=>"100011000",
  22719=>"100010111",
  22720=>"111111100",
  22721=>"110111010",
  22722=>"100011110",
  22723=>"110000010",
  22724=>"001000010",
  22725=>"110000101",
  22726=>"000100101",
  22727=>"000111011",
  22728=>"100000101",
  22729=>"101111101",
  22730=>"000101000",
  22731=>"111001001",
  22732=>"100110000",
  22733=>"001000001",
  22734=>"101011111",
  22735=>"111001111",
  22736=>"000000011",
  22737=>"001101100",
  22738=>"100011110",
  22739=>"000000010",
  22740=>"001101000",
  22741=>"010100010",
  22742=>"101011010",
  22743=>"101100100",
  22744=>"100110000",
  22745=>"111111011",
  22746=>"001111010",
  22747=>"111001100",
  22748=>"100101010",
  22749=>"001110001",
  22750=>"111000111",
  22751=>"001000010",
  22752=>"110011000",
  22753=>"001001100",
  22754=>"001010111",
  22755=>"000100100",
  22756=>"100010110",
  22757=>"010011000",
  22758=>"110000000",
  22759=>"100111111",
  22760=>"010001011",
  22761=>"101011010",
  22762=>"010110111",
  22763=>"001110100",
  22764=>"100100110",
  22765=>"000100110",
  22766=>"001011101",
  22767=>"100001111",
  22768=>"010000110",
  22769=>"011000101",
  22770=>"001000011",
  22771=>"100101001",
  22772=>"111111101",
  22773=>"111000000",
  22774=>"011111001",
  22775=>"010001111",
  22776=>"000000000",
  22777=>"011101111",
  22778=>"100100100",
  22779=>"000011001",
  22780=>"001011001",
  22781=>"000111011",
  22782=>"000110110",
  22783=>"000101000",
  22784=>"000100000",
  22785=>"100001110",
  22786=>"110010010",
  22787=>"100100001",
  22788=>"101101010",
  22789=>"010111110",
  22790=>"111010000",
  22791=>"100001101",
  22792=>"001110011",
  22793=>"100000000",
  22794=>"011010110",
  22795=>"000110010",
  22796=>"011001110",
  22797=>"111101010",
  22798=>"100000110",
  22799=>"000110001",
  22800=>"001101011",
  22801=>"100001000",
  22802=>"011110110",
  22803=>"110001001",
  22804=>"011010110",
  22805=>"000010001",
  22806=>"010001011",
  22807=>"011010011",
  22808=>"011011101",
  22809=>"101101100",
  22810=>"110101000",
  22811=>"011011101",
  22812=>"111011000",
  22813=>"101010001",
  22814=>"010011001",
  22815=>"101101011",
  22816=>"010110000",
  22817=>"101101010",
  22818=>"010110101",
  22819=>"000010010",
  22820=>"010110011",
  22821=>"110000101",
  22822=>"010100000",
  22823=>"110110011",
  22824=>"010010001",
  22825=>"011011010",
  22826=>"111000100",
  22827=>"101101011",
  22828=>"101101111",
  22829=>"010000101",
  22830=>"000000000",
  22831=>"001101110",
  22832=>"101100010",
  22833=>"110111000",
  22834=>"111111111",
  22835=>"001100111",
  22836=>"000000010",
  22837=>"010100001",
  22838=>"111010100",
  22839=>"100101000",
  22840=>"000010111",
  22841=>"111110010",
  22842=>"001111001",
  22843=>"100001011",
  22844=>"111000100",
  22845=>"111000100",
  22846=>"110100101",
  22847=>"110101110",
  22848=>"101101101",
  22849=>"111011101",
  22850=>"111001100",
  22851=>"100000001",
  22852=>"110111111",
  22853=>"111101111",
  22854=>"000010010",
  22855=>"100101100",
  22856=>"010110111",
  22857=>"010110000",
  22858=>"110100000",
  22859=>"111001110",
  22860=>"100011111",
  22861=>"111000011",
  22862=>"110001010",
  22863=>"101010101",
  22864=>"010100111",
  22865=>"000100101",
  22866=>"100110100",
  22867=>"110001001",
  22868=>"010010011",
  22869=>"010111111",
  22870=>"011001100",
  22871=>"111110110",
  22872=>"000010001",
  22873=>"111011010",
  22874=>"000110011",
  22875=>"110110001",
  22876=>"001001100",
  22877=>"111110011",
  22878=>"110011010",
  22879=>"001001001",
  22880=>"100011011",
  22881=>"000001011",
  22882=>"001011001",
  22883=>"000010110",
  22884=>"101001100",
  22885=>"011010111",
  22886=>"010011010",
  22887=>"001011000",
  22888=>"011101101",
  22889=>"010001000",
  22890=>"011001011",
  22891=>"000000001",
  22892=>"101001001",
  22893=>"100100010",
  22894=>"100000011",
  22895=>"101001011",
  22896=>"000010001",
  22897=>"111001000",
  22898=>"010010000",
  22899=>"111010001",
  22900=>"110101100",
  22901=>"111110001",
  22902=>"000111011",
  22903=>"101101101",
  22904=>"000101101",
  22905=>"011011010",
  22906=>"000011001",
  22907=>"111100111",
  22908=>"110011011",
  22909=>"100000111",
  22910=>"011100111",
  22911=>"101100111",
  22912=>"111001010",
  22913=>"000101100",
  22914=>"010110001",
  22915=>"110001000",
  22916=>"101000001",
  22917=>"000101111",
  22918=>"100111111",
  22919=>"000010000",
  22920=>"001011000",
  22921=>"001000000",
  22922=>"110110001",
  22923=>"001110101",
  22924=>"111101100",
  22925=>"110011101",
  22926=>"100111111",
  22927=>"001011011",
  22928=>"100111000",
  22929=>"000001010",
  22930=>"111011001",
  22931=>"100111111",
  22932=>"101001001",
  22933=>"011000010",
  22934=>"010111000",
  22935=>"000111111",
  22936=>"100000010",
  22937=>"100000101",
  22938=>"110011100",
  22939=>"010001110",
  22940=>"100010000",
  22941=>"000011110",
  22942=>"011110000",
  22943=>"011001101",
  22944=>"010000000",
  22945=>"000111101",
  22946=>"011111011",
  22947=>"000000000",
  22948=>"010011000",
  22949=>"001001111",
  22950=>"000111111",
  22951=>"010001110",
  22952=>"111000001",
  22953=>"100001100",
  22954=>"000101010",
  22955=>"110001001",
  22956=>"000000101",
  22957=>"100110110",
  22958=>"010100110",
  22959=>"011010100",
  22960=>"000011000",
  22961=>"111000111",
  22962=>"110000111",
  22963=>"010100001",
  22964=>"111101111",
  22965=>"101110011",
  22966=>"010000010",
  22967=>"011000001",
  22968=>"110100000",
  22969=>"110010110",
  22970=>"001111110",
  22971=>"011110101",
  22972=>"000101100",
  22973=>"100100101",
  22974=>"001101000",
  22975=>"000001011",
  22976=>"000000100",
  22977=>"010011101",
  22978=>"000000110",
  22979=>"100101111",
  22980=>"001111010",
  22981=>"111001010",
  22982=>"000010010",
  22983=>"100010000",
  22984=>"010100010",
  22985=>"000110011",
  22986=>"101010001",
  22987=>"101010011",
  22988=>"000111010",
  22989=>"001001101",
  22990=>"111101110",
  22991=>"100000101",
  22992=>"011010001",
  22993=>"101101010",
  22994=>"001101110",
  22995=>"111110110",
  22996=>"110010110",
  22997=>"000100010",
  22998=>"010000110",
  22999=>"011000000",
  23000=>"011100100",
  23001=>"000110111",
  23002=>"010111000",
  23003=>"110000011",
  23004=>"011010111",
  23005=>"111000110",
  23006=>"101101111",
  23007=>"110111001",
  23008=>"001000011",
  23009=>"110001101",
  23010=>"010101011",
  23011=>"000001101",
  23012=>"010111000",
  23013=>"111100001",
  23014=>"100110111",
  23015=>"000010000",
  23016=>"100000111",
  23017=>"111010101",
  23018=>"000110000",
  23019=>"011001110",
  23020=>"100001101",
  23021=>"000001100",
  23022=>"001000011",
  23023=>"000010010",
  23024=>"011101000",
  23025=>"100001110",
  23026=>"010110110",
  23027=>"010000010",
  23028=>"001111010",
  23029=>"011111110",
  23030=>"111011011",
  23031=>"011001101",
  23032=>"111011101",
  23033=>"011010011",
  23034=>"010010101",
  23035=>"101001100",
  23036=>"000010101",
  23037=>"101110010",
  23038=>"011101111",
  23039=>"001111000",
  23040=>"101110111",
  23041=>"110000101",
  23042=>"000000110",
  23043=>"100010000",
  23044=>"010111011",
  23045=>"001110010",
  23046=>"111111000",
  23047=>"101001010",
  23048=>"000101101",
  23049=>"100010111",
  23050=>"010110101",
  23051=>"000101100",
  23052=>"110111001",
  23053=>"000010000",
  23054=>"000000001",
  23055=>"001011101",
  23056=>"111100110",
  23057=>"000000000",
  23058=>"101111000",
  23059=>"001101100",
  23060=>"011010010",
  23061=>"101110011",
  23062=>"110010011",
  23063=>"111111100",
  23064=>"110010100",
  23065=>"100101101",
  23066=>"001100000",
  23067=>"100101000",
  23068=>"011010100",
  23069=>"001001010",
  23070=>"100111011",
  23071=>"110000011",
  23072=>"000001100",
  23073=>"111111101",
  23074=>"000000111",
  23075=>"010001101",
  23076=>"100100011",
  23077=>"010101011",
  23078=>"101110101",
  23079=>"101100000",
  23080=>"000010000",
  23081=>"111010101",
  23082=>"011111000",
  23083=>"101110011",
  23084=>"010101111",
  23085=>"000010001",
  23086=>"010100100",
  23087=>"001011000",
  23088=>"000011111",
  23089=>"001011001",
  23090=>"100111100",
  23091=>"011101100",
  23092=>"010000000",
  23093=>"111101010",
  23094=>"110011100",
  23095=>"000110001",
  23096=>"101110100",
  23097=>"010111111",
  23098=>"110100000",
  23099=>"100100110",
  23100=>"111010101",
  23101=>"101000000",
  23102=>"100111111",
  23103=>"101100001",
  23104=>"110101010",
  23105=>"010001100",
  23106=>"000010100",
  23107=>"111100011",
  23108=>"010100011",
  23109=>"010100101",
  23110=>"000000000",
  23111=>"100110010",
  23112=>"001000011",
  23113=>"110111011",
  23114=>"010111100",
  23115=>"110100101",
  23116=>"011110110",
  23117=>"011111010",
  23118=>"111110100",
  23119=>"001101010",
  23120=>"110111011",
  23121=>"110001110",
  23122=>"100000101",
  23123=>"011000001",
  23124=>"101001101",
  23125=>"001010011",
  23126=>"110101100",
  23127=>"000001110",
  23128=>"101101011",
  23129=>"000011100",
  23130=>"000001000",
  23131=>"000011101",
  23132=>"001111000",
  23133=>"100001010",
  23134=>"111101101",
  23135=>"011100011",
  23136=>"111010110",
  23137=>"001101000",
  23138=>"101000000",
  23139=>"001001001",
  23140=>"100010010",
  23141=>"000000100",
  23142=>"110101100",
  23143=>"111101001",
  23144=>"110011011",
  23145=>"010101000",
  23146=>"100111010",
  23147=>"010000001",
  23148=>"101100001",
  23149=>"001000011",
  23150=>"001001000",
  23151=>"001001100",
  23152=>"000100100",
  23153=>"001111101",
  23154=>"001110111",
  23155=>"001110011",
  23156=>"100001100",
  23157=>"100001100",
  23158=>"011100110",
  23159=>"010001111",
  23160=>"000110011",
  23161=>"110000000",
  23162=>"001001000",
  23163=>"101111001",
  23164=>"101000000",
  23165=>"011011010",
  23166=>"101111000",
  23167=>"011111001",
  23168=>"100001110",
  23169=>"100100100",
  23170=>"001010110",
  23171=>"101101101",
  23172=>"101001010",
  23173=>"100001110",
  23174=>"110111110",
  23175=>"011110100",
  23176=>"101110100",
  23177=>"011101001",
  23178=>"101001101",
  23179=>"010010000",
  23180=>"010001010",
  23181=>"111111101",
  23182=>"001001010",
  23183=>"110000110",
  23184=>"100110011",
  23185=>"000111111",
  23186=>"111111101",
  23187=>"011001001",
  23188=>"000101010",
  23189=>"101011000",
  23190=>"101100010",
  23191=>"101111101",
  23192=>"110101010",
  23193=>"111111101",
  23194=>"001101010",
  23195=>"011100110",
  23196=>"000110101",
  23197=>"100111001",
  23198=>"011110101",
  23199=>"000001100",
  23200=>"100001111",
  23201=>"000001110",
  23202=>"011111000",
  23203=>"011111111",
  23204=>"001111011",
  23205=>"000011111",
  23206=>"000101100",
  23207=>"000001011",
  23208=>"000011110",
  23209=>"001001100",
  23210=>"011101011",
  23211=>"110010000",
  23212=>"100010000",
  23213=>"001110101",
  23214=>"001101000",
  23215=>"111010110",
  23216=>"001101010",
  23217=>"100001011",
  23218=>"000110111",
  23219=>"101011110",
  23220=>"100100011",
  23221=>"111101111",
  23222=>"110111011",
  23223=>"111101011",
  23224=>"110101001",
  23225=>"011111010",
  23226=>"100101111",
  23227=>"111111100",
  23228=>"100110111",
  23229=>"010110001",
  23230=>"000010101",
  23231=>"101101101",
  23232=>"111001100",
  23233=>"001101100",
  23234=>"101001111",
  23235=>"101101111",
  23236=>"000101001",
  23237=>"010100001",
  23238=>"000110111",
  23239=>"001010000",
  23240=>"011011011",
  23241=>"100001111",
  23242=>"010001110",
  23243=>"001111111",
  23244=>"010000110",
  23245=>"111100101",
  23246=>"100011000",
  23247=>"011100000",
  23248=>"000111001",
  23249=>"110001000",
  23250=>"100100001",
  23251=>"000110100",
  23252=>"111000101",
  23253=>"011111101",
  23254=>"001101110",
  23255=>"010011000",
  23256=>"101110101",
  23257=>"011110000",
  23258=>"000101100",
  23259=>"101001111",
  23260=>"001011010",
  23261=>"011100110",
  23262=>"110010010",
  23263=>"011100001",
  23264=>"110011001",
  23265=>"001111101",
  23266=>"000101010",
  23267=>"001100000",
  23268=>"111011101",
  23269=>"100100010",
  23270=>"111101000",
  23271=>"101110110",
  23272=>"001011010",
  23273=>"111011011",
  23274=>"000000110",
  23275=>"011100010",
  23276=>"011011001",
  23277=>"000011011",
  23278=>"001000010",
  23279=>"101101111",
  23280=>"011110011",
  23281=>"101000111",
  23282=>"010000111",
  23283=>"100010110",
  23284=>"010110111",
  23285=>"110100111",
  23286=>"001110011",
  23287=>"000010000",
  23288=>"100100010",
  23289=>"011111010",
  23290=>"110101000",
  23291=>"000110111",
  23292=>"010001001",
  23293=>"110000110",
  23294=>"001110110",
  23295=>"000111110",
  23296=>"110011100",
  23297=>"011111010",
  23298=>"100111100",
  23299=>"110100111",
  23300=>"100101101",
  23301=>"100011111",
  23302=>"111111001",
  23303=>"001000011",
  23304=>"111101011",
  23305=>"011100001",
  23306=>"100101101",
  23307=>"101010101",
  23308=>"101111001",
  23309=>"111110010",
  23310=>"101110000",
  23311=>"101111111",
  23312=>"000100110",
  23313=>"101000010",
  23314=>"110110000",
  23315=>"011010110",
  23316=>"110000000",
  23317=>"010001000",
  23318=>"111101100",
  23319=>"100111100",
  23320=>"001000001",
  23321=>"010000110",
  23322=>"000111111",
  23323=>"011111010",
  23324=>"001011001",
  23325=>"010010000",
  23326=>"111001011",
  23327=>"000000000",
  23328=>"010110100",
  23329=>"100011001",
  23330=>"100011010",
  23331=>"011100011",
  23332=>"110110000",
  23333=>"110100001",
  23334=>"000010111",
  23335=>"000010001",
  23336=>"110111000",
  23337=>"111001101",
  23338=>"111111000",
  23339=>"011001011",
  23340=>"000010010",
  23341=>"100101011",
  23342=>"000011011",
  23343=>"101010101",
  23344=>"001001110",
  23345=>"100100110",
  23346=>"110110001",
  23347=>"100010000",
  23348=>"000010001",
  23349=>"000100111",
  23350=>"100100010",
  23351=>"000101000",
  23352=>"001010000",
  23353=>"101100110",
  23354=>"001001001",
  23355=>"101010010",
  23356=>"101101001",
  23357=>"111001100",
  23358=>"000000000",
  23359=>"111110001",
  23360=>"010010100",
  23361=>"101101011",
  23362=>"101110111",
  23363=>"000110011",
  23364=>"010100101",
  23365=>"001010111",
  23366=>"111010011",
  23367=>"010000000",
  23368=>"111101011",
  23369=>"011011101",
  23370=>"010110111",
  23371=>"111000111",
  23372=>"110101100",
  23373=>"001101000",
  23374=>"000100001",
  23375=>"010110000",
  23376=>"110000001",
  23377=>"101110100",
  23378=>"000000001",
  23379=>"000110100",
  23380=>"111001111",
  23381=>"010100101",
  23382=>"011100010",
  23383=>"000101101",
  23384=>"001001001",
  23385=>"110111000",
  23386=>"101110011",
  23387=>"001001001",
  23388=>"000000011",
  23389=>"001001010",
  23390=>"101011101",
  23391=>"100101001",
  23392=>"011111101",
  23393=>"001110000",
  23394=>"000011001",
  23395=>"100110101",
  23396=>"100100110",
  23397=>"101001000",
  23398=>"011110000",
  23399=>"111111001",
  23400=>"101011010",
  23401=>"100001000",
  23402=>"110000101",
  23403=>"011011010",
  23404=>"001000000",
  23405=>"010010110",
  23406=>"000010000",
  23407=>"101100100",
  23408=>"110000110",
  23409=>"111011111",
  23410=>"001111001",
  23411=>"010010010",
  23412=>"010111010",
  23413=>"101001100",
  23414=>"111011110",
  23415=>"000111110",
  23416=>"110011110",
  23417=>"110001110",
  23418=>"110110110",
  23419=>"001110010",
  23420=>"001100011",
  23421=>"010010010",
  23422=>"001010110",
  23423=>"111111011",
  23424=>"111110000",
  23425=>"011010111",
  23426=>"110110110",
  23427=>"010010100",
  23428=>"000010001",
  23429=>"001000110",
  23430=>"011001010",
  23431=>"011010100",
  23432=>"100100010",
  23433=>"111011011",
  23434=>"101101110",
  23435=>"011100111",
  23436=>"000010101",
  23437=>"011001100",
  23438=>"100001011",
  23439=>"011101101",
  23440=>"011111100",
  23441=>"111000011",
  23442=>"000010111",
  23443=>"001001000",
  23444=>"001011111",
  23445=>"001111100",
  23446=>"011000001",
  23447=>"101000010",
  23448=>"100100001",
  23449=>"111011010",
  23450=>"000001011",
  23451=>"010110101",
  23452=>"100110101",
  23453=>"111101001",
  23454=>"100010001",
  23455=>"010011000",
  23456=>"001000000",
  23457=>"011111011",
  23458=>"010011111",
  23459=>"010011000",
  23460=>"010011010",
  23461=>"000101111",
  23462=>"110000110",
  23463=>"011001110",
  23464=>"010010001",
  23465=>"000001000",
  23466=>"100110000",
  23467=>"011111110",
  23468=>"100000011",
  23469=>"110010001",
  23470=>"110111100",
  23471=>"000100010",
  23472=>"111011110",
  23473=>"101010000",
  23474=>"100100000",
  23475=>"010100011",
  23476=>"001010001",
  23477=>"000111110",
  23478=>"110111010",
  23479=>"001110110",
  23480=>"111101111",
  23481=>"010000100",
  23482=>"001001000",
  23483=>"010111000",
  23484=>"000101000",
  23485=>"010000000",
  23486=>"100111000",
  23487=>"101011000",
  23488=>"011011101",
  23489=>"101011110",
  23490=>"110011101",
  23491=>"000100010",
  23492=>"101001011",
  23493=>"111111011",
  23494=>"011100111",
  23495=>"101101111",
  23496=>"010011100",
  23497=>"010001111",
  23498=>"011100000",
  23499=>"011101000",
  23500=>"001111101",
  23501=>"101100111",
  23502=>"100101110",
  23503=>"100101111",
  23504=>"111011110",
  23505=>"011011001",
  23506=>"001010110",
  23507=>"110100110",
  23508=>"010001000",
  23509=>"011000100",
  23510=>"101001110",
  23511=>"001010100",
  23512=>"111011101",
  23513=>"011010000",
  23514=>"100000100",
  23515=>"111110010",
  23516=>"110000000",
  23517=>"111100101",
  23518=>"001001101",
  23519=>"010100000",
  23520=>"001010100",
  23521=>"001100100",
  23522=>"001100001",
  23523=>"100011000",
  23524=>"010111010",
  23525=>"100000110",
  23526=>"000111100",
  23527=>"000100000",
  23528=>"000011110",
  23529=>"110110000",
  23530=>"101001000",
  23531=>"000110100",
  23532=>"001100111",
  23533=>"010100001",
  23534=>"011100000",
  23535=>"101111111",
  23536=>"110111101",
  23537=>"010111110",
  23538=>"010110111",
  23539=>"010011011",
  23540=>"110110110",
  23541=>"111110001",
  23542=>"010000101",
  23543=>"101000110",
  23544=>"111110010",
  23545=>"100010010",
  23546=>"001000011",
  23547=>"100101001",
  23548=>"111001010",
  23549=>"011100010",
  23550=>"011101010",
  23551=>"011011111",
  23552=>"110100101",
  23553=>"100010010",
  23554=>"100000011",
  23555=>"100110111",
  23556=>"001110001",
  23557=>"001101011",
  23558=>"010101001",
  23559=>"010010110",
  23560=>"010011011",
  23561=>"010001101",
  23562=>"000110000",
  23563=>"010001101",
  23564=>"010010001",
  23565=>"111100001",
  23566=>"100000000",
  23567=>"100111011",
  23568=>"100011100",
  23569=>"010000001",
  23570=>"000001000",
  23571=>"011000011",
  23572=>"111111011",
  23573=>"100011010",
  23574=>"101110110",
  23575=>"101000001",
  23576=>"110110011",
  23577=>"111010110",
  23578=>"000001100",
  23579=>"011000000",
  23580=>"100000100",
  23581=>"011100111",
  23582=>"011010111",
  23583=>"101010100",
  23584=>"100101010",
  23585=>"100000010",
  23586=>"000000010",
  23587=>"010010010",
  23588=>"101110101",
  23589=>"010101110",
  23590=>"111110000",
  23591=>"010000000",
  23592=>"110000010",
  23593=>"000101001",
  23594=>"011110110",
  23595=>"110010111",
  23596=>"101010001",
  23597=>"010010001",
  23598=>"010110011",
  23599=>"001001101",
  23600=>"110110011",
  23601=>"010010111",
  23602=>"011101100",
  23603=>"010010011",
  23604=>"010011111",
  23605=>"000110010",
  23606=>"001001110",
  23607=>"111101010",
  23608=>"000111011",
  23609=>"111110000",
  23610=>"110111110",
  23611=>"011000111",
  23612=>"100000010",
  23613=>"000000000",
  23614=>"111111001",
  23615=>"111010110",
  23616=>"110011001",
  23617=>"001111000",
  23618=>"101100011",
  23619=>"010011010",
  23620=>"110111001",
  23621=>"101000111",
  23622=>"001101010",
  23623=>"101101010",
  23624=>"010111010",
  23625=>"100100001",
  23626=>"001010010",
  23627=>"001001110",
  23628=>"111100010",
  23629=>"111011011",
  23630=>"011001001",
  23631=>"101011110",
  23632=>"010000010",
  23633=>"111001011",
  23634=>"110111010",
  23635=>"110010001",
  23636=>"100100100",
  23637=>"000000011",
  23638=>"101100101",
  23639=>"001000100",
  23640=>"011000110",
  23641=>"110110000",
  23642=>"000001011",
  23643=>"000000011",
  23644=>"000100101",
  23645=>"100010010",
  23646=>"010101110",
  23647=>"100001001",
  23648=>"011010111",
  23649=>"100000001",
  23650=>"100001101",
  23651=>"001101100",
  23652=>"110110011",
  23653=>"111110010",
  23654=>"101100101",
  23655=>"100000111",
  23656=>"101100011",
  23657=>"001010111",
  23658=>"111000100",
  23659=>"110110000",
  23660=>"000010110",
  23661=>"111000111",
  23662=>"000011000",
  23663=>"101011010",
  23664=>"000101000",
  23665=>"101100111",
  23666=>"011100110",
  23667=>"001110100",
  23668=>"101101010",
  23669=>"101011010",
  23670=>"101100101",
  23671=>"100010100",
  23672=>"110110010",
  23673=>"101011010",
  23674=>"010110010",
  23675=>"001100110",
  23676=>"000000000",
  23677=>"101001010",
  23678=>"101000100",
  23679=>"010100000",
  23680=>"010011111",
  23681=>"101101100",
  23682=>"100000000",
  23683=>"001111000",
  23684=>"100110000",
  23685=>"011011010",
  23686=>"100011001",
  23687=>"111010011",
  23688=>"001101010",
  23689=>"000010011",
  23690=>"010010011",
  23691=>"011101100",
  23692=>"001100110",
  23693=>"001011111",
  23694=>"100100001",
  23695=>"110111110",
  23696=>"110110100",
  23697=>"111000000",
  23698=>"100011111",
  23699=>"001100000",
  23700=>"100111101",
  23701=>"010100010",
  23702=>"000011110",
  23703=>"111001001",
  23704=>"011001100",
  23705=>"001100101",
  23706=>"111111010",
  23707=>"100001000",
  23708=>"000000000",
  23709=>"001011111",
  23710=>"111111110",
  23711=>"110100101",
  23712=>"011110101",
  23713=>"000110010",
  23714=>"100100001",
  23715=>"110001011",
  23716=>"001100011",
  23717=>"110111010",
  23718=>"110100111",
  23719=>"000000000",
  23720=>"111101100",
  23721=>"101001000",
  23722=>"110011011",
  23723=>"100111000",
  23724=>"100001000",
  23725=>"110111010",
  23726=>"001110101",
  23727=>"110110111",
  23728=>"111001100",
  23729=>"001110110",
  23730=>"100000111",
  23731=>"010101010",
  23732=>"000001000",
  23733=>"011010100",
  23734=>"010111111",
  23735=>"010110101",
  23736=>"001110101",
  23737=>"100000010",
  23738=>"100000010",
  23739=>"101010010",
  23740=>"000010000",
  23741=>"100101011",
  23742=>"100001101",
  23743=>"000000000",
  23744=>"110101111",
  23745=>"100011111",
  23746=>"110101011",
  23747=>"010100101",
  23748=>"101001110",
  23749=>"010011000",
  23750=>"101111110",
  23751=>"011100000",
  23752=>"001100110",
  23753=>"011001110",
  23754=>"100101010",
  23755=>"111111010",
  23756=>"001101000",
  23757=>"000000111",
  23758=>"000111001",
  23759=>"000010010",
  23760=>"001000110",
  23761=>"000111010",
  23762=>"011100100",
  23763=>"101001000",
  23764=>"011100111",
  23765=>"000000100",
  23766=>"010010100",
  23767=>"101011101",
  23768=>"101101011",
  23769=>"011111011",
  23770=>"010111010",
  23771=>"011111000",
  23772=>"111100000",
  23773=>"100001101",
  23774=>"010110001",
  23775=>"110111101",
  23776=>"101001000",
  23777=>"011111001",
  23778=>"010110111",
  23779=>"100000101",
  23780=>"101001001",
  23781=>"000101101",
  23782=>"000010010",
  23783=>"110101110",
  23784=>"000101010",
  23785=>"010011100",
  23786=>"100100011",
  23787=>"000010111",
  23788=>"000000110",
  23789=>"000101101",
  23790=>"011111010",
  23791=>"100000101",
  23792=>"110101111",
  23793=>"010011000",
  23794=>"110010010",
  23795=>"101010100",
  23796=>"000010101",
  23797=>"010111110",
  23798=>"101001101",
  23799=>"000111101",
  23800=>"111101110",
  23801=>"011010110",
  23802=>"100111111",
  23803=>"010100101",
  23804=>"011111110",
  23805=>"101000001",
  23806=>"000101000",
  23807=>"110000011",
  23808=>"100111001",
  23809=>"010110001",
  23810=>"101011100",
  23811=>"111000111",
  23812=>"000011110",
  23813=>"100111011",
  23814=>"000011101",
  23815=>"001111000",
  23816=>"111010000",
  23817=>"011110111",
  23818=>"110011110",
  23819=>"100000001",
  23820=>"110101010",
  23821=>"010001100",
  23822=>"001011101",
  23823=>"100010000",
  23824=>"010000111",
  23825=>"001000010",
  23826=>"100110001",
  23827=>"110011100",
  23828=>"101000111",
  23829=>"100111011",
  23830=>"001000110",
  23831=>"100111010",
  23832=>"011101011",
  23833=>"111101111",
  23834=>"010011111",
  23835=>"001010001",
  23836=>"111110000",
  23837=>"010110100",
  23838=>"010100011",
  23839=>"000001000",
  23840=>"011010000",
  23841=>"001111011",
  23842=>"111000011",
  23843=>"000110110",
  23844=>"011100001",
  23845=>"000010000",
  23846=>"101111101",
  23847=>"000000100",
  23848=>"101100101",
  23849=>"101110000",
  23850=>"111010010",
  23851=>"010111110",
  23852=>"101110011",
  23853=>"100010101",
  23854=>"110010111",
  23855=>"100010000",
  23856=>"011010111",
  23857=>"011110000",
  23858=>"010010100",
  23859=>"111010001",
  23860=>"001001110",
  23861=>"000110110",
  23862=>"000001010",
  23863=>"011011011",
  23864=>"111100011",
  23865=>"001010000",
  23866=>"000011000",
  23867=>"100110110",
  23868=>"110101011",
  23869=>"100101010",
  23870=>"101010100",
  23871=>"101011101",
  23872=>"110101111",
  23873=>"011111011",
  23874=>"010100010",
  23875=>"110111001",
  23876=>"101101000",
  23877=>"011100011",
  23878=>"000000110",
  23879=>"000011000",
  23880=>"010100000",
  23881=>"000111001",
  23882=>"001111001",
  23883=>"100010100",
  23884=>"000110011",
  23885=>"010001010",
  23886=>"010111001",
  23887=>"011110011",
  23888=>"001011011",
  23889=>"111011010",
  23890=>"011100010",
  23891=>"001000111",
  23892=>"000010010",
  23893=>"101101010",
  23894=>"001110111",
  23895=>"110000010",
  23896=>"010000001",
  23897=>"001011000",
  23898=>"010110001",
  23899=>"001011000",
  23900=>"101010111",
  23901=>"000010010",
  23902=>"110111000",
  23903=>"000001100",
  23904=>"100111010",
  23905=>"001001101",
  23906=>"111100011",
  23907=>"101101001",
  23908=>"101110100",
  23909=>"101011110",
  23910=>"011100000",
  23911=>"000001110",
  23912=>"011111011",
  23913=>"110001110",
  23914=>"000111011",
  23915=>"111110101",
  23916=>"001101001",
  23917=>"110101010",
  23918=>"111001101",
  23919=>"011000100",
  23920=>"000100000",
  23921=>"001101111",
  23922=>"000100110",
  23923=>"101110010",
  23924=>"000000110",
  23925=>"101110110",
  23926=>"000000010",
  23927=>"000001010",
  23928=>"001100101",
  23929=>"101001011",
  23930=>"111111100",
  23931=>"000010100",
  23932=>"011111111",
  23933=>"110001011",
  23934=>"011000001",
  23935=>"110010111",
  23936=>"111011101",
  23937=>"000100111",
  23938=>"100111110",
  23939=>"111010001",
  23940=>"101010111",
  23941=>"010110100",
  23942=>"101101101",
  23943=>"110011001",
  23944=>"100100001",
  23945=>"110100100",
  23946=>"011110000",
  23947=>"000011001",
  23948=>"111001011",
  23949=>"110011110",
  23950=>"010001101",
  23951=>"010001000",
  23952=>"110101101",
  23953=>"101000111",
  23954=>"011110000",
  23955=>"000000101",
  23956=>"000010110",
  23957=>"010111010",
  23958=>"111110100",
  23959=>"011001001",
  23960=>"001100111",
  23961=>"011110100",
  23962=>"000001011",
  23963=>"010100010",
  23964=>"101111010",
  23965=>"111010001",
  23966=>"100110100",
  23967=>"101110100",
  23968=>"001110111",
  23969=>"100001010",
  23970=>"001101001",
  23971=>"010000010",
  23972=>"100000101",
  23973=>"110001110",
  23974=>"101110101",
  23975=>"110001001",
  23976=>"100011001",
  23977=>"001111001",
  23978=>"000001100",
  23979=>"111101101",
  23980=>"111101001",
  23981=>"000100111",
  23982=>"000110110",
  23983=>"011001000",
  23984=>"010010100",
  23985=>"111001001",
  23986=>"011110001",
  23987=>"001010001",
  23988=>"011010101",
  23989=>"100100010",
  23990=>"001000111",
  23991=>"110101111",
  23992=>"111101011",
  23993=>"001100011",
  23994=>"000000011",
  23995=>"000101000",
  23996=>"001001010",
  23997=>"001000000",
  23998=>"100010111",
  23999=>"111111101",
  24000=>"101111101",
  24001=>"110001011",
  24002=>"111000111",
  24003=>"000100100",
  24004=>"110111000",
  24005=>"000101101",
  24006=>"111110000",
  24007=>"010110111",
  24008=>"111010011",
  24009=>"110111001",
  24010=>"100100111",
  24011=>"111100100",
  24012=>"011100100",
  24013=>"111001110",
  24014=>"111101101",
  24015=>"010100011",
  24016=>"110011001",
  24017=>"111011010",
  24018=>"000100100",
  24019=>"010001100",
  24020=>"111001000",
  24021=>"111100001",
  24022=>"001000000",
  24023=>"101010111",
  24024=>"100111101",
  24025=>"110111000",
  24026=>"111001110",
  24027=>"000110111",
  24028=>"010011001",
  24029=>"101100001",
  24030=>"110011011",
  24031=>"000010111",
  24032=>"100011011",
  24033=>"101010010",
  24034=>"101001110",
  24035=>"011101011",
  24036=>"111001101",
  24037=>"010110101",
  24038=>"011001011",
  24039=>"000111010",
  24040=>"110000111",
  24041=>"011011101",
  24042=>"101101101",
  24043=>"100100001",
  24044=>"001010010",
  24045=>"110100111",
  24046=>"111010101",
  24047=>"010100100",
  24048=>"000001100",
  24049=>"010101110",
  24050=>"001110100",
  24051=>"011010000",
  24052=>"111111110",
  24053=>"111111100",
  24054=>"100000011",
  24055=>"000110100",
  24056=>"001111010",
  24057=>"101101011",
  24058=>"010101011",
  24059=>"010000010",
  24060=>"111100100",
  24061=>"001001101",
  24062=>"000010010",
  24063=>"111001001",
  24064=>"010000101",
  24065=>"010000110",
  24066=>"110011110",
  24067=>"011001111",
  24068=>"000110110",
  24069=>"000100101",
  24070=>"000010100",
  24071=>"111111111",
  24072=>"000001010",
  24073=>"011111111",
  24074=>"101011101",
  24075=>"110001101",
  24076=>"111011110",
  24077=>"101101111",
  24078=>"010101110",
  24079=>"111111010",
  24080=>"010011101",
  24081=>"101111100",
  24082=>"000111001",
  24083=>"111010101",
  24084=>"001000111",
  24085=>"100110101",
  24086=>"100011101",
  24087=>"110011111",
  24088=>"010101110",
  24089=>"010100001",
  24090=>"110111111",
  24091=>"010111010",
  24092=>"101000011",
  24093=>"010010101",
  24094=>"001000000",
  24095=>"110111101",
  24096=>"000100111",
  24097=>"001110001",
  24098=>"110001100",
  24099=>"111001001",
  24100=>"100001111",
  24101=>"101000010",
  24102=>"110010101",
  24103=>"111001101",
  24104=>"001100010",
  24105=>"100111011",
  24106=>"111000100",
  24107=>"110110000",
  24108=>"000000101",
  24109=>"000001001",
  24110=>"000111000",
  24111=>"101010001",
  24112=>"011110010",
  24113=>"011101010",
  24114=>"110111110",
  24115=>"010000100",
  24116=>"001110010",
  24117=>"110001000",
  24118=>"010000100",
  24119=>"000001110",
  24120=>"001010111",
  24121=>"101000111",
  24122=>"000100011",
  24123=>"001111101",
  24124=>"011101000",
  24125=>"001100011",
  24126=>"100111000",
  24127=>"010010110",
  24128=>"100000100",
  24129=>"000000011",
  24130=>"000111011",
  24131=>"010000001",
  24132=>"010011010",
  24133=>"100100100",
  24134=>"100111100",
  24135=>"001000011",
  24136=>"000001010",
  24137=>"110101100",
  24138=>"100100001",
  24139=>"111101011",
  24140=>"111010010",
  24141=>"000000010",
  24142=>"111101110",
  24143=>"011001000",
  24144=>"111010010",
  24145=>"010111111",
  24146=>"100111000",
  24147=>"001000000",
  24148=>"101001001",
  24149=>"011001011",
  24150=>"011101110",
  24151=>"001011001",
  24152=>"001010011",
  24153=>"001011001",
  24154=>"101000110",
  24155=>"000001001",
  24156=>"001000110",
  24157=>"011001000",
  24158=>"110110001",
  24159=>"010100001",
  24160=>"110100011",
  24161=>"000010110",
  24162=>"110000010",
  24163=>"101011001",
  24164=>"111111101",
  24165=>"100000100",
  24166=>"000001100",
  24167=>"001000101",
  24168=>"100011100",
  24169=>"010101001",
  24170=>"100110100",
  24171=>"101011101",
  24172=>"000100110",
  24173=>"001101101",
  24174=>"011001011",
  24175=>"001111010",
  24176=>"000000101",
  24177=>"101100011",
  24178=>"010111111",
  24179=>"011000000",
  24180=>"101001001",
  24181=>"110000101",
  24182=>"011100010",
  24183=>"101001010",
  24184=>"111101001",
  24185=>"011010101",
  24186=>"001111000",
  24187=>"100000000",
  24188=>"000000010",
  24189=>"111111011",
  24190=>"001000110",
  24191=>"110011100",
  24192=>"000101011",
  24193=>"000100101",
  24194=>"111001000",
  24195=>"100011000",
  24196=>"100110100",
  24197=>"000001100",
  24198=>"101100001",
  24199=>"011000010",
  24200=>"011101101",
  24201=>"011100000",
  24202=>"101000011",
  24203=>"101101011",
  24204=>"001111100",
  24205=>"010101111",
  24206=>"000110011",
  24207=>"111011110",
  24208=>"010011110",
  24209=>"101101011",
  24210=>"000010010",
  24211=>"011111101",
  24212=>"101010101",
  24213=>"110101100",
  24214=>"100111101",
  24215=>"000110101",
  24216=>"110011101",
  24217=>"011101000",
  24218=>"011111001",
  24219=>"001111000",
  24220=>"110000000",
  24221=>"000100001",
  24222=>"100100100",
  24223=>"000000011",
  24224=>"001111000",
  24225=>"000001111",
  24226=>"000011101",
  24227=>"001000101",
  24228=>"101011011",
  24229=>"101100111",
  24230=>"111001110",
  24231=>"100000001",
  24232=>"110100101",
  24233=>"110001111",
  24234=>"000000111",
  24235=>"111110101",
  24236=>"001111010",
  24237=>"111011100",
  24238=>"101001010",
  24239=>"111100101",
  24240=>"101111001",
  24241=>"001101111",
  24242=>"001111111",
  24243=>"101011101",
  24244=>"110110000",
  24245=>"110100010",
  24246=>"001100111",
  24247=>"100001111",
  24248=>"010110100",
  24249=>"111110110",
  24250=>"101010100",
  24251=>"011011000",
  24252=>"001001000",
  24253=>"010100010",
  24254=>"000110010",
  24255=>"001011011",
  24256=>"101011011",
  24257=>"001100110",
  24258=>"100010101",
  24259=>"101000101",
  24260=>"110101111",
  24261=>"100101111",
  24262=>"000011101",
  24263=>"100111000",
  24264=>"001110111",
  24265=>"100010010",
  24266=>"010011100",
  24267=>"110110010",
  24268=>"100111110",
  24269=>"010111100",
  24270=>"110111001",
  24271=>"101011011",
  24272=>"101010000",
  24273=>"010100111",
  24274=>"110000110",
  24275=>"100101001",
  24276=>"111110000",
  24277=>"011001010",
  24278=>"001000111",
  24279=>"101101000",
  24280=>"000110101",
  24281=>"100100010",
  24282=>"110011000",
  24283=>"111100010",
  24284=>"100000101",
  24285=>"011000100",
  24286=>"111100110",
  24287=>"110101110",
  24288=>"110101101",
  24289=>"100011111",
  24290=>"101011000",
  24291=>"100100010",
  24292=>"100001101",
  24293=>"100001010",
  24294=>"111111110",
  24295=>"111100010",
  24296=>"110000111",
  24297=>"000001111",
  24298=>"100101111",
  24299=>"011110101",
  24300=>"111110010",
  24301=>"010110010",
  24302=>"100001011",
  24303=>"001100011",
  24304=>"101011010",
  24305=>"111011001",
  24306=>"000111111",
  24307=>"101100101",
  24308=>"011010110",
  24309=>"100001100",
  24310=>"101100010",
  24311=>"001010111",
  24312=>"111101100",
  24313=>"001101011",
  24314=>"101101110",
  24315=>"100101110",
  24316=>"000111000",
  24317=>"111001100",
  24318=>"110011111",
  24319=>"100111000",
  24320=>"010000101",
  24321=>"101010000",
  24322=>"101010101",
  24323=>"010110100",
  24324=>"001111101",
  24325=>"101011001",
  24326=>"011000011",
  24327=>"110010110",
  24328=>"010111101",
  24329=>"101011000",
  24330=>"101001110",
  24331=>"001111011",
  24332=>"100000000",
  24333=>"110100111",
  24334=>"001100000",
  24335=>"101111101",
  24336=>"100010111",
  24337=>"100110000",
  24338=>"010100110",
  24339=>"010110010",
  24340=>"000101110",
  24341=>"000010110",
  24342=>"101101100",
  24343=>"000111101",
  24344=>"100111110",
  24345=>"101000110",
  24346=>"010101111",
  24347=>"101011100",
  24348=>"110011011",
  24349=>"011101001",
  24350=>"000111100",
  24351=>"100010010",
  24352=>"110100011",
  24353=>"101100000",
  24354=>"110010111",
  24355=>"001101111",
  24356=>"010111101",
  24357=>"001001010",
  24358=>"100111001",
  24359=>"100011100",
  24360=>"001101100",
  24361=>"111011110",
  24362=>"001111100",
  24363=>"111001101",
  24364=>"110000110",
  24365=>"000100100",
  24366=>"010011111",
  24367=>"111111110",
  24368=>"011000110",
  24369=>"000000110",
  24370=>"001101011",
  24371=>"011111001",
  24372=>"100111010",
  24373=>"111100111",
  24374=>"101011000",
  24375=>"111101000",
  24376=>"010011000",
  24377=>"101000010",
  24378=>"110010110",
  24379=>"110010110",
  24380=>"100100001",
  24381=>"110100010",
  24382=>"000000111",
  24383=>"011111101",
  24384=>"000100000",
  24385=>"000000111",
  24386=>"111111011",
  24387=>"001010101",
  24388=>"111011000",
  24389=>"001101111",
  24390=>"000011110",
  24391=>"000101001",
  24392=>"010110111",
  24393=>"111111011",
  24394=>"111101001",
  24395=>"010100011",
  24396=>"001010110",
  24397=>"111101011",
  24398=>"001101001",
  24399=>"000001010",
  24400=>"000001010",
  24401=>"001001000",
  24402=>"100110001",
  24403=>"101001101",
  24404=>"011011000",
  24405=>"000111100",
  24406=>"110100011",
  24407=>"011011001",
  24408=>"111011001",
  24409=>"111110001",
  24410=>"111000010",
  24411=>"110011111",
  24412=>"110010011",
  24413=>"100110101",
  24414=>"100000111",
  24415=>"000000010",
  24416=>"011010000",
  24417=>"110010011",
  24418=>"000011110",
  24419=>"001011000",
  24420=>"111100110",
  24421=>"010010111",
  24422=>"001000000",
  24423=>"110000100",
  24424=>"001001010",
  24425=>"101101110",
  24426=>"100000101",
  24427=>"101101110",
  24428=>"001101000",
  24429=>"010010010",
  24430=>"111001100",
  24431=>"011000011",
  24432=>"111001000",
  24433=>"110001100",
  24434=>"000010001",
  24435=>"100100100",
  24436=>"010100000",
  24437=>"011001110",
  24438=>"101111111",
  24439=>"100001001",
  24440=>"000000001",
  24441=>"100010100",
  24442=>"001110111",
  24443=>"101011100",
  24444=>"110011111",
  24445=>"000000000",
  24446=>"000111110",
  24447=>"111110000",
  24448=>"001100101",
  24449=>"000010010",
  24450=>"101110101",
  24451=>"010010000",
  24452=>"001000010",
  24453=>"011111010",
  24454=>"001000101",
  24455=>"100011110",
  24456=>"100111101",
  24457=>"010100010",
  24458=>"111000001",
  24459=>"101000001",
  24460=>"010100011",
  24461=>"000110100",
  24462=>"010100110",
  24463=>"101110100",
  24464=>"100010110",
  24465=>"111000101",
  24466=>"100001111",
  24467=>"011011111",
  24468=>"110111100",
  24469=>"111100010",
  24470=>"110011100",
  24471=>"110010111",
  24472=>"001111010",
  24473=>"000110011",
  24474=>"001100111",
  24475=>"000100000",
  24476=>"011010111",
  24477=>"011110000",
  24478=>"101100101",
  24479=>"011001000",
  24480=>"001000100",
  24481=>"010111100",
  24482=>"101010010",
  24483=>"111101100",
  24484=>"110100001",
  24485=>"000111000",
  24486=>"100000100",
  24487=>"110010110",
  24488=>"111101001",
  24489=>"010101111",
  24490=>"101100001",
  24491=>"000100010",
  24492=>"000100110",
  24493=>"001101000",
  24494=>"101001111",
  24495=>"111010111",
  24496=>"110001111",
  24497=>"101111100",
  24498=>"101111001",
  24499=>"110010010",
  24500=>"110100100",
  24501=>"111110101",
  24502=>"000000101",
  24503=>"101000101",
  24504=>"111001001",
  24505=>"011000000",
  24506=>"010011110",
  24507=>"000101100",
  24508=>"110000101",
  24509=>"101011101",
  24510=>"110100001",
  24511=>"010001111",
  24512=>"110101111",
  24513=>"011111011",
  24514=>"011011000",
  24515=>"000001011",
  24516=>"100111111",
  24517=>"110101111",
  24518=>"001101100",
  24519=>"010011100",
  24520=>"001100011",
  24521=>"000010000",
  24522=>"001000101",
  24523=>"011001100",
  24524=>"000101011",
  24525=>"100100111",
  24526=>"101000001",
  24527=>"001011100",
  24528=>"011100010",
  24529=>"001100110",
  24530=>"001101111",
  24531=>"000101101",
  24532=>"111000001",
  24533=>"011011010",
  24534=>"000111100",
  24535=>"101100101",
  24536=>"001011110",
  24537=>"111001010",
  24538=>"111111100",
  24539=>"010011000",
  24540=>"011111110",
  24541=>"101110111",
  24542=>"111101011",
  24543=>"000010010",
  24544=>"000000000",
  24545=>"111111001",
  24546=>"101110010",
  24547=>"000110100",
  24548=>"010000111",
  24549=>"000011001",
  24550=>"111100111",
  24551=>"010011010",
  24552=>"110100000",
  24553=>"111000000",
  24554=>"010001000",
  24555=>"001100111",
  24556=>"000111010",
  24557=>"000100111",
  24558=>"010110000",
  24559=>"101000101",
  24560=>"111101100",
  24561=>"000100100",
  24562=>"111111101",
  24563=>"111100100",
  24564=>"001001110",
  24565=>"000010110",
  24566=>"100111000",
  24567=>"110110101",
  24568=>"101100011",
  24569=>"110101110",
  24570=>"100100000",
  24571=>"010001111",
  24572=>"100010110",
  24573=>"100100111",
  24574=>"100011110",
  24575=>"000000110",
  24576=>"111000000",
  24577=>"110111110",
  24578=>"000011011",
  24579=>"110111010",
  24580=>"000110101",
  24581=>"010001010",
  24582=>"110111101",
  24583=>"111001011",
  24584=>"111011001",
  24585=>"110110101",
  24586=>"001001101",
  24587=>"100000001",
  24588=>"000101000",
  24589=>"010110101",
  24590=>"101010100",
  24591=>"100100101",
  24592=>"111111011",
  24593=>"001001010",
  24594=>"000001100",
  24595=>"001110110",
  24596=>"001011100",
  24597=>"101000111",
  24598=>"100000100",
  24599=>"000010010",
  24600=>"011011110",
  24601=>"100010111",
  24602=>"010100010",
  24603=>"001011111",
  24604=>"111101111",
  24605=>"011010011",
  24606=>"010010001",
  24607=>"011000001",
  24608=>"101101000",
  24609=>"001110011",
  24610=>"000001010",
  24611=>"000001001",
  24612=>"100101101",
  24613=>"101110101",
  24614=>"100001010",
  24615=>"010100001",
  24616=>"101100011",
  24617=>"111000010",
  24618=>"000011010",
  24619=>"011110100",
  24620=>"110101111",
  24621=>"101000100",
  24622=>"111011010",
  24623=>"011011110",
  24624=>"111000010",
  24625=>"001010111",
  24626=>"101101011",
  24627=>"100100101",
  24628=>"100111011",
  24629=>"011011100",
  24630=>"001010110",
  24631=>"101110010",
  24632=>"001100100",
  24633=>"100001101",
  24634=>"111011000",
  24635=>"101000000",
  24636=>"101000100",
  24637=>"111010101",
  24638=>"010000001",
  24639=>"110011101",
  24640=>"011111011",
  24641=>"111001100",
  24642=>"110110111",
  24643=>"111001101",
  24644=>"011010110",
  24645=>"101100111",
  24646=>"111101001",
  24647=>"000011111",
  24648=>"010101011",
  24649=>"110010000",
  24650=>"111101101",
  24651=>"010111000",
  24652=>"111010001",
  24653=>"011111101",
  24654=>"111000010",
  24655=>"101001111",
  24656=>"001110011",
  24657=>"001011001",
  24658=>"101000010",
  24659=>"101000000",
  24660=>"110000010",
  24661=>"100101000",
  24662=>"110100111",
  24663=>"011000111",
  24664=>"100000111",
  24665=>"110001101",
  24666=>"111011000",
  24667=>"110010011",
  24668=>"100010100",
  24669=>"000001011",
  24670=>"101001000",
  24671=>"011110000",
  24672=>"000001001",
  24673=>"010100101",
  24674=>"001010010",
  24675=>"000100001",
  24676=>"101100001",
  24677=>"111110100",
  24678=>"001001110",
  24679=>"011110010",
  24680=>"101011010",
  24681=>"001011010",
  24682=>"100000001",
  24683=>"011101100",
  24684=>"001011100",
  24685=>"001010100",
  24686=>"101110011",
  24687=>"000010011",
  24688=>"111010101",
  24689=>"010101000",
  24690=>"101000110",
  24691=>"000110110",
  24692=>"110110001",
  24693=>"101100111",
  24694=>"011110111",
  24695=>"001100010",
  24696=>"001110010",
  24697=>"110111000",
  24698=>"011010010",
  24699=>"001000100",
  24700=>"001000010",
  24701=>"010100001",
  24702=>"000001001",
  24703=>"000001011",
  24704=>"000110001",
  24705=>"011010010",
  24706=>"001101000",
  24707=>"101101111",
  24708=>"010011000",
  24709=>"001110110",
  24710=>"000011000",
  24711=>"101000110",
  24712=>"010100101",
  24713=>"101111001",
  24714=>"011010100",
  24715=>"110101010",
  24716=>"000011101",
  24717=>"111010010",
  24718=>"111101111",
  24719=>"101010100",
  24720=>"001110001",
  24721=>"111000110",
  24722=>"111011011",
  24723=>"001001101",
  24724=>"110010001",
  24725=>"111000110",
  24726=>"111011001",
  24727=>"000110101",
  24728=>"111101101",
  24729=>"010001011",
  24730=>"010010011",
  24731=>"100000110",
  24732=>"011100101",
  24733=>"111110110",
  24734=>"001011110",
  24735=>"110111011",
  24736=>"101101100",
  24737=>"000000100",
  24738=>"011100110",
  24739=>"000111100",
  24740=>"100000000",
  24741=>"001011001",
  24742=>"110100000",
  24743=>"000110100",
  24744=>"011110011",
  24745=>"110110101",
  24746=>"011011000",
  24747=>"101110110",
  24748=>"001101010",
  24749=>"011010110",
  24750=>"000011010",
  24751=>"010010110",
  24752=>"110000100",
  24753=>"010000110",
  24754=>"001100100",
  24755=>"001000000",
  24756=>"100000000",
  24757=>"000111011",
  24758=>"100100011",
  24759=>"000000100",
  24760=>"011100111",
  24761=>"000111011",
  24762=>"111110100",
  24763=>"001100010",
  24764=>"011111011",
  24765=>"111110101",
  24766=>"101011101",
  24767=>"001010110",
  24768=>"010010101",
  24769=>"110010011",
  24770=>"001000101",
  24771=>"010100001",
  24772=>"010000111",
  24773=>"101100110",
  24774=>"101010110",
  24775=>"101110111",
  24776=>"101000110",
  24777=>"101000110",
  24778=>"010110000",
  24779=>"110111001",
  24780=>"011111110",
  24781=>"101010011",
  24782=>"001110000",
  24783=>"110100010",
  24784=>"010010010",
  24785=>"001001101",
  24786=>"000001010",
  24787=>"100101000",
  24788=>"010100111",
  24789=>"100011001",
  24790=>"011001001",
  24791=>"000111100",
  24792=>"001110100",
  24793=>"001010000",
  24794=>"100110100",
  24795=>"101101111",
  24796=>"010010101",
  24797=>"100001111",
  24798=>"001001000",
  24799=>"011111101",
  24800=>"111010000",
  24801=>"000001000",
  24802=>"011010000",
  24803=>"010000100",
  24804=>"100001001",
  24805=>"010111001",
  24806=>"101010011",
  24807=>"111110111",
  24808=>"100010110",
  24809=>"010100100",
  24810=>"000100111",
  24811=>"101000111",
  24812=>"100110011",
  24813=>"111110010",
  24814=>"010011100",
  24815=>"010000111",
  24816=>"010101101",
  24817=>"101110110",
  24818=>"110100011",
  24819=>"110010110",
  24820=>"001000001",
  24821=>"111100000",
  24822=>"011000110",
  24823=>"100000111",
  24824=>"011101000",
  24825=>"100011010",
  24826=>"001111001",
  24827=>"000000011",
  24828=>"000100111",
  24829=>"101110010",
  24830=>"111011001",
  24831=>"100101101",
  24832=>"010011111",
  24833=>"111011110",
  24834=>"000101010",
  24835=>"010010101",
  24836=>"100101011",
  24837=>"100001011",
  24838=>"000000010",
  24839=>"100111100",
  24840=>"111110111",
  24841=>"101011101",
  24842=>"011001011",
  24843=>"111101010",
  24844=>"110100011",
  24845=>"111101010",
  24846=>"011111110",
  24847=>"000010011",
  24848=>"111110111",
  24849=>"001001101",
  24850=>"011001010",
  24851=>"100001110",
  24852=>"100111100",
  24853=>"010000010",
  24854=>"010001110",
  24855=>"000101111",
  24856=>"110111000",
  24857=>"111101010",
  24858=>"101010000",
  24859=>"000101110",
  24860=>"101101001",
  24861=>"101100110",
  24862=>"101000010",
  24863=>"000000011",
  24864=>"000100010",
  24865=>"111101011",
  24866=>"011010100",
  24867=>"000011101",
  24868=>"111010001",
  24869=>"010010101",
  24870=>"110011000",
  24871=>"011110110",
  24872=>"111000000",
  24873=>"101011101",
  24874=>"000111111",
  24875=>"001010000",
  24876=>"111001110",
  24877=>"101010000",
  24878=>"000100000",
  24879=>"100011111",
  24880=>"010001111",
  24881=>"000101101",
  24882=>"011001011",
  24883=>"101101101",
  24884=>"111011101",
  24885=>"011001100",
  24886=>"101001011",
  24887=>"110111100",
  24888=>"111010111",
  24889=>"111101110",
  24890=>"110011111",
  24891=>"001010000",
  24892=>"110001100",
  24893=>"111111111",
  24894=>"110011100",
  24895=>"011011010",
  24896=>"010001010",
  24897=>"111101101",
  24898=>"001001000",
  24899=>"010011101",
  24900=>"000100000",
  24901=>"001110101",
  24902=>"010111001",
  24903=>"110101001",
  24904=>"001101010",
  24905=>"000110111",
  24906=>"011001101",
  24907=>"001011100",
  24908=>"000111101",
  24909=>"001010101",
  24910=>"011000011",
  24911=>"001001010",
  24912=>"111001000",
  24913=>"101011000",
  24914=>"000101010",
  24915=>"110010100",
  24916=>"110100011",
  24917=>"011000001",
  24918=>"111000000",
  24919=>"000110101",
  24920=>"010000011",
  24921=>"000010011",
  24922=>"101010000",
  24923=>"000010011",
  24924=>"100001101",
  24925=>"111101100",
  24926=>"100101101",
  24927=>"111101100",
  24928=>"101011110",
  24929=>"000000100",
  24930=>"110010001",
  24931=>"110110101",
  24932=>"111101110",
  24933=>"000011000",
  24934=>"010100101",
  24935=>"010000010",
  24936=>"011001001",
  24937=>"010011001",
  24938=>"101101111",
  24939=>"111001001",
  24940=>"111010000",
  24941=>"001001110",
  24942=>"001011111",
  24943=>"011011001",
  24944=>"111110010",
  24945=>"010001000",
  24946=>"101001000",
  24947=>"100000101",
  24948=>"011100111",
  24949=>"101111110",
  24950=>"001000000",
  24951=>"101110000",
  24952=>"100110011",
  24953=>"000010001",
  24954=>"110000110",
  24955=>"111000000",
  24956=>"011010110",
  24957=>"110001001",
  24958=>"011110111",
  24959=>"111110110",
  24960=>"111001111",
  24961=>"001001110",
  24962=>"000110110",
  24963=>"100100001",
  24964=>"111001000",
  24965=>"000110010",
  24966=>"001000001",
  24967=>"001101001",
  24968=>"000000000",
  24969=>"001100000",
  24970=>"100001001",
  24971=>"011011100",
  24972=>"000000111",
  24973=>"011001011",
  24974=>"101100000",
  24975=>"010011001",
  24976=>"101100101",
  24977=>"010001110",
  24978=>"000000000",
  24979=>"111111110",
  24980=>"100011110",
  24981=>"111000111",
  24982=>"010100001",
  24983=>"111100011",
  24984=>"000010110",
  24985=>"011101100",
  24986=>"111100000",
  24987=>"001011000",
  24988=>"000000000",
  24989=>"000101010",
  24990=>"100011110",
  24991=>"100010101",
  24992=>"000110000",
  24993=>"111100001",
  24994=>"101000110",
  24995=>"111001100",
  24996=>"010010000",
  24997=>"111100111",
  24998=>"011011000",
  24999=>"101000101",
  25000=>"100011010",
  25001=>"001100101",
  25002=>"000100101",
  25003=>"110110110",
  25004=>"110101110",
  25005=>"110001111",
  25006=>"010000101",
  25007=>"101000000",
  25008=>"110011101",
  25009=>"000110001",
  25010=>"010111111",
  25011=>"011000110",
  25012=>"000000101",
  25013=>"000001101",
  25014=>"000111000",
  25015=>"110100001",
  25016=>"010000011",
  25017=>"101100011",
  25018=>"110010110",
  25019=>"001111010",
  25020=>"010110100",
  25021=>"000001011",
  25022=>"000101100",
  25023=>"110011111",
  25024=>"000111111",
  25025=>"100111010",
  25026=>"111100111",
  25027=>"000001100",
  25028=>"100111110",
  25029=>"111111101",
  25030=>"101111110",
  25031=>"000000111",
  25032=>"110101100",
  25033=>"011011110",
  25034=>"110100000",
  25035=>"101000000",
  25036=>"010000100",
  25037=>"100101101",
  25038=>"000001001",
  25039=>"110010100",
  25040=>"101000010",
  25041=>"010001000",
  25042=>"011010010",
  25043=>"000101011",
  25044=>"001001110",
  25045=>"000000001",
  25046=>"001100011",
  25047=>"001001110",
  25048=>"111000111",
  25049=>"111101111",
  25050=>"001001100",
  25051=>"111011000",
  25052=>"101111111",
  25053=>"001011111",
  25054=>"110011111",
  25055=>"111111001",
  25056=>"110001000",
  25057=>"100110100",
  25058=>"011101110",
  25059=>"000000000",
  25060=>"001001101",
  25061=>"001001000",
  25062=>"110100101",
  25063=>"111010101",
  25064=>"111111101",
  25065=>"111100010",
  25066=>"110000010",
  25067=>"101101111",
  25068=>"010101011",
  25069=>"000100011",
  25070=>"001100100",
  25071=>"101100111",
  25072=>"000000000",
  25073=>"100110000",
  25074=>"010100010",
  25075=>"010100001",
  25076=>"110111000",
  25077=>"111010001",
  25078=>"000111010",
  25079=>"110101110",
  25080=>"110101000",
  25081=>"001011101",
  25082=>"110100001",
  25083=>"100011000",
  25084=>"001100001",
  25085=>"101010011",
  25086=>"100000100",
  25087=>"010101100",
  25088=>"110000100",
  25089=>"100100110",
  25090=>"000011101",
  25091=>"000011101",
  25092=>"111111101",
  25093=>"000001010",
  25094=>"010010010",
  25095=>"110100100",
  25096=>"101101110",
  25097=>"001110110",
  25098=>"111001100",
  25099=>"110001101",
  25100=>"001010011",
  25101=>"111110000",
  25102=>"010100000",
  25103=>"100111111",
  25104=>"100001001",
  25105=>"001101111",
  25106=>"111010011",
  25107=>"101001010",
  25108=>"000101001",
  25109=>"110110110",
  25110=>"101111000",
  25111=>"110011010",
  25112=>"000100000",
  25113=>"110110010",
  25114=>"000111100",
  25115=>"010110001",
  25116=>"001111000",
  25117=>"110100100",
  25118=>"100011110",
  25119=>"110101011",
  25120=>"100001000",
  25121=>"101110100",
  25122=>"011000011",
  25123=>"001100100",
  25124=>"111100110",
  25125=>"100111000",
  25126=>"010100011",
  25127=>"110011010",
  25128=>"001010010",
  25129=>"000001101",
  25130=>"111111111",
  25131=>"110010010",
  25132=>"000000101",
  25133=>"110010010",
  25134=>"110011000",
  25135=>"010100100",
  25136=>"001001011",
  25137=>"110111100",
  25138=>"101010111",
  25139=>"110000001",
  25140=>"100110110",
  25141=>"110100110",
  25142=>"010011011",
  25143=>"000111101",
  25144=>"000010011",
  25145=>"110000010",
  25146=>"101111111",
  25147=>"111011101",
  25148=>"100001101",
  25149=>"010010000",
  25150=>"001110011",
  25151=>"100101011",
  25152=>"111111001",
  25153=>"000000101",
  25154=>"001000001",
  25155=>"101000010",
  25156=>"101111010",
  25157=>"110110010",
  25158=>"100010000",
  25159=>"110100111",
  25160=>"100100011",
  25161=>"001101000",
  25162=>"110101100",
  25163=>"011100110",
  25164=>"001110100",
  25165=>"001110011",
  25166=>"001011001",
  25167=>"001001101",
  25168=>"111101111",
  25169=>"101101110",
  25170=>"111101011",
  25171=>"000110110",
  25172=>"101000010",
  25173=>"001001101",
  25174=>"101010110",
  25175=>"111010001",
  25176=>"011100110",
  25177=>"000011001",
  25178=>"001001000",
  25179=>"000000101",
  25180=>"100000100",
  25181=>"000000011",
  25182=>"011000111",
  25183=>"100101001",
  25184=>"000111001",
  25185=>"111010001",
  25186=>"100100100",
  25187=>"101001100",
  25188=>"101111100",
  25189=>"011011001",
  25190=>"100110101",
  25191=>"011111101",
  25192=>"000100001",
  25193=>"011001011",
  25194=>"111011010",
  25195=>"011001001",
  25196=>"010111101",
  25197=>"111000110",
  25198=>"011110000",
  25199=>"001100000",
  25200=>"110101011",
  25201=>"000100100",
  25202=>"010111010",
  25203=>"110110011",
  25204=>"101110010",
  25205=>"101011000",
  25206=>"010010001",
  25207=>"100101100",
  25208=>"011100111",
  25209=>"110000000",
  25210=>"111001110",
  25211=>"100001101",
  25212=>"110100110",
  25213=>"001110000",
  25214=>"010011100",
  25215=>"011011111",
  25216=>"100001101",
  25217=>"101111011",
  25218=>"011011110",
  25219=>"001010110",
  25220=>"111101001",
  25221=>"000110111",
  25222=>"010000000",
  25223=>"000111000",
  25224=>"110011100",
  25225=>"110001110",
  25226=>"010101000",
  25227=>"111101000",
  25228=>"010100010",
  25229=>"111101011",
  25230=>"111011011",
  25231=>"111000000",
  25232=>"111100010",
  25233=>"100110100",
  25234=>"001101100",
  25235=>"110111100",
  25236=>"100010100",
  25237=>"100100101",
  25238=>"111101111",
  25239=>"101010000",
  25240=>"101100001",
  25241=>"110000001",
  25242=>"110010100",
  25243=>"011001101",
  25244=>"001011011",
  25245=>"001001101",
  25246=>"001000101",
  25247=>"001001010",
  25248=>"110101010",
  25249=>"110010010",
  25250=>"110111101",
  25251=>"101001001",
  25252=>"010100111",
  25253=>"001101010",
  25254=>"000011111",
  25255=>"001001100",
  25256=>"101101000",
  25257=>"101110001",
  25258=>"111100111",
  25259=>"111100010",
  25260=>"000010010",
  25261=>"000000001",
  25262=>"010001000",
  25263=>"001000111",
  25264=>"011001011",
  25265=>"111001100",
  25266=>"110111111",
  25267=>"100010000",
  25268=>"010110111",
  25269=>"110111110",
  25270=>"000001110",
  25271=>"100000001",
  25272=>"111001010",
  25273=>"111101110",
  25274=>"100000001",
  25275=>"111111010",
  25276=>"111100001",
  25277=>"000001000",
  25278=>"101000001",
  25279=>"001000000",
  25280=>"100000110",
  25281=>"101100111",
  25282=>"100111010",
  25283=>"000110100",
  25284=>"101100110",
  25285=>"100001010",
  25286=>"000010100",
  25287=>"000011001",
  25288=>"011101011",
  25289=>"111101111",
  25290=>"111111000",
  25291=>"100111010",
  25292=>"111011101",
  25293=>"110000101",
  25294=>"110110101",
  25295=>"000110111",
  25296=>"011000111",
  25297=>"100011100",
  25298=>"110100011",
  25299=>"111101100",
  25300=>"101110110",
  25301=>"000001100",
  25302=>"000011101",
  25303=>"011110000",
  25304=>"101110001",
  25305=>"011000000",
  25306=>"100000000",
  25307=>"001000001",
  25308=>"101000110",
  25309=>"100010011",
  25310=>"000100011",
  25311=>"100111110",
  25312=>"100110111",
  25313=>"101101000",
  25314=>"110100010",
  25315=>"100101111",
  25316=>"101101101",
  25317=>"110111000",
  25318=>"001110100",
  25319=>"110011100",
  25320=>"100110111",
  25321=>"100110111",
  25322=>"100101010",
  25323=>"111110001",
  25324=>"000011111",
  25325=>"100111111",
  25326=>"111010001",
  25327=>"011001011",
  25328=>"100010000",
  25329=>"001011100",
  25330=>"100100101",
  25331=>"000000010",
  25332=>"001011011",
  25333=>"101000110",
  25334=>"011101100",
  25335=>"110111000",
  25336=>"011000001",
  25337=>"001100010",
  25338=>"000000011",
  25339=>"000011000",
  25340=>"101010100",
  25341=>"000001111",
  25342=>"101100001",
  25343=>"110010001",
  25344=>"000000011",
  25345=>"010100101",
  25346=>"111100001",
  25347=>"101010111",
  25348=>"100001110",
  25349=>"001101000",
  25350=>"111111101",
  25351=>"101100101",
  25352=>"100001100",
  25353=>"111001111",
  25354=>"111011000",
  25355=>"001011100",
  25356=>"000001100",
  25357=>"101110001",
  25358=>"000010110",
  25359=>"101111011",
  25360=>"101101111",
  25361=>"101100101",
  25362=>"000000111",
  25363=>"000111110",
  25364=>"100100000",
  25365=>"101000000",
  25366=>"100000100",
  25367=>"100101110",
  25368=>"100011110",
  25369=>"001010011",
  25370=>"101010110",
  25371=>"001011100",
  25372=>"110110100",
  25373=>"010111010",
  25374=>"011010000",
  25375=>"010000100",
  25376=>"100101110",
  25377=>"000111111",
  25378=>"111011000",
  25379=>"010011111",
  25380=>"111001001",
  25381=>"010110110",
  25382=>"001100010",
  25383=>"001111101",
  25384=>"101001101",
  25385=>"101111111",
  25386=>"101100110",
  25387=>"000000001",
  25388=>"101101001",
  25389=>"000000000",
  25390=>"010001001",
  25391=>"100000101",
  25392=>"000000000",
  25393=>"111001111",
  25394=>"001010101",
  25395=>"011111111",
  25396=>"000001101",
  25397=>"010010100",
  25398=>"110110111",
  25399=>"101001000",
  25400=>"110101001",
  25401=>"000101111",
  25402=>"001101101",
  25403=>"100101100",
  25404=>"101110100",
  25405=>"100001000",
  25406=>"111100111",
  25407=>"111011101",
  25408=>"100010001",
  25409=>"100100101",
  25410=>"110010010",
  25411=>"101001101",
  25412=>"100101010",
  25413=>"111100011",
  25414=>"010111101",
  25415=>"110011010",
  25416=>"010011101",
  25417=>"110011110",
  25418=>"001001110",
  25419=>"001001110",
  25420=>"100010101",
  25421=>"111001111",
  25422=>"000110000",
  25423=>"010010101",
  25424=>"010011010",
  25425=>"111011100",
  25426=>"111010011",
  25427=>"011000011",
  25428=>"100101100",
  25429=>"111000011",
  25430=>"011000110",
  25431=>"000000111",
  25432=>"111101010",
  25433=>"001011100",
  25434=>"111011010",
  25435=>"101100100",
  25436=>"100101100",
  25437=>"111100110",
  25438=>"110101101",
  25439=>"000010010",
  25440=>"111110010",
  25441=>"000110011",
  25442=>"110100010",
  25443=>"010111101",
  25444=>"000010110",
  25445=>"000011001",
  25446=>"100110011",
  25447=>"000111011",
  25448=>"110010010",
  25449=>"101100010",
  25450=>"000001110",
  25451=>"011000001",
  25452=>"111011111",
  25453=>"011000110",
  25454=>"000010111",
  25455=>"100000000",
  25456=>"001001011",
  25457=>"011010111",
  25458=>"011100010",
  25459=>"101101010",
  25460=>"110010101",
  25461=>"111100110",
  25462=>"001111000",
  25463=>"111000010",
  25464=>"110110011",
  25465=>"000111000",
  25466=>"001101000",
  25467=>"111001110",
  25468=>"011000000",
  25469=>"000010000",
  25470=>"111111011",
  25471=>"000110101",
  25472=>"000010010",
  25473=>"111010111",
  25474=>"101101000",
  25475=>"010000000",
  25476=>"010000101",
  25477=>"100010000",
  25478=>"011101010",
  25479=>"011100001",
  25480=>"000100010",
  25481=>"001100000",
  25482=>"111000001",
  25483=>"000000001",
  25484=>"011001011",
  25485=>"111010110",
  25486=>"000111011",
  25487=>"110001111",
  25488=>"100011001",
  25489=>"110001100",
  25490=>"000000000",
  25491=>"000010100",
  25492=>"110010111",
  25493=>"001010010",
  25494=>"001101000",
  25495=>"101110011",
  25496=>"110000000",
  25497=>"010010110",
  25498=>"010110111",
  25499=>"111101111",
  25500=>"111010100",
  25501=>"011011010",
  25502=>"100101111",
  25503=>"010000010",
  25504=>"100111111",
  25505=>"100011011",
  25506=>"101011111",
  25507=>"111111111",
  25508=>"010000000",
  25509=>"010010111",
  25510=>"011101011",
  25511=>"011001100",
  25512=>"011110101",
  25513=>"011000100",
  25514=>"100111101",
  25515=>"011001111",
  25516=>"010100011",
  25517=>"001000011",
  25518=>"101111000",
  25519=>"101001100",
  25520=>"011010111",
  25521=>"001101111",
  25522=>"111111100",
  25523=>"101110111",
  25524=>"001101001",
  25525=>"001000110",
  25526=>"110110101",
  25527=>"000010101",
  25528=>"111000100",
  25529=>"000011010",
  25530=>"101001010",
  25531=>"001010101",
  25532=>"011001100",
  25533=>"010111110",
  25534=>"001110010",
  25535=>"000110000",
  25536=>"111000111",
  25537=>"010000010",
  25538=>"001000110",
  25539=>"011110001",
  25540=>"100001110",
  25541=>"110100111",
  25542=>"011010100",
  25543=>"011101011",
  25544=>"000000000",
  25545=>"110011101",
  25546=>"111001100",
  25547=>"101001101",
  25548=>"110001000",
  25549=>"001111011",
  25550=>"011010000",
  25551=>"011011011",
  25552=>"110110000",
  25553=>"011101100",
  25554=>"111010101",
  25555=>"001100001",
  25556=>"010011010",
  25557=>"111000010",
  25558=>"000011101",
  25559=>"110110110",
  25560=>"101101110",
  25561=>"010100001",
  25562=>"010111110",
  25563=>"000000000",
  25564=>"000000000",
  25565=>"110110110",
  25566=>"010110110",
  25567=>"000000101",
  25568=>"110011001",
  25569=>"110101000",
  25570=>"000100011",
  25571=>"110111101",
  25572=>"000000010",
  25573=>"111111101",
  25574=>"000000010",
  25575=>"000001000",
  25576=>"110100001",
  25577=>"001110000",
  25578=>"100111010",
  25579=>"001000110",
  25580=>"100101001",
  25581=>"101110110",
  25582=>"100000110",
  25583=>"100010111",
  25584=>"010100100",
  25585=>"101111010",
  25586=>"101001101",
  25587=>"011010001",
  25588=>"100010111",
  25589=>"111010101",
  25590=>"101011001",
  25591=>"111110111",
  25592=>"101101111",
  25593=>"000111101",
  25594=>"001100011",
  25595=>"010011110",
  25596=>"001000000",
  25597=>"110001101",
  25598=>"011010011",
  25599=>"010110010",
  25600=>"111111000",
  25601=>"111100001",
  25602=>"111111000",
  25603=>"110000100",
  25604=>"000101010",
  25605=>"100101010",
  25606=>"011101100",
  25607=>"000011000",
  25608=>"000001111",
  25609=>"011011000",
  25610=>"010000001",
  25611=>"110111111",
  25612=>"000000111",
  25613=>"100100000",
  25614=>"010001100",
  25615=>"110001110",
  25616=>"011000010",
  25617=>"010100111",
  25618=>"100000100",
  25619=>"100101100",
  25620=>"110110111",
  25621=>"100100100",
  25622=>"100111101",
  25623=>"110101101",
  25624=>"101000100",
  25625=>"110110100",
  25626=>"100110110",
  25627=>"010111100",
  25628=>"110110110",
  25629=>"011011101",
  25630=>"000101101",
  25631=>"110100110",
  25632=>"011001111",
  25633=>"110010100",
  25634=>"110100100",
  25635=>"100000010",
  25636=>"001111100",
  25637=>"010000001",
  25638=>"111010010",
  25639=>"011000010",
  25640=>"010011111",
  25641=>"111101101",
  25642=>"101100111",
  25643=>"101101000",
  25644=>"101101011",
  25645=>"111000011",
  25646=>"100110011",
  25647=>"110110110",
  25648=>"001101110",
  25649=>"111011001",
  25650=>"001011000",
  25651=>"100000100",
  25652=>"111111010",
  25653=>"001110001",
  25654=>"111011111",
  25655=>"111101110",
  25656=>"100000101",
  25657=>"110111010",
  25658=>"000111111",
  25659=>"101001000",
  25660=>"100100110",
  25661=>"000100000",
  25662=>"111010010",
  25663=>"011111100",
  25664=>"111000111",
  25665=>"111110101",
  25666=>"110010000",
  25667=>"100101110",
  25668=>"101111111",
  25669=>"110001011",
  25670=>"011011110",
  25671=>"000101100",
  25672=>"011000011",
  25673=>"110000110",
  25674=>"101111100",
  25675=>"111001111",
  25676=>"110010010",
  25677=>"111101111",
  25678=>"000110111",
  25679=>"110111000",
  25680=>"000011110",
  25681=>"100110101",
  25682=>"111011001",
  25683=>"101000001",
  25684=>"000100110",
  25685=>"110110111",
  25686=>"011011011",
  25687=>"011011000",
  25688=>"000001100",
  25689=>"010000001",
  25690=>"101100100",
  25691=>"101111001",
  25692=>"111111000",
  25693=>"100111110",
  25694=>"001001100",
  25695=>"001001010",
  25696=>"000001101",
  25697=>"110111101",
  25698=>"100010000",
  25699=>"001100011",
  25700=>"101011111",
  25701=>"110111011",
  25702=>"110001100",
  25703=>"101011101",
  25704=>"000101100",
  25705=>"110100000",
  25706=>"101100001",
  25707=>"100100001",
  25708=>"100111011",
  25709=>"000000100",
  25710=>"111111110",
  25711=>"110010010",
  25712=>"110101101",
  25713=>"000101101",
  25714=>"001001000",
  25715=>"110110001",
  25716=>"001001101",
  25717=>"111110111",
  25718=>"010001000",
  25719=>"111101110",
  25720=>"010011001",
  25721=>"000110110",
  25722=>"111100100",
  25723=>"010011000",
  25724=>"111111011",
  25725=>"000110010",
  25726=>"111110110",
  25727=>"010111111",
  25728=>"110111001",
  25729=>"011111100",
  25730=>"010001001",
  25731=>"011100011",
  25732=>"100101011",
  25733=>"011011110",
  25734=>"110111111",
  25735=>"011011010",
  25736=>"001100110",
  25737=>"100111100",
  25738=>"101111010",
  25739=>"010000010",
  25740=>"111101001",
  25741=>"100111100",
  25742=>"011001101",
  25743=>"000100010",
  25744=>"010100000",
  25745=>"101000110",
  25746=>"001110000",
  25747=>"000001100",
  25748=>"000000000",
  25749=>"000100101",
  25750=>"101111000",
  25751=>"100111010",
  25752=>"001011110",
  25753=>"110011000",
  25754=>"011001111",
  25755=>"001101011",
  25756=>"101001100",
  25757=>"011100011",
  25758=>"110101101",
  25759=>"010110001",
  25760=>"110001110",
  25761=>"111001110",
  25762=>"000101011",
  25763=>"100000001",
  25764=>"010110110",
  25765=>"111110000",
  25766=>"000001111",
  25767=>"111001011",
  25768=>"000101001",
  25769=>"100011111",
  25770=>"100001001",
  25771=>"100011011",
  25772=>"010101110",
  25773=>"000011001",
  25774=>"001110000",
  25775=>"001001001",
  25776=>"110001001",
  25777=>"101110110",
  25778=>"110100001",
  25779=>"101101001",
  25780=>"000001010",
  25781=>"000010000",
  25782=>"010011001",
  25783=>"111100101",
  25784=>"110000011",
  25785=>"001001100",
  25786=>"011101111",
  25787=>"101010011",
  25788=>"000101000",
  25789=>"011011111",
  25790=>"001110111",
  25791=>"101000110",
  25792=>"111110011",
  25793=>"110110110",
  25794=>"110000011",
  25795=>"011000011",
  25796=>"011000100",
  25797=>"000101001",
  25798=>"011000110",
  25799=>"111111100",
  25800=>"011101010",
  25801=>"101010010",
  25802=>"111110100",
  25803=>"000110100",
  25804=>"100000011",
  25805=>"111101010",
  25806=>"111101010",
  25807=>"011000000",
  25808=>"011000011",
  25809=>"100110010",
  25810=>"010011100",
  25811=>"000000100",
  25812=>"010011110",
  25813=>"111010100",
  25814=>"100101101",
  25815=>"010111111",
  25816=>"010010111",
  25817=>"100111011",
  25818=>"100111101",
  25819=>"011100101",
  25820=>"100101101",
  25821=>"001001011",
  25822=>"101001111",
  25823=>"000100011",
  25824=>"110101101",
  25825=>"100100111",
  25826=>"100001100",
  25827=>"000101010",
  25828=>"000101001",
  25829=>"110001100",
  25830=>"110110011",
  25831=>"111010010",
  25832=>"011011000",
  25833=>"010010111",
  25834=>"010010110",
  25835=>"000101000",
  25836=>"011001000",
  25837=>"100111011",
  25838=>"110110111",
  25839=>"100000100",
  25840=>"100110000",
  25841=>"000111011",
  25842=>"101001101",
  25843=>"000110110",
  25844=>"100100110",
  25845=>"111100110",
  25846=>"011100011",
  25847=>"111101100",
  25848=>"011110000",
  25849=>"101001101",
  25850=>"100110111",
  25851=>"101111100",
  25852=>"011001011",
  25853=>"101100100",
  25854=>"011111001",
  25855=>"010101010",
  25856=>"110101110",
  25857=>"110110111",
  25858=>"000000000",
  25859=>"011110101",
  25860=>"011000100",
  25861=>"111111000",
  25862=>"111101011",
  25863=>"101110101",
  25864=>"011110111",
  25865=>"101011111",
  25866=>"000101011",
  25867=>"110111010",
  25868=>"000101011",
  25869=>"110101111",
  25870=>"001000011",
  25871=>"011111100",
  25872=>"010010000",
  25873=>"110001001",
  25874=>"111010100",
  25875=>"110101011",
  25876=>"111011000",
  25877=>"011010101",
  25878=>"000110111",
  25879=>"101011000",
  25880=>"000000010",
  25881=>"110100100",
  25882=>"110101011",
  25883=>"111010111",
  25884=>"101111011",
  25885=>"110001011",
  25886=>"100001000",
  25887=>"101011111",
  25888=>"000011010",
  25889=>"100101111",
  25890=>"011101111",
  25891=>"001010011",
  25892=>"001101110",
  25893=>"001101111",
  25894=>"110101100",
  25895=>"010000010",
  25896=>"111011110",
  25897=>"101111101",
  25898=>"010101011",
  25899=>"111110111",
  25900=>"110001010",
  25901=>"111101111",
  25902=>"100101000",
  25903=>"110111001",
  25904=>"110010100",
  25905=>"000110111",
  25906=>"111100110",
  25907=>"111010111",
  25908=>"101101001",
  25909=>"010101110",
  25910=>"111001110",
  25911=>"101110011",
  25912=>"111101011",
  25913=>"001001001",
  25914=>"110110100",
  25915=>"100000000",
  25916=>"111010000",
  25917=>"101111111",
  25918=>"000100100",
  25919=>"111110010",
  25920=>"100010001",
  25921=>"110111101",
  25922=>"010101010",
  25923=>"000000001",
  25924=>"100100011",
  25925=>"100011100",
  25926=>"101110110",
  25927=>"101110000",
  25928=>"000011011",
  25929=>"001010001",
  25930=>"000101000",
  25931=>"000101101",
  25932=>"100010101",
  25933=>"100010100",
  25934=>"111101011",
  25935=>"110111110",
  25936=>"000101001",
  25937=>"101011101",
  25938=>"000001010",
  25939=>"011010110",
  25940=>"011100001",
  25941=>"000111101",
  25942=>"101010110",
  25943=>"010100111",
  25944=>"110110100",
  25945=>"100111101",
  25946=>"000100110",
  25947=>"100011001",
  25948=>"110110010",
  25949=>"100100011",
  25950=>"011111010",
  25951=>"001100110",
  25952=>"011011101",
  25953=>"000110000",
  25954=>"001001011",
  25955=>"101000011",
  25956=>"110011111",
  25957=>"100001011",
  25958=>"000001110",
  25959=>"011001010",
  25960=>"010100011",
  25961=>"011111110",
  25962=>"011000011",
  25963=>"001000100",
  25964=>"000100000",
  25965=>"100111100",
  25966=>"111110101",
  25967=>"011100001",
  25968=>"110100101",
  25969=>"111101100",
  25970=>"100110011",
  25971=>"101110101",
  25972=>"101110111",
  25973=>"001000110",
  25974=>"101010010",
  25975=>"001001111",
  25976=>"010111100",
  25977=>"010010000",
  25978=>"100110110",
  25979=>"100101100",
  25980=>"101101010",
  25981=>"100010111",
  25982=>"100100101",
  25983=>"101100001",
  25984=>"000010001",
  25985=>"110000010",
  25986=>"101001000",
  25987=>"110111001",
  25988=>"010001001",
  25989=>"010101001",
  25990=>"001111110",
  25991=>"101100110",
  25992=>"011100011",
  25993=>"001010000",
  25994=>"110010101",
  25995=>"101100000",
  25996=>"110110100",
  25997=>"110000001",
  25998=>"101101000",
  25999=>"110100111",
  26000=>"000100101",
  26001=>"110110000",
  26002=>"111001000",
  26003=>"010001001",
  26004=>"111010001",
  26005=>"000110100",
  26006=>"100010111",
  26007=>"101110010",
  26008=>"011001111",
  26009=>"111111010",
  26010=>"110011101",
  26011=>"011101111",
  26012=>"000101000",
  26013=>"001111110",
  26014=>"111001101",
  26015=>"011101000",
  26016=>"000101010",
  26017=>"110101010",
  26018=>"111111011",
  26019=>"011110101",
  26020=>"001010011",
  26021=>"000101011",
  26022=>"100100111",
  26023=>"001000110",
  26024=>"001001101",
  26025=>"001101000",
  26026=>"010000101",
  26027=>"001010011",
  26028=>"101101110",
  26029=>"110100100",
  26030=>"000000101",
  26031=>"010111010",
  26032=>"000111100",
  26033=>"100100101",
  26034=>"000110010",
  26035=>"100010011",
  26036=>"011000111",
  26037=>"111110001",
  26038=>"011101111",
  26039=>"100001000",
  26040=>"101110111",
  26041=>"010101010",
  26042=>"110100110",
  26043=>"101111111",
  26044=>"110110100",
  26045=>"100001011",
  26046=>"011001000",
  26047=>"110111000",
  26048=>"101100101",
  26049=>"011010101",
  26050=>"001001010",
  26051=>"010101101",
  26052=>"110101000",
  26053=>"100111111",
  26054=>"000100001",
  26055=>"011011110",
  26056=>"101011010",
  26057=>"101101110",
  26058=>"000100100",
  26059=>"011000100",
  26060=>"111110000",
  26061=>"100000001",
  26062=>"101100011",
  26063=>"110100111",
  26064=>"110010001",
  26065=>"100000100",
  26066=>"110110100",
  26067=>"110110100",
  26068=>"000101001",
  26069=>"010111010",
  26070=>"001101001",
  26071=>"001000100",
  26072=>"001000100",
  26073=>"101111100",
  26074=>"000010101",
  26075=>"011000011",
  26076=>"111011111",
  26077=>"101110011",
  26078=>"011011110",
  26079=>"010111110",
  26080=>"111011011",
  26081=>"010010000",
  26082=>"110000000",
  26083=>"011100111",
  26084=>"010101101",
  26085=>"001101000",
  26086=>"100010011",
  26087=>"111101101",
  26088=>"110000010",
  26089=>"010011110",
  26090=>"111111000",
  26091=>"110101101",
  26092=>"001101010",
  26093=>"100000111",
  26094=>"111111110",
  26095=>"100110000",
  26096=>"100000000",
  26097=>"101001000",
  26098=>"100010000",
  26099=>"011000000",
  26100=>"110011000",
  26101=>"000001010",
  26102=>"011001001",
  26103=>"010010011",
  26104=>"110111010",
  26105=>"001101111",
  26106=>"110001100",
  26107=>"111010110",
  26108=>"101000101",
  26109=>"010000000",
  26110=>"101001111",
  26111=>"000110111",
  26112=>"100111101",
  26113=>"000101101",
  26114=>"000000001",
  26115=>"110111111",
  26116=>"111100100",
  26117=>"000010111",
  26118=>"110111000",
  26119=>"000110111",
  26120=>"111010011",
  26121=>"100010110",
  26122=>"000110000",
  26123=>"100101100",
  26124=>"110111010",
  26125=>"001010111",
  26126=>"000111011",
  26127=>"000101101",
  26128=>"000001011",
  26129=>"011001100",
  26130=>"101110111",
  26131=>"110111000",
  26132=>"100101011",
  26133=>"011000001",
  26134=>"000110101",
  26135=>"100101101",
  26136=>"111110001",
  26137=>"000000110",
  26138=>"111001000",
  26139=>"010011101",
  26140=>"011011011",
  26141=>"010000110",
  26142=>"010000111",
  26143=>"111010111",
  26144=>"001010101",
  26145=>"101111011",
  26146=>"011111101",
  26147=>"110101111",
  26148=>"100100110",
  26149=>"110000101",
  26150=>"111000001",
  26151=>"001010110",
  26152=>"100110100",
  26153=>"100010111",
  26154=>"001000111",
  26155=>"101011011",
  26156=>"110110101",
  26157=>"101001000",
  26158=>"111110111",
  26159=>"101101110",
  26160=>"010000111",
  26161=>"001101111",
  26162=>"011111110",
  26163=>"001000101",
  26164=>"011011110",
  26165=>"100110101",
  26166=>"110001001",
  26167=>"100000000",
  26168=>"011000101",
  26169=>"100100100",
  26170=>"011001011",
  26171=>"100001011",
  26172=>"011001011",
  26173=>"111001100",
  26174=>"010000000",
  26175=>"100110111",
  26176=>"001101101",
  26177=>"101101111",
  26178=>"100001010",
  26179=>"111111010",
  26180=>"100110111",
  26181=>"100100100",
  26182=>"010000101",
  26183=>"100101010",
  26184=>"111010000",
  26185=>"011101100",
  26186=>"000000111",
  26187=>"101111100",
  26188=>"110000100",
  26189=>"110101111",
  26190=>"000100101",
  26191=>"000000100",
  26192=>"100110000",
  26193=>"101011100",
  26194=>"010001110",
  26195=>"111100001",
  26196=>"010111110",
  26197=>"010000101",
  26198=>"100110111",
  26199=>"110101110",
  26200=>"000010100",
  26201=>"000111010",
  26202=>"010000010",
  26203=>"100011101",
  26204=>"111111011",
  26205=>"001010110",
  26206=>"111010110",
  26207=>"000101111",
  26208=>"000001000",
  26209=>"011110011",
  26210=>"101010000",
  26211=>"110101010",
  26212=>"001000101",
  26213=>"011111110",
  26214=>"011111110",
  26215=>"110010101",
  26216=>"111110011",
  26217=>"111010001",
  26218=>"100010001",
  26219=>"110011111",
  26220=>"101111100",
  26221=>"001100101",
  26222=>"110101101",
  26223=>"111111101",
  26224=>"000110101",
  26225=>"101101101",
  26226=>"011011011",
  26227=>"010000000",
  26228=>"110100000",
  26229=>"111101101",
  26230=>"110010010",
  26231=>"000000011",
  26232=>"111011111",
  26233=>"000111000",
  26234=>"000001111",
  26235=>"010110010",
  26236=>"001111101",
  26237=>"101000001",
  26238=>"110110111",
  26239=>"001000101",
  26240=>"010010110",
  26241=>"010111101",
  26242=>"000101001",
  26243=>"000110100",
  26244=>"000000011",
  26245=>"010011101",
  26246=>"110111111",
  26247=>"111001011",
  26248=>"001011001",
  26249=>"000011000",
  26250=>"010000000",
  26251=>"010000100",
  26252=>"110000001",
  26253=>"110101110",
  26254=>"100000010",
  26255=>"101101001",
  26256=>"001001011",
  26257=>"010010101",
  26258=>"100001111",
  26259=>"011100111",
  26260=>"101001110",
  26261=>"001001011",
  26262=>"001101100",
  26263=>"101110010",
  26264=>"101000000",
  26265=>"011011010",
  26266=>"001001010",
  26267=>"010111111",
  26268=>"001010000",
  26269=>"111110110",
  26270=>"101111001",
  26271=>"100101110",
  26272=>"001011100",
  26273=>"110000011",
  26274=>"100011101",
  26275=>"111010101",
  26276=>"001101001",
  26277=>"101100110",
  26278=>"110110110",
  26279=>"110000001",
  26280=>"111100010",
  26281=>"010000111",
  26282=>"100110000",
  26283=>"001000110",
  26284=>"001001011",
  26285=>"101111011",
  26286=>"011010010",
  26287=>"010111101",
  26288=>"000000000",
  26289=>"101101110",
  26290=>"111001110",
  26291=>"011100010",
  26292=>"011010011",
  26293=>"100111100",
  26294=>"010110010",
  26295=>"111101111",
  26296=>"111000001",
  26297=>"010001101",
  26298=>"111101100",
  26299=>"111001001",
  26300=>"010110001",
  26301=>"011000100",
  26302=>"101010010",
  26303=>"110111010",
  26304=>"001101101",
  26305=>"100110100",
  26306=>"011111111",
  26307=>"011101010",
  26308=>"000000000",
  26309=>"101101111",
  26310=>"100110010",
  26311=>"000010111",
  26312=>"011111001",
  26313=>"001101111",
  26314=>"100000011",
  26315=>"111011110",
  26316=>"111110000",
  26317=>"001110000",
  26318=>"000011000",
  26319=>"101110010",
  26320=>"001111011",
  26321=>"111100110",
  26322=>"110100100",
  26323=>"011010011",
  26324=>"111000000",
  26325=>"100111110",
  26326=>"001001011",
  26327=>"011000111",
  26328=>"110010011",
  26329=>"010011111",
  26330=>"100101000",
  26331=>"001010010",
  26332=>"111110000",
  26333=>"100110110",
  26334=>"011001011",
  26335=>"011010001",
  26336=>"100100010",
  26337=>"001100111",
  26338=>"110010001",
  26339=>"101101110",
  26340=>"100100101",
  26341=>"000110001",
  26342=>"010101111",
  26343=>"000000000",
  26344=>"111101011",
  26345=>"001000001",
  26346=>"111000000",
  26347=>"000000010",
  26348=>"011100001",
  26349=>"010100100",
  26350=>"110110000",
  26351=>"110011000",
  26352=>"110110010",
  26353=>"111001001",
  26354=>"111100010",
  26355=>"100000100",
  26356=>"100111110",
  26357=>"001010011",
  26358=>"111111011",
  26359=>"111000101",
  26360=>"110001111",
  26361=>"110101011",
  26362=>"101101010",
  26363=>"001011110",
  26364=>"111000000",
  26365=>"100010111",
  26366=>"110100110",
  26367=>"100110000",
  26368=>"110110110",
  26369=>"011101101",
  26370=>"110010000",
  26371=>"100100011",
  26372=>"010111010",
  26373=>"000101110",
  26374=>"011010010",
  26375=>"110111001",
  26376=>"010011010",
  26377=>"001100001",
  26378=>"111101101",
  26379=>"001010010",
  26380=>"001010101",
  26381=>"110101011",
  26382=>"011000011",
  26383=>"010110001",
  26384=>"110110100",
  26385=>"110011110",
  26386=>"000110000",
  26387=>"110110001",
  26388=>"000111111",
  26389=>"110111011",
  26390=>"000110011",
  26391=>"011110100",
  26392=>"000010001",
  26393=>"111101101",
  26394=>"001000001",
  26395=>"000111101",
  26396=>"010100110",
  26397=>"010001100",
  26398=>"100111111",
  26399=>"101110101",
  26400=>"011001111",
  26401=>"101111111",
  26402=>"011100101",
  26403=>"100100011",
  26404=>"110001111",
  26405=>"110111111",
  26406=>"001101011",
  26407=>"011100000",
  26408=>"010100000",
  26409=>"101001101",
  26410=>"100110000",
  26411=>"010100100",
  26412=>"001101001",
  26413=>"000010100",
  26414=>"111100011",
  26415=>"010110011",
  26416=>"111100011",
  26417=>"100111011",
  26418=>"111000010",
  26419=>"111111011",
  26420=>"010000000",
  26421=>"011001101",
  26422=>"110010100",
  26423=>"010010111",
  26424=>"001010011",
  26425=>"000100000",
  26426=>"011101011",
  26427=>"001001010",
  26428=>"101000101",
  26429=>"011101001",
  26430=>"100110001",
  26431=>"100010011",
  26432=>"001100010",
  26433=>"010011000",
  26434=>"000101100",
  26435=>"111111110",
  26436=>"101011110",
  26437=>"001101110",
  26438=>"001100110",
  26439=>"100100100",
  26440=>"110101111",
  26441=>"011101010",
  26442=>"111001001",
  26443=>"000010010",
  26444=>"100111001",
  26445=>"011000011",
  26446=>"110110111",
  26447=>"100001010",
  26448=>"010111100",
  26449=>"110010001",
  26450=>"010011011",
  26451=>"010010010",
  26452=>"111101100",
  26453=>"110110110",
  26454=>"001101011",
  26455=>"010000110",
  26456=>"010011101",
  26457=>"010001110",
  26458=>"011101010",
  26459=>"000001100",
  26460=>"011010011",
  26461=>"111011001",
  26462=>"010011010",
  26463=>"111111110",
  26464=>"011110000",
  26465=>"101110010",
  26466=>"100010010",
  26467=>"000101101",
  26468=>"001011000",
  26469=>"010001111",
  26470=>"010101111",
  26471=>"010111110",
  26472=>"110101010",
  26473=>"101011000",
  26474=>"110011010",
  26475=>"011000101",
  26476=>"101101100",
  26477=>"101100100",
  26478=>"111111100",
  26479=>"101110010",
  26480=>"011100000",
  26481=>"000010000",
  26482=>"100000010",
  26483=>"000001000",
  26484=>"101111101",
  26485=>"101101000",
  26486=>"101000000",
  26487=>"011001111",
  26488=>"101011011",
  26489=>"000011010",
  26490=>"000101000",
  26491=>"001100011",
  26492=>"010111000",
  26493=>"100110000",
  26494=>"011110111",
  26495=>"110100000",
  26496=>"001111010",
  26497=>"101011000",
  26498=>"111001111",
  26499=>"001101101",
  26500=>"101011100",
  26501=>"000011110",
  26502=>"110110001",
  26503=>"001010110",
  26504=>"010110011",
  26505=>"011010000",
  26506=>"000001011",
  26507=>"000110101",
  26508=>"111111110",
  26509=>"000111000",
  26510=>"110011010",
  26511=>"101011010",
  26512=>"100100100",
  26513=>"100101111",
  26514=>"100100110",
  26515=>"011000101",
  26516=>"100111010",
  26517=>"111010110",
  26518=>"100001110",
  26519=>"000010011",
  26520=>"010011001",
  26521=>"000111101",
  26522=>"100100110",
  26523=>"111101001",
  26524=>"011111001",
  26525=>"101111100",
  26526=>"001001011",
  26527=>"010111110",
  26528=>"111111010",
  26529=>"011010000",
  26530=>"101111001",
  26531=>"100011101",
  26532=>"111001000",
  26533=>"010111110",
  26534=>"011101001",
  26535=>"100011101",
  26536=>"011110110",
  26537=>"111001101",
  26538=>"101111111",
  26539=>"000011101",
  26540=>"101011111",
  26541=>"111110111",
  26542=>"100011101",
  26543=>"111110111",
  26544=>"111001101",
  26545=>"010100000",
  26546=>"010100101",
  26547=>"110100000",
  26548=>"011011011",
  26549=>"101001001",
  26550=>"001001010",
  26551=>"101100100",
  26552=>"010000110",
  26553=>"001111111",
  26554=>"101100110",
  26555=>"011100101",
  26556=>"100011100",
  26557=>"100010010",
  26558=>"110110011",
  26559=>"100100101",
  26560=>"100110111",
  26561=>"001110001",
  26562=>"111011011",
  26563=>"110000001",
  26564=>"101111011",
  26565=>"001001100",
  26566=>"110111110",
  26567=>"001001111",
  26568=>"110101111",
  26569=>"000010011",
  26570=>"010011111",
  26571=>"100001011",
  26572=>"000011111",
  26573=>"110011110",
  26574=>"111110011",
  26575=>"101001100",
  26576=>"011110111",
  26577=>"001100111",
  26578=>"101110000",
  26579=>"001101000",
  26580=>"001001101",
  26581=>"011011110",
  26582=>"101011000",
  26583=>"011001000",
  26584=>"111010010",
  26585=>"111011001",
  26586=>"011010001",
  26587=>"111101011",
  26588=>"110010110",
  26589=>"100001011",
  26590=>"111001001",
  26591=>"111011111",
  26592=>"011001001",
  26593=>"111010001",
  26594=>"111101100",
  26595=>"101010100",
  26596=>"111111110",
  26597=>"110110010",
  26598=>"101010111",
  26599=>"110001000",
  26600=>"111111000",
  26601=>"011011110",
  26602=>"010111010",
  26603=>"100010100",
  26604=>"110100011",
  26605=>"011011110",
  26606=>"111110010",
  26607=>"011001110",
  26608=>"001000100",
  26609=>"011011010",
  26610=>"011010100",
  26611=>"000101101",
  26612=>"110001001",
  26613=>"110111111",
  26614=>"000110110",
  26615=>"100110110",
  26616=>"000100001",
  26617=>"001100110",
  26618=>"011011000",
  26619=>"110111011",
  26620=>"110010110",
  26621=>"010111101",
  26622=>"011101110",
  26623=>"101111111",
  26624=>"101001000",
  26625=>"000110101",
  26626=>"110011010",
  26627=>"101100011",
  26628=>"110001110",
  26629=>"001101011",
  26630=>"111011011",
  26631=>"110110010",
  26632=>"101010100",
  26633=>"000001000",
  26634=>"111111111",
  26635=>"010110001",
  26636=>"111001011",
  26637=>"011110000",
  26638=>"101001010",
  26639=>"001110100",
  26640=>"100011101",
  26641=>"101011100",
  26642=>"001000001",
  26643=>"011001010",
  26644=>"000100110",
  26645=>"000100101",
  26646=>"111101000",
  26647=>"011011000",
  26648=>"111101011",
  26649=>"011011011",
  26650=>"100101100",
  26651=>"011100000",
  26652=>"100011101",
  26653=>"110111110",
  26654=>"100000000",
  26655=>"000100010",
  26656=>"111100111",
  26657=>"001001110",
  26658=>"000011100",
  26659=>"111100000",
  26660=>"001111101",
  26661=>"101001101",
  26662=>"001010100",
  26663=>"111011001",
  26664=>"010010010",
  26665=>"000100110",
  26666=>"000001000",
  26667=>"101011100",
  26668=>"001110100",
  26669=>"001101110",
  26670=>"111111011",
  26671=>"111111110",
  26672=>"111001100",
  26673=>"111100011",
  26674=>"111000110",
  26675=>"000001101",
  26676=>"100101000",
  26677=>"100100001",
  26678=>"100010010",
  26679=>"111111011",
  26680=>"010010000",
  26681=>"101010001",
  26682=>"001101011",
  26683=>"010010000",
  26684=>"111011111",
  26685=>"101111111",
  26686=>"101101010",
  26687=>"100010110",
  26688=>"011000100",
  26689=>"101001011",
  26690=>"111101001",
  26691=>"011000010",
  26692=>"001011011",
  26693=>"111100110",
  26694=>"010000011",
  26695=>"011101011",
  26696=>"000101011",
  26697=>"111100011",
  26698=>"110110011",
  26699=>"000100000",
  26700=>"110111111",
  26701=>"101010000",
  26702=>"111011010",
  26703=>"011011110",
  26704=>"100110000",
  26705=>"101011110",
  26706=>"110000111",
  26707=>"110100110",
  26708=>"010011110",
  26709=>"110000011",
  26710=>"000010110",
  26711=>"000100111",
  26712=>"001110011",
  26713=>"101000101",
  26714=>"000000101",
  26715=>"100001001",
  26716=>"111000111",
  26717=>"100000111",
  26718=>"111101010",
  26719=>"010101101",
  26720=>"111001010",
  26721=>"010011001",
  26722=>"011011010",
  26723=>"001010101",
  26724=>"000000101",
  26725=>"101000000",
  26726=>"111001101",
  26727=>"100111100",
  26728=>"010101110",
  26729=>"011010100",
  26730=>"110010001",
  26731=>"001001100",
  26732=>"111111001",
  26733=>"101011111",
  26734=>"100101110",
  26735=>"011001011",
  26736=>"100010011",
  26737=>"000100001",
  26738=>"111100001",
  26739=>"111111100",
  26740=>"111111110",
  26741=>"010000100",
  26742=>"011101100",
  26743=>"001000110",
  26744=>"110111010",
  26745=>"011010011",
  26746=>"110000110",
  26747=>"001111111",
  26748=>"010101110",
  26749=>"111001110",
  26750=>"000100101",
  26751=>"111001001",
  26752=>"100000011",
  26753=>"001010111",
  26754=>"100100110",
  26755=>"010000110",
  26756=>"010010100",
  26757=>"110111010",
  26758=>"001110001",
  26759=>"000101101",
  26760=>"001101010",
  26761=>"100111000",
  26762=>"111011010",
  26763=>"011101111",
  26764=>"010111010",
  26765=>"110000000",
  26766=>"011000011",
  26767=>"110010011",
  26768=>"111001111",
  26769=>"111111001",
  26770=>"101000010",
  26771=>"101100101",
  26772=>"111010000",
  26773=>"110111000",
  26774=>"110011111",
  26775=>"100100101",
  26776=>"000101111",
  26777=>"010100101",
  26778=>"100001110",
  26779=>"110111100",
  26780=>"001000001",
  26781=>"010000000",
  26782=>"110111001",
  26783=>"101011001",
  26784=>"011000010",
  26785=>"110111111",
  26786=>"010110101",
  26787=>"101010110",
  26788=>"110100011",
  26789=>"010100110",
  26790=>"010101100",
  26791=>"000101100",
  26792=>"000101001",
  26793=>"101001100",
  26794=>"011011000",
  26795=>"000100101",
  26796=>"111101111",
  26797=>"011100010",
  26798=>"000001000",
  26799=>"111010101",
  26800=>"010000010",
  26801=>"111110000",
  26802=>"111101010",
  26803=>"000000000",
  26804=>"011101101",
  26805=>"111011001",
  26806=>"110000000",
  26807=>"010100101",
  26808=>"010110101",
  26809=>"011100011",
  26810=>"000010011",
  26811=>"101111111",
  26812=>"100001000",
  26813=>"101111000",
  26814=>"011010000",
  26815=>"111100111",
  26816=>"001001111",
  26817=>"000111110",
  26818=>"011011010",
  26819=>"111111001",
  26820=>"010100110",
  26821=>"111101011",
  26822=>"011001110",
  26823=>"011001111",
  26824=>"011100101",
  26825=>"000000110",
  26826=>"110110000",
  26827=>"100110100",
  26828=>"110101110",
  26829=>"010111001",
  26830=>"100001011",
  26831=>"001101000",
  26832=>"010011000",
  26833=>"111101101",
  26834=>"001100100",
  26835=>"111011011",
  26836=>"010110001",
  26837=>"000010011",
  26838=>"000001100",
  26839=>"111011100",
  26840=>"111000101",
  26841=>"100100110",
  26842=>"000011001",
  26843=>"111011001",
  26844=>"010111100",
  26845=>"001100010",
  26846=>"010111110",
  26847=>"110010011",
  26848=>"010011011",
  26849=>"011010001",
  26850=>"110100000",
  26851=>"011001001",
  26852=>"010101011",
  26853=>"000000101",
  26854=>"001010011",
  26855=>"010111111",
  26856=>"100110110",
  26857=>"010001010",
  26858=>"000001101",
  26859=>"011001000",
  26860=>"011111000",
  26861=>"010111100",
  26862=>"110100001",
  26863=>"101010000",
  26864=>"111000011",
  26865=>"101001011",
  26866=>"011011101",
  26867=>"000101100",
  26868=>"000101101",
  26869=>"110111111",
  26870=>"101011001",
  26871=>"000001110",
  26872=>"101101001",
  26873=>"000011000",
  26874=>"111111001",
  26875=>"110111011",
  26876=>"001100000",
  26877=>"110011101",
  26878=>"001001000",
  26879=>"111111011",
  26880=>"000011100",
  26881=>"111001110",
  26882=>"010110001",
  26883=>"001111000",
  26884=>"011010110",
  26885=>"101001011",
  26886=>"101000101",
  26887=>"010111000",
  26888=>"001110111",
  26889=>"000001010",
  26890=>"000010000",
  26891=>"010110100",
  26892=>"100010011",
  26893=>"111000101",
  26894=>"011000110",
  26895=>"101001011",
  26896=>"011011111",
  26897=>"100010000",
  26898=>"101100011",
  26899=>"111110101",
  26900=>"011100000",
  26901=>"010001000",
  26902=>"001010110",
  26903=>"000100101",
  26904=>"111010001",
  26905=>"111001010",
  26906=>"000110111",
  26907=>"001100001",
  26908=>"110101011",
  26909=>"110100111",
  26910=>"010011111",
  26911=>"110001100",
  26912=>"001010111",
  26913=>"010110000",
  26914=>"111101000",
  26915=>"100111111",
  26916=>"010101010",
  26917=>"000100010",
  26918=>"110000001",
  26919=>"001101001",
  26920=>"111001111",
  26921=>"000000100",
  26922=>"110101100",
  26923=>"000011100",
  26924=>"100000010",
  26925=>"101101001",
  26926=>"111001001",
  26927=>"001110100",
  26928=>"110101101",
  26929=>"001100100",
  26930=>"110000000",
  26931=>"011111111",
  26932=>"001000100",
  26933=>"001011101",
  26934=>"110100101",
  26935=>"100111000",
  26936=>"100101110",
  26937=>"011100001",
  26938=>"010111000",
  26939=>"011000000",
  26940=>"010001001",
  26941=>"001000100",
  26942=>"100101000",
  26943=>"100000010",
  26944=>"110100011",
  26945=>"101000011",
  26946=>"011011111",
  26947=>"110011011",
  26948=>"110110010",
  26949=>"100111000",
  26950=>"111001000",
  26951=>"011011000",
  26952=>"110001010",
  26953=>"000111010",
  26954=>"001001111",
  26955=>"001101000",
  26956=>"110010000",
  26957=>"110110111",
  26958=>"010110100",
  26959=>"111010011",
  26960=>"110111110",
  26961=>"000110011",
  26962=>"110100011",
  26963=>"111010000",
  26964=>"001110011",
  26965=>"010010111",
  26966=>"100010111",
  26967=>"001010101",
  26968=>"101111011",
  26969=>"100010101",
  26970=>"111100101",
  26971=>"000100110",
  26972=>"101010001",
  26973=>"011011101",
  26974=>"110100100",
  26975=>"010010001",
  26976=>"011001000",
  26977=>"001010010",
  26978=>"010111110",
  26979=>"110001101",
  26980=>"011111011",
  26981=>"011100011",
  26982=>"001001101",
  26983=>"010001011",
  26984=>"000110101",
  26985=>"100111000",
  26986=>"010011111",
  26987=>"001111110",
  26988=>"001000111",
  26989=>"000110010",
  26990=>"100101001",
  26991=>"010011000",
  26992=>"001111111",
  26993=>"110010101",
  26994=>"011111001",
  26995=>"000010001",
  26996=>"100100111",
  26997=>"001101101",
  26998=>"001100101",
  26999=>"010100000",
  27000=>"101010101",
  27001=>"011000110",
  27002=>"011110101",
  27003=>"000110111",
  27004=>"001010110",
  27005=>"010000001",
  27006=>"101101110",
  27007=>"101010011",
  27008=>"011001100",
  27009=>"110100010",
  27010=>"010010100",
  27011=>"100110100",
  27012=>"111110110",
  27013=>"101000001",
  27014=>"011111001",
  27015=>"000010001",
  27016=>"001101001",
  27017=>"001011111",
  27018=>"010010000",
  27019=>"011011110",
  27020=>"000011011",
  27021=>"100101101",
  27022=>"110101100",
  27023=>"100111110",
  27024=>"111010000",
  27025=>"011011011",
  27026=>"111000111",
  27027=>"110000010",
  27028=>"101101100",
  27029=>"000101001",
  27030=>"111011101",
  27031=>"001111011",
  27032=>"100011100",
  27033=>"001011101",
  27034=>"101101001",
  27035=>"000001110",
  27036=>"001111011",
  27037=>"110010101",
  27038=>"101010000",
  27039=>"010110100",
  27040=>"001001001",
  27041=>"000010110",
  27042=>"001101111",
  27043=>"010000001",
  27044=>"100100110",
  27045=>"010010100",
  27046=>"001000000",
  27047=>"101101110",
  27048=>"011011000",
  27049=>"101111011",
  27050=>"001010001",
  27051=>"010011000",
  27052=>"111100101",
  27053=>"011110001",
  27054=>"111111101",
  27055=>"001101110",
  27056=>"000101101",
  27057=>"010001011",
  27058=>"010000010",
  27059=>"111111011",
  27060=>"101110101",
  27061=>"100100100",
  27062=>"000001100",
  27063=>"101011010",
  27064=>"101000110",
  27065=>"101101010",
  27066=>"000100000",
  27067=>"001100100",
  27068=>"111000101",
  27069=>"101100011",
  27070=>"010011111",
  27071=>"110011010",
  27072=>"011000000",
  27073=>"100001111",
  27074=>"011000111",
  27075=>"011110100",
  27076=>"110000001",
  27077=>"000101110",
  27078=>"101100100",
  27079=>"100000000",
  27080=>"010010110",
  27081=>"100110101",
  27082=>"000010111",
  27083=>"010110110",
  27084=>"101010011",
  27085=>"010110011",
  27086=>"001000000",
  27087=>"011010010",
  27088=>"000001011",
  27089=>"000011011",
  27090=>"110100111",
  27091=>"011010011",
  27092=>"011101100",
  27093=>"001010111",
  27094=>"000000101",
  27095=>"011101111",
  27096=>"110000100",
  27097=>"110101101",
  27098=>"110101000",
  27099=>"111011011",
  27100=>"101101011",
  27101=>"000101101",
  27102=>"110101110",
  27103=>"001110110",
  27104=>"000000001",
  27105=>"000010011",
  27106=>"000011011",
  27107=>"110000001",
  27108=>"101111111",
  27109=>"101000111",
  27110=>"110000000",
  27111=>"111000001",
  27112=>"011011101",
  27113=>"110011010",
  27114=>"011100001",
  27115=>"010111111",
  27116=>"001111100",
  27117=>"101001101",
  27118=>"000010001",
  27119=>"001001011",
  27120=>"110100101",
  27121=>"110011100",
  27122=>"111001011",
  27123=>"011101101",
  27124=>"000011001",
  27125=>"111011100",
  27126=>"001000101",
  27127=>"010000000",
  27128=>"010110111",
  27129=>"111111001",
  27130=>"110001000",
  27131=>"111111000",
  27132=>"010111010",
  27133=>"010100111",
  27134=>"111010101",
  27135=>"000010000",
  27136=>"110110111",
  27137=>"010111110",
  27138=>"101110011",
  27139=>"010110101",
  27140=>"011000101",
  27141=>"111010111",
  27142=>"100100001",
  27143=>"001001110",
  27144=>"110100101",
  27145=>"101001010",
  27146=>"001001000",
  27147=>"011010111",
  27148=>"100100000",
  27149=>"000110011",
  27150=>"001001111",
  27151=>"111110100",
  27152=>"001110111",
  27153=>"001111111",
  27154=>"100111100",
  27155=>"101000110",
  27156=>"101010111",
  27157=>"100000011",
  27158=>"010110000",
  27159=>"000011000",
  27160=>"001110100",
  27161=>"011111000",
  27162=>"111011001",
  27163=>"100011101",
  27164=>"001000001",
  27165=>"001000101",
  27166=>"100101101",
  27167=>"100000110",
  27168=>"001100111",
  27169=>"011001000",
  27170=>"110101110",
  27171=>"001010100",
  27172=>"001010111",
  27173=>"101111010",
  27174=>"101111110",
  27175=>"010110101",
  27176=>"001111010",
  27177=>"001000000",
  27178=>"111001110",
  27179=>"111011101",
  27180=>"011111000",
  27181=>"100100100",
  27182=>"000111000",
  27183=>"000000001",
  27184=>"011000011",
  27185=>"001111101",
  27186=>"011000011",
  27187=>"001000111",
  27188=>"000101100",
  27189=>"010000010",
  27190=>"010010101",
  27191=>"010100111",
  27192=>"111101111",
  27193=>"001001011",
  27194=>"100010100",
  27195=>"000110101",
  27196=>"000000111",
  27197=>"000100001",
  27198=>"111011111",
  27199=>"101110100",
  27200=>"000110001",
  27201=>"111100000",
  27202=>"001101111",
  27203=>"101001000",
  27204=>"000001111",
  27205=>"000000100",
  27206=>"011010011",
  27207=>"100001011",
  27208=>"001011000",
  27209=>"110110100",
  27210=>"000100111",
  27211=>"001001101",
  27212=>"111111010",
  27213=>"001000111",
  27214=>"110000111",
  27215=>"110001100",
  27216=>"001110000",
  27217=>"110010100",
  27218=>"011111110",
  27219=>"110011011",
  27220=>"111110010",
  27221=>"000000001",
  27222=>"000000010",
  27223=>"111011100",
  27224=>"000000111",
  27225=>"000000100",
  27226=>"000000000",
  27227=>"101101101",
  27228=>"111001011",
  27229=>"100000011",
  27230=>"101100101",
  27231=>"011010100",
  27232=>"111010100",
  27233=>"010000000",
  27234=>"011010000",
  27235=>"100000011",
  27236=>"010111011",
  27237=>"001110000",
  27238=>"100100011",
  27239=>"000011010",
  27240=>"110010000",
  27241=>"011000111",
  27242=>"100111111",
  27243=>"000100010",
  27244=>"101000010",
  27245=>"100010001",
  27246=>"001110001",
  27247=>"111011111",
  27248=>"011011110",
  27249=>"011001001",
  27250=>"010001110",
  27251=>"000000111",
  27252=>"010000000",
  27253=>"110001000",
  27254=>"011001010",
  27255=>"001111011",
  27256=>"000001000",
  27257=>"001101011",
  27258=>"000111000",
  27259=>"000100110",
  27260=>"001101100",
  27261=>"001011000",
  27262=>"111010000",
  27263=>"110001101",
  27264=>"111000101",
  27265=>"111100111",
  27266=>"011011011",
  27267=>"110010000",
  27268=>"001000111",
  27269=>"010100101",
  27270=>"110100011",
  27271=>"100110110",
  27272=>"011101110",
  27273=>"011110111",
  27274=>"010100100",
  27275=>"100100110",
  27276=>"010011111",
  27277=>"010101000",
  27278=>"101001001",
  27279=>"011000100",
  27280=>"111011111",
  27281=>"011101000",
  27282=>"011011101",
  27283=>"000000101",
  27284=>"010110101",
  27285=>"110100111",
  27286=>"001100000",
  27287=>"000001100",
  27288=>"110100101",
  27289=>"110010001",
  27290=>"000010101",
  27291=>"110110101",
  27292=>"011111111",
  27293=>"010101011",
  27294=>"101011000",
  27295=>"001100011",
  27296=>"111111111",
  27297=>"011000100",
  27298=>"011001010",
  27299=>"110111011",
  27300=>"000011101",
  27301=>"011001111",
  27302=>"011001001",
  27303=>"011111111",
  27304=>"001101111",
  27305=>"001011001",
  27306=>"000000001",
  27307=>"111011110",
  27308=>"110101000",
  27309=>"101010111",
  27310=>"011110000",
  27311=>"110011000",
  27312=>"101011001",
  27313=>"001000100",
  27314=>"000010001",
  27315=>"001001011",
  27316=>"000100001",
  27317=>"001000000",
  27318=>"010100111",
  27319=>"000000010",
  27320=>"101101110",
  27321=>"101101101",
  27322=>"010100001",
  27323=>"101100010",
  27324=>"000110010",
  27325=>"011011011",
  27326=>"000001001",
  27327=>"010111100",
  27328=>"100011100",
  27329=>"010000110",
  27330=>"010101111",
  27331=>"100110110",
  27332=>"110100001",
  27333=>"001000110",
  27334=>"111100001",
  27335=>"101001011",
  27336=>"110010000",
  27337=>"010000011",
  27338=>"101001000",
  27339=>"100101111",
  27340=>"110111010",
  27341=>"000110001",
  27342=>"010101111",
  27343=>"011111010",
  27344=>"010011000",
  27345=>"011100110",
  27346=>"110010110",
  27347=>"101000111",
  27348=>"001100101",
  27349=>"011000111",
  27350=>"001101100",
  27351=>"111110000",
  27352=>"111001011",
  27353=>"111010110",
  27354=>"110100101",
  27355=>"110010100",
  27356=>"000000110",
  27357=>"000100010",
  27358=>"010000111",
  27359=>"110000100",
  27360=>"001110000",
  27361=>"110001100",
  27362=>"111011011",
  27363=>"101110001",
  27364=>"101101111",
  27365=>"001011000",
  27366=>"100001000",
  27367=>"011001010",
  27368=>"111111100",
  27369=>"011001001",
  27370=>"110101001",
  27371=>"001100000",
  27372=>"110001110",
  27373=>"011000001",
  27374=>"011100110",
  27375=>"111100010",
  27376=>"010001010",
  27377=>"101010100",
  27378=>"001011110",
  27379=>"110011001",
  27380=>"000111111",
  27381=>"011011001",
  27382=>"100110101",
  27383=>"111100011",
  27384=>"001100110",
  27385=>"111101101",
  27386=>"100111000",
  27387=>"111101011",
  27388=>"100001110",
  27389=>"101001011",
  27390=>"000001111",
  27391=>"111011000",
  27392=>"000011110",
  27393=>"100101101",
  27394=>"100110011",
  27395=>"010010001",
  27396=>"011101001",
  27397=>"100000111",
  27398=>"111101101",
  27399=>"101111000",
  27400=>"111101111",
  27401=>"101101111",
  27402=>"010110101",
  27403=>"000111011",
  27404=>"110111011",
  27405=>"111110111",
  27406=>"000010110",
  27407=>"011101110",
  27408=>"000011100",
  27409=>"001001001",
  27410=>"100101000",
  27411=>"100000110",
  27412=>"000010111",
  27413=>"110110101",
  27414=>"010110101",
  27415=>"110011100",
  27416=>"101011111",
  27417=>"001011011",
  27418=>"000010110",
  27419=>"011101100",
  27420=>"001101100",
  27421=>"110011101",
  27422=>"000011001",
  27423=>"110000000",
  27424=>"000111011",
  27425=>"111001111",
  27426=>"001011010",
  27427=>"011101011",
  27428=>"101111101",
  27429=>"010100100",
  27430=>"111010100",
  27431=>"101101001",
  27432=>"011001101",
  27433=>"000101001",
  27434=>"010011111",
  27435=>"010110101",
  27436=>"101110110",
  27437=>"110110111",
  27438=>"001111010",
  27439=>"011001010",
  27440=>"010110111",
  27441=>"101111111",
  27442=>"000000001",
  27443=>"001100010",
  27444=>"001101011",
  27445=>"001001101",
  27446=>"001010100",
  27447=>"010110011",
  27448=>"100000010",
  27449=>"000011011",
  27450=>"010111100",
  27451=>"000000101",
  27452=>"000001010",
  27453=>"011100111",
  27454=>"010101101",
  27455=>"011110000",
  27456=>"101111101",
  27457=>"011001011",
  27458=>"110010111",
  27459=>"010000000",
  27460=>"101001011",
  27461=>"111111110",
  27462=>"010111000",
  27463=>"101011101",
  27464=>"101101100",
  27465=>"010111110",
  27466=>"000110000",
  27467=>"011111000",
  27468=>"000110100",
  27469=>"110100100",
  27470=>"010110110",
  27471=>"101011010",
  27472=>"001011110",
  27473=>"100001011",
  27474=>"010111011",
  27475=>"000111000",
  27476=>"010010001",
  27477=>"011101011",
  27478=>"010101010",
  27479=>"100010011",
  27480=>"001011011",
  27481=>"110100010",
  27482=>"100110101",
  27483=>"011111000",
  27484=>"001101001",
  27485=>"101011000",
  27486=>"101110000",
  27487=>"010101100",
  27488=>"110000100",
  27489=>"111000001",
  27490=>"011000110",
  27491=>"111001111",
  27492=>"100101000",
  27493=>"000111101",
  27494=>"001110010",
  27495=>"100110110",
  27496=>"100110011",
  27497=>"101111011",
  27498=>"100010010",
  27499=>"100001111",
  27500=>"110011000",
  27501=>"011111010",
  27502=>"001110000",
  27503=>"100000101",
  27504=>"010111010",
  27505=>"100100101",
  27506=>"101011011",
  27507=>"001110010",
  27508=>"111001001",
  27509=>"011001000",
  27510=>"111100100",
  27511=>"001000001",
  27512=>"001010001",
  27513=>"100110111",
  27514=>"111111001",
  27515=>"100101011",
  27516=>"001011001",
  27517=>"111100100",
  27518=>"011011000",
  27519=>"011100011",
  27520=>"010101000",
  27521=>"110011110",
  27522=>"111111010",
  27523=>"011111111",
  27524=>"110100100",
  27525=>"110101000",
  27526=>"011111001",
  27527=>"101110010",
  27528=>"011101100",
  27529=>"000111101",
  27530=>"111101100",
  27531=>"010011011",
  27532=>"111100010",
  27533=>"001100011",
  27534=>"001100111",
  27535=>"011000000",
  27536=>"000101001",
  27537=>"111010000",
  27538=>"000011010",
  27539=>"010101101",
  27540=>"010010100",
  27541=>"011101111",
  27542=>"111001001",
  27543=>"010100001",
  27544=>"001100010",
  27545=>"011010011",
  27546=>"100100011",
  27547=>"011001000",
  27548=>"110011110",
  27549=>"111010111",
  27550=>"100010011",
  27551=>"011000111",
  27552=>"001001000",
  27553=>"001000001",
  27554=>"011001110",
  27555=>"001010100",
  27556=>"101111000",
  27557=>"111110010",
  27558=>"110100101",
  27559=>"100011011",
  27560=>"001010100",
  27561=>"000111011",
  27562=>"000010010",
  27563=>"100001010",
  27564=>"011001001",
  27565=>"000001010",
  27566=>"100000100",
  27567=>"001111001",
  27568=>"110010111",
  27569=>"101001001",
  27570=>"110111101",
  27571=>"111100101",
  27572=>"110111010",
  27573=>"110110110",
  27574=>"101011111",
  27575=>"101101010",
  27576=>"011001011",
  27577=>"011100100",
  27578=>"001001100",
  27579=>"111110101",
  27580=>"001110111",
  27581=>"101010010",
  27582=>"011001101",
  27583=>"111001011",
  27584=>"101000001",
  27585=>"001100011",
  27586=>"000000101",
  27587=>"000101111",
  27588=>"000100001",
  27589=>"110111011",
  27590=>"011110010",
  27591=>"100100011",
  27592=>"011110010",
  27593=>"110111111",
  27594=>"010101000",
  27595=>"001011000",
  27596=>"000111011",
  27597=>"100110010",
  27598=>"011000111",
  27599=>"110001001",
  27600=>"100101110",
  27601=>"000100001",
  27602=>"100011010",
  27603=>"000110100",
  27604=>"000110101",
  27605=>"011101111",
  27606=>"110100010",
  27607=>"110111010",
  27608=>"111010000",
  27609=>"001101101",
  27610=>"001000001",
  27611=>"010001001",
  27612=>"001110110",
  27613=>"000110010",
  27614=>"001000101",
  27615=>"001010010",
  27616=>"100101010",
  27617=>"110000101",
  27618=>"000110100",
  27619=>"001000100",
  27620=>"011001001",
  27621=>"011101001",
  27622=>"101111101",
  27623=>"111010100",
  27624=>"001111011",
  27625=>"010111010",
  27626=>"000101101",
  27627=>"000001110",
  27628=>"111011100",
  27629=>"001000000",
  27630=>"001001111",
  27631=>"011111100",
  27632=>"110110101",
  27633=>"001011100",
  27634=>"110101010",
  27635=>"111000111",
  27636=>"100101001",
  27637=>"011110100",
  27638=>"010111001",
  27639=>"111010100",
  27640=>"010100011",
  27641=>"000110011",
  27642=>"101111101",
  27643=>"110001011",
  27644=>"001110000",
  27645=>"001100100",
  27646=>"110110111",
  27647=>"111111010",
  27648=>"110000001",
  27649=>"101011111",
  27650=>"010110111",
  27651=>"000010000",
  27652=>"010110110",
  27653=>"101000001",
  27654=>"110010111",
  27655=>"100101000",
  27656=>"010000000",
  27657=>"101111101",
  27658=>"010001000",
  27659=>"000100111",
  27660=>"000110100",
  27661=>"000101001",
  27662=>"010000001",
  27663=>"110001010",
  27664=>"110000001",
  27665=>"110110110",
  27666=>"101100001",
  27667=>"111110010",
  27668=>"111110001",
  27669=>"001100010",
  27670=>"110110110",
  27671=>"011011000",
  27672=>"010101111",
  27673=>"100100000",
  27674=>"001111000",
  27675=>"000101001",
  27676=>"111000000",
  27677=>"111010111",
  27678=>"001001000",
  27679=>"100001000",
  27680=>"011100000",
  27681=>"001011110",
  27682=>"111111100",
  27683=>"101010100",
  27684=>"011011111",
  27685=>"000000111",
  27686=>"111110010",
  27687=>"110011111",
  27688=>"110110100",
  27689=>"000110111",
  27690=>"101011010",
  27691=>"010111001",
  27692=>"010101111",
  27693=>"110010011",
  27694=>"101000011",
  27695=>"001001111",
  27696=>"011100111",
  27697=>"011011111",
  27698=>"101110111",
  27699=>"010111100",
  27700=>"001001101",
  27701=>"000010011",
  27702=>"001100000",
  27703=>"101101100",
  27704=>"010001011",
  27705=>"010000001",
  27706=>"101111010",
  27707=>"010000000",
  27708=>"100010000",
  27709=>"101111101",
  27710=>"010110100",
  27711=>"000001111",
  27712=>"100001111",
  27713=>"100010110",
  27714=>"100001110",
  27715=>"111111100",
  27716=>"001010000",
  27717=>"011010101",
  27718=>"110100101",
  27719=>"011000001",
  27720=>"101101010",
  27721=>"010100001",
  27722=>"101111001",
  27723=>"111001000",
  27724=>"100011110",
  27725=>"001110100",
  27726=>"010000110",
  27727=>"010001011",
  27728=>"001111101",
  27729=>"111111010",
  27730=>"011110001",
  27731=>"110111000",
  27732=>"111010000",
  27733=>"110111110",
  27734=>"110011101",
  27735=>"101000101",
  27736=>"111011011",
  27737=>"110010101",
  27738=>"000111111",
  27739=>"000000111",
  27740=>"010000110",
  27741=>"000011110",
  27742=>"010000101",
  27743=>"110110000",
  27744=>"100100011",
  27745=>"101001001",
  27746=>"110011111",
  27747=>"011010110",
  27748=>"110000100",
  27749=>"110100110",
  27750=>"011111000",
  27751=>"111001000",
  27752=>"000000110",
  27753=>"000010101",
  27754=>"000101000",
  27755=>"011000100",
  27756=>"001100101",
  27757=>"101110101",
  27758=>"100110110",
  27759=>"111011100",
  27760=>"000100000",
  27761=>"011111010",
  27762=>"100101001",
  27763=>"000001111",
  27764=>"000001100",
  27765=>"001110110",
  27766=>"100000101",
  27767=>"010010001",
  27768=>"011100100",
  27769=>"111011001",
  27770=>"110000000",
  27771=>"110000010",
  27772=>"001000000",
  27773=>"010011111",
  27774=>"101100000",
  27775=>"011110000",
  27776=>"010010001",
  27777=>"010001101",
  27778=>"101110110",
  27779=>"101000100",
  27780=>"100011010",
  27781=>"100011010",
  27782=>"101000100",
  27783=>"010001110",
  27784=>"100110101",
  27785=>"001101100",
  27786=>"111100011",
  27787=>"001111100",
  27788=>"101110011",
  27789=>"001111111",
  27790=>"000000101",
  27791=>"010011100",
  27792=>"111011101",
  27793=>"000111100",
  27794=>"100111010",
  27795=>"100000111",
  27796=>"100000000",
  27797=>"000010010",
  27798=>"001001100",
  27799=>"101111001",
  27800=>"111111001",
  27801=>"101101010",
  27802=>"011101001",
  27803=>"001100010",
  27804=>"000110111",
  27805=>"010101110",
  27806=>"010111001",
  27807=>"111100001",
  27808=>"011001111",
  27809=>"000000100",
  27810=>"011000001",
  27811=>"011010101",
  27812=>"010001110",
  27813=>"000010101",
  27814=>"001110010",
  27815=>"110000100",
  27816=>"101000001",
  27817=>"100100101",
  27818=>"111010010",
  27819=>"111011111",
  27820=>"000010011",
  27821=>"101101000",
  27822=>"010111010",
  27823=>"010010011",
  27824=>"110001000",
  27825=>"100110101",
  27826=>"111010010",
  27827=>"111111010",
  27828=>"000001000",
  27829=>"100011100",
  27830=>"011001000",
  27831=>"100011111",
  27832=>"001001111",
  27833=>"011110111",
  27834=>"101000001",
  27835=>"101100010",
  27836=>"001100101",
  27837=>"111101001",
  27838=>"110111001",
  27839=>"010010111",
  27840=>"111111000",
  27841=>"011000110",
  27842=>"000000000",
  27843=>"100101111",
  27844=>"001110011",
  27845=>"010111001",
  27846=>"110101101",
  27847=>"011000111",
  27848=>"011011101",
  27849=>"001010010",
  27850=>"000010110",
  27851=>"010000111",
  27852=>"001010111",
  27853=>"101000001",
  27854=>"001100101",
  27855=>"100010000",
  27856=>"011000101",
  27857=>"110100001",
  27858=>"100111001",
  27859=>"111110101",
  27860=>"110111100",
  27861=>"111111110",
  27862=>"011000100",
  27863=>"010110111",
  27864=>"110011000",
  27865=>"000111110",
  27866=>"100010110",
  27867=>"101001111",
  27868=>"000110101",
  27869=>"111110011",
  27870=>"100001010",
  27871=>"101100101",
  27872=>"101110011",
  27873=>"001100010",
  27874=>"111011010",
  27875=>"000010110",
  27876=>"010001110",
  27877=>"101101101",
  27878=>"000010000",
  27879=>"011101001",
  27880=>"001001001",
  27881=>"111110100",
  27882=>"100100110",
  27883=>"011010100",
  27884=>"000001011",
  27885=>"100100000",
  27886=>"010100110",
  27887=>"110111101",
  27888=>"101110110",
  27889=>"101010111",
  27890=>"000101101",
  27891=>"101111001",
  27892=>"001101100",
  27893=>"011010100",
  27894=>"000110000",
  27895=>"100001101",
  27896=>"000111110",
  27897=>"001111111",
  27898=>"001110001",
  27899=>"010100001",
  27900=>"101000011",
  27901=>"111001010",
  27902=>"001001000",
  27903=>"000101011",
  27904=>"111010110",
  27905=>"100110011",
  27906=>"111110101",
  27907=>"000011100",
  27908=>"111111100",
  27909=>"001111110",
  27910=>"100011011",
  27911=>"001010010",
  27912=>"000000000",
  27913=>"010000110",
  27914=>"001100101",
  27915=>"010011001",
  27916=>"001011100",
  27917=>"010100000",
  27918=>"011010111",
  27919=>"001000000",
  27920=>"110100110",
  27921=>"010000010",
  27922=>"000010011",
  27923=>"111101001",
  27924=>"000000010",
  27925=>"010101110",
  27926=>"111111011",
  27927=>"010110110",
  27928=>"101011100",
  27929=>"001111110",
  27930=>"010011011",
  27931=>"010101110",
  27932=>"011111011",
  27933=>"000100110",
  27934=>"011000001",
  27935=>"111000010",
  27936=>"000100011",
  27937=>"010100001",
  27938=>"111110101",
  27939=>"001101100",
  27940=>"100111100",
  27941=>"010110111",
  27942=>"101101000",
  27943=>"000101110",
  27944=>"110110011",
  27945=>"000100011",
  27946=>"000100010",
  27947=>"111101011",
  27948=>"000101101",
  27949=>"011001110",
  27950=>"111000001",
  27951=>"101001101",
  27952=>"101010000",
  27953=>"010010010",
  27954=>"100001010",
  27955=>"101101010",
  27956=>"111000010",
  27957=>"101110110",
  27958=>"011000000",
  27959=>"010100010",
  27960=>"101000000",
  27961=>"111110001",
  27962=>"101000010",
  27963=>"101010100",
  27964=>"010001101",
  27965=>"111110101",
  27966=>"010001000",
  27967=>"111111010",
  27968=>"000001110",
  27969=>"011110001",
  27970=>"100011110",
  27971=>"001111110",
  27972=>"111010100",
  27973=>"110101111",
  27974=>"100111000",
  27975=>"011010010",
  27976=>"101100011",
  27977=>"000000110",
  27978=>"000100011",
  27979=>"100111110",
  27980=>"101001011",
  27981=>"110101010",
  27982=>"101111011",
  27983=>"000011101",
  27984=>"111001001",
  27985=>"011011001",
  27986=>"011101011",
  27987=>"101110101",
  27988=>"011110100",
  27989=>"100001101",
  27990=>"000101011",
  27991=>"100001101",
  27992=>"011111110",
  27993=>"000010111",
  27994=>"101100100",
  27995=>"001011100",
  27996=>"101110010",
  27997=>"110000111",
  27998=>"110001000",
  27999=>"101110011",
  28000=>"101110110",
  28001=>"010010000",
  28002=>"101011010",
  28003=>"000010110",
  28004=>"110001101",
  28005=>"110000110",
  28006=>"001110111",
  28007=>"001010000",
  28008=>"011010001",
  28009=>"011111100",
  28010=>"101101010",
  28011=>"010100100",
  28012=>"100111110",
  28013=>"001111010",
  28014=>"101011111",
  28015=>"100101000",
  28016=>"111010000",
  28017=>"011000010",
  28018=>"101100101",
  28019=>"001111101",
  28020=>"101101000",
  28021=>"011111110",
  28022=>"100010010",
  28023=>"100010011",
  28024=>"110101111",
  28025=>"100111100",
  28026=>"010000010",
  28027=>"001111010",
  28028=>"010100110",
  28029=>"011100111",
  28030=>"100000010",
  28031=>"000001010",
  28032=>"101010001",
  28033=>"001101001",
  28034=>"101011111",
  28035=>"101100111",
  28036=>"010110111",
  28037=>"001000000",
  28038=>"100111111",
  28039=>"100100000",
  28040=>"110100100",
  28041=>"101000101",
  28042=>"010010101",
  28043=>"101000011",
  28044=>"111000000",
  28045=>"001101011",
  28046=>"000001101",
  28047=>"011000101",
  28048=>"010110011",
  28049=>"010100100",
  28050=>"101010011",
  28051=>"110111111",
  28052=>"000100111",
  28053=>"010110000",
  28054=>"101001011",
  28055=>"110010110",
  28056=>"100110101",
  28057=>"111000000",
  28058=>"110010101",
  28059=>"110010101",
  28060=>"001000000",
  28061=>"001101000",
  28062=>"001001111",
  28063=>"111010000",
  28064=>"000111101",
  28065=>"010010000",
  28066=>"011000010",
  28067=>"000001100",
  28068=>"111010000",
  28069=>"001110001",
  28070=>"001001110",
  28071=>"110101000",
  28072=>"001011101",
  28073=>"001000100",
  28074=>"100111101",
  28075=>"110110000",
  28076=>"000000011",
  28077=>"000000101",
  28078=>"000011001",
  28079=>"101000111",
  28080=>"010010000",
  28081=>"011101010",
  28082=>"100110101",
  28083=>"110101001",
  28084=>"001010101",
  28085=>"110111001",
  28086=>"010100100",
  28087=>"101011110",
  28088=>"011101000",
  28089=>"000001010",
  28090=>"100100000",
  28091=>"010101101",
  28092=>"001000001",
  28093=>"110001000",
  28094=>"110000010",
  28095=>"100011110",
  28096=>"100000100",
  28097=>"101101001",
  28098=>"011001110",
  28099=>"110100011",
  28100=>"001100100",
  28101=>"001000010",
  28102=>"010101001",
  28103=>"100011101",
  28104=>"100010011",
  28105=>"001110100",
  28106=>"110011110",
  28107=>"110110101",
  28108=>"101111011",
  28109=>"101110000",
  28110=>"100111101",
  28111=>"111110011",
  28112=>"010111101",
  28113=>"101001010",
  28114=>"001101101",
  28115=>"100110101",
  28116=>"000101100",
  28117=>"101010000",
  28118=>"000101011",
  28119=>"000010110",
  28120=>"011000001",
  28121=>"000101001",
  28122=>"111110100",
  28123=>"000101011",
  28124=>"010001000",
  28125=>"000101111",
  28126=>"110010001",
  28127=>"110100111",
  28128=>"011011111",
  28129=>"101100001",
  28130=>"110001100",
  28131=>"000100001",
  28132=>"001011110",
  28133=>"000111100",
  28134=>"111011110",
  28135=>"101111010",
  28136=>"011011110",
  28137=>"101010010",
  28138=>"001101010",
  28139=>"100010100",
  28140=>"111010001",
  28141=>"100101101",
  28142=>"001001010",
  28143=>"111101000",
  28144=>"011000101",
  28145=>"101110011",
  28146=>"001111111",
  28147=>"011100011",
  28148=>"110000110",
  28149=>"111010001",
  28150=>"100001100",
  28151=>"011000101",
  28152=>"000000000",
  28153=>"111001100",
  28154=>"101110101",
  28155=>"011101010",
  28156=>"110101111",
  28157=>"000110010",
  28158=>"100000100",
  28159=>"100100010",
  28160=>"000110000",
  28161=>"111101100",
  28162=>"000000100",
  28163=>"100010010",
  28164=>"111100010",
  28165=>"001001110",
  28166=>"110101111",
  28167=>"000011100",
  28168=>"011000001",
  28169=>"000000111",
  28170=>"110000010",
  28171=>"001000011",
  28172=>"010100100",
  28173=>"100010111",
  28174=>"000010100",
  28175=>"011011011",
  28176=>"100110001",
  28177=>"101000010",
  28178=>"101110110",
  28179=>"011010100",
  28180=>"110101111",
  28181=>"010010000",
  28182=>"001001010",
  28183=>"110101000",
  28184=>"111110100",
  28185=>"001111100",
  28186=>"111100011",
  28187=>"101001001",
  28188=>"111100001",
  28189=>"011000000",
  28190=>"000001101",
  28191=>"111101100",
  28192=>"110111001",
  28193=>"101010010",
  28194=>"101000001",
  28195=>"111111111",
  28196=>"111111110",
  28197=>"101110000",
  28198=>"011101100",
  28199=>"100010101",
  28200=>"111101101",
  28201=>"010101101",
  28202=>"100010011",
  28203=>"110110001",
  28204=>"001011011",
  28205=>"000000001",
  28206=>"011111000",
  28207=>"011101101",
  28208=>"110010111",
  28209=>"100101000",
  28210=>"101111011",
  28211=>"010100111",
  28212=>"001001010",
  28213=>"110011000",
  28214=>"111111001",
  28215=>"001010110",
  28216=>"111101011",
  28217=>"110011010",
  28218=>"111101001",
  28219=>"001000011",
  28220=>"001101100",
  28221=>"000001111",
  28222=>"110000000",
  28223=>"010010011",
  28224=>"101011000",
  28225=>"011110110",
  28226=>"011001110",
  28227=>"010001011",
  28228=>"011011110",
  28229=>"011111101",
  28230=>"011111110",
  28231=>"011110110",
  28232=>"111111110",
  28233=>"011001111",
  28234=>"001011010",
  28235=>"000101000",
  28236=>"110000110",
  28237=>"001110100",
  28238=>"011000110",
  28239=>"001101001",
  28240=>"010001111",
  28241=>"010011001",
  28242=>"001011101",
  28243=>"000000010",
  28244=>"110110101",
  28245=>"000000011",
  28246=>"110111011",
  28247=>"000101111",
  28248=>"101111000",
  28249=>"101101001",
  28250=>"000101111",
  28251=>"011000101",
  28252=>"000110111",
  28253=>"001100001",
  28254=>"010100010",
  28255=>"111111111",
  28256=>"000110101",
  28257=>"011101010",
  28258=>"100111001",
  28259=>"000001101",
  28260=>"001101101",
  28261=>"111010010",
  28262=>"101011111",
  28263=>"000100101",
  28264=>"011000000",
  28265=>"001101000",
  28266=>"011000010",
  28267=>"100010000",
  28268=>"001010110",
  28269=>"101001111",
  28270=>"110010110",
  28271=>"100011111",
  28272=>"010100001",
  28273=>"100000111",
  28274=>"001001100",
  28275=>"001101010",
  28276=>"101100111",
  28277=>"100011001",
  28278=>"110100100",
  28279=>"110101101",
  28280=>"011110000",
  28281=>"001001000",
  28282=>"010111010",
  28283=>"100100100",
  28284=>"001010010",
  28285=>"111101000",
  28286=>"001000010",
  28287=>"101010111",
  28288=>"001101111",
  28289=>"100100010",
  28290=>"010111110",
  28291=>"100100100",
  28292=>"000001001",
  28293=>"100100010",
  28294=>"111010001",
  28295=>"101001110",
  28296=>"001110110",
  28297=>"010011000",
  28298=>"001001010",
  28299=>"100110010",
  28300=>"001001111",
  28301=>"011100101",
  28302=>"100000010",
  28303=>"111101001",
  28304=>"011100100",
  28305=>"111110110",
  28306=>"110101011",
  28307=>"111111011",
  28308=>"001101110",
  28309=>"110111110",
  28310=>"100100011",
  28311=>"010101101",
  28312=>"111001001",
  28313=>"100001011",
  28314=>"111101001",
  28315=>"100011110",
  28316=>"001000100",
  28317=>"100101000",
  28318=>"100110110",
  28319=>"110000100",
  28320=>"100011000",
  28321=>"010000001",
  28322=>"111110110",
  28323=>"110010010",
  28324=>"011010010",
  28325=>"101101011",
  28326=>"111010011",
  28327=>"100100011",
  28328=>"101010100",
  28329=>"011011101",
  28330=>"010011101",
  28331=>"111001010",
  28332=>"001001011",
  28333=>"010111000",
  28334=>"111110000",
  28335=>"011110100",
  28336=>"001000000",
  28337=>"000000111",
  28338=>"000000010",
  28339=>"101100100",
  28340=>"011111000",
  28341=>"001010000",
  28342=>"110001101",
  28343=>"010110001",
  28344=>"010011100",
  28345=>"011100101",
  28346=>"111110010",
  28347=>"011010010",
  28348=>"011011010",
  28349=>"000001101",
  28350=>"000100000",
  28351=>"001111001",
  28352=>"000010011",
  28353=>"111001110",
  28354=>"000011000",
  28355=>"111001011",
  28356=>"110100111",
  28357=>"110110101",
  28358=>"101010101",
  28359=>"010010100",
  28360=>"010001111",
  28361=>"011001101",
  28362=>"010101101",
  28363=>"101001010",
  28364=>"010001100",
  28365=>"110100111",
  28366=>"101010100",
  28367=>"101111111",
  28368=>"111111111",
  28369=>"000101101",
  28370=>"101111111",
  28371=>"000000010",
  28372=>"111110011",
  28373=>"100000010",
  28374=>"110101001",
  28375=>"101001101",
  28376=>"000001011",
  28377=>"111011001",
  28378=>"000001101",
  28379=>"100010110",
  28380=>"000001010",
  28381=>"111110101",
  28382=>"001010001",
  28383=>"111000010",
  28384=>"111000100",
  28385=>"000100010",
  28386=>"110111110",
  28387=>"111011110",
  28388=>"011111000",
  28389=>"111111000",
  28390=>"111000110",
  28391=>"000101011",
  28392=>"000110011",
  28393=>"010111010",
  28394=>"110001011",
  28395=>"001011000",
  28396=>"001011000",
  28397=>"010011011",
  28398=>"001101001",
  28399=>"111100101",
  28400=>"110011010",
  28401=>"000000111",
  28402=>"101011111",
  28403=>"111101100",
  28404=>"000110101",
  28405=>"001111001",
  28406=>"010110101",
  28407=>"001001001",
  28408=>"101100010",
  28409=>"000101011",
  28410=>"101001110",
  28411=>"100010001",
  28412=>"000001001",
  28413=>"001100001",
  28414=>"010010110",
  28415=>"001111010",
  28416=>"101110100",
  28417=>"110000111",
  28418=>"011011010",
  28419=>"000001100",
  28420=>"001001010",
  28421=>"101100111",
  28422=>"010111001",
  28423=>"101101101",
  28424=>"010101101",
  28425=>"100010110",
  28426=>"110010000",
  28427=>"110100110",
  28428=>"101001111",
  28429=>"001011001",
  28430=>"011111001",
  28431=>"010100011",
  28432=>"010011111",
  28433=>"000101000",
  28434=>"100000111",
  28435=>"001000001",
  28436=>"011101110",
  28437=>"100100001",
  28438=>"111011000",
  28439=>"010110011",
  28440=>"010001101",
  28441=>"000100110",
  28442=>"010101011",
  28443=>"111010101",
  28444=>"010010111",
  28445=>"101100011",
  28446=>"100010010",
  28447=>"111101000",
  28448=>"000101001",
  28449=>"101111000",
  28450=>"100001010",
  28451=>"010011011",
  28452=>"101101011",
  28453=>"101000000",
  28454=>"001111111",
  28455=>"000011111",
  28456=>"011000000",
  28457=>"011111001",
  28458=>"000001011",
  28459=>"110111100",
  28460=>"101010110",
  28461=>"101001010",
  28462=>"110010100",
  28463=>"101100000",
  28464=>"101011101",
  28465=>"101110001",
  28466=>"110100000",
  28467=>"111111111",
  28468=>"001001001",
  28469=>"100010101",
  28470=>"011011100",
  28471=>"011100111",
  28472=>"011001010",
  28473=>"101001010",
  28474=>"011001101",
  28475=>"110000100",
  28476=>"011010000",
  28477=>"110111000",
  28478=>"110101010",
  28479=>"011101110",
  28480=>"110001101",
  28481=>"111110111",
  28482=>"111100010",
  28483=>"110000111",
  28484=>"000100101",
  28485=>"110110011",
  28486=>"101000100",
  28487=>"111111110",
  28488=>"100100011",
  28489=>"000010111",
  28490=>"101110110",
  28491=>"001100010",
  28492=>"010000101",
  28493=>"000111011",
  28494=>"100111101",
  28495=>"111010001",
  28496=>"010000111",
  28497=>"001011011",
  28498=>"100101001",
  28499=>"010111011",
  28500=>"001010011",
  28501=>"000101010",
  28502=>"001101101",
  28503=>"101100110",
  28504=>"110000110",
  28505=>"100101001",
  28506=>"011011101",
  28507=>"000110100",
  28508=>"110010010",
  28509=>"110000000",
  28510=>"100000110",
  28511=>"100000001",
  28512=>"101110001",
  28513=>"101101000",
  28514=>"101100000",
  28515=>"010001100",
  28516=>"011101001",
  28517=>"010101001",
  28518=>"100000111",
  28519=>"001101010",
  28520=>"000111000",
  28521=>"101111000",
  28522=>"011101100",
  28523=>"011010110",
  28524=>"101101010",
  28525=>"001000001",
  28526=>"000001011",
  28527=>"000110000",
  28528=>"111111100",
  28529=>"001111000",
  28530=>"011100011",
  28531=>"011000000",
  28532=>"010011111",
  28533=>"110011011",
  28534=>"011000000",
  28535=>"111110000",
  28536=>"001111001",
  28537=>"100111011",
  28538=>"110001011",
  28539=>"111111111",
  28540=>"011010001",
  28541=>"000011000",
  28542=>"000110010",
  28543=>"000111111",
  28544=>"110110110",
  28545=>"100001010",
  28546=>"000100001",
  28547=>"010010111",
  28548=>"101001111",
  28549=>"010100100",
  28550=>"101111111",
  28551=>"100100001",
  28552=>"010111001",
  28553=>"000011100",
  28554=>"001000011",
  28555=>"100000111",
  28556=>"000010110",
  28557=>"101110110",
  28558=>"010100011",
  28559=>"011001010",
  28560=>"101101111",
  28561=>"110010011",
  28562=>"110000010",
  28563=>"101100100",
  28564=>"010001010",
  28565=>"111001110",
  28566=>"110111101",
  28567=>"101011010",
  28568=>"001110101",
  28569=>"011110110",
  28570=>"101111000",
  28571=>"100100010",
  28572=>"100100011",
  28573=>"111101111",
  28574=>"001110010",
  28575=>"000110001",
  28576=>"010000100",
  28577=>"000100000",
  28578=>"101011011",
  28579=>"100101010",
  28580=>"010010110",
  28581=>"101010110",
  28582=>"100000101",
  28583=>"101010011",
  28584=>"001101011",
  28585=>"110101110",
  28586=>"010101100",
  28587=>"100111000",
  28588=>"010101000",
  28589=>"000101101",
  28590=>"010100101",
  28591=>"100011000",
  28592=>"010000001",
  28593=>"001111101",
  28594=>"011010011",
  28595=>"100001011",
  28596=>"110010110",
  28597=>"010110101",
  28598=>"101101100",
  28599=>"101100100",
  28600=>"100101101",
  28601=>"110010011",
  28602=>"001000110",
  28603=>"011111011",
  28604=>"001011000",
  28605=>"011110100",
  28606=>"000000100",
  28607=>"000010010",
  28608=>"111000000",
  28609=>"010110001",
  28610=>"100011000",
  28611=>"001001101",
  28612=>"000011111",
  28613=>"111000111",
  28614=>"011000010",
  28615=>"100111111",
  28616=>"000000011",
  28617=>"000011011",
  28618=>"000101001",
  28619=>"111110010",
  28620=>"100011110",
  28621=>"000000101",
  28622=>"101001010",
  28623=>"010101110",
  28624=>"100010001",
  28625=>"101000000",
  28626=>"110011010",
  28627=>"111000011",
  28628=>"010010000",
  28629=>"111101011",
  28630=>"101000000",
  28631=>"001000010",
  28632=>"110001100",
  28633=>"100001111",
  28634=>"110001011",
  28635=>"101110011",
  28636=>"010100011",
  28637=>"110110110",
  28638=>"100110011",
  28639=>"010000010",
  28640=>"110010101",
  28641=>"101011001",
  28642=>"000010100",
  28643=>"000000111",
  28644=>"101100001",
  28645=>"010101011",
  28646=>"011010101",
  28647=>"101001011",
  28648=>"000001100",
  28649=>"101001011",
  28650=>"101010100",
  28651=>"100010101",
  28652=>"011101110",
  28653=>"001110100",
  28654=>"110001010",
  28655=>"100010100",
  28656=>"110111110",
  28657=>"100100000",
  28658=>"000101010",
  28659=>"000100111",
  28660=>"011001100",
  28661=>"000010110",
  28662=>"111110000",
  28663=>"001000111",
  28664=>"111111001",
  28665=>"000011001",
  28666=>"000010010",
  28667=>"110001111",
  28668=>"101001110",
  28669=>"000101111",
  28670=>"010101101",
  28671=>"001111101",
  28672=>"111111010",
  28673=>"111111110",
  28674=>"000011111",
  28675=>"111111100",
  28676=>"000100011",
  28677=>"110101111",
  28678=>"001101010",
  28679=>"101001110",
  28680=>"011011111",
  28681=>"100111101",
  28682=>"011111010",
  28683=>"000011010",
  28684=>"101000000",
  28685=>"011101010",
  28686=>"000101111",
  28687=>"011110011",
  28688=>"001111111",
  28689=>"011101010",
  28690=>"100111001",
  28691=>"101010101",
  28692=>"001011011",
  28693=>"001110111",
  28694=>"100110010",
  28695=>"000000000",
  28696=>"110000100",
  28697=>"101110101",
  28698=>"111111001",
  28699=>"110001100",
  28700=>"001001001",
  28701=>"011000010",
  28702=>"110111100",
  28703=>"100001100",
  28704=>"011111011",
  28705=>"011011001",
  28706=>"001011110",
  28707=>"100110001",
  28708=>"111011111",
  28709=>"011100101",
  28710=>"101110011",
  28711=>"111110010",
  28712=>"111001000",
  28713=>"010001100",
  28714=>"110000011",
  28715=>"110100111",
  28716=>"101101010",
  28717=>"000001011",
  28718=>"010111101",
  28719=>"110001001",
  28720=>"101011110",
  28721=>"011001100",
  28722=>"010100111",
  28723=>"101111010",
  28724=>"100001010",
  28725=>"110011011",
  28726=>"101001001",
  28727=>"011111100",
  28728=>"001100100",
  28729=>"011000000",
  28730=>"100001111",
  28731=>"111101111",
  28732=>"001001001",
  28733=>"100101011",
  28734=>"101000011",
  28735=>"111010010",
  28736=>"001111101",
  28737=>"100001011",
  28738=>"101110001",
  28739=>"101110100",
  28740=>"010111001",
  28741=>"011011101",
  28742=>"000110001",
  28743=>"000001100",
  28744=>"011010100",
  28745=>"111100111",
  28746=>"111111100",
  28747=>"111000110",
  28748=>"111101001",
  28749=>"011010111",
  28750=>"110000101",
  28751=>"000111000",
  28752=>"100010111",
  28753=>"100101100",
  28754=>"100000011",
  28755=>"110010011",
  28756=>"000000110",
  28757=>"000101101",
  28758=>"001101110",
  28759=>"111101011",
  28760=>"111111011",
  28761=>"010001101",
  28762=>"110110100",
  28763=>"100110101",
  28764=>"100111101",
  28765=>"000001001",
  28766=>"011100110",
  28767=>"010110000",
  28768=>"000100101",
  28769=>"111011011",
  28770=>"101110000",
  28771=>"000001001",
  28772=>"110011001",
  28773=>"110011010",
  28774=>"011101010",
  28775=>"101100010",
  28776=>"010010101",
  28777=>"011111101",
  28778=>"000011000",
  28779=>"111110010",
  28780=>"001011010",
  28781=>"101000001",
  28782=>"010011100",
  28783=>"110100111",
  28784=>"110001110",
  28785=>"110110100",
  28786=>"011101111",
  28787=>"001011101",
  28788=>"011011011",
  28789=>"101011111",
  28790=>"001100100",
  28791=>"111000100",
  28792=>"001111010",
  28793=>"010010111",
  28794=>"111001101",
  28795=>"100110001",
  28796=>"101000010",
  28797=>"010111111",
  28798=>"110110101",
  28799=>"011110001",
  28800=>"111011010",
  28801=>"101001111",
  28802=>"101100001",
  28803=>"111010010",
  28804=>"110110100",
  28805=>"011100101",
  28806=>"010010001",
  28807=>"101110110",
  28808=>"000011010",
  28809=>"110010101",
  28810=>"101010011",
  28811=>"011011001",
  28812=>"011000110",
  28813=>"100110100",
  28814=>"101110000",
  28815=>"010010100",
  28816=>"011110111",
  28817=>"000100011",
  28818=>"001000100",
  28819=>"000100111",
  28820=>"111111110",
  28821=>"101100110",
  28822=>"001111011",
  28823=>"001101001",
  28824=>"011011010",
  28825=>"001111000",
  28826=>"101010011",
  28827=>"011010110",
  28828=>"111010100",
  28829=>"100111100",
  28830=>"011110011",
  28831=>"010000001",
  28832=>"001011110",
  28833=>"101000101",
  28834=>"110111100",
  28835=>"001101110",
  28836=>"011010101",
  28837=>"101001110",
  28838=>"110011110",
  28839=>"111001000",
  28840=>"001110101",
  28841=>"000000100",
  28842=>"001010001",
  28843=>"100010000",
  28844=>"001100110",
  28845=>"100110100",
  28846=>"100001011",
  28847=>"110010110",
  28848=>"001011000",
  28849=>"111001111",
  28850=>"101110100",
  28851=>"101000101",
  28852=>"111011101",
  28853=>"001101111",
  28854=>"111101111",
  28855=>"110100011",
  28856=>"100100000",
  28857=>"110000101",
  28858=>"111110111",
  28859=>"110111101",
  28860=>"001010101",
  28861=>"000110111",
  28862=>"111100101",
  28863=>"011100001",
  28864=>"000000100",
  28865=>"011000000",
  28866=>"111101111",
  28867=>"110110010",
  28868=>"011010111",
  28869=>"001101011",
  28870=>"111010111",
  28871=>"101000111",
  28872=>"100111101",
  28873=>"001010101",
  28874=>"010010110",
  28875=>"100101100",
  28876=>"010000110",
  28877=>"100101110",
  28878=>"000111111",
  28879=>"001011011",
  28880=>"100100111",
  28881=>"110011001",
  28882=>"100000011",
  28883=>"111111101",
  28884=>"101110110",
  28885=>"111011011",
  28886=>"101111100",
  28887=>"100001010",
  28888=>"110101010",
  28889=>"110100010",
  28890=>"010001111",
  28891=>"011100101",
  28892=>"110110011",
  28893=>"101001000",
  28894=>"001100110",
  28895=>"000111010",
  28896=>"111111010",
  28897=>"101100101",
  28898=>"011010010",
  28899=>"011101110",
  28900=>"100100110",
  28901=>"010110100",
  28902=>"011001110",
  28903=>"100000010",
  28904=>"010101001",
  28905=>"000011010",
  28906=>"111011001",
  28907=>"111100010",
  28908=>"011100110",
  28909=>"110111111",
  28910=>"000101001",
  28911=>"101000000",
  28912=>"001111110",
  28913=>"101111101",
  28914=>"010011111",
  28915=>"101111101",
  28916=>"000011001",
  28917=>"011010000",
  28918=>"000110001",
  28919=>"010111000",
  28920=>"001000111",
  28921=>"010010011",
  28922=>"000001101",
  28923=>"000001110",
  28924=>"101001000",
  28925=>"111101111",
  28926=>"111100111",
  28927=>"001100111",
  28928=>"010000000",
  28929=>"111101111",
  28930=>"011101111",
  28931=>"111101001",
  28932=>"011111110",
  28933=>"001001101",
  28934=>"001100011",
  28935=>"111101111",
  28936=>"001010001",
  28937=>"101000100",
  28938=>"011111101",
  28939=>"000110101",
  28940=>"010100111",
  28941=>"111101110",
  28942=>"010111110",
  28943=>"101111100",
  28944=>"010111100",
  28945=>"000001101",
  28946=>"010000011",
  28947=>"111111100",
  28948=>"101001010",
  28949=>"101110001",
  28950=>"001110110",
  28951=>"111001110",
  28952=>"110011111",
  28953=>"011001101",
  28954=>"010010111",
  28955=>"110001000",
  28956=>"011011011",
  28957=>"111111100",
  28958=>"110010011",
  28959=>"101100111",
  28960=>"111010000",
  28961=>"000100011",
  28962=>"001110010",
  28963=>"010000011",
  28964=>"000110100",
  28965=>"101000010",
  28966=>"001111010",
  28967=>"001110101",
  28968=>"011001010",
  28969=>"000110111",
  28970=>"011011010",
  28971=>"010111100",
  28972=>"110111100",
  28973=>"111110000",
  28974=>"000010010",
  28975=>"001111101",
  28976=>"110100100",
  28977=>"000111010",
  28978=>"001100001",
  28979=>"011101010",
  28980=>"100111100",
  28981=>"110101110",
  28982=>"110100100",
  28983=>"000011000",
  28984=>"100011010",
  28985=>"111101011",
  28986=>"001110100",
  28987=>"000011001",
  28988=>"011001001",
  28989=>"101110101",
  28990=>"101111011",
  28991=>"011100101",
  28992=>"000001100",
  28993=>"100110110",
  28994=>"101001011",
  28995=>"110101100",
  28996=>"111111111",
  28997=>"100111101",
  28998=>"001000101",
  28999=>"011001101",
  29000=>"010100001",
  29001=>"110101111",
  29002=>"101011000",
  29003=>"101110000",
  29004=>"111011111",
  29005=>"011001011",
  29006=>"111001010",
  29007=>"100001011",
  29008=>"101110011",
  29009=>"111010111",
  29010=>"111010000",
  29011=>"011000111",
  29012=>"101011100",
  29013=>"101100001",
  29014=>"000110011",
  29015=>"111001000",
  29016=>"010100011",
  29017=>"001000000",
  29018=>"001101101",
  29019=>"000011110",
  29020=>"010101010",
  29021=>"110101110",
  29022=>"000001011",
  29023=>"000001101",
  29024=>"010000010",
  29025=>"010010111",
  29026=>"000011000",
  29027=>"010111010",
  29028=>"001000010",
  29029=>"000000010",
  29030=>"100000100",
  29031=>"101100110",
  29032=>"111001000",
  29033=>"100110010",
  29034=>"010000011",
  29035=>"001000011",
  29036=>"010000010",
  29037=>"010101101",
  29038=>"001010001",
  29039=>"100110011",
  29040=>"000010100",
  29041=>"000000010",
  29042=>"001000111",
  29043=>"111001110",
  29044=>"000100101",
  29045=>"100111111",
  29046=>"000000100",
  29047=>"100001001",
  29048=>"001011110",
  29049=>"010101011",
  29050=>"111111110",
  29051=>"110011001",
  29052=>"000101000",
  29053=>"111101011",
  29054=>"110001111",
  29055=>"100010000",
  29056=>"111100010",
  29057=>"110011010",
  29058=>"010000011",
  29059=>"001100000",
  29060=>"000100011",
  29061=>"100000011",
  29062=>"010000111",
  29063=>"000011000",
  29064=>"001001100",
  29065=>"000110010",
  29066=>"010001111",
  29067=>"000001111",
  29068=>"110101101",
  29069=>"101111001",
  29070=>"100110101",
  29071=>"101011111",
  29072=>"011110011",
  29073=>"101111111",
  29074=>"111001011",
  29075=>"100010011",
  29076=>"001111001",
  29077=>"011110111",
  29078=>"100010000",
  29079=>"011111101",
  29080=>"010010001",
  29081=>"000100110",
  29082=>"011111111",
  29083=>"100011010",
  29084=>"101010111",
  29085=>"110100000",
  29086=>"000111010",
  29087=>"110001001",
  29088=>"000100100",
  29089=>"001110101",
  29090=>"001000000",
  29091=>"011110000",
  29092=>"100100111",
  29093=>"111110010",
  29094=>"011111000",
  29095=>"010000001",
  29096=>"101001011",
  29097=>"000111111",
  29098=>"000001100",
  29099=>"111101111",
  29100=>"100011000",
  29101=>"000100110",
  29102=>"100001110",
  29103=>"101111000",
  29104=>"101011000",
  29105=>"101101000",
  29106=>"000011001",
  29107=>"001000011",
  29108=>"000011111",
  29109=>"100010101",
  29110=>"000011010",
  29111=>"101000100",
  29112=>"110111110",
  29113=>"100111110",
  29114=>"111100111",
  29115=>"101111000",
  29116=>"011001100",
  29117=>"011001100",
  29118=>"110001010",
  29119=>"111000111",
  29120=>"101111100",
  29121=>"110111010",
  29122=>"101100010",
  29123=>"101001011",
  29124=>"111101101",
  29125=>"001000000",
  29126=>"101010100",
  29127=>"000000101",
  29128=>"001100111",
  29129=>"000010000",
  29130=>"111100011",
  29131=>"001010011",
  29132=>"001001110",
  29133=>"101011010",
  29134=>"101101111",
  29135=>"100111110",
  29136=>"101110110",
  29137=>"101111110",
  29138=>"101000011",
  29139=>"101101101",
  29140=>"100111111",
  29141=>"111010111",
  29142=>"000110011",
  29143=>"000101100",
  29144=>"011010010",
  29145=>"000011000",
  29146=>"111000110",
  29147=>"110000111",
  29148=>"010111101",
  29149=>"001001001",
  29150=>"111110000",
  29151=>"001010110",
  29152=>"010011001",
  29153=>"110010110",
  29154=>"110001111",
  29155=>"100001101",
  29156=>"001011011",
  29157=>"010000000",
  29158=>"001111111",
  29159=>"001000011",
  29160=>"111001001",
  29161=>"110011010",
  29162=>"000111110",
  29163=>"111101100",
  29164=>"011101001",
  29165=>"110110011",
  29166=>"111010100",
  29167=>"001001011",
  29168=>"100111111",
  29169=>"000110001",
  29170=>"010110100",
  29171=>"100000111",
  29172=>"111011111",
  29173=>"111000010",
  29174=>"111010000",
  29175=>"011000101",
  29176=>"110010100",
  29177=>"110111110",
  29178=>"110010000",
  29179=>"111011111",
  29180=>"011101101",
  29181=>"111000000",
  29182=>"110000101",
  29183=>"110100100",
  29184=>"100111010",
  29185=>"000111110",
  29186=>"110100000",
  29187=>"010000000",
  29188=>"101110101",
  29189=>"110110111",
  29190=>"000000010",
  29191=>"111100011",
  29192=>"011011111",
  29193=>"011100011",
  29194=>"111101010",
  29195=>"110011000",
  29196=>"011001111",
  29197=>"001011100",
  29198=>"000110111",
  29199=>"010110100",
  29200=>"101101001",
  29201=>"001010000",
  29202=>"100111011",
  29203=>"111100110",
  29204=>"001000111",
  29205=>"100010010",
  29206=>"011100111",
  29207=>"100001000",
  29208=>"000000100",
  29209=>"010010110",
  29210=>"011111010",
  29211=>"101011010",
  29212=>"100101011",
  29213=>"011000011",
  29214=>"111011100",
  29215=>"110111110",
  29216=>"100000010",
  29217=>"100001000",
  29218=>"000010001",
  29219=>"000000010",
  29220=>"000100110",
  29221=>"101001010",
  29222=>"111011000",
  29223=>"101000011",
  29224=>"100100101",
  29225=>"000110001",
  29226=>"000001001",
  29227=>"101000010",
  29228=>"100111101",
  29229=>"101101011",
  29230=>"100101101",
  29231=>"111111100",
  29232=>"010010101",
  29233=>"110100100",
  29234=>"100010101",
  29235=>"101011101",
  29236=>"010011010",
  29237=>"100001110",
  29238=>"101101101",
  29239=>"011111111",
  29240=>"010101110",
  29241=>"010010000",
  29242=>"010100100",
  29243=>"111000111",
  29244=>"110110101",
  29245=>"000100001",
  29246=>"000010001",
  29247=>"101111110",
  29248=>"100111010",
  29249=>"100011101",
  29250=>"001001001",
  29251=>"110010010",
  29252=>"011000111",
  29253=>"001111011",
  29254=>"011111111",
  29255=>"001001000",
  29256=>"011100111",
  29257=>"110100010",
  29258=>"011011100",
  29259=>"001001001",
  29260=>"000010000",
  29261=>"110101101",
  29262=>"101100111",
  29263=>"000000001",
  29264=>"111110100",
  29265=>"101011010",
  29266=>"001110100",
  29267=>"001111010",
  29268=>"111110000",
  29269=>"010111011",
  29270=>"110110110",
  29271=>"010101001",
  29272=>"000111100",
  29273=>"011100000",
  29274=>"111011101",
  29275=>"000101001",
  29276=>"101101100",
  29277=>"000000000",
  29278=>"111111110",
  29279=>"111111100",
  29280=>"100000110",
  29281=>"100010011",
  29282=>"111001100",
  29283=>"011111000",
  29284=>"010010110",
  29285=>"100111001",
  29286=>"011011100",
  29287=>"000110101",
  29288=>"011001101",
  29289=>"111111000",
  29290=>"101110110",
  29291=>"011011100",
  29292=>"000101100",
  29293=>"001110011",
  29294=>"011100000",
  29295=>"010010011",
  29296=>"001110111",
  29297=>"111111101",
  29298=>"001010110",
  29299=>"100111001",
  29300=>"100101110",
  29301=>"110011011",
  29302=>"000001000",
  29303=>"001101010",
  29304=>"001011100",
  29305=>"101000101",
  29306=>"101011110",
  29307=>"101101111",
  29308=>"011000000",
  29309=>"110110110",
  29310=>"011001100",
  29311=>"101110110",
  29312=>"000011100",
  29313=>"010011100",
  29314=>"101101111",
  29315=>"100010010",
  29316=>"011011111",
  29317=>"111111110",
  29318=>"101010111",
  29319=>"001001110",
  29320=>"100111111",
  29321=>"010001000",
  29322=>"110010001",
  29323=>"100101001",
  29324=>"110001010",
  29325=>"000111000",
  29326=>"111011000",
  29327=>"001101111",
  29328=>"011011000",
  29329=>"010100111",
  29330=>"100101000",
  29331=>"111101000",
  29332=>"100001000",
  29333=>"111000000",
  29334=>"001010000",
  29335=>"101001010",
  29336=>"010100111",
  29337=>"111011100",
  29338=>"101011101",
  29339=>"111110010",
  29340=>"001101101",
  29341=>"001001111",
  29342=>"010001111",
  29343=>"010001001",
  29344=>"011010100",
  29345=>"110101101",
  29346=>"101101001",
  29347=>"111101111",
  29348=>"011111101",
  29349=>"010110100",
  29350=>"000001110",
  29351=>"101110001",
  29352=>"010111110",
  29353=>"100111110",
  29354=>"011000010",
  29355=>"000100111",
  29356=>"111110001",
  29357=>"111100111",
  29358=>"011001110",
  29359=>"110001001",
  29360=>"001001010",
  29361=>"011011001",
  29362=>"011011000",
  29363=>"000011101",
  29364=>"101100110",
  29365=>"011011000",
  29366=>"110111011",
  29367=>"110010111",
  29368=>"001111001",
  29369=>"101000000",
  29370=>"100000111",
  29371=>"100111101",
  29372=>"011110010",
  29373=>"010011010",
  29374=>"100100101",
  29375=>"110001000",
  29376=>"001000110",
  29377=>"010011010",
  29378=>"111000110",
  29379=>"010011001",
  29380=>"001110111",
  29381=>"100100001",
  29382=>"101001101",
  29383=>"101110001",
  29384=>"000110010",
  29385=>"101111010",
  29386=>"100011010",
  29387=>"000111011",
  29388=>"000010000",
  29389=>"011110110",
  29390=>"001101001",
  29391=>"101110010",
  29392=>"100001000",
  29393=>"001110101",
  29394=>"101100001",
  29395=>"101101000",
  29396=>"011000111",
  29397=>"011110001",
  29398=>"001111110",
  29399=>"101100010",
  29400=>"000001100",
  29401=>"011110010",
  29402=>"001111000",
  29403=>"111000101",
  29404=>"100001110",
  29405=>"111100111",
  29406=>"110100000",
  29407=>"100100100",
  29408=>"000000000",
  29409=>"001010011",
  29410=>"111101000",
  29411=>"110010010",
  29412=>"000100110",
  29413=>"001000110",
  29414=>"000011111",
  29415=>"101011000",
  29416=>"010100000",
  29417=>"010010011",
  29418=>"011001110",
  29419=>"101111000",
  29420=>"010000011",
  29421=>"101111010",
  29422=>"011110101",
  29423=>"001010101",
  29424=>"101101110",
  29425=>"001101110",
  29426=>"100111110",
  29427=>"010010100",
  29428=>"010100010",
  29429=>"001001111",
  29430=>"000110011",
  29431=>"001111101",
  29432=>"110010100",
  29433=>"110010111",
  29434=>"111001011",
  29435=>"101001101",
  29436=>"001000110",
  29437=>"001001011",
  29438=>"010111100",
  29439=>"111001111",
  29440=>"001001001",
  29441=>"000110011",
  29442=>"000010110",
  29443=>"111111001",
  29444=>"011000000",
  29445=>"110110100",
  29446=>"000011010",
  29447=>"100001000",
  29448=>"111001011",
  29449=>"111010001",
  29450=>"100001010",
  29451=>"010110101",
  29452=>"000010110",
  29453=>"011011111",
  29454=>"000100100",
  29455=>"110001100",
  29456=>"101010001",
  29457=>"101001101",
  29458=>"000100100",
  29459=>"101100001",
  29460=>"111101000",
  29461=>"100100010",
  29462=>"011101111",
  29463=>"100101011",
  29464=>"000000001",
  29465=>"000001001",
  29466=>"011011001",
  29467=>"111001100",
  29468=>"011101110",
  29469=>"011100001",
  29470=>"100100000",
  29471=>"011111001",
  29472=>"110001110",
  29473=>"000011011",
  29474=>"110101011",
  29475=>"010000010",
  29476=>"001011111",
  29477=>"001000001",
  29478=>"000111000",
  29479=>"001010011",
  29480=>"001011111",
  29481=>"011110010",
  29482=>"110001000",
  29483=>"000001100",
  29484=>"100000101",
  29485=>"101101001",
  29486=>"110110001",
  29487=>"100010100",
  29488=>"000011011",
  29489=>"011110110",
  29490=>"000011001",
  29491=>"000110000",
  29492=>"101101111",
  29493=>"110011011",
  29494=>"001010001",
  29495=>"010010000",
  29496=>"010111001",
  29497=>"101111010",
  29498=>"011001100",
  29499=>"011000101",
  29500=>"100100010",
  29501=>"101011101",
  29502=>"000100001",
  29503=>"001010000",
  29504=>"100101100",
  29505=>"001011000",
  29506=>"100111111",
  29507=>"101000000",
  29508=>"111000011",
  29509=>"001011110",
  29510=>"000110110",
  29511=>"111010101",
  29512=>"000000100",
  29513=>"001001100",
  29514=>"101000100",
  29515=>"010100001",
  29516=>"000010001",
  29517=>"110010101",
  29518=>"010000011",
  29519=>"110000110",
  29520=>"110110100",
  29521=>"000100110",
  29522=>"000000010",
  29523=>"000001011",
  29524=>"110110111",
  29525=>"010001101",
  29526=>"111011000",
  29527=>"010101101",
  29528=>"011100101",
  29529=>"001011101",
  29530=>"111110010",
  29531=>"010000111",
  29532=>"011111011",
  29533=>"001010010",
  29534=>"000001101",
  29535=>"001101010",
  29536=>"001110101",
  29537=>"001111100",
  29538=>"100000011",
  29539=>"111010011",
  29540=>"000000010",
  29541=>"001010101",
  29542=>"110000011",
  29543=>"001100110",
  29544=>"000001101",
  29545=>"101111001",
  29546=>"000010111",
  29547=>"101011101",
  29548=>"100000000",
  29549=>"001000001",
  29550=>"100100100",
  29551=>"010000111",
  29552=>"110001110",
  29553=>"001100000",
  29554=>"010110001",
  29555=>"000000011",
  29556=>"110111111",
  29557=>"111101010",
  29558=>"010000011",
  29559=>"110010011",
  29560=>"101100111",
  29561=>"010000101",
  29562=>"110100110",
  29563=>"101100110",
  29564=>"100001110",
  29565=>"011011000",
  29566=>"101111101",
  29567=>"100000011",
  29568=>"101011111",
  29569=>"000010011",
  29570=>"100100000",
  29571=>"101100001",
  29572=>"100001011",
  29573=>"010010011",
  29574=>"001001111",
  29575=>"110100000",
  29576=>"100000010",
  29577=>"010111011",
  29578=>"011110101",
  29579=>"001000100",
  29580=>"001001010",
  29581=>"111110011",
  29582=>"011010100",
  29583=>"000100100",
  29584=>"111001101",
  29585=>"100110111",
  29586=>"010101101",
  29587=>"111000011",
  29588=>"101000100",
  29589=>"010111000",
  29590=>"100100101",
  29591=>"000101110",
  29592=>"010011011",
  29593=>"010000100",
  29594=>"101101101",
  29595=>"110110101",
  29596=>"100000110",
  29597=>"101001111",
  29598=>"111001101",
  29599=>"000010100",
  29600=>"100011100",
  29601=>"011001010",
  29602=>"110110010",
  29603=>"000100010",
  29604=>"000010001",
  29605=>"111111111",
  29606=>"000001100",
  29607=>"011101011",
  29608=>"100101111",
  29609=>"010111000",
  29610=>"110101010",
  29611=>"011010000",
  29612=>"110100010",
  29613=>"000010000",
  29614=>"100100011",
  29615=>"000101011",
  29616=>"011011111",
  29617=>"110000111",
  29618=>"110100101",
  29619=>"100001000",
  29620=>"000101011",
  29621=>"000100001",
  29622=>"101111000",
  29623=>"111010010",
  29624=>"111011110",
  29625=>"100110110",
  29626=>"010010000",
  29627=>"011011101",
  29628=>"010010000",
  29629=>"111111111",
  29630=>"001111110",
  29631=>"100001100",
  29632=>"001100111",
  29633=>"011110101",
  29634=>"000001000",
  29635=>"000010000",
  29636=>"101001000",
  29637=>"011111101",
  29638=>"110101101",
  29639=>"001011010",
  29640=>"101001111",
  29641=>"111000101",
  29642=>"011100100",
  29643=>"100100011",
  29644=>"110000100",
  29645=>"001101100",
  29646=>"010001000",
  29647=>"101000000",
  29648=>"101000100",
  29649=>"000000111",
  29650=>"000010011",
  29651=>"000101110",
  29652=>"110000001",
  29653=>"010000000",
  29654=>"010001000",
  29655=>"010011000",
  29656=>"000110000",
  29657=>"111000000",
  29658=>"001000000",
  29659=>"001000101",
  29660=>"100000100",
  29661=>"010111010",
  29662=>"001001010",
  29663=>"000001000",
  29664=>"001110110",
  29665=>"100100010",
  29666=>"000010110",
  29667=>"001111000",
  29668=>"100110000",
  29669=>"011101111",
  29670=>"001101011",
  29671=>"000111111",
  29672=>"000000010",
  29673=>"010101011",
  29674=>"001101001",
  29675=>"000100100",
  29676=>"010011000",
  29677=>"011001100",
  29678=>"101001100",
  29679=>"110011001",
  29680=>"010000000",
  29681=>"100011110",
  29682=>"110100010",
  29683=>"101110011",
  29684=>"011111011",
  29685=>"110110001",
  29686=>"001001110",
  29687=>"010101011",
  29688=>"000010010",
  29689=>"011011000",
  29690=>"010000110",
  29691=>"100000110",
  29692=>"001101111",
  29693=>"011011001",
  29694=>"001011101",
  29695=>"011011010",
  29696=>"010000000",
  29697=>"111100111",
  29698=>"011111101",
  29699=>"000000000",
  29700=>"111010001",
  29701=>"000000011",
  29702=>"100011101",
  29703=>"111101001",
  29704=>"110110100",
  29705=>"100111101",
  29706=>"011001110",
  29707=>"100011001",
  29708=>"011001101",
  29709=>"001110100",
  29710=>"111010111",
  29711=>"000010001",
  29712=>"011100101",
  29713=>"000110101",
  29714=>"101111010",
  29715=>"000110100",
  29716=>"000001011",
  29717=>"111111001",
  29718=>"001111110",
  29719=>"001101011",
  29720=>"001011001",
  29721=>"000010100",
  29722=>"000101001",
  29723=>"000000000",
  29724=>"111010100",
  29725=>"001111111",
  29726=>"001111001",
  29727=>"001001010",
  29728=>"011001000",
  29729=>"010110011",
  29730=>"001000011",
  29731=>"111000000",
  29732=>"000011011",
  29733=>"101110100",
  29734=>"100000011",
  29735=>"111111100",
  29736=>"110100001",
  29737=>"010110111",
  29738=>"001000010",
  29739=>"111110011",
  29740=>"011000010",
  29741=>"000111111",
  29742=>"001011110",
  29743=>"010100111",
  29744=>"001001001",
  29745=>"110101100",
  29746=>"001001001",
  29747=>"111100011",
  29748=>"101101011",
  29749=>"110001000",
  29750=>"110101000",
  29751=>"110001011",
  29752=>"101111011",
  29753=>"110111101",
  29754=>"111100111",
  29755=>"000000110",
  29756=>"110010101",
  29757=>"000111001",
  29758=>"100000111",
  29759=>"101001010",
  29760=>"000011000",
  29761=>"011101010",
  29762=>"110010011",
  29763=>"110101110",
  29764=>"010011110",
  29765=>"101010001",
  29766=>"101011110",
  29767=>"011011101",
  29768=>"000001000",
  29769=>"010101000",
  29770=>"111111101",
  29771=>"010100011",
  29772=>"101101011",
  29773=>"110011011",
  29774=>"101000000",
  29775=>"010110111",
  29776=>"100110100",
  29777=>"001010100",
  29778=>"100100100",
  29779=>"101101111",
  29780=>"101111011",
  29781=>"010000100",
  29782=>"110111100",
  29783=>"001010001",
  29784=>"000010011",
  29785=>"111101001",
  29786=>"111110101",
  29787=>"100110010",
  29788=>"100001000",
  29789=>"000010011",
  29790=>"111001010",
  29791=>"100010000",
  29792=>"001001111",
  29793=>"110001011",
  29794=>"101001000",
  29795=>"011111001",
  29796=>"110000000",
  29797=>"100110000",
  29798=>"000110001",
  29799=>"011010111",
  29800=>"101011001",
  29801=>"010101111",
  29802=>"000101100",
  29803=>"000110100",
  29804=>"101010100",
  29805=>"000000000",
  29806=>"000000000",
  29807=>"010001010",
  29808=>"110010011",
  29809=>"001001000",
  29810=>"000011100",
  29811=>"010111111",
  29812=>"000010110",
  29813=>"111000100",
  29814=>"100011001",
  29815=>"011101010",
  29816=>"101011110",
  29817=>"101000001",
  29818=>"011111010",
  29819=>"101011001",
  29820=>"010011111",
  29821=>"100001001",
  29822=>"000001011",
  29823=>"111101000",
  29824=>"110110001",
  29825=>"000111100",
  29826=>"111011001",
  29827=>"111001101",
  29828=>"000010000",
  29829=>"101110101",
  29830=>"100000001",
  29831=>"010011010",
  29832=>"001111011",
  29833=>"011010010",
  29834=>"110101101",
  29835=>"001011001",
  29836=>"100010011",
  29837=>"000010101",
  29838=>"000001110",
  29839=>"011010100",
  29840=>"001111011",
  29841=>"001110110",
  29842=>"010100101",
  29843=>"101100100",
  29844=>"110101110",
  29845=>"000101000",
  29846=>"010111011",
  29847=>"110111011",
  29848=>"101010010",
  29849=>"010011111",
  29850=>"101010011",
  29851=>"111111111",
  29852=>"011100110",
  29853=>"111101000",
  29854=>"010110011",
  29855=>"110000100",
  29856=>"001001011",
  29857=>"011100110",
  29858=>"001110000",
  29859=>"101101001",
  29860=>"011111001",
  29861=>"100100000",
  29862=>"101110101",
  29863=>"010011011",
  29864=>"101010111",
  29865=>"101010111",
  29866=>"000110100",
  29867=>"100010000",
  29868=>"100010010",
  29869=>"001110011",
  29870=>"110101101",
  29871=>"011101110",
  29872=>"101110110",
  29873=>"110101111",
  29874=>"010111110",
  29875=>"011010011",
  29876=>"000000001",
  29877=>"001010000",
  29878=>"011011110",
  29879=>"110111111",
  29880=>"101110010",
  29881=>"101000110",
  29882=>"011111001",
  29883=>"110111110",
  29884=>"100111101",
  29885=>"011101001",
  29886=>"100010111",
  29887=>"111101000",
  29888=>"100000011",
  29889=>"011010110",
  29890=>"111101011",
  29891=>"100010101",
  29892=>"100001111",
  29893=>"111110100",
  29894=>"110100001",
  29895=>"101110100",
  29896=>"110010100",
  29897=>"101110110",
  29898=>"001000111",
  29899=>"010100010",
  29900=>"011111111",
  29901=>"111010010",
  29902=>"010010111",
  29903=>"010010011",
  29904=>"101000011",
  29905=>"011000100",
  29906=>"001001010",
  29907=>"000011101",
  29908=>"011111001",
  29909=>"000110001",
  29910=>"100010000",
  29911=>"101000001",
  29912=>"001011011",
  29913=>"010001000",
  29914=>"010000101",
  29915=>"101110100",
  29916=>"010000000",
  29917=>"101000000",
  29918=>"101100010",
  29919=>"110100111",
  29920=>"101011001",
  29921=>"110011001",
  29922=>"011000001",
  29923=>"010000010",
  29924=>"100111000",
  29925=>"101111111",
  29926=>"111011111",
  29927=>"111111111",
  29928=>"111001100",
  29929=>"111100110",
  29930=>"101110111",
  29931=>"010111010",
  29932=>"000001110",
  29933=>"001010010",
  29934=>"011000101",
  29935=>"100010000",
  29936=>"000100010",
  29937=>"111100111",
  29938=>"001110010",
  29939=>"110110101",
  29940=>"110001001",
  29941=>"010110111",
  29942=>"110101000",
  29943=>"010110011",
  29944=>"111101011",
  29945=>"111001101",
  29946=>"001011110",
  29947=>"010100101",
  29948=>"111100011",
  29949=>"111100110",
  29950=>"011110010",
  29951=>"111000101",
  29952=>"110010000",
  29953=>"111100010",
  29954=>"001011010",
  29955=>"110000111",
  29956=>"000110110",
  29957=>"010000011",
  29958=>"111000000",
  29959=>"111110111",
  29960=>"000101010",
  29961=>"011011010",
  29962=>"101011101",
  29963=>"100010101",
  29964=>"111110001",
  29965=>"001011001",
  29966=>"111010101",
  29967=>"010001100",
  29968=>"100101000",
  29969=>"111011001",
  29970=>"011000001",
  29971=>"100100011",
  29972=>"110010010",
  29973=>"011100000",
  29974=>"101100110",
  29975=>"011011000",
  29976=>"101010101",
  29977=>"011110111",
  29978=>"111111100",
  29979=>"001011100",
  29980=>"011101100",
  29981=>"010011011",
  29982=>"101000100",
  29983=>"110011011",
  29984=>"111010000",
  29985=>"000111001",
  29986=>"101110100",
  29987=>"000100011",
  29988=>"100110100",
  29989=>"010100010",
  29990=>"011110111",
  29991=>"101100111",
  29992=>"001000000",
  29993=>"100000000",
  29994=>"011011111",
  29995=>"100000011",
  29996=>"001000111",
  29997=>"101010110",
  29998=>"101000101",
  29999=>"010101111",
  30000=>"100001001",
  30001=>"101010000",
  30002=>"000011110",
  30003=>"001010101",
  30004=>"001011011",
  30005=>"001110111",
  30006=>"100011010",
  30007=>"000110000",
  30008=>"000111111",
  30009=>"000100001",
  30010=>"000101001",
  30011=>"111110011",
  30012=>"111101001",
  30013=>"001000101",
  30014=>"101010001",
  30015=>"110101111",
  30016=>"000110010",
  30017=>"111011111",
  30018=>"100101001",
  30019=>"101101111",
  30020=>"000111110",
  30021=>"000111001",
  30022=>"110100100",
  30023=>"000000001",
  30024=>"011110011",
  30025=>"111010010",
  30026=>"100011111",
  30027=>"101110000",
  30028=>"100001001",
  30029=>"110101110",
  30030=>"000011110",
  30031=>"000111111",
  30032=>"110101000",
  30033=>"100110010",
  30034=>"111101111",
  30035=>"001101111",
  30036=>"110010001",
  30037=>"001000011",
  30038=>"101000110",
  30039=>"010011011",
  30040=>"111111000",
  30041=>"001011001",
  30042=>"001101110",
  30043=>"111000010",
  30044=>"000000100",
  30045=>"010001000",
  30046=>"110111100",
  30047=>"100100101",
  30048=>"000010110",
  30049=>"110000000",
  30050=>"010011100",
  30051=>"001011011",
  30052=>"010101100",
  30053=>"011000110",
  30054=>"011000001",
  30055=>"100011001",
  30056=>"000101010",
  30057=>"000101110",
  30058=>"110111110",
  30059=>"011011111",
  30060=>"010010111",
  30061=>"110111111",
  30062=>"000011001",
  30063=>"110100011",
  30064=>"001010100",
  30065=>"001100001",
  30066=>"111101001",
  30067=>"001011101",
  30068=>"111010000",
  30069=>"011010000",
  30070=>"111110010",
  30071=>"010011011",
  30072=>"101000101",
  30073=>"111000000",
  30074=>"101101001",
  30075=>"011101000",
  30076=>"001000011",
  30077=>"001010001",
  30078=>"001100111",
  30079=>"110101101",
  30080=>"101111101",
  30081=>"110111010",
  30082=>"100000100",
  30083=>"000001101",
  30084=>"111011000",
  30085=>"000010101",
  30086=>"100111010",
  30087=>"010000101",
  30088=>"001001011",
  30089=>"000101001",
  30090=>"011100100",
  30091=>"101110011",
  30092=>"000000010",
  30093=>"011001011",
  30094=>"111010000",
  30095=>"000110011",
  30096=>"101101001",
  30097=>"111010101",
  30098=>"101010011",
  30099=>"011001101",
  30100=>"000100101",
  30101=>"001110111",
  30102=>"010010100",
  30103=>"010011000",
  30104=>"001000001",
  30105=>"111010010",
  30106=>"100111010",
  30107=>"001101010",
  30108=>"100010001",
  30109=>"011000100",
  30110=>"101101100",
  30111=>"100111001",
  30112=>"000010101",
  30113=>"010001000",
  30114=>"010000000",
  30115=>"111100011",
  30116=>"111101011",
  30117=>"111111000",
  30118=>"101000000",
  30119=>"110011001",
  30120=>"100011011",
  30121=>"001110011",
  30122=>"100000011",
  30123=>"111101111",
  30124=>"101111111",
  30125=>"011011011",
  30126=>"110011100",
  30127=>"101010001",
  30128=>"010001101",
  30129=>"010000111",
  30130=>"101101101",
  30131=>"110100100",
  30132=>"100011100",
  30133=>"000010110",
  30134=>"100100010",
  30135=>"000111110",
  30136=>"100110110",
  30137=>"110111010",
  30138=>"011010101",
  30139=>"011000100",
  30140=>"010111011",
  30141=>"110101111",
  30142=>"111111000",
  30143=>"111111110",
  30144=>"110000000",
  30145=>"001111110",
  30146=>"000110010",
  30147=>"101110000",
  30148=>"010111101",
  30149=>"010100111",
  30150=>"111111111",
  30151=>"001001101",
  30152=>"100001010",
  30153=>"011011011",
  30154=>"100101010",
  30155=>"011001000",
  30156=>"100111110",
  30157=>"101110111",
  30158=>"010101000",
  30159=>"101101100",
  30160=>"110000000",
  30161=>"010101011",
  30162=>"001011100",
  30163=>"100101100",
  30164=>"011011111",
  30165=>"000100111",
  30166=>"100110111",
  30167=>"110011001",
  30168=>"010000011",
  30169=>"111100011",
  30170=>"011000010",
  30171=>"110010100",
  30172=>"010011001",
  30173=>"011101000",
  30174=>"000001001",
  30175=>"000110111",
  30176=>"010001010",
  30177=>"110010011",
  30178=>"001111100",
  30179=>"110100000",
  30180=>"000001001",
  30181=>"111111111",
  30182=>"001100000",
  30183=>"101110111",
  30184=>"001101010",
  30185=>"111010101",
  30186=>"001000101",
  30187=>"001111000",
  30188=>"101000001",
  30189=>"111010101",
  30190=>"001101001",
  30191=>"010011011",
  30192=>"111001110",
  30193=>"001101000",
  30194=>"011111100",
  30195=>"110001100",
  30196=>"101101010",
  30197=>"000001100",
  30198=>"111110010",
  30199=>"010000010",
  30200=>"000010111",
  30201=>"001100000",
  30202=>"000000000",
  30203=>"110010011",
  30204=>"100111001",
  30205=>"110010110",
  30206=>"000110111",
  30207=>"001000111",
  30208=>"010011000",
  30209=>"001110011",
  30210=>"011000100",
  30211=>"110100110",
  30212=>"110100110",
  30213=>"111101111",
  30214=>"101001111",
  30215=>"100011011",
  30216=>"111001111",
  30217=>"010011101",
  30218=>"011011011",
  30219=>"010100000",
  30220=>"101010001",
  30221=>"110101000",
  30222=>"110110011",
  30223=>"110111011",
  30224=>"111111101",
  30225=>"000111001",
  30226=>"000110001",
  30227=>"111100011",
  30228=>"101010101",
  30229=>"101010011",
  30230=>"110111101",
  30231=>"000101110",
  30232=>"011100110",
  30233=>"110101111",
  30234=>"011111010",
  30235=>"101100101",
  30236=>"011010101",
  30237=>"100000100",
  30238=>"101111010",
  30239=>"100110010",
  30240=>"011110011",
  30241=>"111101011",
  30242=>"010001101",
  30243=>"110011001",
  30244=>"011010100",
  30245=>"111011010",
  30246=>"011001010",
  30247=>"011101110",
  30248=>"111100101",
  30249=>"111000100",
  30250=>"011111100",
  30251=>"011000000",
  30252=>"001110101",
  30253=>"110001010",
  30254=>"101001111",
  30255=>"010010010",
  30256=>"010100110",
  30257=>"011001010",
  30258=>"111001011",
  30259=>"010101100",
  30260=>"010011011",
  30261=>"111000001",
  30262=>"111000111",
  30263=>"110010010",
  30264=>"111010000",
  30265=>"001011101",
  30266=>"010101011",
  30267=>"000000110",
  30268=>"000110111",
  30269=>"000101100",
  30270=>"111010111",
  30271=>"110111100",
  30272=>"001000011",
  30273=>"111110010",
  30274=>"000101101",
  30275=>"010010010",
  30276=>"000110011",
  30277=>"001010000",
  30278=>"010000000",
  30279=>"000000101",
  30280=>"111101100",
  30281=>"111001101",
  30282=>"110110101",
  30283=>"110111111",
  30284=>"000011011",
  30285=>"111111111",
  30286=>"001101110",
  30287=>"000001010",
  30288=>"001001111",
  30289=>"111111100",
  30290=>"100111100",
  30291=>"110010110",
  30292=>"101000101",
  30293=>"100010110",
  30294=>"100011000",
  30295=>"011001110",
  30296=>"111011010",
  30297=>"101111010",
  30298=>"100100110",
  30299=>"110101010",
  30300=>"100010100",
  30301=>"010100011",
  30302=>"010110101",
  30303=>"111011111",
  30304=>"110110111",
  30305=>"010110110",
  30306=>"011100000",
  30307=>"100011000",
  30308=>"100011101",
  30309=>"100101010",
  30310=>"011011001",
  30311=>"110110110",
  30312=>"100000100",
  30313=>"110000101",
  30314=>"111101110",
  30315=>"011011111",
  30316=>"010110010",
  30317=>"011010000",
  30318=>"110110111",
  30319=>"000110111",
  30320=>"011000101",
  30321=>"000001110",
  30322=>"010110110",
  30323=>"111011111",
  30324=>"011011000",
  30325=>"100000110",
  30326=>"011011101",
  30327=>"011111101",
  30328=>"101101000",
  30329=>"101101101",
  30330=>"011101000",
  30331=>"001111101",
  30332=>"110111101",
  30333=>"011101111",
  30334=>"000100001",
  30335=>"100110111",
  30336=>"001010110",
  30337=>"000011001",
  30338=>"010011100",
  30339=>"111000110",
  30340=>"100010001",
  30341=>"001010011",
  30342=>"100010100",
  30343=>"111001010",
  30344=>"111110101",
  30345=>"111110010",
  30346=>"010111000",
  30347=>"110111000",
  30348=>"000010110",
  30349=>"011001000",
  30350=>"011100100",
  30351=>"011001101",
  30352=>"001010011",
  30353=>"100011100",
  30354=>"100011111",
  30355=>"010100001",
  30356=>"110000001",
  30357=>"111111010",
  30358=>"000100100",
  30359=>"001110110",
  30360=>"000000101",
  30361=>"101001100",
  30362=>"100000010",
  30363=>"010101001",
  30364=>"101101110",
  30365=>"100100100",
  30366=>"010111101",
  30367=>"011000110",
  30368=>"111101111",
  30369=>"010101011",
  30370=>"111101101",
  30371=>"110101111",
  30372=>"011111111",
  30373=>"101111111",
  30374=>"011101000",
  30375=>"110101011",
  30376=>"111101000",
  30377=>"101001000",
  30378=>"001001111",
  30379=>"011101010",
  30380=>"110001010",
  30381=>"000101001",
  30382=>"011111111",
  30383=>"000001111",
  30384=>"000001111",
  30385=>"000000000",
  30386=>"110000100",
  30387=>"101011000",
  30388=>"101010100",
  30389=>"010000010",
  30390=>"011101101",
  30391=>"100111101",
  30392=>"000000110",
  30393=>"010001001",
  30394=>"011101001",
  30395=>"100111110",
  30396=>"111001111",
  30397=>"111011010",
  30398=>"011000001",
  30399=>"011001100",
  30400=>"001001010",
  30401=>"001010010",
  30402=>"101110011",
  30403=>"001110100",
  30404=>"001000010",
  30405=>"000110000",
  30406=>"100111110",
  30407=>"000111111",
  30408=>"010101100",
  30409=>"111111110",
  30410=>"001010100",
  30411=>"000010110",
  30412=>"011101111",
  30413=>"000100001",
  30414=>"100011001",
  30415=>"011110000",
  30416=>"100110001",
  30417=>"010001100",
  30418=>"010100111",
  30419=>"010110111",
  30420=>"111011000",
  30421=>"000000100",
  30422=>"100101101",
  30423=>"010111110",
  30424=>"001001010",
  30425=>"011100101",
  30426=>"100111100",
  30427=>"100011100",
  30428=>"010110010",
  30429=>"001101010",
  30430=>"111100101",
  30431=>"111110001",
  30432=>"100000110",
  30433=>"100011001",
  30434=>"000111111",
  30435=>"111111111",
  30436=>"101001011",
  30437=>"111110110",
  30438=>"101001110",
  30439=>"101001000",
  30440=>"111010000",
  30441=>"101110001",
  30442=>"001110010",
  30443=>"101010100",
  30444=>"000101011",
  30445=>"101111000",
  30446=>"111111110",
  30447=>"001010101",
  30448=>"110111100",
  30449=>"011100001",
  30450=>"010001010",
  30451=>"011110111",
  30452=>"101111010",
  30453=>"100000110",
  30454=>"011100011",
  30455=>"011100100",
  30456=>"111000110",
  30457=>"111011001",
  30458=>"101000101",
  30459=>"001000001",
  30460=>"011011011",
  30461=>"010101110",
  30462=>"110010011",
  30463=>"011011000",
  30464=>"100011110",
  30465=>"010011100",
  30466=>"101110100",
  30467=>"011110000",
  30468=>"010100011",
  30469=>"010110010",
  30470=>"100110001",
  30471=>"010010010",
  30472=>"011011111",
  30473=>"110001010",
  30474=>"101110111",
  30475=>"111001101",
  30476=>"010011010",
  30477=>"100010111",
  30478=>"000010100",
  30479=>"001011111",
  30480=>"010111111",
  30481=>"011110010",
  30482=>"010100011",
  30483=>"100010110",
  30484=>"001111100",
  30485=>"111111101",
  30486=>"010100011",
  30487=>"000000101",
  30488=>"110111101",
  30489=>"001100101",
  30490=>"100100101",
  30491=>"001101110",
  30492=>"110110101",
  30493=>"110011100",
  30494=>"000100101",
  30495=>"101000101",
  30496=>"111111111",
  30497=>"000000101",
  30498=>"101001110",
  30499=>"011110101",
  30500=>"011001010",
  30501=>"010000101",
  30502=>"101101110",
  30503=>"001110101",
  30504=>"111111011",
  30505=>"110110111",
  30506=>"100001101",
  30507=>"011000110",
  30508=>"000010000",
  30509=>"001001010",
  30510=>"000011011",
  30511=>"011110001",
  30512=>"001110111",
  30513=>"001111111",
  30514=>"010000011",
  30515=>"000001111",
  30516=>"000010001",
  30517=>"001000010",
  30518=>"000010011",
  30519=>"110001001",
  30520=>"110100001",
  30521=>"011100011",
  30522=>"101001101",
  30523=>"101010000",
  30524=>"011000101",
  30525=>"110101111",
  30526=>"011110010",
  30527=>"101000101",
  30528=>"001100111",
  30529=>"001001100",
  30530=>"110011101",
  30531=>"001100110",
  30532=>"110101100",
  30533=>"011111111",
  30534=>"011111100",
  30535=>"101000011",
  30536=>"011011001",
  30537=>"101000000",
  30538=>"000000010",
  30539=>"110101101",
  30540=>"111001000",
  30541=>"101010010",
  30542=>"100011111",
  30543=>"000111111",
  30544=>"111011000",
  30545=>"010100110",
  30546=>"111101101",
  30547=>"010000111",
  30548=>"100101000",
  30549=>"011011101",
  30550=>"101101101",
  30551=>"000011011",
  30552=>"100111111",
  30553=>"011111100",
  30554=>"100001101",
  30555=>"011000000",
  30556=>"010011110",
  30557=>"111100111",
  30558=>"111111111",
  30559=>"011101011",
  30560=>"011100101",
  30561=>"110001011",
  30562=>"000010011",
  30563=>"010101011",
  30564=>"000001100",
  30565=>"001000111",
  30566=>"111000001",
  30567=>"001110000",
  30568=>"111010000",
  30569=>"011001110",
  30570=>"100100110",
  30571=>"110101111",
  30572=>"100001100",
  30573=>"110110101",
  30574=>"000011011",
  30575=>"000000000",
  30576=>"101001011",
  30577=>"111010100",
  30578=>"010110011",
  30579=>"111101110",
  30580=>"101111101",
  30581=>"010011000",
  30582=>"110101011",
  30583=>"100100111",
  30584=>"001110010",
  30585=>"001101111",
  30586=>"101011001",
  30587=>"101001001",
  30588=>"001100100",
  30589=>"011010111",
  30590=>"100100110",
  30591=>"100111110",
  30592=>"000110001",
  30593=>"111011000",
  30594=>"110111001",
  30595=>"011000100",
  30596=>"110100111",
  30597=>"111100000",
  30598=>"001011111",
  30599=>"000001001",
  30600=>"010100101",
  30601=>"101110111",
  30602=>"001000010",
  30603=>"111100111",
  30604=>"011101100",
  30605=>"011100000",
  30606=>"010111001",
  30607=>"111000101",
  30608=>"111011111",
  30609=>"101010001",
  30610=>"000001110",
  30611=>"110111011",
  30612=>"110000010",
  30613=>"001001100",
  30614=>"110101110",
  30615=>"000011100",
  30616=>"101001110",
  30617=>"011101100",
  30618=>"111011111",
  30619=>"001001100",
  30620=>"111000100",
  30621=>"111101110",
  30622=>"010111111",
  30623=>"111101010",
  30624=>"100101010",
  30625=>"001111100",
  30626=>"011000001",
  30627=>"110101101",
  30628=>"111001110",
  30629=>"001010110",
  30630=>"100100110",
  30631=>"110010110",
  30632=>"010101110",
  30633=>"000010111",
  30634=>"100000110",
  30635=>"110000100",
  30636=>"011010100",
  30637=>"000100011",
  30638=>"110111000",
  30639=>"010000001",
  30640=>"110111010",
  30641=>"001011010",
  30642=>"011010100",
  30643=>"111111101",
  30644=>"110100000",
  30645=>"011000100",
  30646=>"001001001",
  30647=>"100011001",
  30648=>"111111001",
  30649=>"100001111",
  30650=>"000011110",
  30651=>"001111000",
  30652=>"011110110",
  30653=>"110001111",
  30654=>"000011101",
  30655=>"011111111",
  30656=>"111011101",
  30657=>"000001100",
  30658=>"000110110",
  30659=>"111001110",
  30660=>"011011111",
  30661=>"110011110",
  30662=>"101110101",
  30663=>"001110011",
  30664=>"011110110",
  30665=>"011110100",
  30666=>"000000111",
  30667=>"101101011",
  30668=>"011100011",
  30669=>"011110110",
  30670=>"000000011",
  30671=>"011101011",
  30672=>"101011010",
  30673=>"001011110",
  30674=>"111110111",
  30675=>"010001001",
  30676=>"010010000",
  30677=>"011011100",
  30678=>"011101011",
  30679=>"110100111",
  30680=>"011101000",
  30681=>"100100011",
  30682=>"110110000",
  30683=>"110100010",
  30684=>"101011011",
  30685=>"001101001",
  30686=>"001101110",
  30687=>"100000100",
  30688=>"111010010",
  30689=>"110000010",
  30690=>"111000000",
  30691=>"000001011",
  30692=>"010000101",
  30693=>"100001000",
  30694=>"001011110",
  30695=>"101000101",
  30696=>"001000101",
  30697=>"101000111",
  30698=>"101111101",
  30699=>"010011011",
  30700=>"001101000",
  30701=>"110000000",
  30702=>"001000100",
  30703=>"001100101",
  30704=>"100101110",
  30705=>"010100011",
  30706=>"111100001",
  30707=>"111000110",
  30708=>"011011101",
  30709=>"000101110",
  30710=>"000100110",
  30711=>"100001101",
  30712=>"010101101",
  30713=>"001110111",
  30714=>"100000001",
  30715=>"001111111",
  30716=>"000010000",
  30717=>"001101111",
  30718=>"010010000",
  30719=>"001011011",
  30720=>"110100101",
  30721=>"110000110",
  30722=>"011011100",
  30723=>"000010010",
  30724=>"100100011",
  30725=>"000000010",
  30726=>"100010011",
  30727=>"001100000",
  30728=>"001010001",
  30729=>"000100100",
  30730=>"010000111",
  30731=>"101111111",
  30732=>"111000000",
  30733=>"111110010",
  30734=>"110000101",
  30735=>"110110001",
  30736=>"111001100",
  30737=>"000011100",
  30738=>"100010100",
  30739=>"110111001",
  30740=>"100001111",
  30741=>"101111000",
  30742=>"111111111",
  30743=>"011011100",
  30744=>"011001101",
  30745=>"110100101",
  30746=>"111000010",
  30747=>"100001110",
  30748=>"110101100",
  30749=>"110110010",
  30750=>"110111001",
  30751=>"010000100",
  30752=>"111111100",
  30753=>"110000101",
  30754=>"001101010",
  30755=>"000100010",
  30756=>"101100111",
  30757=>"100101110",
  30758=>"100000100",
  30759=>"000001101",
  30760=>"100000100",
  30761=>"110110011",
  30762=>"111010010",
  30763=>"101101101",
  30764=>"001001011",
  30765=>"111000111",
  30766=>"011010000",
  30767=>"101101110",
  30768=>"110001000",
  30769=>"001011011",
  30770=>"101100011",
  30771=>"110001011",
  30772=>"011000000",
  30773=>"000010101",
  30774=>"110000000",
  30775=>"000111101",
  30776=>"100011111",
  30777=>"011100011",
  30778=>"010010001",
  30779=>"001011101",
  30780=>"010010111",
  30781=>"011010101",
  30782=>"110011000",
  30783=>"010000100",
  30784=>"100111010",
  30785=>"001000001",
  30786=>"000010100",
  30787=>"001110101",
  30788=>"111000110",
  30789=>"101101110",
  30790=>"111011011",
  30791=>"010100101",
  30792=>"110110101",
  30793=>"000111001",
  30794=>"000000000",
  30795=>"010010001",
  30796=>"100010001",
  30797=>"010101100",
  30798=>"110100000",
  30799=>"101001000",
  30800=>"010010110",
  30801=>"000011101",
  30802=>"010100110",
  30803=>"101100010",
  30804=>"110011001",
  30805=>"001001111",
  30806=>"110100001",
  30807=>"111001001",
  30808=>"001101110",
  30809=>"001100010",
  30810=>"111111110",
  30811=>"001101100",
  30812=>"001010010",
  30813=>"100011000",
  30814=>"101111001",
  30815=>"111101110",
  30816=>"000000011",
  30817=>"001111100",
  30818=>"010110110",
  30819=>"000000001",
  30820=>"101101001",
  30821=>"111111010",
  30822=>"011111111",
  30823=>"100110100",
  30824=>"110001001",
  30825=>"101110100",
  30826=>"111011000",
  30827=>"110101011",
  30828=>"010111100",
  30829=>"000100111",
  30830=>"101000000",
  30831=>"100101100",
  30832=>"110100001",
  30833=>"011001001",
  30834=>"001100110",
  30835=>"111001011",
  30836=>"001100011",
  30837=>"011100110",
  30838=>"001111011",
  30839=>"101101100",
  30840=>"011011111",
  30841=>"010011001",
  30842=>"101011010",
  30843=>"101111111",
  30844=>"010010001",
  30845=>"011010100",
  30846=>"101010111",
  30847=>"000010110",
  30848=>"100000011",
  30849=>"010111011",
  30850=>"110001110",
  30851=>"001011100",
  30852=>"000111111",
  30853=>"010101110",
  30854=>"011011011",
  30855=>"111000010",
  30856=>"110000010",
  30857=>"011001010",
  30858=>"010111110",
  30859=>"010011100",
  30860=>"001101101",
  30861=>"000110101",
  30862=>"100101110",
  30863=>"110111101",
  30864=>"110001110",
  30865=>"101100001",
  30866=>"100010111",
  30867=>"011101001",
  30868=>"001110010",
  30869=>"110000110",
  30870=>"000111110",
  30871=>"010011000",
  30872=>"010111000",
  30873=>"101100001",
  30874=>"110000010",
  30875=>"011101101",
  30876=>"111111111",
  30877=>"011011110",
  30878=>"101001010",
  30879=>"110100111",
  30880=>"110110001",
  30881=>"011001011",
  30882=>"111010010",
  30883=>"000001011",
  30884=>"001000111",
  30885=>"011011010",
  30886=>"001010000",
  30887=>"000010011",
  30888=>"010000101",
  30889=>"011011001",
  30890=>"010111100",
  30891=>"101111001",
  30892=>"000100101",
  30893=>"010111011",
  30894=>"101000110",
  30895=>"100100001",
  30896=>"011000010",
  30897=>"010110100",
  30898=>"010000001",
  30899=>"010111101",
  30900=>"000110101",
  30901=>"001011110",
  30902=>"011010010",
  30903=>"000111010",
  30904=>"001000111",
  30905=>"111000001",
  30906=>"110011111",
  30907=>"000110111",
  30908=>"111100000",
  30909=>"011001000",
  30910=>"000111010",
  30911=>"101000101",
  30912=>"000010011",
  30913=>"000110011",
  30914=>"110001110",
  30915=>"000011000",
  30916=>"110001000",
  30917=>"111101100",
  30918=>"010001111",
  30919=>"100010010",
  30920=>"000111111",
  30921=>"001000000",
  30922=>"000011011",
  30923=>"101111011",
  30924=>"110101001",
  30925=>"100111110",
  30926=>"010000000",
  30927=>"100111101",
  30928=>"000000100",
  30929=>"011101100",
  30930=>"000110100",
  30931=>"111100111",
  30932=>"010000001",
  30933=>"011010011",
  30934=>"001101110",
  30935=>"101011100",
  30936=>"100000011",
  30937=>"110101101",
  30938=>"010001011",
  30939=>"111110000",
  30940=>"001010011",
  30941=>"001110011",
  30942=>"000000001",
  30943=>"101100000",
  30944=>"010001111",
  30945=>"000110010",
  30946=>"111101010",
  30947=>"110000010",
  30948=>"110011110",
  30949=>"101111001",
  30950=>"110110010",
  30951=>"101111000",
  30952=>"110010101",
  30953=>"000000101",
  30954=>"010000000",
  30955=>"111010010",
  30956=>"110101100",
  30957=>"101000111",
  30958=>"101001100",
  30959=>"001111101",
  30960=>"110110010",
  30961=>"001100100",
  30962=>"101101111",
  30963=>"001011000",
  30964=>"011000000",
  30965=>"011111100",
  30966=>"100000010",
  30967=>"111110101",
  30968=>"111101100",
  30969=>"111001010",
  30970=>"111111101",
  30971=>"011101000",
  30972=>"000010010",
  30973=>"100010101",
  30974=>"000111111",
  30975=>"101100110",
  30976=>"010110101",
  30977=>"011101100",
  30978=>"101011000",
  30979=>"000000000",
  30980=>"000000110",
  30981=>"101001000",
  30982=>"001010101",
  30983=>"101111101",
  30984=>"111000010",
  30985=>"111000011",
  30986=>"001000001",
  30987=>"111110000",
  30988=>"110100010",
  30989=>"111010010",
  30990=>"110010110",
  30991=>"000001101",
  30992=>"111001110",
  30993=>"010010111",
  30994=>"011001110",
  30995=>"111011010",
  30996=>"111111100",
  30997=>"110110001",
  30998=>"110100011",
  30999=>"011000101",
  31000=>"101001101",
  31001=>"101001110",
  31002=>"111001100",
  31003=>"101110000",
  31004=>"010010011",
  31005=>"001111000",
  31006=>"101001001",
  31007=>"010001010",
  31008=>"000101001",
  31009=>"111010110",
  31010=>"110110101",
  31011=>"010110000",
  31012=>"101000000",
  31013=>"010111101",
  31014=>"110000001",
  31015=>"000111000",
  31016=>"001101110",
  31017=>"101101001",
  31018=>"001010001",
  31019=>"101010100",
  31020=>"000110000",
  31021=>"001110101",
  31022=>"110101100",
  31023=>"100011010",
  31024=>"101001100",
  31025=>"111110111",
  31026=>"010111101",
  31027=>"100100001",
  31028=>"000010010",
  31029=>"100011101",
  31030=>"001110110",
  31031=>"011101111",
  31032=>"110101100",
  31033=>"110011101",
  31034=>"101011111",
  31035=>"010100101",
  31036=>"011111110",
  31037=>"011011110",
  31038=>"000111001",
  31039=>"100111101",
  31040=>"000000011",
  31041=>"101111110",
  31042=>"010011000",
  31043=>"110111000",
  31044=>"001000111",
  31045=>"110000110",
  31046=>"000010010",
  31047=>"111110010",
  31048=>"010001100",
  31049=>"011000011",
  31050=>"011101001",
  31051=>"001010000",
  31052=>"010011010",
  31053=>"001011101",
  31054=>"001110010",
  31055=>"000011010",
  31056=>"000010010",
  31057=>"111001000",
  31058=>"010001000",
  31059=>"000110111",
  31060=>"101110100",
  31061=>"111011101",
  31062=>"011100011",
  31063=>"011000111",
  31064=>"101000000",
  31065=>"110100000",
  31066=>"100111110",
  31067=>"101000011",
  31068=>"111111000",
  31069=>"000101100",
  31070=>"111010101",
  31071=>"010100111",
  31072=>"110101010",
  31073=>"010010011",
  31074=>"000011001",
  31075=>"011001001",
  31076=>"101011101",
  31077=>"000011010",
  31078=>"000101000",
  31079=>"010111111",
  31080=>"011110011",
  31081=>"001110111",
  31082=>"110011010",
  31083=>"100010100",
  31084=>"100101100",
  31085=>"101001100",
  31086=>"110100101",
  31087=>"100000100",
  31088=>"010111000",
  31089=>"011100111",
  31090=>"011010011",
  31091=>"111101000",
  31092=>"101000101",
  31093=>"001100111",
  31094=>"011111010",
  31095=>"110010011",
  31096=>"111001110",
  31097=>"010011001",
  31098=>"110010001",
  31099=>"101111101",
  31100=>"111101100",
  31101=>"111110110",
  31102=>"010010100",
  31103=>"110000000",
  31104=>"101010101",
  31105=>"001010010",
  31106=>"101110001",
  31107=>"001100100",
  31108=>"000101000",
  31109=>"111110000",
  31110=>"110101110",
  31111=>"000110011",
  31112=>"110001001",
  31113=>"010011101",
  31114=>"111010001",
  31115=>"101100111",
  31116=>"010000011",
  31117=>"010100111",
  31118=>"111110101",
  31119=>"101110001",
  31120=>"100011100",
  31121=>"110011110",
  31122=>"001001101",
  31123=>"101010101",
  31124=>"110100001",
  31125=>"001100000",
  31126=>"000000000",
  31127=>"000011001",
  31128=>"000010111",
  31129=>"000010000",
  31130=>"001100101",
  31131=>"110101101",
  31132=>"001101111",
  31133=>"000001010",
  31134=>"111110100",
  31135=>"101001100",
  31136=>"011100011",
  31137=>"010010101",
  31138=>"011100010",
  31139=>"000000000",
  31140=>"111101000",
  31141=>"001100111",
  31142=>"100000111",
  31143=>"100011011",
  31144=>"010100001",
  31145=>"110110001",
  31146=>"011011000",
  31147=>"000011010",
  31148=>"100110011",
  31149=>"110001001",
  31150=>"011110100",
  31151=>"011011101",
  31152=>"100100110",
  31153=>"100110010",
  31154=>"000110101",
  31155=>"100011000",
  31156=>"001100000",
  31157=>"110100100",
  31158=>"011001001",
  31159=>"000011001",
  31160=>"010011101",
  31161=>"101001000",
  31162=>"111001011",
  31163=>"111000111",
  31164=>"000001001",
  31165=>"100000101",
  31166=>"000010100",
  31167=>"111111001",
  31168=>"101011101",
  31169=>"010000000",
  31170=>"000001111",
  31171=>"011110100",
  31172=>"010001000",
  31173=>"000010101",
  31174=>"110000101",
  31175=>"101101000",
  31176=>"001011001",
  31177=>"111001100",
  31178=>"010000101",
  31179=>"101101010",
  31180=>"000111100",
  31181=>"100101100",
  31182=>"001011110",
  31183=>"011001001",
  31184=>"010110101",
  31185=>"101101001",
  31186=>"010100000",
  31187=>"001000001",
  31188=>"110000000",
  31189=>"011101001",
  31190=>"111000001",
  31191=>"111101110",
  31192=>"100000001",
  31193=>"111010010",
  31194=>"001010001",
  31195=>"111011010",
  31196=>"110011110",
  31197=>"010100011",
  31198=>"011010010",
  31199=>"101011110",
  31200=>"010001011",
  31201=>"010001110",
  31202=>"001010011",
  31203=>"001011011",
  31204=>"011011001",
  31205=>"111001110",
  31206=>"010000110",
  31207=>"000001101",
  31208=>"011010101",
  31209=>"110000100",
  31210=>"000000010",
  31211=>"001011001",
  31212=>"000001001",
  31213=>"110110101",
  31214=>"011110100",
  31215=>"101011111",
  31216=>"100111101",
  31217=>"000111100",
  31218=>"001011101",
  31219=>"101011010",
  31220=>"000011101",
  31221=>"000001111",
  31222=>"111100010",
  31223=>"101110101",
  31224=>"011111111",
  31225=>"001100111",
  31226=>"110101100",
  31227=>"101111000",
  31228=>"101110111",
  31229=>"000001000",
  31230=>"010111000",
  31231=>"000001010",
  31232=>"011111101",
  31233=>"000101100",
  31234=>"010111111",
  31235=>"000100000",
  31236=>"011000011",
  31237=>"101100011",
  31238=>"111011010",
  31239=>"010100101",
  31240=>"100001100",
  31241=>"001110100",
  31242=>"101100011",
  31243=>"011110000",
  31244=>"001001101",
  31245=>"010001101",
  31246=>"111010110",
  31247=>"000100010",
  31248=>"000100011",
  31249=>"111000000",
  31250=>"001001000",
  31251=>"101000100",
  31252=>"101101111",
  31253=>"011011000",
  31254=>"010011010",
  31255=>"101001110",
  31256=>"101011110",
  31257=>"111001111",
  31258=>"000011001",
  31259=>"110101000",
  31260=>"100011100",
  31261=>"001001111",
  31262=>"111001101",
  31263=>"110011011",
  31264=>"011010100",
  31265=>"110001110",
  31266=>"000001100",
  31267=>"011011101",
  31268=>"111111111",
  31269=>"110100110",
  31270=>"011100100",
  31271=>"000110001",
  31272=>"101110011",
  31273=>"000011000",
  31274=>"101011001",
  31275=>"111111001",
  31276=>"100010100",
  31277=>"101100001",
  31278=>"110101000",
  31279=>"001000001",
  31280=>"101010010",
  31281=>"001000000",
  31282=>"011001100",
  31283=>"111001000",
  31284=>"110110000",
  31285=>"111001101",
  31286=>"111110001",
  31287=>"101010010",
  31288=>"000110010",
  31289=>"111101110",
  31290=>"100010000",
  31291=>"100010010",
  31292=>"110111110",
  31293=>"001001001",
  31294=>"011100110",
  31295=>"001011011",
  31296=>"010111011",
  31297=>"011101110",
  31298=>"111111000",
  31299=>"011011101",
  31300=>"100000000",
  31301=>"100010110",
  31302=>"100001001",
  31303=>"011010001",
  31304=>"001011111",
  31305=>"100111000",
  31306=>"001110100",
  31307=>"100010100",
  31308=>"100011111",
  31309=>"111010010",
  31310=>"000101000",
  31311=>"101101001",
  31312=>"101101010",
  31313=>"110011101",
  31314=>"000101101",
  31315=>"100001110",
  31316=>"001011000",
  31317=>"011000100",
  31318=>"011001011",
  31319=>"011001001",
  31320=>"111001111",
  31321=>"101001110",
  31322=>"011011001",
  31323=>"100100100",
  31324=>"011111110",
  31325=>"000100000",
  31326=>"100100110",
  31327=>"100100001",
  31328=>"001010110",
  31329=>"001010001",
  31330=>"101110111",
  31331=>"101101110",
  31332=>"110111011",
  31333=>"101010011",
  31334=>"001111110",
  31335=>"001100011",
  31336=>"001111101",
  31337=>"101111101",
  31338=>"100111111",
  31339=>"011001100",
  31340=>"100011110",
  31341=>"001011011",
  31342=>"100111010",
  31343=>"100000000",
  31344=>"000011010",
  31345=>"101000011",
  31346=>"000101001",
  31347=>"110110000",
  31348=>"111100110",
  31349=>"011111001",
  31350=>"110001111",
  31351=>"110101100",
  31352=>"100111101",
  31353=>"000001001",
  31354=>"111001100",
  31355=>"110001000",
  31356=>"011100010",
  31357=>"001110100",
  31358=>"110111010",
  31359=>"110011110",
  31360=>"010011110",
  31361=>"111011111",
  31362=>"010111011",
  31363=>"010011101",
  31364=>"111010110",
  31365=>"001110101",
  31366=>"101011111",
  31367=>"011101100",
  31368=>"100001110",
  31369=>"011010111",
  31370=>"100010000",
  31371=>"011111011",
  31372=>"111011100",
  31373=>"100111100",
  31374=>"100001100",
  31375=>"101100100",
  31376=>"010010001",
  31377=>"111110011",
  31378=>"111101111",
  31379=>"001001000",
  31380=>"110110111",
  31381=>"111001100",
  31382=>"110101111",
  31383=>"110110000",
  31384=>"011011010",
  31385=>"010010010",
  31386=>"101110111",
  31387=>"010011100",
  31388=>"110111110",
  31389=>"010011100",
  31390=>"111000000",
  31391=>"000111000",
  31392=>"011001001",
  31393=>"101011101",
  31394=>"000010101",
  31395=>"011101111",
  31396=>"110011011",
  31397=>"011010010",
  31398=>"001110100",
  31399=>"000010001",
  31400=>"111110111",
  31401=>"010001111",
  31402=>"110001010",
  31403=>"111110010",
  31404=>"011111001",
  31405=>"011110001",
  31406=>"011111101",
  31407=>"000000101",
  31408=>"101001100",
  31409=>"111110001",
  31410=>"110110001",
  31411=>"001111110",
  31412=>"000110001",
  31413=>"010001101",
  31414=>"100000000",
  31415=>"111011100",
  31416=>"110000001",
  31417=>"011010010",
  31418=>"000110110",
  31419=>"001000100",
  31420=>"111000000",
  31421=>"010100010",
  31422=>"010011111",
  31423=>"110000110",
  31424=>"001000000",
  31425=>"101100111",
  31426=>"001100001",
  31427=>"011101110",
  31428=>"110000111",
  31429=>"100101000",
  31430=>"000010100",
  31431=>"100100000",
  31432=>"000000011",
  31433=>"001010111",
  31434=>"110001101",
  31435=>"100000111",
  31436=>"100001000",
  31437=>"100010111",
  31438=>"011001010",
  31439=>"111111110",
  31440=>"001101000",
  31441=>"100011111",
  31442=>"101101110",
  31443=>"110101101",
  31444=>"000110010",
  31445=>"010000001",
  31446=>"001110111",
  31447=>"101010101",
  31448=>"011110100",
  31449=>"100001011",
  31450=>"111000111",
  31451=>"110001010",
  31452=>"011001011",
  31453=>"000010111",
  31454=>"110000000",
  31455=>"010110010",
  31456=>"000111000",
  31457=>"000101000",
  31458=>"101111100",
  31459=>"111001110",
  31460=>"010101100",
  31461=>"110010100",
  31462=>"000110000",
  31463=>"010000110",
  31464=>"011000010",
  31465=>"111101101",
  31466=>"000001100",
  31467=>"010101000",
  31468=>"000111101",
  31469=>"001000011",
  31470=>"001010011",
  31471=>"101110110",
  31472=>"001011001",
  31473=>"010001101",
  31474=>"010101110",
  31475=>"011000100",
  31476=>"110010110",
  31477=>"111001101",
  31478=>"011110001",
  31479=>"111001110",
  31480=>"100010100",
  31481=>"010111001",
  31482=>"011001011",
  31483=>"111111011",
  31484=>"001010100",
  31485=>"111011010",
  31486=>"110101001",
  31487=>"001110101",
  31488=>"010100011",
  31489=>"001101101",
  31490=>"111010001",
  31491=>"000001111",
  31492=>"100111001",
  31493=>"100011101",
  31494=>"000110011",
  31495=>"001100100",
  31496=>"101001101",
  31497=>"100001000",
  31498=>"111010100",
  31499=>"111100010",
  31500=>"011001101",
  31501=>"011100101",
  31502=>"101011110",
  31503=>"000011111",
  31504=>"110011001",
  31505=>"000000000",
  31506=>"111001011",
  31507=>"000001011",
  31508=>"110110100",
  31509=>"101100101",
  31510=>"100011110",
  31511=>"101000110",
  31512=>"010101100",
  31513=>"100111010",
  31514=>"010001111",
  31515=>"001000011",
  31516=>"110100001",
  31517=>"001100010",
  31518=>"101100000",
  31519=>"111001000",
  31520=>"010011101",
  31521=>"110000101",
  31522=>"101001111",
  31523=>"111100001",
  31524=>"110111110",
  31525=>"010011000",
  31526=>"001111111",
  31527=>"011111001",
  31528=>"001100010",
  31529=>"011010110",
  31530=>"101111111",
  31531=>"011010110",
  31532=>"010011110",
  31533=>"010001000",
  31534=>"100010000",
  31535=>"010010000",
  31536=>"010001100",
  31537=>"000101011",
  31538=>"011100111",
  31539=>"001110100",
  31540=>"001100110",
  31541=>"111101000",
  31542=>"101010101",
  31543=>"000110101",
  31544=>"100000111",
  31545=>"101111100",
  31546=>"101111010",
  31547=>"001000100",
  31548=>"100110110",
  31549=>"101100001",
  31550=>"001111111",
  31551=>"101001011",
  31552=>"000010000",
  31553=>"100101010",
  31554=>"111001000",
  31555=>"011111100",
  31556=>"110001100",
  31557=>"010000011",
  31558=>"001000010",
  31559=>"110111110",
  31560=>"000001110",
  31561=>"011111110",
  31562=>"101010001",
  31563=>"101010000",
  31564=>"100101111",
  31565=>"011011010",
  31566=>"110101011",
  31567=>"101111000",
  31568=>"010110100",
  31569=>"000110001",
  31570=>"110100101",
  31571=>"001000001",
  31572=>"010000110",
  31573=>"111010101",
  31574=>"110011101",
  31575=>"010001001",
  31576=>"011011000",
  31577=>"111001111",
  31578=>"001011010",
  31579=>"010000111",
  31580=>"011101101",
  31581=>"010101111",
  31582=>"010011101",
  31583=>"010100100",
  31584=>"110000111",
  31585=>"100011001",
  31586=>"001001101",
  31587=>"111011100",
  31588=>"110001010",
  31589=>"011001110",
  31590=>"000001100",
  31591=>"111110010",
  31592=>"001101010",
  31593=>"001110010",
  31594=>"111100001",
  31595=>"001110111",
  31596=>"100110110",
  31597=>"010101000",
  31598=>"100110111",
  31599=>"100011111",
  31600=>"000001001",
  31601=>"110100110",
  31602=>"111110010",
  31603=>"101101110",
  31604=>"101010001",
  31605=>"001100001",
  31606=>"100101010",
  31607=>"001111101",
  31608=>"001100101",
  31609=>"111001100",
  31610=>"011100000",
  31611=>"010101001",
  31612=>"111001110",
  31613=>"110001110",
  31614=>"000000100",
  31615=>"000011000",
  31616=>"100111111",
  31617=>"111111000",
  31618=>"000111100",
  31619=>"100110110",
  31620=>"110010011",
  31621=>"110101111",
  31622=>"010100000",
  31623=>"100011000",
  31624=>"100111110",
  31625=>"001000011",
  31626=>"100010000",
  31627=>"110000010",
  31628=>"001000010",
  31629=>"101111111",
  31630=>"101110101",
  31631=>"100111111",
  31632=>"010110000",
  31633=>"110110000",
  31634=>"100001000",
  31635=>"010110011",
  31636=>"111011110",
  31637=>"011101100",
  31638=>"011110111",
  31639=>"100100101",
  31640=>"010011101",
  31641=>"010101000",
  31642=>"011010000",
  31643=>"101100111",
  31644=>"000010110",
  31645=>"100000111",
  31646=>"001011101",
  31647=>"101110111",
  31648=>"100011101",
  31649=>"010111001",
  31650=>"110111000",
  31651=>"001000110",
  31652=>"001000110",
  31653=>"100011111",
  31654=>"100011010",
  31655=>"111110000",
  31656=>"001000011",
  31657=>"100001010",
  31658=>"010011111",
  31659=>"111001011",
  31660=>"000101101",
  31661=>"011011010",
  31662=>"011111111",
  31663=>"111110111",
  31664=>"001011011",
  31665=>"111110111",
  31666=>"010010101",
  31667=>"011100111",
  31668=>"110011101",
  31669=>"111110011",
  31670=>"011001010",
  31671=>"010100101",
  31672=>"101111010",
  31673=>"010000000",
  31674=>"100011001",
  31675=>"100000010",
  31676=>"011101101",
  31677=>"000001000",
  31678=>"100111101",
  31679=>"000010011",
  31680=>"101000111",
  31681=>"000110011",
  31682=>"101000110",
  31683=>"110100101",
  31684=>"111001011",
  31685=>"110011110",
  31686=>"000001110",
  31687=>"010000010",
  31688=>"100010111",
  31689=>"010101111",
  31690=>"101011100",
  31691=>"100000000",
  31692=>"001001101",
  31693=>"100111001",
  31694=>"011010000",
  31695=>"111101100",
  31696=>"001011101",
  31697=>"111001000",
  31698=>"111110100",
  31699=>"011101011",
  31700=>"100011001",
  31701=>"010000001",
  31702=>"011101110",
  31703=>"001001011",
  31704=>"100100011",
  31705=>"011101100",
  31706=>"010000101",
  31707=>"100000100",
  31708=>"100011000",
  31709=>"011100111",
  31710=>"101011100",
  31711=>"000101110",
  31712=>"111001101",
  31713=>"000001011",
  31714=>"000010100",
  31715=>"001001001",
  31716=>"000000110",
  31717=>"111001111",
  31718=>"111000100",
  31719=>"111001011",
  31720=>"111101111",
  31721=>"011111011",
  31722=>"110001100",
  31723=>"111100001",
  31724=>"100000001",
  31725=>"111001101",
  31726=>"010111000",
  31727=>"110100101",
  31728=>"011110100",
  31729=>"011001010",
  31730=>"001011100",
  31731=>"001100100",
  31732=>"011100001",
  31733=>"110011000",
  31734=>"001100000",
  31735=>"000100011",
  31736=>"110111110",
  31737=>"001111100",
  31738=>"111001101",
  31739=>"010010000",
  31740=>"110000100",
  31741=>"111110011",
  31742=>"111000101",
  31743=>"101001000",
  31744=>"100110001",
  31745=>"101011111",
  31746=>"100101111",
  31747=>"001111010",
  31748=>"001010011",
  31749=>"111100101",
  31750=>"010101101",
  31751=>"100010100",
  31752=>"011100111",
  31753=>"111110111",
  31754=>"001001000",
  31755=>"001000101",
  31756=>"110111001",
  31757=>"100001011",
  31758=>"110110111",
  31759=>"111011111",
  31760=>"100111101",
  31761=>"101100101",
  31762=>"011111101",
  31763=>"010010100",
  31764=>"001011011",
  31765=>"010011010",
  31766=>"000000110",
  31767=>"010101100",
  31768=>"100111011",
  31769=>"100111011",
  31770=>"000011100",
  31771=>"001110110",
  31772=>"011100011",
  31773=>"011011111",
  31774=>"010000010",
  31775=>"000010010",
  31776=>"000100101",
  31777=>"110000010",
  31778=>"100101010",
  31779=>"010100010",
  31780=>"011001110",
  31781=>"101001010",
  31782=>"001100101",
  31783=>"101011010",
  31784=>"101100111",
  31785=>"000100110",
  31786=>"010011011",
  31787=>"111111110",
  31788=>"101110010",
  31789=>"110011000",
  31790=>"001011100",
  31791=>"111010000",
  31792=>"010001000",
  31793=>"001001011",
  31794=>"110000000",
  31795=>"101110100",
  31796=>"011100010",
  31797=>"011010000",
  31798=>"001110001",
  31799=>"100110100",
  31800=>"011001111",
  31801=>"000111001",
  31802=>"100100101",
  31803=>"100001100",
  31804=>"101111000",
  31805=>"011100000",
  31806=>"000010001",
  31807=>"010111100",
  31808=>"010101000",
  31809=>"000100100",
  31810=>"111001010",
  31811=>"100011000",
  31812=>"010100011",
  31813=>"111001101",
  31814=>"110110100",
  31815=>"101001011",
  31816=>"001100111",
  31817=>"000100001",
  31818=>"100000110",
  31819=>"000001111",
  31820=>"010111011",
  31821=>"010011000",
  31822=>"111001110",
  31823=>"110011110",
  31824=>"001101011",
  31825=>"111001110",
  31826=>"111000010",
  31827=>"100101111",
  31828=>"110111010",
  31829=>"110110111",
  31830=>"110000100",
  31831=>"000111100",
  31832=>"100011110",
  31833=>"000001010",
  31834=>"100000100",
  31835=>"000010100",
  31836=>"010000001",
  31837=>"011000000",
  31838=>"001001011",
  31839=>"101000111",
  31840=>"000011000",
  31841=>"011100000",
  31842=>"010110101",
  31843=>"010000011",
  31844=>"010010000",
  31845=>"000110110",
  31846=>"010110011",
  31847=>"000001111",
  31848=>"111001100",
  31849=>"101000000",
  31850=>"000111001",
  31851=>"110010011",
  31852=>"111011010",
  31853=>"110001000",
  31854=>"101101110",
  31855=>"010011010",
  31856=>"001010011",
  31857=>"100010010",
  31858=>"101011011",
  31859=>"011111000",
  31860=>"000001011",
  31861=>"100111100",
  31862=>"110101011",
  31863=>"101010111",
  31864=>"011001001",
  31865=>"111000010",
  31866=>"010110101",
  31867=>"011100111",
  31868=>"010110011",
  31869=>"111010011",
  31870=>"111011100",
  31871=>"011001110",
  31872=>"001101001",
  31873=>"011000001",
  31874=>"100010101",
  31875=>"010101100",
  31876=>"001010100",
  31877=>"000001110",
  31878=>"110110000",
  31879=>"101011110",
  31880=>"001110011",
  31881=>"100101011",
  31882=>"010111010",
  31883=>"111000000",
  31884=>"101000110",
  31885=>"001001100",
  31886=>"000000110",
  31887=>"001011001",
  31888=>"011001000",
  31889=>"100001001",
  31890=>"101011000",
  31891=>"101001011",
  31892=>"010110100",
  31893=>"111101001",
  31894=>"111101000",
  31895=>"111111101",
  31896=>"111000101",
  31897=>"101101011",
  31898=>"010010101",
  31899=>"001001100",
  31900=>"000101111",
  31901=>"111001100",
  31902=>"101111011",
  31903=>"110110001",
  31904=>"101110000",
  31905=>"011011001",
  31906=>"000001100",
  31907=>"001001100",
  31908=>"010010000",
  31909=>"000111001",
  31910=>"111010110",
  31911=>"011110001",
  31912=>"011011111",
  31913=>"011011011",
  31914=>"001110000",
  31915=>"111100110",
  31916=>"100010001",
  31917=>"000111001",
  31918=>"110010111",
  31919=>"000111101",
  31920=>"000011100",
  31921=>"101010100",
  31922=>"000111001",
  31923=>"101100110",
  31924=>"011101111",
  31925=>"000000100",
  31926=>"101000010",
  31927=>"101111100",
  31928=>"001001011",
  31929=>"100000001",
  31930=>"100111110",
  31931=>"101111100",
  31932=>"011001111",
  31933=>"111011111",
  31934=>"000011111",
  31935=>"000111010",
  31936=>"101111011",
  31937=>"000100000",
  31938=>"011110001",
  31939=>"011011001",
  31940=>"000101101",
  31941=>"011100101",
  31942=>"101011000",
  31943=>"100000110",
  31944=>"111010100",
  31945=>"010000011",
  31946=>"100000001",
  31947=>"011000110",
  31948=>"010110000",
  31949=>"000010011",
  31950=>"000101010",
  31951=>"101000001",
  31952=>"101111011",
  31953=>"111101000",
  31954=>"000101000",
  31955=>"011101010",
  31956=>"111101000",
  31957=>"000111111",
  31958=>"000101011",
  31959=>"111011101",
  31960=>"100100010",
  31961=>"101111101",
  31962=>"001000111",
  31963=>"001100101",
  31964=>"001000011",
  31965=>"111100001",
  31966=>"111110111",
  31967=>"001110001",
  31968=>"001000000",
  31969=>"010110100",
  31970=>"011111100",
  31971=>"100000101",
  31972=>"110101001",
  31973=>"000111110",
  31974=>"000100111",
  31975=>"000010011",
  31976=>"010100110",
  31977=>"001001111",
  31978=>"010110100",
  31979=>"101011001",
  31980=>"111100010",
  31981=>"010010111",
  31982=>"000000011",
  31983=>"101111011",
  31984=>"001100010",
  31985=>"001000000",
  31986=>"101100100",
  31987=>"001010011",
  31988=>"000100110",
  31989=>"101101100",
  31990=>"110101101",
  31991=>"100010001",
  31992=>"101010000",
  31993=>"101101101",
  31994=>"111100011",
  31995=>"000010010",
  31996=>"001111111",
  31997=>"101011010",
  31998=>"011000111",
  31999=>"111100010",
  32000=>"100100110",
  32001=>"011111010",
  32002=>"111111100",
  32003=>"101100100",
  32004=>"111000010",
  32005=>"110101100",
  32006=>"010001001",
  32007=>"110011010",
  32008=>"110111110",
  32009=>"110100001",
  32010=>"010011000",
  32011=>"100000001",
  32012=>"110001100",
  32013=>"110110001",
  32014=>"100000000",
  32015=>"000111010",
  32016=>"100100001",
  32017=>"001000000",
  32018=>"100010110",
  32019=>"000111111",
  32020=>"100100010",
  32021=>"111110010",
  32022=>"011100000",
  32023=>"001000011",
  32024=>"110000101",
  32025=>"001011011",
  32026=>"010011001",
  32027=>"011001001",
  32028=>"011011000",
  32029=>"000010111",
  32030=>"001010111",
  32031=>"010001101",
  32032=>"111000001",
  32033=>"110001000",
  32034=>"100000110",
  32035=>"100001001",
  32036=>"010000111",
  32037=>"001011111",
  32038=>"011001010",
  32039=>"010010000",
  32040=>"100010011",
  32041=>"001100010",
  32042=>"111000101",
  32043=>"110001100",
  32044=>"010111101",
  32045=>"001100000",
  32046=>"111011011",
  32047=>"010110111",
  32048=>"111011110",
  32049=>"001110110",
  32050=>"001011100",
  32051=>"101010001",
  32052=>"000001100",
  32053=>"011001000",
  32054=>"100101111",
  32055=>"111111000",
  32056=>"100000000",
  32057=>"000001001",
  32058=>"111110000",
  32059=>"001001111",
  32060=>"000101101",
  32061=>"000011101",
  32062=>"001100010",
  32063=>"010110011",
  32064=>"101111111",
  32065=>"111101011",
  32066=>"001000001",
  32067=>"000001000",
  32068=>"000001110",
  32069=>"011010011",
  32070=>"110011100",
  32071=>"000001101",
  32072=>"110100101",
  32073=>"101000101",
  32074=>"101000111",
  32075=>"001001111",
  32076=>"010000101",
  32077=>"100110110",
  32078=>"100011001",
  32079=>"111100001",
  32080=>"100010010",
  32081=>"000001110",
  32082=>"010110100",
  32083=>"101100101",
  32084=>"001110101",
  32085=>"010000011",
  32086=>"011100100",
  32087=>"101100001",
  32088=>"010111010",
  32089=>"000011110",
  32090=>"111111100",
  32091=>"100100100",
  32092=>"100100101",
  32093=>"001110011",
  32094=>"001000100",
  32095=>"111111000",
  32096=>"001010010",
  32097=>"111010001",
  32098=>"001111010",
  32099=>"001100110",
  32100=>"111101111",
  32101=>"010110100",
  32102=>"010101011",
  32103=>"000100111",
  32104=>"010010011",
  32105=>"001001111",
  32106=>"000111010",
  32107=>"110001100",
  32108=>"011111000",
  32109=>"011110010",
  32110=>"011111011",
  32111=>"110011000",
  32112=>"111110110",
  32113=>"101001100",
  32114=>"111000010",
  32115=>"110010110",
  32116=>"001001000",
  32117=>"000010001",
  32118=>"110110011",
  32119=>"010001011",
  32120=>"011000101",
  32121=>"110001100",
  32122=>"100011011",
  32123=>"101000000",
  32124=>"011011010",
  32125=>"100101000",
  32126=>"110100111",
  32127=>"101001000",
  32128=>"000011111",
  32129=>"110010011",
  32130=>"001101011",
  32131=>"000000011",
  32132=>"000000100",
  32133=>"111100011",
  32134=>"000001001",
  32135=>"000110000",
  32136=>"111011001",
  32137=>"110111111",
  32138=>"111000000",
  32139=>"000000011",
  32140=>"101100010",
  32141=>"111011000",
  32142=>"001110000",
  32143=>"000100110",
  32144=>"001111101",
  32145=>"101101101",
  32146=>"101011010",
  32147=>"111000111",
  32148=>"000010001",
  32149=>"000101101",
  32150=>"110100110",
  32151=>"111001001",
  32152=>"110010111",
  32153=>"011101111",
  32154=>"010101011",
  32155=>"001101001",
  32156=>"001100101",
  32157=>"111010000",
  32158=>"100110110",
  32159=>"011001000",
  32160=>"110011111",
  32161=>"100011010",
  32162=>"000111110",
  32163=>"000100001",
  32164=>"000101101",
  32165=>"100011010",
  32166=>"000001110",
  32167=>"101100101",
  32168=>"001110010",
  32169=>"001100010",
  32170=>"100000001",
  32171=>"011011110",
  32172=>"010010001",
  32173=>"110011010",
  32174=>"100101111",
  32175=>"000100010",
  32176=>"101011100",
  32177=>"100100111",
  32178=>"000101010",
  32179=>"000010000",
  32180=>"011001000",
  32181=>"110100101",
  32182=>"000010110",
  32183=>"010110001",
  32184=>"011111001",
  32185=>"110001110",
  32186=>"011000100",
  32187=>"101000000",
  32188=>"110100100",
  32189=>"010000000",
  32190=>"101011011",
  32191=>"110111000",
  32192=>"001100000",
  32193=>"001001101",
  32194=>"110100001",
  32195=>"010010111",
  32196=>"001110110",
  32197=>"111100111",
  32198=>"101010110",
  32199=>"010100100",
  32200=>"100011101",
  32201=>"111010001",
  32202=>"101000000",
  32203=>"010111010",
  32204=>"010010010",
  32205=>"101011011",
  32206=>"011001010",
  32207=>"001000110",
  32208=>"010000110",
  32209=>"110011111",
  32210=>"101011110",
  32211=>"100010110",
  32212=>"010010001",
  32213=>"001010011",
  32214=>"010111110",
  32215=>"111010001",
  32216=>"011011100",
  32217=>"000101110",
  32218=>"100100101",
  32219=>"001100000",
  32220=>"000111101",
  32221=>"101010110",
  32222=>"111010010",
  32223=>"101100011",
  32224=>"011001001",
  32225=>"111010110",
  32226=>"011011000",
  32227=>"000111000",
  32228=>"011010101",
  32229=>"111101111",
  32230=>"110111001",
  32231=>"110101001",
  32232=>"101111011",
  32233=>"010010111",
  32234=>"010110111",
  32235=>"101011011",
  32236=>"000101001",
  32237=>"010000000",
  32238=>"111010000",
  32239=>"011111010",
  32240=>"000110111",
  32241=>"000010000",
  32242=>"001101001",
  32243=>"010010110",
  32244=>"101001011",
  32245=>"111000111",
  32246=>"100111010",
  32247=>"111101000",
  32248=>"011111111",
  32249=>"101101110",
  32250=>"010111001",
  32251=>"011011100",
  32252=>"011011100",
  32253=>"111000001",
  32254=>"111010010",
  32255=>"010000101",
  32256=>"101101001",
  32257=>"100001011",
  32258=>"100101001",
  32259=>"000110111",
  32260=>"011010101",
  32261=>"010100001",
  32262=>"000000000",
  32263=>"110101000",
  32264=>"111000100",
  32265=>"001011010",
  32266=>"000100010",
  32267=>"001011000",
  32268=>"010111110",
  32269=>"001111011",
  32270=>"101101111",
  32271=>"111101010",
  32272=>"000010100",
  32273=>"001001010",
  32274=>"111101001",
  32275=>"101000001",
  32276=>"110011101",
  32277=>"101101111",
  32278=>"000110110",
  32279=>"101111110",
  32280=>"010111111",
  32281=>"001100001",
  32282=>"001111101",
  32283=>"001011111",
  32284=>"000010011",
  32285=>"010100110",
  32286=>"101101011",
  32287=>"100111110",
  32288=>"011010110",
  32289=>"100010001",
  32290=>"000101110",
  32291=>"001011110",
  32292=>"000100100",
  32293=>"110111001",
  32294=>"100001010",
  32295=>"100010001",
  32296=>"111111001",
  32297=>"110000010",
  32298=>"010111100",
  32299=>"111010010",
  32300=>"010100101",
  32301=>"110000010",
  32302=>"010110111",
  32303=>"000101001",
  32304=>"010110010",
  32305=>"001001110",
  32306=>"001110111",
  32307=>"111110011",
  32308=>"011100111",
  32309=>"011110000",
  32310=>"001101011",
  32311=>"100000000",
  32312=>"001100011",
  32313=>"010110010",
  32314=>"010100011",
  32315=>"001000001",
  32316=>"000010000",
  32317=>"101010111",
  32318=>"111111110",
  32319=>"100000111",
  32320=>"111100111",
  32321=>"001010100",
  32322=>"011010010",
  32323=>"011101100",
  32324=>"001000110",
  32325=>"011100010",
  32326=>"110011110",
  32327=>"000100110",
  32328=>"101111000",
  32329=>"011000000",
  32330=>"001010101",
  32331=>"000001010",
  32332=>"111100111",
  32333=>"010011000",
  32334=>"011100000",
  32335=>"010010010",
  32336=>"111111111",
  32337=>"100110110",
  32338=>"101100100",
  32339=>"001100010",
  32340=>"100011011",
  32341=>"000100101",
  32342=>"000011101",
  32343=>"010011011",
  32344=>"000110100",
  32345=>"101100111",
  32346=>"000000011",
  32347=>"010100001",
  32348=>"010111001",
  32349=>"000000001",
  32350=>"110010000",
  32351=>"100111001",
  32352=>"111111101",
  32353=>"010001010",
  32354=>"001000101",
  32355=>"000001000",
  32356=>"001100111",
  32357=>"000000101",
  32358=>"011100100",
  32359=>"111100111",
  32360=>"000000101",
  32361=>"011011011",
  32362=>"111111010",
  32363=>"111011110",
  32364=>"110100101",
  32365=>"011100100",
  32366=>"011011110",
  32367=>"100100100",
  32368=>"110110010",
  32369=>"001100110",
  32370=>"011100001",
  32371=>"000001101",
  32372=>"011101010",
  32373=>"010011010",
  32374=>"110100100",
  32375=>"101111000",
  32376=>"010111101",
  32377=>"101100111",
  32378=>"011101100",
  32379=>"100000000",
  32380=>"000011110",
  32381=>"101011101",
  32382=>"101000101",
  32383=>"110010110",
  32384=>"001000000",
  32385=>"100100110",
  32386=>"000100100",
  32387=>"000101101",
  32388=>"010011000",
  32389=>"101000010",
  32390=>"111010101",
  32391=>"011010001",
  32392=>"010000101",
  32393=>"101011000",
  32394=>"010100000",
  32395=>"100101000",
  32396=>"100101010",
  32397=>"111110011",
  32398=>"011010111",
  32399=>"000011100",
  32400=>"111111110",
  32401=>"111001011",
  32402=>"000110000",
  32403=>"011001000",
  32404=>"111100011",
  32405=>"011100001",
  32406=>"101011000",
  32407=>"110000101",
  32408=>"010100110",
  32409=>"100111101",
  32410=>"100101000",
  32411=>"001101001",
  32412=>"001001111",
  32413=>"011100110",
  32414=>"101101111",
  32415=>"100000010",
  32416=>"011110101",
  32417=>"101001011",
  32418=>"101101111",
  32419=>"010100000",
  32420=>"111010111",
  32421=>"000000010",
  32422=>"110010110",
  32423=>"110101011",
  32424=>"000111001",
  32425=>"000100100",
  32426=>"000010000",
  32427=>"010101001",
  32428=>"101011111",
  32429=>"010011110",
  32430=>"001111111",
  32431=>"011011111",
  32432=>"010011101",
  32433=>"001101111",
  32434=>"111100001",
  32435=>"011111111",
  32436=>"010100010",
  32437=>"000001010",
  32438=>"111111111",
  32439=>"011001011",
  32440=>"101101011",
  32441=>"010010100",
  32442=>"011001101",
  32443=>"111100111",
  32444=>"100000111",
  32445=>"000011110",
  32446=>"010010010",
  32447=>"110010101",
  32448=>"110111010",
  32449=>"011001110",
  32450=>"100011100",
  32451=>"110010110",
  32452=>"010010010",
  32453=>"010010000",
  32454=>"011101011",
  32455=>"000001110",
  32456=>"110000001",
  32457=>"111011111",
  32458=>"010110101",
  32459=>"100010010",
  32460=>"101100100",
  32461=>"111000100",
  32462=>"111111110",
  32463=>"100111001",
  32464=>"110101001",
  32465=>"111011000",
  32466=>"010110111",
  32467=>"100011010",
  32468=>"000111110",
  32469=>"001111100",
  32470=>"001111101",
  32471=>"100110010",
  32472=>"000111011",
  32473=>"011010011",
  32474=>"011011000",
  32475=>"101101111",
  32476=>"001110111",
  32477=>"101010000",
  32478=>"111000100",
  32479=>"110011100",
  32480=>"000110001",
  32481=>"100000000",
  32482=>"001110100",
  32483=>"101101100",
  32484=>"000011100",
  32485=>"010011101",
  32486=>"000111000",
  32487=>"001001101",
  32488=>"110111001",
  32489=>"010010100",
  32490=>"011101110",
  32491=>"100000010",
  32492=>"000110110",
  32493=>"001001111",
  32494=>"110101011",
  32495=>"001000111",
  32496=>"111011001",
  32497=>"101100011",
  32498=>"111101001",
  32499=>"101011101",
  32500=>"101000110",
  32501=>"001001111",
  32502=>"111111001",
  32503=>"101000010",
  32504=>"010010000",
  32505=>"000011100",
  32506=>"011111111",
  32507=>"010001001",
  32508=>"001111111",
  32509=>"001110011",
  32510=>"100101101",
  32511=>"100011001",
  32512=>"000110011",
  32513=>"111011000",
  32514=>"000010000",
  32515=>"010111111",
  32516=>"010001111",
  32517=>"010110100",
  32518=>"101100100",
  32519=>"010110111",
  32520=>"100000110",
  32521=>"110101110",
  32522=>"110001101",
  32523=>"000111011",
  32524=>"101110000",
  32525=>"100101100",
  32526=>"010010010",
  32527=>"101110110",
  32528=>"011001000",
  32529=>"010001001",
  32530=>"010001010",
  32531=>"111111110",
  32532=>"110110101",
  32533=>"111111000",
  32534=>"111100100",
  32535=>"101111011",
  32536=>"000101101",
  32537=>"101111010",
  32538=>"100001100",
  32539=>"110111110",
  32540=>"110000010",
  32541=>"110000001",
  32542=>"001100111",
  32543=>"010000000",
  32544=>"110011110",
  32545=>"101011000",
  32546=>"100000100",
  32547=>"110111111",
  32548=>"010001101",
  32549=>"110100101",
  32550=>"011000011",
  32551=>"011010110",
  32552=>"010101110",
  32553=>"111110111",
  32554=>"100100111",
  32555=>"001000101",
  32556=>"100101000",
  32557=>"110110110",
  32558=>"100101111",
  32559=>"010010000",
  32560=>"110000111",
  32561=>"011111100",
  32562=>"010011010",
  32563=>"001101000",
  32564=>"101100011",
  32565=>"011001001",
  32566=>"000111110",
  32567=>"001101010",
  32568=>"001000001",
  32569=>"111001111",
  32570=>"101010100",
  32571=>"100110110",
  32572=>"011101101",
  32573=>"001110101",
  32574=>"110100000",
  32575=>"000110111",
  32576=>"010010000",
  32577=>"010011010",
  32578=>"010110001",
  32579=>"000000011",
  32580=>"010000001",
  32581=>"000110010",
  32582=>"011111010",
  32583=>"001001111",
  32584=>"000001100",
  32585=>"001000100",
  32586=>"010000001",
  32587=>"100101000",
  32588=>"100100111",
  32589=>"101000010",
  32590=>"011010111",
  32591=>"111100100",
  32592=>"010110111",
  32593=>"100010001",
  32594=>"101110011",
  32595=>"001010111",
  32596=>"101111000",
  32597=>"000011110",
  32598=>"001110001",
  32599=>"110111011",
  32600=>"011111011",
  32601=>"110011100",
  32602=>"110110100",
  32603=>"010111001",
  32604=>"011000001",
  32605=>"100100111",
  32606=>"110001110",
  32607=>"101000111",
  32608=>"111110010",
  32609=>"011011011",
  32610=>"000111100",
  32611=>"011011000",
  32612=>"010011000",
  32613=>"101010011",
  32614=>"000101111",
  32615=>"000111001",
  32616=>"100000000",
  32617=>"001110101",
  32618=>"010111010",
  32619=>"011110111",
  32620=>"001110100",
  32621=>"011100000",
  32622=>"100000101",
  32623=>"101010001",
  32624=>"000101100",
  32625=>"111101010",
  32626=>"000100101",
  32627=>"000010101",
  32628=>"011100010",
  32629=>"011010010",
  32630=>"101111000",
  32631=>"111100111",
  32632=>"010110110",
  32633=>"100000000",
  32634=>"100011001",
  32635=>"011101010",
  32636=>"000100010",
  32637=>"000111111",
  32638=>"100101001",
  32639=>"101010011",
  32640=>"000110000",
  32641=>"100001010",
  32642=>"000011111",
  32643=>"010001101",
  32644=>"000001000",
  32645=>"010001101",
  32646=>"100100010",
  32647=>"010101001",
  32648=>"000100101",
  32649=>"011010000",
  32650=>"110011111",
  32651=>"000000110",
  32652=>"010100101",
  32653=>"111110111",
  32654=>"000001100",
  32655=>"000101111",
  32656=>"001111011",
  32657=>"100111011",
  32658=>"100110111",
  32659=>"110011011",
  32660=>"101010000",
  32661=>"001100110",
  32662=>"010001000",
  32663=>"110010000",
  32664=>"010111110",
  32665=>"010011110",
  32666=>"011101110",
  32667=>"011101000",
  32668=>"010010000",
  32669=>"011010001",
  32670=>"100110001",
  32671=>"100000101",
  32672=>"110111000",
  32673=>"101100111",
  32674=>"110011111",
  32675=>"100100111",
  32676=>"100010000",
  32677=>"101001000",
  32678=>"011010100",
  32679=>"100100100",
  32680=>"010000000",
  32681=>"001101000",
  32682=>"111110100",
  32683=>"001001110",
  32684=>"010101111",
  32685=>"101111110",
  32686=>"110101001",
  32687=>"000001101",
  32688=>"011100100",
  32689=>"011111001",
  32690=>"000000001",
  32691=>"101011111",
  32692=>"101011001",
  32693=>"100100001",
  32694=>"010010011",
  32695=>"010010111",
  32696=>"011010110",
  32697=>"111110100",
  32698=>"110010011",
  32699=>"011100100",
  32700=>"011010000",
  32701=>"100011110",
  32702=>"111011011",
  32703=>"000110001",
  32704=>"110101100",
  32705=>"111101100",
  32706=>"000011010",
  32707=>"010001011",
  32708=>"101010000",
  32709=>"101010010",
  32710=>"110001000",
  32711=>"111110011",
  32712=>"110000011",
  32713=>"010110111",
  32714=>"111110000",
  32715=>"111101010",
  32716=>"000010011",
  32717=>"010011110",
  32718=>"010011000",
  32719=>"001010100",
  32720=>"010101000",
  32721=>"101001010",
  32722=>"111011111",
  32723=>"001010000",
  32724=>"101010111",
  32725=>"111111011",
  32726=>"010111110",
  32727=>"000100000",
  32728=>"001000111",
  32729=>"101000101",
  32730=>"011111010",
  32731=>"000110001",
  32732=>"011001010",
  32733=>"100000001",
  32734=>"100011110",
  32735=>"110110001",
  32736=>"000010110",
  32737=>"101000101",
  32738=>"000100110",
  32739=>"100001110",
  32740=>"100000011",
  32741=>"011111111",
  32742=>"101101110",
  32743=>"001100110",
  32744=>"010011111",
  32745=>"101011110",
  32746=>"111111111",
  32747=>"000110010",
  32748=>"101110001",
  32749=>"111110100",
  32750=>"011100011",
  32751=>"111110111",
  32752=>"110111000",
  32753=>"101001001",
  32754=>"011111101",
  32755=>"100110111",
  32756=>"000000111",
  32757=>"100101101",
  32758=>"011010100",
  32759=>"011101000",
  32760=>"110100111",
  32761=>"111011001",
  32762=>"011010001",
  32763=>"011011100",
  32764=>"111010010",
  32765=>"000100111",
  32766=>"010100001",
  32767=>"000010001",
  32768=>"111111000",
  32769=>"011111011",
  32770=>"100000100",
  32771=>"100101011",
  32772=>"100101101",
  32773=>"011101010",
  32774=>"011000100",
  32775=>"000000001",
  32776=>"110011010",
  32777=>"001001010",
  32778=>"010100011",
  32779=>"110100110",
  32780=>"011011001",
  32781=>"001000000",
  32782=>"000110100",
  32783=>"101001000",
  32784=>"111111010",
  32785=>"010000000",
  32786=>"010100110",
  32787=>"010111000",
  32788=>"011001001",
  32789=>"101110001",
  32790=>"111100010",
  32791=>"100000000",
  32792=>"100001010",
  32793=>"111110001",
  32794=>"110101001",
  32795=>"110011101",
  32796=>"000100111",
  32797=>"100010110",
  32798=>"001001100",
  32799=>"010001111",
  32800=>"100001011",
  32801=>"010101111",
  32802=>"011011011",
  32803=>"101100011",
  32804=>"010100011",
  32805=>"101111101",
  32806=>"001001111",
  32807=>"101000100",
  32808=>"001101111",
  32809=>"000001000",
  32810=>"000001110",
  32811=>"000010000",
  32812=>"010100001",
  32813=>"111111011",
  32814=>"110101001",
  32815=>"010100000",
  32816=>"111001110",
  32817=>"001011111",
  32818=>"011001001",
  32819=>"001000010",
  32820=>"110001011",
  32821=>"100111110",
  32822=>"000000111",
  32823=>"001101001",
  32824=>"100001010",
  32825=>"000010111",
  32826=>"111111111",
  32827=>"100101001",
  32828=>"111011110",
  32829=>"010111011",
  32830=>"110101111",
  32831=>"011011100",
  32832=>"111111100",
  32833=>"000110000",
  32834=>"100010011",
  32835=>"101011100",
  32836=>"100000001",
  32837=>"010101110",
  32838=>"111111010",
  32839=>"111001100",
  32840=>"110001110",
  32841=>"010000000",
  32842=>"111110011",
  32843=>"101101011",
  32844=>"010011010",
  32845=>"101110101",
  32846=>"011111111",
  32847=>"011100100",
  32848=>"100000100",
  32849=>"011100111",
  32850=>"001011101",
  32851=>"100011101",
  32852=>"010010010",
  32853=>"001110011",
  32854=>"010010000",
  32855=>"000110110",
  32856=>"100110101",
  32857=>"001110010",
  32858=>"010001101",
  32859=>"111110101",
  32860=>"001100101",
  32861=>"011011100",
  32862=>"010000011",
  32863=>"010011110",
  32864=>"001010101",
  32865=>"011101111",
  32866=>"111100000",
  32867=>"000001001",
  32868=>"001001010",
  32869=>"111111001",
  32870=>"111011001",
  32871=>"000110010",
  32872=>"010011000",
  32873=>"110000101",
  32874=>"011010011",
  32875=>"100010100",
  32876=>"001010010",
  32877=>"011001001",
  32878=>"011111010",
  32879=>"000100000",
  32880=>"000000001",
  32881=>"011011100",
  32882=>"011100011",
  32883=>"111011001",
  32884=>"010001001",
  32885=>"100111111",
  32886=>"110001111",
  32887=>"011001111",
  32888=>"110010011",
  32889=>"100101100",
  32890=>"101011000",
  32891=>"110110011",
  32892=>"001001110",
  32893=>"010101110",
  32894=>"110000001",
  32895=>"101111000",
  32896=>"011000101",
  32897=>"100101000",
  32898=>"010011100",
  32899=>"101110001",
  32900=>"110101101",
  32901=>"000010111",
  32902=>"010101010",
  32903=>"100000110",
  32904=>"011101001",
  32905=>"000000010",
  32906=>"010001001",
  32907=>"111010010",
  32908=>"001010111",
  32909=>"100010011",
  32910=>"001101101",
  32911=>"011001010",
  32912=>"000011010",
  32913=>"101000000",
  32914=>"001101100",
  32915=>"011101100",
  32916=>"110110111",
  32917=>"010100110",
  32918=>"011111011",
  32919=>"000100100",
  32920=>"010000010",
  32921=>"110101010",
  32922=>"111111101",
  32923=>"111111101",
  32924=>"111100010",
  32925=>"000000001",
  32926=>"110011101",
  32927=>"100011110",
  32928=>"011100001",
  32929=>"011011001",
  32930=>"001010011",
  32931=>"101101101",
  32932=>"000111111",
  32933=>"000100101",
  32934=>"110101000",
  32935=>"101111100",
  32936=>"100100111",
  32937=>"101011111",
  32938=>"000001110",
  32939=>"110000100",
  32940=>"110100010",
  32941=>"110101000",
  32942=>"101010001",
  32943=>"111110101",
  32944=>"000000110",
  32945=>"111111000",
  32946=>"100110111",
  32947=>"001100000",
  32948=>"000010100",
  32949=>"000101010",
  32950=>"101000000",
  32951=>"100010100",
  32952=>"011101101",
  32953=>"011110001",
  32954=>"110001011",
  32955=>"100110101",
  32956=>"010001111",
  32957=>"001100011",
  32958=>"000110011",
  32959=>"100111100",
  32960=>"111000001",
  32961=>"100011101",
  32962=>"000101011",
  32963=>"011001011",
  32964=>"111000111",
  32965=>"010010111",
  32966=>"110011000",
  32967=>"101111101",
  32968=>"110111110",
  32969=>"000111001",
  32970=>"111001001",
  32971=>"111111000",
  32972=>"001110100",
  32973=>"101100111",
  32974=>"011000000",
  32975=>"111110111",
  32976=>"101110011",
  32977=>"000101110",
  32978=>"010110011",
  32979=>"100011011",
  32980=>"001111100",
  32981=>"001101000",
  32982=>"011100010",
  32983=>"011010111",
  32984=>"100100001",
  32985=>"001100111",
  32986=>"100111110",
  32987=>"111001010",
  32988=>"111011011",
  32989=>"000011011",
  32990=>"110110000",
  32991=>"000100010",
  32992=>"111001101",
  32993=>"101001110",
  32994=>"100101001",
  32995=>"000100100",
  32996=>"100111001",
  32997=>"111111010",
  32998=>"100101011",
  32999=>"011000011",
  33000=>"101111010",
  33001=>"001010000",
  33002=>"100110110",
  33003=>"100100011",
  33004=>"001001001",
  33005=>"010111000",
  33006=>"000110100",
  33007=>"110111111",
  33008=>"100001100",
  33009=>"010101000",
  33010=>"101000000",
  33011=>"011110101",
  33012=>"111101000",
  33013=>"111001000",
  33014=>"010000111",
  33015=>"110000011",
  33016=>"101010001",
  33017=>"100010000",
  33018=>"011110011",
  33019=>"110110000",
  33020=>"101100100",
  33021=>"101101000",
  33022=>"011100110",
  33023=>"000000010",
  33024=>"010001101",
  33025=>"010011111",
  33026=>"001011100",
  33027=>"101000111",
  33028=>"101101110",
  33029=>"001000010",
  33030=>"000000001",
  33031=>"100000101",
  33032=>"111111100",
  33033=>"011010110",
  33034=>"000111011",
  33035=>"110001110",
  33036=>"001010111",
  33037=>"001011111",
  33038=>"010001011",
  33039=>"101000101",
  33040=>"000111110",
  33041=>"101000100",
  33042=>"110010111",
  33043=>"010101110",
  33044=>"101000111",
  33045=>"110000011",
  33046=>"010011000",
  33047=>"101101100",
  33048=>"010100011",
  33049=>"001110000",
  33050=>"100101101",
  33051=>"001000100",
  33052=>"001000101",
  33053=>"000000001",
  33054=>"010100010",
  33055=>"011001110",
  33056=>"100100111",
  33057=>"001011101",
  33058=>"011110101",
  33059=>"011010011",
  33060=>"010101110",
  33061=>"011010100",
  33062=>"110010010",
  33063=>"000101001",
  33064=>"111100001",
  33065=>"111000000",
  33066=>"110011000",
  33067=>"111100101",
  33068=>"110001110",
  33069=>"001110110",
  33070=>"101110011",
  33071=>"001110011",
  33072=>"011000010",
  33073=>"110100000",
  33074=>"110101110",
  33075=>"000000000",
  33076=>"010100111",
  33077=>"010101001",
  33078=>"011111011",
  33079=>"100001110",
  33080=>"111101111",
  33081=>"011100100",
  33082=>"110011111",
  33083=>"111110100",
  33084=>"010110110",
  33085=>"001111110",
  33086=>"111001110",
  33087=>"001100001",
  33088=>"011100111",
  33089=>"111110001",
  33090=>"100001100",
  33091=>"001011101",
  33092=>"101010010",
  33093=>"110010101",
  33094=>"000100000",
  33095=>"101111001",
  33096=>"111101000",
  33097=>"111100110",
  33098=>"001001111",
  33099=>"100111011",
  33100=>"101011011",
  33101=>"001101111",
  33102=>"101000110",
  33103=>"001000001",
  33104=>"100000011",
  33105=>"110101111",
  33106=>"111111101",
  33107=>"100111001",
  33108=>"101000101",
  33109=>"011010110",
  33110=>"110110100",
  33111=>"010001011",
  33112=>"000000011",
  33113=>"001100010",
  33114=>"010100010",
  33115=>"101110011",
  33116=>"001010100",
  33117=>"000011110",
  33118=>"110010011",
  33119=>"011011100",
  33120=>"001000011",
  33121=>"010110110",
  33122=>"011001001",
  33123=>"001100010",
  33124=>"111001111",
  33125=>"011000000",
  33126=>"101010001",
  33127=>"111100101",
  33128=>"001010101",
  33129=>"000101110",
  33130=>"011110011",
  33131=>"100011000",
  33132=>"101011100",
  33133=>"001101101",
  33134=>"111011101",
  33135=>"010101010",
  33136=>"000001100",
  33137=>"001101010",
  33138=>"001010110",
  33139=>"111101010",
  33140=>"000010011",
  33141=>"111000101",
  33142=>"110010010",
  33143=>"100100010",
  33144=>"000001011",
  33145=>"010000011",
  33146=>"011100101",
  33147=>"011000011",
  33148=>"101000111",
  33149=>"110101010",
  33150=>"100010100",
  33151=>"101011100",
  33152=>"001111110",
  33153=>"011000010",
  33154=>"010010100",
  33155=>"000101010",
  33156=>"000011000",
  33157=>"101011111",
  33158=>"101111100",
  33159=>"111111110",
  33160=>"001100101",
  33161=>"010001100",
  33162=>"100011100",
  33163=>"110001011",
  33164=>"011110001",
  33165=>"100101000",
  33166=>"110110000",
  33167=>"100011011",
  33168=>"011001001",
  33169=>"010000001",
  33170=>"000011000",
  33171=>"101011010",
  33172=>"100100110",
  33173=>"010101101",
  33174=>"111110010",
  33175=>"111111011",
  33176=>"011001101",
  33177=>"110001011",
  33178=>"011001100",
  33179=>"000001100",
  33180=>"100011100",
  33181=>"001101110",
  33182=>"000010111",
  33183=>"011000111",
  33184=>"101111110",
  33185=>"001000110",
  33186=>"101111110",
  33187=>"101111010",
  33188=>"101101110",
  33189=>"101101100",
  33190=>"011010110",
  33191=>"111000011",
  33192=>"101001000",
  33193=>"100010010",
  33194=>"001000000",
  33195=>"000101011",
  33196=>"110110111",
  33197=>"111000111",
  33198=>"111000101",
  33199=>"111100111",
  33200=>"011111111",
  33201=>"110000000",
  33202=>"101111001",
  33203=>"010010011",
  33204=>"111111001",
  33205=>"111001011",
  33206=>"100010000",
  33207=>"110011000",
  33208=>"100000010",
  33209=>"000110001",
  33210=>"110001010",
  33211=>"001100010",
  33212=>"111101101",
  33213=>"001000011",
  33214=>"001001001",
  33215=>"110100111",
  33216=>"111000001",
  33217=>"110111000",
  33218=>"011100001",
  33219=>"000110000",
  33220=>"111000100",
  33221=>"101001100",
  33222=>"000000100",
  33223=>"101011110",
  33224=>"010001010",
  33225=>"100111001",
  33226=>"111100011",
  33227=>"111000111",
  33228=>"000101001",
  33229=>"001000111",
  33230=>"101101101",
  33231=>"010101011",
  33232=>"011110101",
  33233=>"110100001",
  33234=>"111001100",
  33235=>"000000101",
  33236=>"011100001",
  33237=>"010110100",
  33238=>"110101100",
  33239=>"000111010",
  33240=>"111110110",
  33241=>"010100000",
  33242=>"001101111",
  33243=>"101011101",
  33244=>"000010100",
  33245=>"001111011",
  33246=>"011101111",
  33247=>"000011100",
  33248=>"101000111",
  33249=>"000001000",
  33250=>"111100101",
  33251=>"010100000",
  33252=>"100110000",
  33253=>"100000110",
  33254=>"100110111",
  33255=>"000110010",
  33256=>"010111011",
  33257=>"000011101",
  33258=>"011101100",
  33259=>"011011100",
  33260=>"001010101",
  33261=>"110111110",
  33262=>"000000111",
  33263=>"101010001",
  33264=>"001111001",
  33265=>"100011101",
  33266=>"101011001",
  33267=>"000100101",
  33268=>"000110000",
  33269=>"111001100",
  33270=>"110101101",
  33271=>"111101101",
  33272=>"101111001",
  33273=>"111011101",
  33274=>"011111111",
  33275=>"001010101",
  33276=>"001001000",
  33277=>"111001010",
  33278=>"101000010",
  33279=>"011000011",
  33280=>"110000110",
  33281=>"011010001",
  33282=>"111000110",
  33283=>"011010001",
  33284=>"011111000",
  33285=>"110110010",
  33286=>"000110001",
  33287=>"100111101",
  33288=>"010110000",
  33289=>"000101011",
  33290=>"000001001",
  33291=>"011111000",
  33292=>"000110011",
  33293=>"111011111",
  33294=>"001100100",
  33295=>"111111010",
  33296=>"111001110",
  33297=>"010001000",
  33298=>"001111011",
  33299=>"010100100",
  33300=>"011101100",
  33301=>"001011111",
  33302=>"110101010",
  33303=>"010110000",
  33304=>"001010100",
  33305=>"101001011",
  33306=>"011011001",
  33307=>"111001100",
  33308=>"001001101",
  33309=>"011010110",
  33310=>"101010010",
  33311=>"011110010",
  33312=>"001010011",
  33313=>"100000100",
  33314=>"101000010",
  33315=>"001110110",
  33316=>"101100000",
  33317=>"111110011",
  33318=>"100101100",
  33319=>"001011001",
  33320=>"101100110",
  33321=>"111011110",
  33322=>"111111111",
  33323=>"000011011",
  33324=>"100110100",
  33325=>"001110110",
  33326=>"000010001",
  33327=>"000110000",
  33328=>"101000000",
  33329=>"101110011",
  33330=>"101000111",
  33331=>"000101110",
  33332=>"100101000",
  33333=>"101001011",
  33334=>"111110000",
  33335=>"100101011",
  33336=>"111000111",
  33337=>"100101111",
  33338=>"100000110",
  33339=>"000001101",
  33340=>"001111000",
  33341=>"010100000",
  33342=>"000101000",
  33343=>"101111001",
  33344=>"101111100",
  33345=>"101111001",
  33346=>"111111100",
  33347=>"010011001",
  33348=>"110010111",
  33349=>"010011110",
  33350=>"010100011",
  33351=>"100100100",
  33352=>"011110100",
  33353=>"111010111",
  33354=>"110110100",
  33355=>"000100000",
  33356=>"100001101",
  33357=>"010110001",
  33358=>"100101110",
  33359=>"101101100",
  33360=>"010010010",
  33361=>"011011010",
  33362=>"011011101",
  33363=>"111101011",
  33364=>"010000011",
  33365=>"010000101",
  33366=>"100000001",
  33367=>"000100011",
  33368=>"110100000",
  33369=>"001011100",
  33370=>"010010000",
  33371=>"000100010",
  33372=>"001111010",
  33373=>"010001001",
  33374=>"110011010",
  33375=>"010000101",
  33376=>"011110110",
  33377=>"101111111",
  33378=>"101000010",
  33379=>"111101110",
  33380=>"111010100",
  33381=>"111100010",
  33382=>"010110100",
  33383=>"010000010",
  33384=>"010110101",
  33385=>"001111010",
  33386=>"000110011",
  33387=>"111100111",
  33388=>"001011111",
  33389=>"010000101",
  33390=>"000100010",
  33391=>"111011011",
  33392=>"000100011",
  33393=>"011010110",
  33394=>"100011110",
  33395=>"111110110",
  33396=>"000110000",
  33397=>"101011001",
  33398=>"100000110",
  33399=>"010110000",
  33400=>"011011011",
  33401=>"001001100",
  33402=>"101100110",
  33403=>"000110001",
  33404=>"111001001",
  33405=>"000010010",
  33406=>"110110100",
  33407=>"010101101",
  33408=>"000010000",
  33409=>"001110001",
  33410=>"100101000",
  33411=>"110101001",
  33412=>"001111011",
  33413=>"011010001",
  33414=>"001101101",
  33415=>"000011111",
  33416=>"110000011",
  33417=>"000011101",
  33418=>"110001100",
  33419=>"001011000",
  33420=>"101100101",
  33421=>"011001110",
  33422=>"001111111",
  33423=>"000001011",
  33424=>"011001000",
  33425=>"100001100",
  33426=>"100110101",
  33427=>"010101110",
  33428=>"011111100",
  33429=>"110011101",
  33430=>"010100101",
  33431=>"111101100",
  33432=>"010110001",
  33433=>"111010100",
  33434=>"101110010",
  33435=>"101010100",
  33436=>"010111011",
  33437=>"000100000",
  33438=>"001000101",
  33439=>"000000001",
  33440=>"001110101",
  33441=>"001010010",
  33442=>"111111100",
  33443=>"110101111",
  33444=>"011101100",
  33445=>"010100101",
  33446=>"010011011",
  33447=>"001011011",
  33448=>"001101000",
  33449=>"010001011",
  33450=>"101110101",
  33451=>"011010110",
  33452=>"011010000",
  33453=>"000001110",
  33454=>"101100000",
  33455=>"101101011",
  33456=>"101001010",
  33457=>"101001110",
  33458=>"001011010",
  33459=>"001111010",
  33460=>"000011011",
  33461=>"011011100",
  33462=>"001101001",
  33463=>"010001000",
  33464=>"010110001",
  33465=>"111010001",
  33466=>"010100000",
  33467=>"100010101",
  33468=>"110111110",
  33469=>"111010100",
  33470=>"111100010",
  33471=>"101100110",
  33472=>"111101111",
  33473=>"110001100",
  33474=>"111000010",
  33475=>"110101100",
  33476=>"010101011",
  33477=>"000001001",
  33478=>"111000000",
  33479=>"010000000",
  33480=>"000001011",
  33481=>"100111110",
  33482=>"011110000",
  33483=>"010111111",
  33484=>"011111010",
  33485=>"010110010",
  33486=>"110111000",
  33487=>"100100001",
  33488=>"101010000",
  33489=>"101010011",
  33490=>"110010001",
  33491=>"011000101",
  33492=>"011110010",
  33493=>"001011111",
  33494=>"101010111",
  33495=>"101111001",
  33496=>"111101110",
  33497=>"000010101",
  33498=>"010111111",
  33499=>"011101001",
  33500=>"110001000",
  33501=>"111110101",
  33502=>"110000001",
  33503=>"111011110",
  33504=>"001011100",
  33505=>"110100010",
  33506=>"011100111",
  33507=>"011111000",
  33508=>"011011100",
  33509=>"011111110",
  33510=>"101110000",
  33511=>"010110001",
  33512=>"101111101",
  33513=>"111110100",
  33514=>"111000110",
  33515=>"111111010",
  33516=>"011110101",
  33517=>"110110110",
  33518=>"111011100",
  33519=>"101100000",
  33520=>"101010111",
  33521=>"101000001",
  33522=>"101010111",
  33523=>"000010101",
  33524=>"010011001",
  33525=>"000010010",
  33526=>"010000010",
  33527=>"110010010",
  33528=>"100100110",
  33529=>"010110110",
  33530=>"001110100",
  33531=>"000000111",
  33532=>"110110001",
  33533=>"001101111",
  33534=>"111000010",
  33535=>"000011010",
  33536=>"101101011",
  33537=>"001101001",
  33538=>"010110110",
  33539=>"101001110",
  33540=>"000001111",
  33541=>"010001000",
  33542=>"101110110",
  33543=>"101110000",
  33544=>"101011011",
  33545=>"100110110",
  33546=>"001010010",
  33547=>"010000010",
  33548=>"101110111",
  33549=>"111011100",
  33550=>"000111111",
  33551=>"011010000",
  33552=>"010011111",
  33553=>"011110111",
  33554=>"000000011",
  33555=>"011010010",
  33556=>"011011111",
  33557=>"110110101",
  33558=>"011110111",
  33559=>"101010100",
  33560=>"000011000",
  33561=>"000000101",
  33562=>"111110110",
  33563=>"010100100",
  33564=>"101110001",
  33565=>"101011011",
  33566=>"000011000",
  33567=>"000101001",
  33568=>"011101101",
  33569=>"111010111",
  33570=>"001111111",
  33571=>"111001001",
  33572=>"000001100",
  33573=>"100001001",
  33574=>"000110101",
  33575=>"011111101",
  33576=>"110010100",
  33577=>"000111010",
  33578=>"011110000",
  33579=>"000001101",
  33580=>"111110010",
  33581=>"110001110",
  33582=>"101101001",
  33583=>"010111111",
  33584=>"110010110",
  33585=>"001101001",
  33586=>"100100101",
  33587=>"010111000",
  33588=>"111010100",
  33589=>"101000101",
  33590=>"111010000",
  33591=>"010011110",
  33592=>"011010001",
  33593=>"001111100",
  33594=>"001000011",
  33595=>"100001011",
  33596=>"000000001",
  33597=>"101100001",
  33598=>"000001110",
  33599=>"100110111",
  33600=>"110110111",
  33601=>"011111010",
  33602=>"111001111",
  33603=>"100111000",
  33604=>"101011110",
  33605=>"110111101",
  33606=>"111000101",
  33607=>"010101000",
  33608=>"110010001",
  33609=>"100111101",
  33610=>"010111001",
  33611=>"101001000",
  33612=>"011011001",
  33613=>"101101111",
  33614=>"100011011",
  33615=>"100001100",
  33616=>"100101111",
  33617=>"011000001",
  33618=>"101001000",
  33619=>"000011100",
  33620=>"101101111",
  33621=>"111110010",
  33622=>"000010110",
  33623=>"100101011",
  33624=>"101010001",
  33625=>"011010110",
  33626=>"100111001",
  33627=>"101101101",
  33628=>"100011101",
  33629=>"111001101",
  33630=>"111111010",
  33631=>"000011010",
  33632=>"010110001",
  33633=>"001111000",
  33634=>"101110011",
  33635=>"101001100",
  33636=>"011111110",
  33637=>"011010011",
  33638=>"011011100",
  33639=>"001101110",
  33640=>"110010111",
  33641=>"001011111",
  33642=>"111101010",
  33643=>"010101000",
  33644=>"000001111",
  33645=>"000011011",
  33646=>"101001001",
  33647=>"101111111",
  33648=>"010000010",
  33649=>"011001010",
  33650=>"111011100",
  33651=>"001001111",
  33652=>"000011010",
  33653=>"111101100",
  33654=>"101111100",
  33655=>"000100001",
  33656=>"001010001",
  33657=>"001010000",
  33658=>"101001010",
  33659=>"100001110",
  33660=>"010010000",
  33661=>"101001111",
  33662=>"111101110",
  33663=>"010010100",
  33664=>"010011110",
  33665=>"011001101",
  33666=>"100010111",
  33667=>"110010111",
  33668=>"001010000",
  33669=>"110011110",
  33670=>"100101110",
  33671=>"101100001",
  33672=>"101011111",
  33673=>"001100011",
  33674=>"110101100",
  33675=>"110100100",
  33676=>"111101011",
  33677=>"100011110",
  33678=>"010011001",
  33679=>"100111111",
  33680=>"001011101",
  33681=>"110111100",
  33682=>"000011011",
  33683=>"010010101",
  33684=>"110101111",
  33685=>"111001101",
  33686=>"101000110",
  33687=>"011001011",
  33688=>"111010000",
  33689=>"001010101",
  33690=>"010000100",
  33691=>"000010100",
  33692=>"000100100",
  33693=>"011010110",
  33694=>"111011111",
  33695=>"011101111",
  33696=>"010110110",
  33697=>"000101000",
  33698=>"100010000",
  33699=>"100001010",
  33700=>"111000000",
  33701=>"000101011",
  33702=>"001011100",
  33703=>"010010000",
  33704=>"000011100",
  33705=>"111000000",
  33706=>"100000011",
  33707=>"011100000",
  33708=>"100010100",
  33709=>"001001000",
  33710=>"110110000",
  33711=>"100101000",
  33712=>"001000000",
  33713=>"000101101",
  33714=>"111100010",
  33715=>"110010101",
  33716=>"011011101",
  33717=>"111010111",
  33718=>"110011111",
  33719=>"110111100",
  33720=>"100000000",
  33721=>"101011110",
  33722=>"001001010",
  33723=>"100000010",
  33724=>"001001001",
  33725=>"000011000",
  33726=>"100001101",
  33727=>"111010110",
  33728=>"110001111",
  33729=>"101000010",
  33730=>"101101100",
  33731=>"111001011",
  33732=>"000001011",
  33733=>"110011111",
  33734=>"101001000",
  33735=>"111000110",
  33736=>"111001000",
  33737=>"100000001",
  33738=>"110100110",
  33739=>"001011010",
  33740=>"101001010",
  33741=>"011000010",
  33742=>"101110101",
  33743=>"101111001",
  33744=>"000110011",
  33745=>"101110110",
  33746=>"100010010",
  33747=>"100101000",
  33748=>"000111110",
  33749=>"001011111",
  33750=>"100001110",
  33751=>"000001000",
  33752=>"000000000",
  33753=>"001110000",
  33754=>"110101111",
  33755=>"100001011",
  33756=>"111011011",
  33757=>"111111000",
  33758=>"101111001",
  33759=>"100000011",
  33760=>"100000001",
  33761=>"000000010",
  33762=>"110001100",
  33763=>"101101010",
  33764=>"010001010",
  33765=>"111001010",
  33766=>"110110101",
  33767=>"110100010",
  33768=>"011111010",
  33769=>"011010010",
  33770=>"000101110",
  33771=>"100010000",
  33772=>"111101111",
  33773=>"101101110",
  33774=>"101100010",
  33775=>"110000000",
  33776=>"101111001",
  33777=>"001010011",
  33778=>"000000101",
  33779=>"001000110",
  33780=>"110110010",
  33781=>"011101011",
  33782=>"010100111",
  33783=>"000000011",
  33784=>"011101010",
  33785=>"000000000",
  33786=>"111010010",
  33787=>"000010110",
  33788=>"110100001",
  33789=>"011100010",
  33790=>"110001000",
  33791=>"001001001",
  33792=>"000000000",
  33793=>"100000001",
  33794=>"111010000",
  33795=>"010101010",
  33796=>"110111001",
  33797=>"011110000",
  33798=>"101000101",
  33799=>"101101110",
  33800=>"101011000",
  33801=>"100001000",
  33802=>"111110010",
  33803=>"110000110",
  33804=>"001001110",
  33805=>"111110000",
  33806=>"011100101",
  33807=>"001001011",
  33808=>"000001011",
  33809=>"110111001",
  33810=>"100010001",
  33811=>"110010101",
  33812=>"100110000",
  33813=>"011011001",
  33814=>"110001110",
  33815=>"010001110",
  33816=>"100100110",
  33817=>"010001010",
  33818=>"101001010",
  33819=>"100011110",
  33820=>"001001000",
  33821=>"010001000",
  33822=>"111011011",
  33823=>"011011000",
  33824=>"001010100",
  33825=>"000111111",
  33826=>"101001100",
  33827=>"101100010",
  33828=>"010011100",
  33829=>"000010101",
  33830=>"001110000",
  33831=>"101000000",
  33832=>"000110100",
  33833=>"101100001",
  33834=>"011011110",
  33835=>"100111001",
  33836=>"111010100",
  33837=>"101101101",
  33838=>"011111100",
  33839=>"100100101",
  33840=>"101001001",
  33841=>"111110001",
  33842=>"100111001",
  33843=>"010111111",
  33844=>"011110001",
  33845=>"100110011",
  33846=>"110110101",
  33847=>"100001010",
  33848=>"100001001",
  33849=>"101010101",
  33850=>"110000001",
  33851=>"111100111",
  33852=>"101000100",
  33853=>"001010001",
  33854=>"110010011",
  33855=>"000011101",
  33856=>"011011111",
  33857=>"000101011",
  33858=>"001111011",
  33859=>"011000110",
  33860=>"110010010",
  33861=>"010101100",
  33862=>"001100011",
  33863=>"110011001",
  33864=>"101011111",
  33865=>"001000001",
  33866=>"100010100",
  33867=>"100101000",
  33868=>"100110101",
  33869=>"110111110",
  33870=>"011100110",
  33871=>"011101101",
  33872=>"000010000",
  33873=>"000001011",
  33874=>"000010001",
  33875=>"000100001",
  33876=>"000100111",
  33877=>"110001110",
  33878=>"111001111",
  33879=>"101100010",
  33880=>"011001100",
  33881=>"001001011",
  33882=>"001011001",
  33883=>"000010000",
  33884=>"000110110",
  33885=>"101011000",
  33886=>"111100010",
  33887=>"000010110",
  33888=>"001010101",
  33889=>"100001011",
  33890=>"001011101",
  33891=>"100100111",
  33892=>"110011001",
  33893=>"001000110",
  33894=>"100000010",
  33895=>"001010110",
  33896=>"100100111",
  33897=>"100111000",
  33898=>"101101110",
  33899=>"100110001",
  33900=>"010001001",
  33901=>"011000001",
  33902=>"010001101",
  33903=>"000010111",
  33904=>"000010000",
  33905=>"110100011",
  33906=>"100011111",
  33907=>"001100000",
  33908=>"111111101",
  33909=>"000000010",
  33910=>"110011011",
  33911=>"101001110",
  33912=>"110011011",
  33913=>"111111101",
  33914=>"000001100",
  33915=>"011001111",
  33916=>"011000011",
  33917=>"000101101",
  33918=>"001011000",
  33919=>"000100110",
  33920=>"000001100",
  33921=>"110011000",
  33922=>"000000100",
  33923=>"110000111",
  33924=>"010001011",
  33925=>"110111000",
  33926=>"001000101",
  33927=>"111100101",
  33928=>"001010010",
  33929=>"011111000",
  33930=>"010000101",
  33931=>"101011011",
  33932=>"000100100",
  33933=>"100001011",
  33934=>"001101101",
  33935=>"100000001",
  33936=>"111111110",
  33937=>"101111110",
  33938=>"011000110",
  33939=>"111000111",
  33940=>"110111101",
  33941=>"110100000",
  33942=>"111110011",
  33943=>"110100101",
  33944=>"010111001",
  33945=>"011101010",
  33946=>"101010101",
  33947=>"110101100",
  33948=>"011000010",
  33949=>"110110101",
  33950=>"010110100",
  33951=>"111010110",
  33952=>"110010001",
  33953=>"001000000",
  33954=>"000110111",
  33955=>"111000010",
  33956=>"001011110",
  33957=>"000000110",
  33958=>"000011100",
  33959=>"100111110",
  33960=>"011111000",
  33961=>"000110110",
  33962=>"100001001",
  33963=>"110101111",
  33964=>"010101110",
  33965=>"101000100",
  33966=>"010110000",
  33967=>"101111101",
  33968=>"011010010",
  33969=>"011101010",
  33970=>"001011000",
  33971=>"101000000",
  33972=>"100011011",
  33973=>"111011101",
  33974=>"100000100",
  33975=>"000100000",
  33976=>"011001100",
  33977=>"011100001",
  33978=>"001110100",
  33979=>"001100101",
  33980=>"000001101",
  33981=>"000010010",
  33982=>"000111000",
  33983=>"100100001",
  33984=>"100100110",
  33985=>"001110001",
  33986=>"111110011",
  33987=>"111110101",
  33988=>"001001010",
  33989=>"011010100",
  33990=>"111111100",
  33991=>"110001110",
  33992=>"110001100",
  33993=>"001001111",
  33994=>"000011101",
  33995=>"101101101",
  33996=>"111000000",
  33997=>"110110100",
  33998=>"110110001",
  33999=>"101001010",
  34000=>"001101000",
  34001=>"001011010",
  34002=>"001110000",
  34003=>"110100000",
  34004=>"001111111",
  34005=>"000100111",
  34006=>"100011000",
  34007=>"100000111",
  34008=>"010111101",
  34009=>"001011011",
  34010=>"010010111",
  34011=>"111110000",
  34012=>"100100000",
  34013=>"111011111",
  34014=>"000100000",
  34015=>"101101010",
  34016=>"000110101",
  34017=>"011010010",
  34018=>"100011111",
  34019=>"011110110",
  34020=>"110101011",
  34021=>"100000100",
  34022=>"001001110",
  34023=>"110111010",
  34024=>"100111101",
  34025=>"111001000",
  34026=>"010110110",
  34027=>"101001101",
  34028=>"011010010",
  34029=>"100000010",
  34030=>"001101010",
  34031=>"011010111",
  34032=>"011111011",
  34033=>"101010001",
  34034=>"110000111",
  34035=>"100000001",
  34036=>"110100110",
  34037=>"111001111",
  34038=>"000110001",
  34039=>"000000000",
  34040=>"011010001",
  34041=>"111111100",
  34042=>"111100100",
  34043=>"110110100",
  34044=>"000001010",
  34045=>"010000010",
  34046=>"110101101",
  34047=>"110000101",
  34048=>"110010111",
  34049=>"110101011",
  34050=>"000101101",
  34051=>"001101001",
  34052=>"011001101",
  34053=>"111101100",
  34054=>"001011110",
  34055=>"010110111",
  34056=>"010101111",
  34057=>"110101011",
  34058=>"001000011",
  34059=>"100101100",
  34060=>"001011110",
  34061=>"011010000",
  34062=>"011011111",
  34063=>"101100100",
  34064=>"011001001",
  34065=>"111000110",
  34066=>"011100110",
  34067=>"101110101",
  34068=>"000111001",
  34069=>"111100100",
  34070=>"100011111",
  34071=>"000001011",
  34072=>"101111011",
  34073=>"001101011",
  34074=>"100110111",
  34075=>"011011001",
  34076=>"011100101",
  34077=>"001101110",
  34078=>"011100010",
  34079=>"011001010",
  34080=>"000000111",
  34081=>"110011110",
  34082=>"000011011",
  34083=>"011000011",
  34084=>"001100111",
  34085=>"111011010",
  34086=>"110111110",
  34087=>"101100001",
  34088=>"101010010",
  34089=>"111100101",
  34090=>"111011100",
  34091=>"110100100",
  34092=>"111001110",
  34093=>"111111111",
  34094=>"101100000",
  34095=>"100101101",
  34096=>"101000110",
  34097=>"100011011",
  34098=>"100110010",
  34099=>"000001001",
  34100=>"000110100",
  34101=>"100011111",
  34102=>"110000110",
  34103=>"010000100",
  34104=>"101111110",
  34105=>"001100001",
  34106=>"010111110",
  34107=>"000111000",
  34108=>"100101111",
  34109=>"111101111",
  34110=>"010100011",
  34111=>"110110111",
  34112=>"001000010",
  34113=>"110001011",
  34114=>"001111110",
  34115=>"000010101",
  34116=>"101000011",
  34117=>"010010100",
  34118=>"001000110",
  34119=>"000100110",
  34120=>"011011110",
  34121=>"011010101",
  34122=>"100001000",
  34123=>"111110100",
  34124=>"100101101",
  34125=>"000001101",
  34126=>"101011111",
  34127=>"001101100",
  34128=>"100100010",
  34129=>"111011011",
  34130=>"100010010",
  34131=>"110111100",
  34132=>"001111100",
  34133=>"101000110",
  34134=>"101110000",
  34135=>"101011001",
  34136=>"111100010",
  34137=>"100101000",
  34138=>"001100101",
  34139=>"110010000",
  34140=>"110001001",
  34141=>"010110111",
  34142=>"101011000",
  34143=>"000010011",
  34144=>"000100000",
  34145=>"011110110",
  34146=>"000111011",
  34147=>"001000001",
  34148=>"101111110",
  34149=>"000011100",
  34150=>"000000010",
  34151=>"101011010",
  34152=>"011011101",
  34153=>"001110011",
  34154=>"001011100",
  34155=>"000011101",
  34156=>"110100100",
  34157=>"001111011",
  34158=>"001101000",
  34159=>"000100111",
  34160=>"101000101",
  34161=>"111000011",
  34162=>"100000010",
  34163=>"010110111",
  34164=>"101111101",
  34165=>"001101111",
  34166=>"101101110",
  34167=>"011110100",
  34168=>"001000011",
  34169=>"100100011",
  34170=>"111110011",
  34171=>"100011101",
  34172=>"100101110",
  34173=>"010011101",
  34174=>"011011111",
  34175=>"101100110",
  34176=>"010101100",
  34177=>"101100011",
  34178=>"010110110",
  34179=>"110001010",
  34180=>"100001100",
  34181=>"001100100",
  34182=>"111001001",
  34183=>"110101010",
  34184=>"010011101",
  34185=>"000001001",
  34186=>"100001000",
  34187=>"011010001",
  34188=>"110000100",
  34189=>"011101111",
  34190=>"011100000",
  34191=>"011001010",
  34192=>"001110110",
  34193=>"000101000",
  34194=>"100111011",
  34195=>"111011001",
  34196=>"111001010",
  34197=>"001010011",
  34198=>"001011100",
  34199=>"100011111",
  34200=>"111111111",
  34201=>"100000100",
  34202=>"100010101",
  34203=>"110100000",
  34204=>"010101110",
  34205=>"001011010",
  34206=>"000000110",
  34207=>"001101001",
  34208=>"110100000",
  34209=>"000001111",
  34210=>"100111110",
  34211=>"111100100",
  34212=>"110011110",
  34213=>"101010100",
  34214=>"111110000",
  34215=>"000110010",
  34216=>"001001010",
  34217=>"110001001",
  34218=>"110110101",
  34219=>"001010100",
  34220=>"000001100",
  34221=>"101011011",
  34222=>"111110010",
  34223=>"001110000",
  34224=>"110011011",
  34225=>"110000000",
  34226=>"000011010",
  34227=>"010010101",
  34228=>"000000011",
  34229=>"001000111",
  34230=>"111100100",
  34231=>"010110100",
  34232=>"001110100",
  34233=>"110101011",
  34234=>"000111101",
  34235=>"101101100",
  34236=>"111000010",
  34237=>"000111010",
  34238=>"000101101",
  34239=>"011001111",
  34240=>"011101001",
  34241=>"000000011",
  34242=>"011111110",
  34243=>"010000100",
  34244=>"100000101",
  34245=>"110001000",
  34246=>"100010000",
  34247=>"000011001",
  34248=>"101010011",
  34249=>"001101101",
  34250=>"011011101",
  34251=>"110100000",
  34252=>"110100010",
  34253=>"010110101",
  34254=>"101010000",
  34255=>"111111010",
  34256=>"010111011",
  34257=>"000000110",
  34258=>"011111110",
  34259=>"111100110",
  34260=>"111101100",
  34261=>"001001001",
  34262=>"110001111",
  34263=>"010010000",
  34264=>"011011001",
  34265=>"101110101",
  34266=>"111011111",
  34267=>"101100010",
  34268=>"001000110",
  34269=>"000111111",
  34270=>"111001000",
  34271=>"110010000",
  34272=>"001011010",
  34273=>"010110000",
  34274=>"101000010",
  34275=>"110010011",
  34276=>"010110111",
  34277=>"010110011",
  34278=>"010001010",
  34279=>"110100110",
  34280=>"011010000",
  34281=>"000111110",
  34282=>"101000001",
  34283=>"000100001",
  34284=>"100001010",
  34285=>"110101100",
  34286=>"000000100",
  34287=>"010000110",
  34288=>"111010011",
  34289=>"010001101",
  34290=>"110010100",
  34291=>"011101111",
  34292=>"111000010",
  34293=>"001100001",
  34294=>"001101000",
  34295=>"111101001",
  34296=>"111111010",
  34297=>"011011100",
  34298=>"011110010",
  34299=>"000011100",
  34300=>"110111000",
  34301=>"111001100",
  34302=>"010000001",
  34303=>"100011001",
  34304=>"011111110",
  34305=>"001000000",
  34306=>"101100110",
  34307=>"000000101",
  34308=>"111110001",
  34309=>"110001010",
  34310=>"111111010",
  34311=>"011010101",
  34312=>"110011001",
  34313=>"000001011",
  34314=>"011111101",
  34315=>"010010011",
  34316=>"101110000",
  34317=>"101010000",
  34318=>"100000101",
  34319=>"101000001",
  34320=>"100110010",
  34321=>"110011101",
  34322=>"000111100",
  34323=>"100100110",
  34324=>"001001110",
  34325=>"010100100",
  34326=>"101111001",
  34327=>"101101110",
  34328=>"001000111",
  34329=>"010010110",
  34330=>"111101010",
  34331=>"001011011",
  34332=>"011011000",
  34333=>"111100000",
  34334=>"010011100",
  34335=>"100011011",
  34336=>"101110110",
  34337=>"101000100",
  34338=>"000101010",
  34339=>"111111011",
  34340=>"011001111",
  34341=>"000011111",
  34342=>"111110111",
  34343=>"010011100",
  34344=>"011010100",
  34345=>"111101011",
  34346=>"000010101",
  34347=>"100101011",
  34348=>"001001111",
  34349=>"010001001",
  34350=>"000010001",
  34351=>"010101111",
  34352=>"101010110",
  34353=>"110001000",
  34354=>"101001101",
  34355=>"100001010",
  34356=>"001011100",
  34357=>"001100111",
  34358=>"000010001",
  34359=>"010000000",
  34360=>"110001100",
  34361=>"010101001",
  34362=>"111010000",
  34363=>"101010000",
  34364=>"000000100",
  34365=>"100000100",
  34366=>"010011111",
  34367=>"001000110",
  34368=>"110101111",
  34369=>"000100010",
  34370=>"001110111",
  34371=>"100101011",
  34372=>"110101000",
  34373=>"001100100",
  34374=>"110011111",
  34375=>"010110000",
  34376=>"111111011",
  34377=>"001101100",
  34378=>"001001000",
  34379=>"000101011",
  34380=>"000001000",
  34381=>"000010011",
  34382=>"011000100",
  34383=>"101100110",
  34384=>"000011000",
  34385=>"111011010",
  34386=>"010100111",
  34387=>"111000000",
  34388=>"011000110",
  34389=>"110101110",
  34390=>"001100001",
  34391=>"111010111",
  34392=>"011000101",
  34393=>"010011111",
  34394=>"001111110",
  34395=>"001001100",
  34396=>"000100011",
  34397=>"100101010",
  34398=>"110001100",
  34399=>"100111010",
  34400=>"000001111",
  34401=>"101001111",
  34402=>"000001111",
  34403=>"111101001",
  34404=>"101111000",
  34405=>"111010110",
  34406=>"100010110",
  34407=>"111001111",
  34408=>"110001010",
  34409=>"001100111",
  34410=>"111010111",
  34411=>"000100110",
  34412=>"111001011",
  34413=>"110001100",
  34414=>"110001100",
  34415=>"101001100",
  34416=>"110001101",
  34417=>"000110100",
  34418=>"011111011",
  34419=>"010100110",
  34420=>"001011011",
  34421=>"101010100",
  34422=>"111101100",
  34423=>"010000010",
  34424=>"010111111",
  34425=>"010111000",
  34426=>"111011011",
  34427=>"111000001",
  34428=>"010100111",
  34429=>"101111001",
  34430=>"000000100",
  34431=>"110001111",
  34432=>"000000101",
  34433=>"111000010",
  34434=>"011011101",
  34435=>"001000101",
  34436=>"001110111",
  34437=>"100101111",
  34438=>"101011011",
  34439=>"111101101",
  34440=>"111001000",
  34441=>"001111000",
  34442=>"101110011",
  34443=>"100110000",
  34444=>"001011100",
  34445=>"100111101",
  34446=>"001111011",
  34447=>"011010111",
  34448=>"010111000",
  34449=>"001100010",
  34450=>"011010100",
  34451=>"000011111",
  34452=>"000111011",
  34453=>"001011111",
  34454=>"001110111",
  34455=>"100010100",
  34456=>"010010101",
  34457=>"000110101",
  34458=>"111100111",
  34459=>"100101001",
  34460=>"001000101",
  34461=>"000000011",
  34462=>"000100001",
  34463=>"100110011",
  34464=>"101110000",
  34465=>"010111111",
  34466=>"011110101",
  34467=>"010101101",
  34468=>"000100100",
  34469=>"111011001",
  34470=>"000100001",
  34471=>"100000100",
  34472=>"001111010",
  34473=>"010101010",
  34474=>"001110111",
  34475=>"100000010",
  34476=>"000011010",
  34477=>"001010111",
  34478=>"011101011",
  34479=>"111110001",
  34480=>"100001101",
  34481=>"100100000",
  34482=>"001000000",
  34483=>"000000001",
  34484=>"001100010",
  34485=>"111111110",
  34486=>"010010000",
  34487=>"010010110",
  34488=>"000101000",
  34489=>"010011011",
  34490=>"001110010",
  34491=>"011111010",
  34492=>"110000010",
  34493=>"010100000",
  34494=>"001111100",
  34495=>"000100010",
  34496=>"011011010",
  34497=>"111100111",
  34498=>"000011001",
  34499=>"010101111",
  34500=>"110100110",
  34501=>"010000000",
  34502=>"011001010",
  34503=>"111100110",
  34504=>"100011000",
  34505=>"100000110",
  34506=>"100111101",
  34507=>"101110001",
  34508=>"111000001",
  34509=>"001111111",
  34510=>"110000100",
  34511=>"100101011",
  34512=>"110100000",
  34513=>"000001011",
  34514=>"010011111",
  34515=>"100110101",
  34516=>"111011000",
  34517=>"100110100",
  34518=>"011011101",
  34519=>"010111101",
  34520=>"111001100",
  34521=>"001011000",
  34522=>"010000010",
  34523=>"110111011",
  34524=>"101000101",
  34525=>"111101001",
  34526=>"101100101",
  34527=>"011010010",
  34528=>"010001101",
  34529=>"000001010",
  34530=>"110101011",
  34531=>"111001001",
  34532=>"001000010",
  34533=>"100001100",
  34534=>"001001111",
  34535=>"000010100",
  34536=>"001000000",
  34537=>"101110010",
  34538=>"011010101",
  34539=>"011000011",
  34540=>"001101000",
  34541=>"011110100",
  34542=>"110010100",
  34543=>"101001100",
  34544=>"110010111",
  34545=>"000001101",
  34546=>"101111100",
  34547=>"000001001",
  34548=>"000011110",
  34549=>"111001101",
  34550=>"110110111",
  34551=>"101011100",
  34552=>"011100111",
  34553=>"111101100",
  34554=>"000111001",
  34555=>"110101100",
  34556=>"011111110",
  34557=>"100010000",
  34558=>"001000001",
  34559=>"110001000",
  34560=>"101110011",
  34561=>"101011111",
  34562=>"111111110",
  34563=>"100010110",
  34564=>"111010011",
  34565=>"100110011",
  34566=>"000001001",
  34567=>"101110100",
  34568=>"110111001",
  34569=>"010111001",
  34570=>"011101101",
  34571=>"101001010",
  34572=>"000010110",
  34573=>"000101100",
  34574=>"011011110",
  34575=>"101011100",
  34576=>"110100011",
  34577=>"000000001",
  34578=>"011000001",
  34579=>"110110010",
  34580=>"111010101",
  34581=>"000011101",
  34582=>"100111011",
  34583=>"011111100",
  34584=>"100010010",
  34585=>"100101000",
  34586=>"000110101",
  34587=>"011110010",
  34588=>"010011111",
  34589=>"011110001",
  34590=>"010010011",
  34591=>"010010101",
  34592=>"101000001",
  34593=>"100110100",
  34594=>"101100111",
  34595=>"110100011",
  34596=>"010001011",
  34597=>"001001100",
  34598=>"100110101",
  34599=>"010010001",
  34600=>"000111011",
  34601=>"001101011",
  34602=>"010010011",
  34603=>"000000001",
  34604=>"011110100",
  34605=>"000000110",
  34606=>"111110111",
  34607=>"011101101",
  34608=>"111001100",
  34609=>"111101100",
  34610=>"000100001",
  34611=>"101011001",
  34612=>"010010010",
  34613=>"101110111",
  34614=>"000110100",
  34615=>"101000110",
  34616=>"011010110",
  34617=>"101011000",
  34618=>"101001111",
  34619=>"000000001",
  34620=>"100001100",
  34621=>"010001100",
  34622=>"001101010",
  34623=>"001000100",
  34624=>"010100000",
  34625=>"001010101",
  34626=>"101011111",
  34627=>"011001111",
  34628=>"000000011",
  34629=>"011100001",
  34630=>"010011010",
  34631=>"111110100",
  34632=>"000000001",
  34633=>"011110001",
  34634=>"001010010",
  34635=>"000100001",
  34636=>"001100100",
  34637=>"010110110",
  34638=>"001001011",
  34639=>"111001010",
  34640=>"101000001",
  34641=>"111011100",
  34642=>"001011111",
  34643=>"111001111",
  34644=>"000011101",
  34645=>"111000110",
  34646=>"101100000",
  34647=>"100101101",
  34648=>"101001000",
  34649=>"001100110",
  34650=>"011011101",
  34651=>"100110101",
  34652=>"111111101",
  34653=>"110111011",
  34654=>"110010100",
  34655=>"001101100",
  34656=>"100011010",
  34657=>"000000011",
  34658=>"000100001",
  34659=>"000001110",
  34660=>"010100000",
  34661=>"000011011",
  34662=>"000001111",
  34663=>"111011111",
  34664=>"000101000",
  34665=>"010111000",
  34666=>"110111011",
  34667=>"110010101",
  34668=>"110111111",
  34669=>"101010011",
  34670=>"111010111",
  34671=>"000010000",
  34672=>"000100100",
  34673=>"101101110",
  34674=>"101110010",
  34675=>"111111011",
  34676=>"101100100",
  34677=>"001000001",
  34678=>"111100000",
  34679=>"011101100",
  34680=>"000111001",
  34681=>"110111101",
  34682=>"010001111",
  34683=>"110011000",
  34684=>"000001110",
  34685=>"111010100",
  34686=>"000000100",
  34687=>"001000101",
  34688=>"101000100",
  34689=>"000100000",
  34690=>"110101000",
  34691=>"101001101",
  34692=>"000000000",
  34693=>"011101101",
  34694=>"110000111",
  34695=>"011101101",
  34696=>"111011001",
  34697=>"000011000",
  34698=>"100000100",
  34699=>"100011001",
  34700=>"100111100",
  34701=>"101001101",
  34702=>"000000100",
  34703=>"110011000",
  34704=>"111100110",
  34705=>"101101100",
  34706=>"010000010",
  34707=>"101010110",
  34708=>"101101100",
  34709=>"111111000",
  34710=>"001000100",
  34711=>"110000100",
  34712=>"010000000",
  34713=>"000010011",
  34714=>"011111110",
  34715=>"011101011",
  34716=>"011100001",
  34717=>"001110111",
  34718=>"001000010",
  34719=>"100011000",
  34720=>"110101010",
  34721=>"011001110",
  34722=>"110000011",
  34723=>"111011101",
  34724=>"000000110",
  34725=>"101101111",
  34726=>"010010111",
  34727=>"001111010",
  34728=>"011000000",
  34729=>"101000111",
  34730=>"101100011",
  34731=>"010000010",
  34732=>"000110001",
  34733=>"010010000",
  34734=>"000000100",
  34735=>"110000010",
  34736=>"100000111",
  34737=>"111010110",
  34738=>"101001100",
  34739=>"101100010",
  34740=>"110110011",
  34741=>"000111101",
  34742=>"110100101",
  34743=>"110001110",
  34744=>"100110000",
  34745=>"001100110",
  34746=>"001001100",
  34747=>"110110100",
  34748=>"001100110",
  34749=>"101010010",
  34750=>"011001010",
  34751=>"011100111",
  34752=>"110010000",
  34753=>"100101111",
  34754=>"111101101",
  34755=>"001100001",
  34756=>"111100001",
  34757=>"111001000",
  34758=>"100111001",
  34759=>"000111111",
  34760=>"000011011",
  34761=>"110111100",
  34762=>"001100100",
  34763=>"100110010",
  34764=>"001011110",
  34765=>"101101110",
  34766=>"111111111",
  34767=>"001011101",
  34768=>"010101101",
  34769=>"111111100",
  34770=>"100001100",
  34771=>"000000100",
  34772=>"000011010",
  34773=>"110010000",
  34774=>"111001110",
  34775=>"001011110",
  34776=>"100001001",
  34777=>"111011110",
  34778=>"110011101",
  34779=>"000100010",
  34780=>"001100101",
  34781=>"001001100",
  34782=>"101011111",
  34783=>"110010011",
  34784=>"100111000",
  34785=>"000110001",
  34786=>"010110000",
  34787=>"101100110",
  34788=>"010100010",
  34789=>"111111000",
  34790=>"001010000",
  34791=>"101001011",
  34792=>"000011000",
  34793=>"110010100",
  34794=>"000001101",
  34795=>"101010010",
  34796=>"011000110",
  34797=>"100011010",
  34798=>"011001010",
  34799=>"011011001",
  34800=>"010110111",
  34801=>"101010101",
  34802=>"101110100",
  34803=>"001100110",
  34804=>"111010011",
  34805=>"110000010",
  34806=>"010111010",
  34807=>"101111000",
  34808=>"100011001",
  34809=>"111000010",
  34810=>"101101101",
  34811=>"000100110",
  34812=>"010010011",
  34813=>"100101000",
  34814=>"011100000",
  34815=>"100110000",
  34816=>"000011101",
  34817=>"011111010",
  34818=>"010101000",
  34819=>"100011110",
  34820=>"001000101",
  34821=>"101110001",
  34822=>"001100011",
  34823=>"100111011",
  34824=>"010000110",
  34825=>"011010001",
  34826=>"000111010",
  34827=>"111001011",
  34828=>"001001100",
  34829=>"111011111",
  34830=>"110000011",
  34831=>"101000010",
  34832=>"010001011",
  34833=>"000111000",
  34834=>"100010101",
  34835=>"000111000",
  34836=>"001111101",
  34837=>"111001001",
  34838=>"011010101",
  34839=>"000101000",
  34840=>"001000000",
  34841=>"101010000",
  34842=>"011000111",
  34843=>"001110010",
  34844=>"011110000",
  34845=>"100001110",
  34846=>"101000011",
  34847=>"010000111",
  34848=>"001000001",
  34849=>"010001011",
  34850=>"011111001",
  34851=>"001001001",
  34852=>"011111000",
  34853=>"101101111",
  34854=>"011100000",
  34855=>"001010000",
  34856=>"110000001",
  34857=>"110011111",
  34858=>"000110001",
  34859=>"100000011",
  34860=>"111001100",
  34861=>"110010001",
  34862=>"100101001",
  34863=>"000100100",
  34864=>"001110100",
  34865=>"001101110",
  34866=>"010001111",
  34867=>"111000110",
  34868=>"100010101",
  34869=>"100000110",
  34870=>"110111011",
  34871=>"000000001",
  34872=>"100110111",
  34873=>"101100010",
  34874=>"111100001",
  34875=>"010010101",
  34876=>"000011111",
  34877=>"011010001",
  34878=>"110001011",
  34879=>"111100101",
  34880=>"001011100",
  34881=>"000110101",
  34882=>"101000010",
  34883=>"011001000",
  34884=>"101100100",
  34885=>"100011000",
  34886=>"011101111",
  34887=>"111010100",
  34888=>"010011000",
  34889=>"101111110",
  34890=>"001001010",
  34891=>"001011011",
  34892=>"011010111",
  34893=>"110101100",
  34894=>"101100111",
  34895=>"010100110",
  34896=>"011100101",
  34897=>"111101100",
  34898=>"100000100",
  34899=>"000011000",
  34900=>"000110111",
  34901=>"100100011",
  34902=>"011111100",
  34903=>"100010100",
  34904=>"000100001",
  34905=>"000000111",
  34906=>"010000111",
  34907=>"010010010",
  34908=>"110000111",
  34909=>"000100111",
  34910=>"000000100",
  34911=>"110111110",
  34912=>"011111011",
  34913=>"010100000",
  34914=>"001111111",
  34915=>"111111101",
  34916=>"011001111",
  34917=>"000000000",
  34918=>"110100100",
  34919=>"000010000",
  34920=>"010010001",
  34921=>"110011110",
  34922=>"110101011",
  34923=>"101001011",
  34924=>"111111100",
  34925=>"010011110",
  34926=>"100010011",
  34927=>"100010000",
  34928=>"100010000",
  34929=>"011100100",
  34930=>"001010111",
  34931=>"100010101",
  34932=>"111001010",
  34933=>"011010001",
  34934=>"010010110",
  34935=>"100100111",
  34936=>"111100000",
  34937=>"010101001",
  34938=>"010110001",
  34939=>"100110000",
  34940=>"101100101",
  34941=>"111101001",
  34942=>"010110001",
  34943=>"010000010",
  34944=>"111010000",
  34945=>"001110011",
  34946=>"010011001",
  34947=>"100010001",
  34948=>"111101001",
  34949=>"100010100",
  34950=>"000001110",
  34951=>"111101010",
  34952=>"000101010",
  34953=>"000111110",
  34954=>"000000000",
  34955=>"000111111",
  34956=>"000101100",
  34957=>"100101000",
  34958=>"111110100",
  34959=>"111000000",
  34960=>"100011111",
  34961=>"010111000",
  34962=>"101110011",
  34963=>"001001001",
  34964=>"110000111",
  34965=>"001100101",
  34966=>"000010000",
  34967=>"101101001",
  34968=>"011000011",
  34969=>"010101000",
  34970=>"001100101",
  34971=>"001000111",
  34972=>"010010100",
  34973=>"111000000",
  34974=>"111011111",
  34975=>"111010101",
  34976=>"001000001",
  34977=>"011100110",
  34978=>"111001100",
  34979=>"001001101",
  34980=>"010111110",
  34981=>"111011001",
  34982=>"101001100",
  34983=>"011010110",
  34984=>"111110110",
  34985=>"110011011",
  34986=>"011001101",
  34987=>"001111000",
  34988=>"111111010",
  34989=>"111110101",
  34990=>"000000111",
  34991=>"101010000",
  34992=>"101100111",
  34993=>"001101110",
  34994=>"010000111",
  34995=>"010000000",
  34996=>"100010101",
  34997=>"001110001",
  34998=>"010011000",
  34999=>"101010010",
  35000=>"011001000",
  35001=>"000010100",
  35002=>"100000000",
  35003=>"011110011",
  35004=>"111000110",
  35005=>"010010010",
  35006=>"100111000",
  35007=>"010101111",
  35008=>"010010110",
  35009=>"110000001",
  35010=>"001111000",
  35011=>"101000110",
  35012=>"101000001",
  35013=>"001010000",
  35014=>"000101101",
  35015=>"110110110",
  35016=>"011000001",
  35017=>"101101111",
  35018=>"101111100",
  35019=>"111001101",
  35020=>"100001101",
  35021=>"111001000",
  35022=>"010010001",
  35023=>"011110000",
  35024=>"111111100",
  35025=>"100000101",
  35026=>"101000000",
  35027=>"111000110",
  35028=>"010100101",
  35029=>"101100111",
  35030=>"000111101",
  35031=>"110100111",
  35032=>"010110100",
  35033=>"000100100",
  35034=>"000001101",
  35035=>"101000101",
  35036=>"001101011",
  35037=>"110101000",
  35038=>"000000111",
  35039=>"110110000",
  35040=>"110100110",
  35041=>"010001101",
  35042=>"010111110",
  35043=>"101010010",
  35044=>"111111001",
  35045=>"101000110",
  35046=>"001111011",
  35047=>"000111101",
  35048=>"000010100",
  35049=>"011000011",
  35050=>"110001100",
  35051=>"110001001",
  35052=>"011001001",
  35053=>"100100010",
  35054=>"010000100",
  35055=>"000011001",
  35056=>"100111011",
  35057=>"111100000",
  35058=>"000011010",
  35059=>"011011011",
  35060=>"011110111",
  35061=>"111110001",
  35062=>"101010110",
  35063=>"101001000",
  35064=>"010100101",
  35065=>"100101000",
  35066=>"101001110",
  35067=>"010001001",
  35068=>"010010110",
  35069=>"011000001",
  35070=>"100111010",
  35071=>"000010001",
  35072=>"010111100",
  35073=>"001111111",
  35074=>"101101011",
  35075=>"001000111",
  35076=>"111110101",
  35077=>"001110111",
  35078=>"000011111",
  35079=>"101100101",
  35080=>"110110110",
  35081=>"101010110",
  35082=>"110000000",
  35083=>"001000000",
  35084=>"011110100",
  35085=>"101011101",
  35086=>"100101010",
  35087=>"001111111",
  35088=>"000010000",
  35089=>"110100101",
  35090=>"111111101",
  35091=>"010101001",
  35092=>"011100110",
  35093=>"011100011",
  35094=>"011001101",
  35095=>"000111010",
  35096=>"100101101",
  35097=>"110100000",
  35098=>"010001110",
  35099=>"101110110",
  35100=>"101000010",
  35101=>"100110010",
  35102=>"110001110",
  35103=>"010000111",
  35104=>"100000000",
  35105=>"100001001",
  35106=>"001000001",
  35107=>"101001100",
  35108=>"011001001",
  35109=>"111110000",
  35110=>"111111001",
  35111=>"100011111",
  35112=>"000111101",
  35113=>"111101010",
  35114=>"000001101",
  35115=>"010110110",
  35116=>"101000101",
  35117=>"011001011",
  35118=>"001101011",
  35119=>"111100111",
  35120=>"100001100",
  35121=>"111001011",
  35122=>"101011001",
  35123=>"110111111",
  35124=>"111101111",
  35125=>"000001000",
  35126=>"111101010",
  35127=>"110111100",
  35128=>"000000011",
  35129=>"010101000",
  35130=>"000010000",
  35131=>"000110001",
  35132=>"000011000",
  35133=>"011011110",
  35134=>"001101101",
  35135=>"101110101",
  35136=>"001110011",
  35137=>"111011110",
  35138=>"000001101",
  35139=>"011101110",
  35140=>"000001101",
  35141=>"010000101",
  35142=>"101000000",
  35143=>"010100100",
  35144=>"001010101",
  35145=>"100010000",
  35146=>"011101111",
  35147=>"010111010",
  35148=>"001101011",
  35149=>"010101111",
  35150=>"011000011",
  35151=>"000001000",
  35152=>"011010011",
  35153=>"110110100",
  35154=>"010111000",
  35155=>"001000010",
  35156=>"111011000",
  35157=>"010110011",
  35158=>"110100101",
  35159=>"100110111",
  35160=>"001110010",
  35161=>"011011011",
  35162=>"100011110",
  35163=>"110011000",
  35164=>"110110101",
  35165=>"100111101",
  35166=>"000011001",
  35167=>"000101001",
  35168=>"001111001",
  35169=>"101001101",
  35170=>"010101111",
  35171=>"001000101",
  35172=>"100001011",
  35173=>"001101001",
  35174=>"101111110",
  35175=>"111101010",
  35176=>"111011010",
  35177=>"010011010",
  35178=>"011010101",
  35179=>"000111000",
  35180=>"010110000",
  35181=>"001101001",
  35182=>"000010010",
  35183=>"110000111",
  35184=>"001100000",
  35185=>"000100100",
  35186=>"011000011",
  35187=>"100110111",
  35188=>"101101000",
  35189=>"110001100",
  35190=>"001110001",
  35191=>"010000100",
  35192=>"001101101",
  35193=>"100100100",
  35194=>"100110011",
  35195=>"110011111",
  35196=>"000000010",
  35197=>"111111101",
  35198=>"000111000",
  35199=>"110001101",
  35200=>"101011000",
  35201=>"000001101",
  35202=>"111000010",
  35203=>"101000011",
  35204=>"100101110",
  35205=>"001100101",
  35206=>"101011100",
  35207=>"100110000",
  35208=>"000110000",
  35209=>"111111101",
  35210=>"111110011",
  35211=>"000100011",
  35212=>"001101010",
  35213=>"010100100",
  35214=>"111111100",
  35215=>"010010111",
  35216=>"011010110",
  35217=>"100000111",
  35218=>"100111011",
  35219=>"100011001",
  35220=>"111110110",
  35221=>"110101100",
  35222=>"100000000",
  35223=>"010010101",
  35224=>"011110000",
  35225=>"011010000",
  35226=>"100111010",
  35227=>"011100001",
  35228=>"100001100",
  35229=>"010001100",
  35230=>"110011111",
  35231=>"001011001",
  35232=>"001000111",
  35233=>"010001001",
  35234=>"111101001",
  35235=>"100100000",
  35236=>"010001011",
  35237=>"011001101",
  35238=>"110100101",
  35239=>"111111110",
  35240=>"101010011",
  35241=>"100101110",
  35242=>"000010101",
  35243=>"101110100",
  35244=>"000100100",
  35245=>"010110001",
  35246=>"010001001",
  35247=>"111110000",
  35248=>"101011000",
  35249=>"110000111",
  35250=>"100010010",
  35251=>"101000110",
  35252=>"110000111",
  35253=>"000001011",
  35254=>"010001101",
  35255=>"110111101",
  35256=>"101000100",
  35257=>"111110001",
  35258=>"100111010",
  35259=>"010110110",
  35260=>"111110110",
  35261=>"111101111",
  35262=>"100111110",
  35263=>"100001001",
  35264=>"010011010",
  35265=>"000100011",
  35266=>"011000110",
  35267=>"111010010",
  35268=>"011101110",
  35269=>"111110001",
  35270=>"000111011",
  35271=>"010010000",
  35272=>"010011001",
  35273=>"010010011",
  35274=>"011001100",
  35275=>"111011000",
  35276=>"000010100",
  35277=>"101111010",
  35278=>"100101111",
  35279=>"011000000",
  35280=>"110011101",
  35281=>"000001100",
  35282=>"011111110",
  35283=>"110010011",
  35284=>"001110000",
  35285=>"101000000",
  35286=>"101101000",
  35287=>"010000111",
  35288=>"000100101",
  35289=>"000000000",
  35290=>"111111011",
  35291=>"011001001",
  35292=>"010010001",
  35293=>"101010000",
  35294=>"000000010",
  35295=>"101110010",
  35296=>"100010010",
  35297=>"111101000",
  35298=>"000000100",
  35299=>"001011001",
  35300=>"001101101",
  35301=>"000101010",
  35302=>"110111011",
  35303=>"111000000",
  35304=>"011001010",
  35305=>"010011100",
  35306=>"000100111",
  35307=>"111100001",
  35308=>"010000001",
  35309=>"011000110",
  35310=>"010111000",
  35311=>"101100000",
  35312=>"111000011",
  35313=>"111010011",
  35314=>"111010000",
  35315=>"000100001",
  35316=>"110111010",
  35317=>"001000001",
  35318=>"010001001",
  35319=>"111000101",
  35320=>"000011010",
  35321=>"111001100",
  35322=>"101010100",
  35323=>"000101110",
  35324=>"010000110",
  35325=>"100111001",
  35326=>"100100111",
  35327=>"000001111",
  35328=>"110101001",
  35329=>"110100111",
  35330=>"111000011",
  35331=>"011011101",
  35332=>"011000001",
  35333=>"111000111",
  35334=>"101000011",
  35335=>"100011010",
  35336=>"000010101",
  35337=>"001001111",
  35338=>"010010011",
  35339=>"111001011",
  35340=>"011000100",
  35341=>"001001000",
  35342=>"101001000",
  35343=>"011100101",
  35344=>"100010011",
  35345=>"001010001",
  35346=>"010100001",
  35347=>"111011101",
  35348=>"101001111",
  35349=>"001100000",
  35350=>"001110000",
  35351=>"010101101",
  35352=>"010011110",
  35353=>"010110010",
  35354=>"101110110",
  35355=>"101010100",
  35356=>"101111001",
  35357=>"110100011",
  35358=>"010000101",
  35359=>"000000011",
  35360=>"101010001",
  35361=>"000100100",
  35362=>"010001001",
  35363=>"111011000",
  35364=>"100000111",
  35365=>"111101011",
  35366=>"010000111",
  35367=>"110110111",
  35368=>"000010100",
  35369=>"111111111",
  35370=>"110110001",
  35371=>"000111010",
  35372=>"111000110",
  35373=>"011001001",
  35374=>"001010110",
  35375=>"001110011",
  35376=>"111100111",
  35377=>"010100110",
  35378=>"000011011",
  35379=>"010000001",
  35380=>"000010011",
  35381=>"111001011",
  35382=>"010010101",
  35383=>"001111100",
  35384=>"000101000",
  35385=>"010110000",
  35386=>"101001011",
  35387=>"011110110",
  35388=>"011111100",
  35389=>"001000111",
  35390=>"110001001",
  35391=>"000011011",
  35392=>"000000110",
  35393=>"111001010",
  35394=>"111000001",
  35395=>"011001110",
  35396=>"001100111",
  35397=>"101110101",
  35398=>"000001001",
  35399=>"110001111",
  35400=>"011111001",
  35401=>"111111010",
  35402=>"010010010",
  35403=>"010011110",
  35404=>"001000111",
  35405=>"000000001",
  35406=>"001001000",
  35407=>"010100000",
  35408=>"010110000",
  35409=>"010010110",
  35410=>"001011110",
  35411=>"101000100",
  35412=>"001110111",
  35413=>"000010000",
  35414=>"100001100",
  35415=>"011010001",
  35416=>"000011101",
  35417=>"001100111",
  35418=>"001011000",
  35419=>"001110011",
  35420=>"011010001",
  35421=>"100010000",
  35422=>"000101010",
  35423=>"011110100",
  35424=>"010101011",
  35425=>"000100000",
  35426=>"000000000",
  35427=>"101001001",
  35428=>"001111001",
  35429=>"100100011",
  35430=>"100111101",
  35431=>"010010100",
  35432=>"111110111",
  35433=>"100100000",
  35434=>"101111011",
  35435=>"110100010",
  35436=>"101110101",
  35437=>"000010101",
  35438=>"110010111",
  35439=>"101100011",
  35440=>"101100011",
  35441=>"100000001",
  35442=>"101001111",
  35443=>"111001110",
  35444=>"001110001",
  35445=>"110100000",
  35446=>"100111011",
  35447=>"011010010",
  35448=>"000111000",
  35449=>"001111000",
  35450=>"010100100",
  35451=>"111100001",
  35452=>"100011010",
  35453=>"110110110",
  35454=>"111000101",
  35455=>"101100111",
  35456=>"011000111",
  35457=>"111010011",
  35458=>"101001011",
  35459=>"011011101",
  35460=>"001110001",
  35461=>"000111000",
  35462=>"000111111",
  35463=>"000100000",
  35464=>"100111111",
  35465=>"100101000",
  35466=>"010110111",
  35467=>"111100011",
  35468=>"101011000",
  35469=>"010000010",
  35470=>"111010011",
  35471=>"010010110",
  35472=>"110000000",
  35473=>"000010001",
  35474=>"101001010",
  35475=>"000101101",
  35476=>"001110100",
  35477=>"110000001",
  35478=>"111101011",
  35479=>"101010000",
  35480=>"111000111",
  35481=>"010001000",
  35482=>"001110101",
  35483=>"011000011",
  35484=>"110010110",
  35485=>"111111011",
  35486=>"111011000",
  35487=>"100101000",
  35488=>"001011001",
  35489=>"110001011",
  35490=>"110000101",
  35491=>"101110101",
  35492=>"000110101",
  35493=>"000110110",
  35494=>"001101111",
  35495=>"001011111",
  35496=>"110011000",
  35497=>"010010001",
  35498=>"010101010",
  35499=>"100110001",
  35500=>"111011010",
  35501=>"001000011",
  35502=>"000001100",
  35503=>"001000111",
  35504=>"110111111",
  35505=>"000110000",
  35506=>"101000000",
  35507=>"001111011",
  35508=>"000101000",
  35509=>"000100011",
  35510=>"110100011",
  35511=>"011101001",
  35512=>"000100001",
  35513=>"110000010",
  35514=>"111111001",
  35515=>"111100111",
  35516=>"011101011",
  35517=>"101000111",
  35518=>"111010001",
  35519=>"000010010",
  35520=>"100111101",
  35521=>"100110110",
  35522=>"001100101",
  35523=>"100000110",
  35524=>"000001101",
  35525=>"101011101",
  35526=>"100001011",
  35527=>"000010011",
  35528=>"111101010",
  35529=>"101001100",
  35530=>"011110001",
  35531=>"101000011",
  35532=>"110111000",
  35533=>"011101101",
  35534=>"000010000",
  35535=>"010000101",
  35536=>"110100010",
  35537=>"100110110",
  35538=>"101000010",
  35539=>"111010111",
  35540=>"110110001",
  35541=>"001101011",
  35542=>"001110001",
  35543=>"100010111",
  35544=>"100101111",
  35545=>"100000100",
  35546=>"111101000",
  35547=>"010011111",
  35548=>"101010001",
  35549=>"110101000",
  35550=>"010101110",
  35551=>"101010011",
  35552=>"000101000",
  35553=>"011010111",
  35554=>"000110100",
  35555=>"110101101",
  35556=>"001100110",
  35557=>"011100110",
  35558=>"011000001",
  35559=>"010101100",
  35560=>"010000000",
  35561=>"110001100",
  35562=>"000101010",
  35563=>"011110101",
  35564=>"010100100",
  35565=>"101001010",
  35566=>"011010100",
  35567=>"100001101",
  35568=>"010111111",
  35569=>"100100111",
  35570=>"010011010",
  35571=>"110111011",
  35572=>"101011000",
  35573=>"001001001",
  35574=>"111111110",
  35575=>"110100010",
  35576=>"110001101",
  35577=>"010010001",
  35578=>"101101100",
  35579=>"101000001",
  35580=>"001110011",
  35581=>"000001111",
  35582=>"110100001",
  35583=>"110100010",
  35584=>"111000100",
  35585=>"000010101",
  35586=>"110110100",
  35587=>"010000010",
  35588=>"011101111",
  35589=>"000011111",
  35590=>"100001010",
  35591=>"110101010",
  35592=>"100010000",
  35593=>"010011111",
  35594=>"001111101",
  35595=>"101110000",
  35596=>"010000101",
  35597=>"010000101",
  35598=>"001111011",
  35599=>"100011000",
  35600=>"010110011",
  35601=>"000010010",
  35602=>"010000001",
  35603=>"011001000",
  35604=>"111100101",
  35605=>"111010001",
  35606=>"100011000",
  35607=>"100001101",
  35608=>"100111011",
  35609=>"101000111",
  35610=>"101110111",
  35611=>"010010000",
  35612=>"000000111",
  35613=>"010101101",
  35614=>"100111110",
  35615=>"011001001",
  35616=>"000101000",
  35617=>"100001010",
  35618=>"011111000",
  35619=>"100010101",
  35620=>"100110100",
  35621=>"110111101",
  35622=>"100000111",
  35623=>"010011010",
  35624=>"111100111",
  35625=>"110101110",
  35626=>"010000001",
  35627=>"111011111",
  35628=>"111111001",
  35629=>"101000000",
  35630=>"000001111",
  35631=>"110101110",
  35632=>"000110000",
  35633=>"001111000",
  35634=>"001010000",
  35635=>"000101100",
  35636=>"100011010",
  35637=>"101001111",
  35638=>"000000101",
  35639=>"001110000",
  35640=>"111110011",
  35641=>"000110100",
  35642=>"001110100",
  35643=>"111110001",
  35644=>"111011000",
  35645=>"001101110",
  35646=>"111110001",
  35647=>"001110011",
  35648=>"100110010",
  35649=>"000111010",
  35650=>"111011011",
  35651=>"110011000",
  35652=>"111111111",
  35653=>"000110111",
  35654=>"000010101",
  35655=>"010101110",
  35656=>"100010101",
  35657=>"111100000",
  35658=>"000001101",
  35659=>"001110101",
  35660=>"001000011",
  35661=>"001010000",
  35662=>"100010000",
  35663=>"001101110",
  35664=>"010100110",
  35665=>"101011100",
  35666=>"101111101",
  35667=>"000000100",
  35668=>"010001110",
  35669=>"000010001",
  35670=>"101010000",
  35671=>"011011000",
  35672=>"101111011",
  35673=>"110000001",
  35674=>"100110000",
  35675=>"011101000",
  35676=>"100001111",
  35677=>"110101111",
  35678=>"100101010",
  35679=>"100101001",
  35680=>"110110100",
  35681=>"000011010",
  35682=>"110100000",
  35683=>"000110000",
  35684=>"000111010",
  35685=>"110111100",
  35686=>"010011111",
  35687=>"000011110",
  35688=>"001001000",
  35689=>"111101101",
  35690=>"000101000",
  35691=>"110110100",
  35692=>"010000010",
  35693=>"011101001",
  35694=>"100010110",
  35695=>"101011101",
  35696=>"011010011",
  35697=>"011111001",
  35698=>"011111011",
  35699=>"001010000",
  35700=>"100011111",
  35701=>"011011100",
  35702=>"111001110",
  35703=>"010001000",
  35704=>"001011010",
  35705=>"101110111",
  35706=>"010011100",
  35707=>"111111110",
  35708=>"001010010",
  35709=>"100001001",
  35710=>"010100111",
  35711=>"010111100",
  35712=>"000100110",
  35713=>"100001010",
  35714=>"000011000",
  35715=>"010010111",
  35716=>"011000011",
  35717=>"001000001",
  35718=>"000100011",
  35719=>"100001010",
  35720=>"101001010",
  35721=>"000000001",
  35722=>"100101010",
  35723=>"010000111",
  35724=>"010101110",
  35725=>"000101010",
  35726=>"001100101",
  35727=>"100110011",
  35728=>"010010110",
  35729=>"100101011",
  35730=>"100000100",
  35731=>"100001011",
  35732=>"101001011",
  35733=>"011111001",
  35734=>"000001010",
  35735=>"011101101",
  35736=>"011011111",
  35737=>"010001101",
  35738=>"001001010",
  35739=>"000000100",
  35740=>"001111101",
  35741=>"010111110",
  35742=>"011100010",
  35743=>"011100010",
  35744=>"010101001",
  35745=>"110010001",
  35746=>"000000000",
  35747=>"110100000",
  35748=>"110000101",
  35749=>"001110011",
  35750=>"001110010",
  35751=>"010111000",
  35752=>"011010010",
  35753=>"010100010",
  35754=>"011101111",
  35755=>"111101011",
  35756=>"100000000",
  35757=>"010000000",
  35758=>"011111100",
  35759=>"100000101",
  35760=>"110011111",
  35761=>"111101000",
  35762=>"010001010",
  35763=>"110111111",
  35764=>"000010110",
  35765=>"110000111",
  35766=>"001110101",
  35767=>"111000100",
  35768=>"100100001",
  35769=>"010000100",
  35770=>"011000111",
  35771=>"001010110",
  35772=>"110000100",
  35773=>"000011101",
  35774=>"010111101",
  35775=>"110000101",
  35776=>"010011101",
  35777=>"011010010",
  35778=>"001110111",
  35779=>"001100110",
  35780=>"000010110",
  35781=>"000100011",
  35782=>"010101010",
  35783=>"111001100",
  35784=>"010110111",
  35785=>"010110011",
  35786=>"111110101",
  35787=>"011000101",
  35788=>"110000111",
  35789=>"001011010",
  35790=>"010100111",
  35791=>"001001001",
  35792=>"001101111",
  35793=>"011110011",
  35794=>"000010111",
  35795=>"101001111",
  35796=>"010000111",
  35797=>"001011101",
  35798=>"001111010",
  35799=>"001011111",
  35800=>"101110101",
  35801=>"010000111",
  35802=>"110111001",
  35803=>"001000111",
  35804=>"010101101",
  35805=>"011100011",
  35806=>"100100000",
  35807=>"100001001",
  35808=>"000000110",
  35809=>"001000010",
  35810=>"000111011",
  35811=>"000110010",
  35812=>"010010101",
  35813=>"000010011",
  35814=>"111010011",
  35815=>"111010101",
  35816=>"000101001",
  35817=>"100100011",
  35818=>"001010000",
  35819=>"111011010",
  35820=>"111100110",
  35821=>"001010111",
  35822=>"011111101",
  35823=>"100000111",
  35824=>"000001010",
  35825=>"000000001",
  35826=>"110000110",
  35827=>"111010001",
  35828=>"110001100",
  35829=>"111100100",
  35830=>"101110100",
  35831=>"100100000",
  35832=>"001111000",
  35833=>"100101111",
  35834=>"101110010",
  35835=>"111111011",
  35836=>"010010110",
  35837=>"000101011",
  35838=>"011101111",
  35839=>"000100101",
  35840=>"011001101",
  35841=>"011001011",
  35842=>"100111110",
  35843=>"010010101",
  35844=>"010000100",
  35845=>"011001010",
  35846=>"100001011",
  35847=>"101011000",
  35848=>"010100110",
  35849=>"111011010",
  35850=>"001110110",
  35851=>"000101010",
  35852=>"000000011",
  35853=>"011011001",
  35854=>"100110100",
  35855=>"111000110",
  35856=>"100101011",
  35857=>"010010100",
  35858=>"100110100",
  35859=>"101001110",
  35860=>"000111010",
  35861=>"000101011",
  35862=>"011100011",
  35863=>"001111011",
  35864=>"100110001",
  35865=>"011110011",
  35866=>"110000111",
  35867=>"110000000",
  35868=>"111000110",
  35869=>"111001111",
  35870=>"010101000",
  35871=>"100100001",
  35872=>"101010101",
  35873=>"010111010",
  35874=>"110011100",
  35875=>"011111111",
  35876=>"101011101",
  35877=>"001001100",
  35878=>"101100000",
  35879=>"110111011",
  35880=>"010111111",
  35881=>"110111001",
  35882=>"111001000",
  35883=>"000111111",
  35884=>"100111100",
  35885=>"000111100",
  35886=>"000111010",
  35887=>"110100011",
  35888=>"101100000",
  35889=>"000101001",
  35890=>"111000000",
  35891=>"100100001",
  35892=>"100110001",
  35893=>"000111100",
  35894=>"110001011",
  35895=>"110101110",
  35896=>"101101111",
  35897=>"001100100",
  35898=>"001001111",
  35899=>"101101110",
  35900=>"111000011",
  35901=>"111011001",
  35902=>"110100101",
  35903=>"111110101",
  35904=>"101010001",
  35905=>"101011000",
  35906=>"111111000",
  35907=>"010011001",
  35908=>"100010110",
  35909=>"101101110",
  35910=>"010000101",
  35911=>"011110010",
  35912=>"110000101",
  35913=>"000100110",
  35914=>"001011000",
  35915=>"110010011",
  35916=>"101000000",
  35917=>"100000100",
  35918=>"101010011",
  35919=>"000111111",
  35920=>"100010000",
  35921=>"111100111",
  35922=>"101011010",
  35923=>"110000010",
  35924=>"101101000",
  35925=>"101101100",
  35926=>"001110111",
  35927=>"011100000",
  35928=>"101010010",
  35929=>"110011101",
  35930=>"000001110",
  35931=>"001111001",
  35932=>"111000100",
  35933=>"000010011",
  35934=>"001111111",
  35935=>"001110011",
  35936=>"111000101",
  35937=>"011011110",
  35938=>"001000101",
  35939=>"000110001",
  35940=>"001010011",
  35941=>"111101100",
  35942=>"101101011",
  35943=>"101010000",
  35944=>"001001101",
  35945=>"100000111",
  35946=>"000010010",
  35947=>"001001010",
  35948=>"111101111",
  35949=>"101011110",
  35950=>"010000111",
  35951=>"110000001",
  35952=>"100011000",
  35953=>"000001110",
  35954=>"111000010",
  35955=>"100110110",
  35956=>"001110100",
  35957=>"101100101",
  35958=>"110001110",
  35959=>"000111110",
  35960=>"110101100",
  35961=>"010111110",
  35962=>"011110111",
  35963=>"001000100",
  35964=>"101100010",
  35965=>"010001111",
  35966=>"110111000",
  35967=>"100101110",
  35968=>"100000000",
  35969=>"001101001",
  35970=>"011000100",
  35971=>"010110011",
  35972=>"001101000",
  35973=>"100101010",
  35974=>"000100111",
  35975=>"011101010",
  35976=>"010111011",
  35977=>"000010101",
  35978=>"101000101",
  35979=>"110100110",
  35980=>"101100101",
  35981=>"010010111",
  35982=>"010001100",
  35983=>"100010000",
  35984=>"001011011",
  35985=>"001001001",
  35986=>"010010010",
  35987=>"000000011",
  35988=>"001001111",
  35989=>"101101100",
  35990=>"111011001",
  35991=>"110100100",
  35992=>"000110001",
  35993=>"011011110",
  35994=>"000010110",
  35995=>"101000010",
  35996=>"000101110",
  35997=>"010100010",
  35998=>"001010000",
  35999=>"000011000",
  36000=>"010100000",
  36001=>"111110111",
  36002=>"110000100",
  36003=>"110100010",
  36004=>"001110010",
  36005=>"100100100",
  36006=>"001010000",
  36007=>"110000110",
  36008=>"001011101",
  36009=>"100100011",
  36010=>"010110010",
  36011=>"110001000",
  36012=>"101111110",
  36013=>"100100111",
  36014=>"011000110",
  36015=>"101000011",
  36016=>"011011000",
  36017=>"101000011",
  36018=>"011011001",
  36019=>"000000011",
  36020=>"101110101",
  36021=>"001111001",
  36022=>"111100011",
  36023=>"011101101",
  36024=>"110110110",
  36025=>"101111110",
  36026=>"110110010",
  36027=>"011100100",
  36028=>"011101011",
  36029=>"000000110",
  36030=>"100000100",
  36031=>"100010101",
  36032=>"101100110",
  36033=>"100010011",
  36034=>"001100111",
  36035=>"101100101",
  36036=>"010100101",
  36037=>"001110111",
  36038=>"101000000",
  36039=>"111100110",
  36040=>"001101101",
  36041=>"110011001",
  36042=>"000100010",
  36043=>"111010101",
  36044=>"101001000",
  36045=>"111101100",
  36046=>"011101110",
  36047=>"101011001",
  36048=>"000100000",
  36049=>"011110111",
  36050=>"100011101",
  36051=>"000011101",
  36052=>"111001110",
  36053=>"101101101",
  36054=>"110001010",
  36055=>"110011010",
  36056=>"100111101",
  36057=>"101111110",
  36058=>"011110011",
  36059=>"101111111",
  36060=>"000110100",
  36061=>"100101000",
  36062=>"100101000",
  36063=>"101000100",
  36064=>"000010110",
  36065=>"101011111",
  36066=>"111011000",
  36067=>"011001111",
  36068=>"100111100",
  36069=>"001101011",
  36070=>"011111001",
  36071=>"001110011",
  36072=>"110010000",
  36073=>"001100000",
  36074=>"110111011",
  36075=>"101110110",
  36076=>"010011101",
  36077=>"011010010",
  36078=>"111101011",
  36079=>"000101011",
  36080=>"110110100",
  36081=>"000000010",
  36082=>"010001010",
  36083=>"101010110",
  36084=>"111001000",
  36085=>"110000101",
  36086=>"101101000",
  36087=>"001000100",
  36088=>"111111011",
  36089=>"101011010",
  36090=>"111001111",
  36091=>"100000010",
  36092=>"101010010",
  36093=>"011000111",
  36094=>"111110110",
  36095=>"011011011",
  36096=>"000001010",
  36097=>"101010111",
  36098=>"101000111",
  36099=>"110101110",
  36100=>"111000000",
  36101=>"101001100",
  36102=>"001011100",
  36103=>"100010100",
  36104=>"000001011",
  36105=>"000010011",
  36106=>"010010110",
  36107=>"110110001",
  36108=>"111110111",
  36109=>"101110101",
  36110=>"111011001",
  36111=>"111010111",
  36112=>"100101010",
  36113=>"110010011",
  36114=>"100110101",
  36115=>"111010000",
  36116=>"010000011",
  36117=>"011011011",
  36118=>"001011110",
  36119=>"101000101",
  36120=>"101101001",
  36121=>"110001010",
  36122=>"111010011",
  36123=>"111101110",
  36124=>"010010101",
  36125=>"000001010",
  36126=>"100011000",
  36127=>"110001101",
  36128=>"111010001",
  36129=>"100001010",
  36130=>"000000000",
  36131=>"010110110",
  36132=>"010111011",
  36133=>"000001100",
  36134=>"011011110",
  36135=>"111011010",
  36136=>"000000100",
  36137=>"000100111",
  36138=>"001100100",
  36139=>"011011111",
  36140=>"110100010",
  36141=>"001000010",
  36142=>"000001011",
  36143=>"101110110",
  36144=>"010101101",
  36145=>"110101011",
  36146=>"010010100",
  36147=>"111110100",
  36148=>"000011110",
  36149=>"001001111",
  36150=>"001001111",
  36151=>"010111101",
  36152=>"010111011",
  36153=>"000100010",
  36154=>"000110001",
  36155=>"111001010",
  36156=>"101000101",
  36157=>"101010001",
  36158=>"110111101",
  36159=>"111111111",
  36160=>"001000000",
  36161=>"101110110",
  36162=>"001010011",
  36163=>"111011000",
  36164=>"110101101",
  36165=>"110010000",
  36166=>"100010100",
  36167=>"110100011",
  36168=>"111011000",
  36169=>"100010000",
  36170=>"100110011",
  36171=>"010010000",
  36172=>"110001010",
  36173=>"001111011",
  36174=>"011011100",
  36175=>"010111110",
  36176=>"010101110",
  36177=>"100111110",
  36178=>"011010101",
  36179=>"100110100",
  36180=>"100000011",
  36181=>"110010101",
  36182=>"011001010",
  36183=>"000101100",
  36184=>"010101001",
  36185=>"000100100",
  36186=>"011001011",
  36187=>"110101111",
  36188=>"101100110",
  36189=>"111010000",
  36190=>"100001000",
  36191=>"100110000",
  36192=>"100111000",
  36193=>"101110001",
  36194=>"111101101",
  36195=>"010001111",
  36196=>"000111011",
  36197=>"110011111",
  36198=>"111110100",
  36199=>"000110000",
  36200=>"011011011",
  36201=>"110111001",
  36202=>"111000000",
  36203=>"110010101",
  36204=>"001111110",
  36205=>"100011011",
  36206=>"001110000",
  36207=>"110111000",
  36208=>"011000111",
  36209=>"011101101",
  36210=>"100010000",
  36211=>"110010101",
  36212=>"101101001",
  36213=>"011010011",
  36214=>"100111010",
  36215=>"011010110",
  36216=>"001011010",
  36217=>"010100000",
  36218=>"100010001",
  36219=>"010101000",
  36220=>"101011100",
  36221=>"100001011",
  36222=>"001011101",
  36223=>"111110111",
  36224=>"101110101",
  36225=>"100011010",
  36226=>"111001000",
  36227=>"011101111",
  36228=>"111000011",
  36229=>"111110110",
  36230=>"011000110",
  36231=>"000101000",
  36232=>"110000011",
  36233=>"101001101",
  36234=>"101011001",
  36235=>"011100100",
  36236=>"011100001",
  36237=>"011111101",
  36238=>"010000001",
  36239=>"111100110",
  36240=>"111010000",
  36241=>"100000111",
  36242=>"110100000",
  36243=>"101000111",
  36244=>"011010100",
  36245=>"000110011",
  36246=>"101010000",
  36247=>"001100110",
  36248=>"110010110",
  36249=>"111000010",
  36250=>"010100001",
  36251=>"101110111",
  36252=>"100101100",
  36253=>"000010000",
  36254=>"011011011",
  36255=>"001000000",
  36256=>"100000000",
  36257=>"010000111",
  36258=>"010101111",
  36259=>"010000110",
  36260=>"001010111",
  36261=>"100010111",
  36262=>"011011010",
  36263=>"111101100",
  36264=>"001010001",
  36265=>"011000001",
  36266=>"111011011",
  36267=>"001110011",
  36268=>"010000111",
  36269=>"011000100",
  36270=>"001010001",
  36271=>"010000000",
  36272=>"100000001",
  36273=>"001010010",
  36274=>"011110010",
  36275=>"011101111",
  36276=>"000100011",
  36277=>"111000110",
  36278=>"110001011",
  36279=>"111110111",
  36280=>"011011011",
  36281=>"111101111",
  36282=>"010100101",
  36283=>"000001101",
  36284=>"111011000",
  36285=>"100010111",
  36286=>"101001110",
  36287=>"110010100",
  36288=>"110001010",
  36289=>"110111101",
  36290=>"110101101",
  36291=>"000111001",
  36292=>"110011010",
  36293=>"110100010",
  36294=>"011111111",
  36295=>"010000110",
  36296=>"100011011",
  36297=>"010110000",
  36298=>"101110000",
  36299=>"111101101",
  36300=>"010001011",
  36301=>"110111110",
  36302=>"000000000",
  36303=>"001000000",
  36304=>"010110001",
  36305=>"011011001",
  36306=>"001111010",
  36307=>"101001000",
  36308=>"100010110",
  36309=>"100011011",
  36310=>"101011101",
  36311=>"001010100",
  36312=>"111110010",
  36313=>"000110100",
  36314=>"010001000",
  36315=>"011010010",
  36316=>"110110111",
  36317=>"010011001",
  36318=>"100000111",
  36319=>"011011010",
  36320=>"001010000",
  36321=>"000001001",
  36322=>"001001010",
  36323=>"011100101",
  36324=>"011100001",
  36325=>"101110101",
  36326=>"101011111",
  36327=>"110100110",
  36328=>"101110010",
  36329=>"000101100",
  36330=>"110110001",
  36331=>"000110000",
  36332=>"000011111",
  36333=>"110011001",
  36334=>"100010111",
  36335=>"100011111",
  36336=>"011000010",
  36337=>"011100011",
  36338=>"000001011",
  36339=>"100100000",
  36340=>"110010111",
  36341=>"111111011",
  36342=>"000100011",
  36343=>"111010011",
  36344=>"100101101",
  36345=>"101001100",
  36346=>"001101000",
  36347=>"110001101",
  36348=>"111111111",
  36349=>"101100100",
  36350=>"111010011",
  36351=>"101111111",
  36352=>"000101110",
  36353=>"110000101",
  36354=>"010101101",
  36355=>"011001011",
  36356=>"111111111",
  36357=>"110011110",
  36358=>"000100100",
  36359=>"000001001",
  36360=>"000000101",
  36361=>"101101000",
  36362=>"000010101",
  36363=>"001100010",
  36364=>"110010111",
  36365=>"100111001",
  36366=>"101111010",
  36367=>"011101100",
  36368=>"000011011",
  36369=>"111000011",
  36370=>"000010010",
  36371=>"011011111",
  36372=>"100000111",
  36373=>"110101011",
  36374=>"100100110",
  36375=>"001111011",
  36376=>"111010000",
  36377=>"110101101",
  36378=>"010110110",
  36379=>"000011011",
  36380=>"100001010",
  36381=>"000011010",
  36382=>"101110011",
  36383=>"101111111",
  36384=>"001010011",
  36385=>"001111110",
  36386=>"011011001",
  36387=>"111101110",
  36388=>"110010000",
  36389=>"110010011",
  36390=>"010110011",
  36391=>"000011100",
  36392=>"101001000",
  36393=>"010010011",
  36394=>"100101011",
  36395=>"111011111",
  36396=>"110111110",
  36397=>"101110011",
  36398=>"010011010",
  36399=>"010101011",
  36400=>"111010001",
  36401=>"011111000",
  36402=>"000001110",
  36403=>"010001110",
  36404=>"011100110",
  36405=>"111101100",
  36406=>"101100101",
  36407=>"100000000",
  36408=>"000000010",
  36409=>"111101100",
  36410=>"101010101",
  36411=>"111111110",
  36412=>"000101000",
  36413=>"001011001",
  36414=>"011110100",
  36415=>"101110001",
  36416=>"100010110",
  36417=>"011000011",
  36418=>"000110011",
  36419=>"111010101",
  36420=>"111101101",
  36421=>"101111111",
  36422=>"011100111",
  36423=>"101101000",
  36424=>"111101011",
  36425=>"010110001",
  36426=>"100111101",
  36427=>"011111011",
  36428=>"111000100",
  36429=>"000001111",
  36430=>"010000101",
  36431=>"010010100",
  36432=>"010000000",
  36433=>"010001001",
  36434=>"111100111",
  36435=>"000110010",
  36436=>"001000000",
  36437=>"010000101",
  36438=>"001100000",
  36439=>"001011000",
  36440=>"110010110",
  36441=>"101100011",
  36442=>"101100011",
  36443=>"011000000",
  36444=>"011111111",
  36445=>"101011100",
  36446=>"011111110",
  36447=>"101010110",
  36448=>"001111111",
  36449=>"000111011",
  36450=>"011001101",
  36451=>"010110100",
  36452=>"111001000",
  36453=>"011000101",
  36454=>"101111100",
  36455=>"011110011",
  36456=>"111001011",
  36457=>"000011101",
  36458=>"100101110",
  36459=>"001100101",
  36460=>"110101100",
  36461=>"011101110",
  36462=>"110110011",
  36463=>"010101011",
  36464=>"000100011",
  36465=>"100101011",
  36466=>"111011100",
  36467=>"011011100",
  36468=>"001001001",
  36469=>"101111001",
  36470=>"110101100",
  36471=>"011010111",
  36472=>"100111101",
  36473=>"001001101",
  36474=>"001111100",
  36475=>"001110010",
  36476=>"110111000",
  36477=>"111001011",
  36478=>"001000000",
  36479=>"110111001",
  36480=>"011011101",
  36481=>"111010101",
  36482=>"001010011",
  36483=>"010011010",
  36484=>"101000011",
  36485=>"001000000",
  36486=>"111101111",
  36487=>"000111001",
  36488=>"000011011",
  36489=>"001001010",
  36490=>"010100011",
  36491=>"100111110",
  36492=>"001111101",
  36493=>"111100000",
  36494=>"000010000",
  36495=>"010010111",
  36496=>"100110110",
  36497=>"100001010",
  36498=>"100101100",
  36499=>"000000100",
  36500=>"110110111",
  36501=>"010010010",
  36502=>"000111100",
  36503=>"110001111",
  36504=>"110011000",
  36505=>"010111001",
  36506=>"111110000",
  36507=>"100000000",
  36508=>"111111000",
  36509=>"111000001",
  36510=>"100001111",
  36511=>"010101101",
  36512=>"001010110",
  36513=>"101100100",
  36514=>"010000010",
  36515=>"010011000",
  36516=>"101011011",
  36517=>"111100101",
  36518=>"110010101",
  36519=>"010010100",
  36520=>"000111110",
  36521=>"111111101",
  36522=>"010010101",
  36523=>"100101101",
  36524=>"111111110",
  36525=>"000100100",
  36526=>"101111111",
  36527=>"111011101",
  36528=>"110000110",
  36529=>"111011001",
  36530=>"111001000",
  36531=>"010010001",
  36532=>"110101011",
  36533=>"010001011",
  36534=>"110001101",
  36535=>"011110101",
  36536=>"110000111",
  36537=>"010000010",
  36538=>"011111110",
  36539=>"001101011",
  36540=>"100010110",
  36541=>"100001001",
  36542=>"000101100",
  36543=>"001010101",
  36544=>"111001011",
  36545=>"000110010",
  36546=>"001001111",
  36547=>"001101111",
  36548=>"111000010",
  36549=>"011011000",
  36550=>"101100001",
  36551=>"111101101",
  36552=>"010000110",
  36553=>"000000011",
  36554=>"101111011",
  36555=>"100100110",
  36556=>"000011101",
  36557=>"000000100",
  36558=>"111111001",
  36559=>"000100011",
  36560=>"101010011",
  36561=>"110101011",
  36562=>"001111100",
  36563=>"111100011",
  36564=>"010001010",
  36565=>"100010001",
  36566=>"000000000",
  36567=>"011101010",
  36568=>"000010000",
  36569=>"001010011",
  36570=>"000101111",
  36571=>"000101110",
  36572=>"110011010",
  36573=>"000010000",
  36574=>"101111101",
  36575=>"110110101",
  36576=>"000110010",
  36577=>"111011100",
  36578=>"011001100",
  36579=>"010101000",
  36580=>"100111001",
  36581=>"000110111",
  36582=>"111110010",
  36583=>"011011001",
  36584=>"010110111",
  36585=>"001011001",
  36586=>"110110000",
  36587=>"011100100",
  36588=>"110011010",
  36589=>"101011011",
  36590=>"111011111",
  36591=>"011001000",
  36592=>"101001000",
  36593=>"111011011",
  36594=>"100001010",
  36595=>"101101100",
  36596=>"000000000",
  36597=>"111110101",
  36598=>"000111011",
  36599=>"010010111",
  36600=>"110111010",
  36601=>"001111011",
  36602=>"111110101",
  36603=>"011101100",
  36604=>"100011111",
  36605=>"110100111",
  36606=>"010111000",
  36607=>"001001111",
  36608=>"011111110",
  36609=>"100111100",
  36610=>"111010000",
  36611=>"011111110",
  36612=>"001101101",
  36613=>"011111000",
  36614=>"011000010",
  36615=>"111011100",
  36616=>"110000111",
  36617=>"101001101",
  36618=>"010011011",
  36619=>"101001101",
  36620=>"101111111",
  36621=>"010111100",
  36622=>"000101111",
  36623=>"010011100",
  36624=>"110011111",
  36625=>"001010001",
  36626=>"010100001",
  36627=>"101111101",
  36628=>"011001000",
  36629=>"010110011",
  36630=>"010000010",
  36631=>"111000000",
  36632=>"101100101",
  36633=>"111110110",
  36634=>"110011000",
  36635=>"100100100",
  36636=>"111111001",
  36637=>"010010110",
  36638=>"000011111",
  36639=>"101101001",
  36640=>"000100010",
  36641=>"001010111",
  36642=>"011100111",
  36643=>"011011000",
  36644=>"101111101",
  36645=>"111100100",
  36646=>"010101100",
  36647=>"000101000",
  36648=>"111110011",
  36649=>"101111101",
  36650=>"111100010",
  36651=>"000000011",
  36652=>"100111100",
  36653=>"000101011",
  36654=>"101101110",
  36655=>"011100101",
  36656=>"111111111",
  36657=>"001011111",
  36658=>"100010000",
  36659=>"010011010",
  36660=>"010001010",
  36661=>"001000000",
  36662=>"100100111",
  36663=>"101001101",
  36664=>"000000001",
  36665=>"010101010",
  36666=>"100100111",
  36667=>"000000001",
  36668=>"101100001",
  36669=>"000110110",
  36670=>"101111111",
  36671=>"000111010",
  36672=>"110110000",
  36673=>"011000111",
  36674=>"100100110",
  36675=>"000000100",
  36676=>"101000011",
  36677=>"011100011",
  36678=>"101111110",
  36679=>"100001101",
  36680=>"001110111",
  36681=>"101111000",
  36682=>"000000100",
  36683=>"001000101",
  36684=>"010110000",
  36685=>"011011101",
  36686=>"111000100",
  36687=>"101100100",
  36688=>"000100010",
  36689=>"101110100",
  36690=>"101001010",
  36691=>"001111000",
  36692=>"000100100",
  36693=>"010111101",
  36694=>"100111000",
  36695=>"010111111",
  36696=>"011111111",
  36697=>"101011000",
  36698=>"011101110",
  36699=>"010010000",
  36700=>"101001111",
  36701=>"101001011",
  36702=>"111101101",
  36703=>"010110001",
  36704=>"111011110",
  36705=>"010110111",
  36706=>"000011000",
  36707=>"011001000",
  36708=>"100000001",
  36709=>"010101100",
  36710=>"101010000",
  36711=>"101000001",
  36712=>"111001001",
  36713=>"111000110",
  36714=>"000100100",
  36715=>"111101101",
  36716=>"100001001",
  36717=>"001001000",
  36718=>"100000100",
  36719=>"011000100",
  36720=>"011011111",
  36721=>"101010111",
  36722=>"011010001",
  36723=>"001010001",
  36724=>"001001100",
  36725=>"110111100",
  36726=>"010111001",
  36727=>"101000110",
  36728=>"000000011",
  36729=>"110011100",
  36730=>"010001001",
  36731=>"011010101",
  36732=>"000000001",
  36733=>"001111011",
  36734=>"101101010",
  36735=>"101110001",
  36736=>"011101110",
  36737=>"110011111",
  36738=>"000101110",
  36739=>"111100011",
  36740=>"011001100",
  36741=>"001011001",
  36742=>"011010101",
  36743=>"000010101",
  36744=>"011001000",
  36745=>"011111101",
  36746=>"100000100",
  36747=>"011001001",
  36748=>"010011001",
  36749=>"011011000",
  36750=>"000000111",
  36751=>"111110100",
  36752=>"011010100",
  36753=>"001010010",
  36754=>"111100100",
  36755=>"011001100",
  36756=>"010000110",
  36757=>"101000100",
  36758=>"000101111",
  36759=>"011101100",
  36760=>"000000001",
  36761=>"010101101",
  36762=>"111001011",
  36763=>"000010000",
  36764=>"110010011",
  36765=>"111101010",
  36766=>"111110100",
  36767=>"100010101",
  36768=>"111010000",
  36769=>"111111101",
  36770=>"110110010",
  36771=>"000001111",
  36772=>"011011010",
  36773=>"100000101",
  36774=>"111101010",
  36775=>"010111001",
  36776=>"101100000",
  36777=>"001011101",
  36778=>"111110100",
  36779=>"111111111",
  36780=>"000110100",
  36781=>"001011111",
  36782=>"000100001",
  36783=>"100101110",
  36784=>"011011010",
  36785=>"101010111",
  36786=>"110011001",
  36787=>"101010110",
  36788=>"111010010",
  36789=>"111100101",
  36790=>"110001010",
  36791=>"011101011",
  36792=>"111101110",
  36793=>"100111100",
  36794=>"101111100",
  36795=>"011100000",
  36796=>"111000111",
  36797=>"011100101",
  36798=>"011000101",
  36799=>"001100001",
  36800=>"010000011",
  36801=>"011100101",
  36802=>"001110110",
  36803=>"001110000",
  36804=>"111110000",
  36805=>"001111100",
  36806=>"100001000",
  36807=>"101101110",
  36808=>"101000101",
  36809=>"010110001",
  36810=>"100000000",
  36811=>"100011101",
  36812=>"011001001",
  36813=>"101010100",
  36814=>"101001001",
  36815=>"001100101",
  36816=>"111101011",
  36817=>"011100010",
  36818=>"001101000",
  36819=>"111000110",
  36820=>"101001101",
  36821=>"000000001",
  36822=>"001001100",
  36823=>"010101000",
  36824=>"000000000",
  36825=>"001100111",
  36826=>"110011010",
  36827=>"010010111",
  36828=>"101100101",
  36829=>"101110000",
  36830=>"111011011",
  36831=>"010010001",
  36832=>"011010100",
  36833=>"000001010",
  36834=>"100010101",
  36835=>"100011010",
  36836=>"011010101",
  36837=>"100001100",
  36838=>"101100111",
  36839=>"101110110",
  36840=>"000000100",
  36841=>"101000010",
  36842=>"011100101",
  36843=>"111101000",
  36844=>"001111100",
  36845=>"101001001",
  36846=>"001011011",
  36847=>"011001111",
  36848=>"111101111",
  36849=>"010110111",
  36850=>"001100110",
  36851=>"111001110",
  36852=>"101010000",
  36853=>"101000100",
  36854=>"110111111",
  36855=>"010110001",
  36856=>"110101110",
  36857=>"110010001",
  36858=>"101010001",
  36859=>"011110011",
  36860=>"101101101",
  36861=>"111100011",
  36862=>"010011011",
  36863=>"110001101",
  36864=>"111100111",
  36865=>"010100000",
  36866=>"111101111",
  36867=>"111101000",
  36868=>"111011110",
  36869=>"101111100",
  36870=>"001010010",
  36871=>"010000000",
  36872=>"011010011",
  36873=>"100100100",
  36874=>"011010101",
  36875=>"101001101",
  36876=>"100100001",
  36877=>"110010000",
  36878=>"110011010",
  36879=>"010110111",
  36880=>"011000110",
  36881=>"100000111",
  36882=>"001101000",
  36883=>"010001100",
  36884=>"000000100",
  36885=>"111101010",
  36886=>"110000010",
  36887=>"001001010",
  36888=>"100110000",
  36889=>"010111000",
  36890=>"000110101",
  36891=>"011101101",
  36892=>"010010000",
  36893=>"000111100",
  36894=>"011000111",
  36895=>"111010100",
  36896=>"010001110",
  36897=>"011101001",
  36898=>"101110101",
  36899=>"000011101",
  36900=>"011101111",
  36901=>"110100100",
  36902=>"000111110",
  36903=>"101110010",
  36904=>"000000010",
  36905=>"010010111",
  36906=>"111000110",
  36907=>"001000000",
  36908=>"000110001",
  36909=>"001010010",
  36910=>"110110111",
  36911=>"101111111",
  36912=>"111100001",
  36913=>"111100111",
  36914=>"010011100",
  36915=>"010111110",
  36916=>"001000000",
  36917=>"011010100",
  36918=>"010000010",
  36919=>"001111101",
  36920=>"100011010",
  36921=>"111100010",
  36922=>"000011010",
  36923=>"101100110",
  36924=>"010111001",
  36925=>"001101111",
  36926=>"000111111",
  36927=>"100110101",
  36928=>"000000101",
  36929=>"101101001",
  36930=>"100101100",
  36931=>"010001000",
  36932=>"111100001",
  36933=>"001000000",
  36934=>"011010111",
  36935=>"010001010",
  36936=>"101001111",
  36937=>"000101000",
  36938=>"111101011",
  36939=>"111001110",
  36940=>"001100001",
  36941=>"100001100",
  36942=>"101000101",
  36943=>"110111110",
  36944=>"001101100",
  36945=>"000111000",
  36946=>"010010001",
  36947=>"011100010",
  36948=>"010011000",
  36949=>"001001101",
  36950=>"111101101",
  36951=>"011011110",
  36952=>"101011001",
  36953=>"000000101",
  36954=>"101001110",
  36955=>"000101010",
  36956=>"011100000",
  36957=>"001010001",
  36958=>"100011001",
  36959=>"101000001",
  36960=>"010001010",
  36961=>"011101110",
  36962=>"111010111",
  36963=>"011001001",
  36964=>"100011100",
  36965=>"101010100",
  36966=>"100001000",
  36967=>"111110001",
  36968=>"000111001",
  36969=>"111011010",
  36970=>"001001001",
  36971=>"001010100",
  36972=>"000000101",
  36973=>"111011100",
  36974=>"100011010",
  36975=>"111010011",
  36976=>"111001100",
  36977=>"101101000",
  36978=>"100011001",
  36979=>"010011010",
  36980=>"011010100",
  36981=>"111010000",
  36982=>"100000010",
  36983=>"100111110",
  36984=>"001001100",
  36985=>"010000111",
  36986=>"000011010",
  36987=>"010110100",
  36988=>"001001000",
  36989=>"111110110",
  36990=>"010001100",
  36991=>"001101001",
  36992=>"010110001",
  36993=>"110111101",
  36994=>"001001011",
  36995=>"000001110",
  36996=>"010001000",
  36997=>"101011010",
  36998=>"001011100",
  36999=>"111011110",
  37000=>"000000010",
  37001=>"011010000",
  37002=>"001000101",
  37003=>"110010100",
  37004=>"011000011",
  37005=>"010111001",
  37006=>"101010000",
  37007=>"011001101",
  37008=>"000010110",
  37009=>"001111110",
  37010=>"100010100",
  37011=>"100101001",
  37012=>"010010100",
  37013=>"010110111",
  37014=>"011001110",
  37015=>"111100010",
  37016=>"101111000",
  37017=>"110011101",
  37018=>"011111001",
  37019=>"000110011",
  37020=>"000111111",
  37021=>"000010001",
  37022=>"110000111",
  37023=>"100101110",
  37024=>"111110000",
  37025=>"001110000",
  37026=>"111010010",
  37027=>"110111101",
  37028=>"111010011",
  37029=>"010101001",
  37030=>"000000101",
  37031=>"010001010",
  37032=>"011000001",
  37033=>"011010111",
  37034=>"110001000",
  37035=>"100010111",
  37036=>"000000010",
  37037=>"100010100",
  37038=>"111100011",
  37039=>"100001000",
  37040=>"001010011",
  37041=>"001000011",
  37042=>"000100010",
  37043=>"100001111",
  37044=>"010111101",
  37045=>"011111001",
  37046=>"111101110",
  37047=>"000010000",
  37048=>"001100011",
  37049=>"001010101",
  37050=>"000011010",
  37051=>"000101101",
  37052=>"111111111",
  37053=>"101001000",
  37054=>"000011111",
  37055=>"000010111",
  37056=>"101001000",
  37057=>"111011100",
  37058=>"000010010",
  37059=>"101100010",
  37060=>"010000111",
  37061=>"110010000",
  37062=>"110101101",
  37063=>"000110100",
  37064=>"001110000",
  37065=>"000000101",
  37066=>"001001100",
  37067=>"101101101",
  37068=>"111010100",
  37069=>"110001000",
  37070=>"110011001",
  37071=>"101001101",
  37072=>"111001111",
  37073=>"011011111",
  37074=>"001011010",
  37075=>"010101110",
  37076=>"001111110",
  37077=>"110011010",
  37078=>"000001110",
  37079=>"011110111",
  37080=>"011100011",
  37081=>"110001111",
  37082=>"101011010",
  37083=>"000001101",
  37084=>"011111001",
  37085=>"000010100",
  37086=>"011100111",
  37087=>"100001000",
  37088=>"111011111",
  37089=>"011110000",
  37090=>"101000000",
  37091=>"001000011",
  37092=>"011110110",
  37093=>"001100000",
  37094=>"011100011",
  37095=>"100001011",
  37096=>"000001001",
  37097=>"010110110",
  37098=>"101111101",
  37099=>"001110011",
  37100=>"110101110",
  37101=>"100111100",
  37102=>"011001110",
  37103=>"010110000",
  37104=>"110000100",
  37105=>"011111111",
  37106=>"110010010",
  37107=>"111000010",
  37108=>"001101001",
  37109=>"000000101",
  37110=>"111011111",
  37111=>"110001101",
  37112=>"010001111",
  37113=>"101100101",
  37114=>"001001110",
  37115=>"010000100",
  37116=>"000011111",
  37117=>"101101000",
  37118=>"001000110",
  37119=>"111001101",
  37120=>"000011111",
  37121=>"100100111",
  37122=>"011011101",
  37123=>"110100010",
  37124=>"100101000",
  37125=>"001111111",
  37126=>"111111101",
  37127=>"001101110",
  37128=>"010001010",
  37129=>"010011101",
  37130=>"001100010",
  37131=>"010110000",
  37132=>"010110101",
  37133=>"110001001",
  37134=>"001110100",
  37135=>"011010000",
  37136=>"000011010",
  37137=>"100101101",
  37138=>"110010010",
  37139=>"101101111",
  37140=>"111011000",
  37141=>"010010101",
  37142=>"011100001",
  37143=>"010110011",
  37144=>"100000001",
  37145=>"100001010",
  37146=>"100010000",
  37147=>"101000101",
  37148=>"110010101",
  37149=>"111100100",
  37150=>"011010000",
  37151=>"011100010",
  37152=>"111000000",
  37153=>"000100010",
  37154=>"011000001",
  37155=>"101110001",
  37156=>"111111100",
  37157=>"001010100",
  37158=>"110101000",
  37159=>"101011011",
  37160=>"001000110",
  37161=>"010110111",
  37162=>"110101011",
  37163=>"000111110",
  37164=>"101111000",
  37165=>"011111111",
  37166=>"011000111",
  37167=>"000001001",
  37168=>"100010000",
  37169=>"100110000",
  37170=>"011111000",
  37171=>"100101010",
  37172=>"111001111",
  37173=>"000110100",
  37174=>"111111000",
  37175=>"001000011",
  37176=>"001110101",
  37177=>"100010111",
  37178=>"100101110",
  37179=>"011110111",
  37180=>"100100011",
  37181=>"001001010",
  37182=>"001111000",
  37183=>"100001101",
  37184=>"110111101",
  37185=>"011100001",
  37186=>"110001011",
  37187=>"111100010",
  37188=>"101110000",
  37189=>"111000011",
  37190=>"101101111",
  37191=>"010011001",
  37192=>"010101110",
  37193=>"000000000",
  37194=>"111011100",
  37195=>"111101100",
  37196=>"011110100",
  37197=>"000010000",
  37198=>"111010101",
  37199=>"011000000",
  37200=>"001101010",
  37201=>"111101000",
  37202=>"100001110",
  37203=>"101000100",
  37204=>"000101110",
  37205=>"101111010",
  37206=>"000011010",
  37207=>"011000010",
  37208=>"001000101",
  37209=>"111010101",
  37210=>"001100010",
  37211=>"000001010",
  37212=>"010010101",
  37213=>"111001101",
  37214=>"111111000",
  37215=>"110100001",
  37216=>"001011010",
  37217=>"110101011",
  37218=>"111110000",
  37219=>"010001010",
  37220=>"110011100",
  37221=>"111000010",
  37222=>"101100101",
  37223=>"101100010",
  37224=>"011000111",
  37225=>"000010111",
  37226=>"001000101",
  37227=>"010011110",
  37228=>"011100011",
  37229=>"110100111",
  37230=>"100010001",
  37231=>"001011000",
  37232=>"011011011",
  37233=>"101010101",
  37234=>"010011101",
  37235=>"110111101",
  37236=>"101010011",
  37237=>"000001001",
  37238=>"111101011",
  37239=>"100101001",
  37240=>"010011001",
  37241=>"010101101",
  37242=>"001101111",
  37243=>"000110000",
  37244=>"110010111",
  37245=>"110101110",
  37246=>"011000011",
  37247=>"111000010",
  37248=>"110111111",
  37249=>"111101011",
  37250=>"101100001",
  37251=>"101111110",
  37252=>"110100001",
  37253=>"010001111",
  37254=>"000010101",
  37255=>"111110011",
  37256=>"011000111",
  37257=>"001111010",
  37258=>"011011111",
  37259=>"110011000",
  37260=>"100010011",
  37261=>"110110010",
  37262=>"001100000",
  37263=>"110101111",
  37264=>"111011101",
  37265=>"110001101",
  37266=>"010111100",
  37267=>"111011010",
  37268=>"100011110",
  37269=>"111010001",
  37270=>"000010001",
  37271=>"000011111",
  37272=>"101010100",
  37273=>"011001001",
  37274=>"111010111",
  37275=>"011101000",
  37276=>"101010110",
  37277=>"101010010",
  37278=>"101001000",
  37279=>"101001000",
  37280=>"000000011",
  37281=>"110000111",
  37282=>"111011100",
  37283=>"101100011",
  37284=>"001001001",
  37285=>"000010111",
  37286=>"000100111",
  37287=>"001111010",
  37288=>"110101000",
  37289=>"010101001",
  37290=>"011111010",
  37291=>"001001111",
  37292=>"010000001",
  37293=>"001101001",
  37294=>"000110001",
  37295=>"110100001",
  37296=>"011111000",
  37297=>"011101000",
  37298=>"100000101",
  37299=>"000000000",
  37300=>"011111010",
  37301=>"110001010",
  37302=>"001000001",
  37303=>"000111001",
  37304=>"100101000",
  37305=>"111000001",
  37306=>"011110011",
  37307=>"110011111",
  37308=>"110101110",
  37309=>"010111111",
  37310=>"010110100",
  37311=>"011010111",
  37312=>"000001101",
  37313=>"111111001",
  37314=>"001111010",
  37315=>"001011010",
  37316=>"011001110",
  37317=>"111001110",
  37318=>"110101111",
  37319=>"011010001",
  37320=>"100011110",
  37321=>"001001011",
  37322=>"111000111",
  37323=>"010100111",
  37324=>"101110110",
  37325=>"010001110",
  37326=>"111110101",
  37327=>"101001010",
  37328=>"011001000",
  37329=>"001110000",
  37330=>"101101011",
  37331=>"011110100",
  37332=>"001000111",
  37333=>"010000100",
  37334=>"110001011",
  37335=>"000111101",
  37336=>"110100110",
  37337=>"100010000",
  37338=>"000000000",
  37339=>"100100011",
  37340=>"001010111",
  37341=>"000000111",
  37342=>"010000100",
  37343=>"000111101",
  37344=>"101101100",
  37345=>"110100111",
  37346=>"001111111",
  37347=>"000101111",
  37348=>"010010101",
  37349=>"100110000",
  37350=>"110101001",
  37351=>"001011100",
  37352=>"101001010",
  37353=>"111010100",
  37354=>"000001000",
  37355=>"111011100",
  37356=>"101100011",
  37357=>"011100001",
  37358=>"100100000",
  37359=>"000010110",
  37360=>"001111111",
  37361=>"010101101",
  37362=>"000010001",
  37363=>"001111100",
  37364=>"001000111",
  37365=>"011000100",
  37366=>"111101010",
  37367=>"111011100",
  37368=>"010100100",
  37369=>"010110000",
  37370=>"010111111",
  37371=>"111110010",
  37372=>"011101110",
  37373=>"100111100",
  37374=>"010001101",
  37375=>"001110110",
  37376=>"000000011",
  37377=>"110000010",
  37378=>"011110110",
  37379=>"100011011",
  37380=>"111011010",
  37381=>"000101100",
  37382=>"100010000",
  37383=>"001111101",
  37384=>"001111110",
  37385=>"000110010",
  37386=>"000101100",
  37387=>"010011101",
  37388=>"000000000",
  37389=>"011010110",
  37390=>"000110110",
  37391=>"111111100",
  37392=>"001010010",
  37393=>"001111100",
  37394=>"101010010",
  37395=>"100011110",
  37396=>"000001000",
  37397=>"010010000",
  37398=>"111100101",
  37399=>"011101110",
  37400=>"010011011",
  37401=>"001110110",
  37402=>"010010100",
  37403=>"011010001",
  37404=>"011110111",
  37405=>"010001011",
  37406=>"100111011",
  37407=>"101111110",
  37408=>"011101110",
  37409=>"101110110",
  37410=>"001110111",
  37411=>"000100011",
  37412=>"010011000",
  37413=>"010100101",
  37414=>"110111110",
  37415=>"001101010",
  37416=>"101010011",
  37417=>"101001111",
  37418=>"100100101",
  37419=>"010101000",
  37420=>"111000010",
  37421=>"111001010",
  37422=>"000000111",
  37423=>"010101111",
  37424=>"111110101",
  37425=>"011100010",
  37426=>"000000000",
  37427=>"010000101",
  37428=>"000111000",
  37429=>"000001100",
  37430=>"011011110",
  37431=>"011110100",
  37432=>"011101011",
  37433=>"010111101",
  37434=>"011100110",
  37435=>"100000110",
  37436=>"111101001",
  37437=>"011011110",
  37438=>"010101111",
  37439=>"110100100",
  37440=>"011000110",
  37441=>"000000111",
  37442=>"011010111",
  37443=>"100010011",
  37444=>"010001100",
  37445=>"010011110",
  37446=>"101100000",
  37447=>"001010001",
  37448=>"111111010",
  37449=>"011101100",
  37450=>"011010111",
  37451=>"110001111",
  37452=>"001110011",
  37453=>"000001010",
  37454=>"011101100",
  37455=>"101110000",
  37456=>"111110100",
  37457=>"001000001",
  37458=>"001101110",
  37459=>"001111000",
  37460=>"110110111",
  37461=>"001110010",
  37462=>"111011000",
  37463=>"110010111",
  37464=>"011011101",
  37465=>"000010110",
  37466=>"010010100",
  37467=>"010101101",
  37468=>"101001000",
  37469=>"000011011",
  37470=>"111101001",
  37471=>"011101000",
  37472=>"100011000",
  37473=>"101110010",
  37474=>"010100111",
  37475=>"110111010",
  37476=>"111011101",
  37477=>"011010100",
  37478=>"000010011",
  37479=>"111000101",
  37480=>"100001111",
  37481=>"110111100",
  37482=>"111111111",
  37483=>"011110111",
  37484=>"100111101",
  37485=>"001000011",
  37486=>"011110111",
  37487=>"110101111",
  37488=>"101011110",
  37489=>"101111110",
  37490=>"010111001",
  37491=>"010101100",
  37492=>"101111000",
  37493=>"100101000",
  37494=>"110110000",
  37495=>"101100000",
  37496=>"100110111",
  37497=>"001101001",
  37498=>"000100011",
  37499=>"111010011",
  37500=>"101010001",
  37501=>"101011010",
  37502=>"001100000",
  37503=>"101111010",
  37504=>"011111011",
  37505=>"000000000",
  37506=>"111101011",
  37507=>"011101010",
  37508=>"010100101",
  37509=>"010111110",
  37510=>"100110000",
  37511=>"100000111",
  37512=>"000110100",
  37513=>"000010011",
  37514=>"011010000",
  37515=>"110110111",
  37516=>"011000000",
  37517=>"111011000",
  37518=>"111101011",
  37519=>"000101110",
  37520=>"001000110",
  37521=>"001101100",
  37522=>"111110011",
  37523=>"011010010",
  37524=>"110100001",
  37525=>"010001011",
  37526=>"000100011",
  37527=>"101110100",
  37528=>"001100010",
  37529=>"110000111",
  37530=>"001010110",
  37531=>"111010110",
  37532=>"000111011",
  37533=>"111010110",
  37534=>"010001011",
  37535=>"111110011",
  37536=>"011001111",
  37537=>"011111101",
  37538=>"000011101",
  37539=>"000011110",
  37540=>"101010101",
  37541=>"011000111",
  37542=>"110011010",
  37543=>"111100111",
  37544=>"110101100",
  37545=>"001111000",
  37546=>"110001100",
  37547=>"010011010",
  37548=>"000001001",
  37549=>"110000001",
  37550=>"011100101",
  37551=>"101111110",
  37552=>"000011011",
  37553=>"100100110",
  37554=>"110111011",
  37555=>"001001111",
  37556=>"101001000",
  37557=>"111100100",
  37558=>"111111000",
  37559=>"101111001",
  37560=>"011001000",
  37561=>"111100010",
  37562=>"110111100",
  37563=>"110010100",
  37564=>"100110010",
  37565=>"110011110",
  37566=>"000010111",
  37567=>"110010010",
  37568=>"010011000",
  37569=>"110000110",
  37570=>"000000001",
  37571=>"000001001",
  37572=>"100000110",
  37573=>"001000111",
  37574=>"111000011",
  37575=>"011010000",
  37576=>"110111100",
  37577=>"011001011",
  37578=>"000010111",
  37579=>"100010010",
  37580=>"100000111",
  37581=>"101111010",
  37582=>"000000110",
  37583=>"111111110",
  37584=>"011101000",
  37585=>"001011101",
  37586=>"010000111",
  37587=>"111100010",
  37588=>"000101111",
  37589=>"001000111",
  37590=>"111100100",
  37591=>"000110001",
  37592=>"101000011",
  37593=>"011011100",
  37594=>"001111100",
  37595=>"000000110",
  37596=>"110000001",
  37597=>"100011110",
  37598=>"010001101",
  37599=>"010010101",
  37600=>"000100011",
  37601=>"101110111",
  37602=>"011111000",
  37603=>"001100101",
  37604=>"000110011",
  37605=>"101010001",
  37606=>"110011111",
  37607=>"000011000",
  37608=>"010001010",
  37609=>"011010010",
  37610=>"011011001",
  37611=>"101001000",
  37612=>"011010011",
  37613=>"101111010",
  37614=>"010111111",
  37615=>"100001000",
  37616=>"110111100",
  37617=>"011101000",
  37618=>"000111001",
  37619=>"110010101",
  37620=>"000000010",
  37621=>"000000000",
  37622=>"100000111",
  37623=>"000110001",
  37624=>"011011101",
  37625=>"011100110",
  37626=>"110110110",
  37627=>"001000110",
  37628=>"000011011",
  37629=>"011110100",
  37630=>"000010011",
  37631=>"000001100",
  37632=>"010100010",
  37633=>"111111111",
  37634=>"011100110",
  37635=>"011100010",
  37636=>"110011101",
  37637=>"110111010",
  37638=>"001101011",
  37639=>"100110000",
  37640=>"100100111",
  37641=>"111101110",
  37642=>"000110011",
  37643=>"110110100",
  37644=>"111100001",
  37645=>"001001100",
  37646=>"110100111",
  37647=>"011001001",
  37648=>"011000110",
  37649=>"101000100",
  37650=>"010101110",
  37651=>"110000001",
  37652=>"001110100",
  37653=>"101000101",
  37654=>"000010100",
  37655=>"000011101",
  37656=>"011010011",
  37657=>"100010010",
  37658=>"000111000",
  37659=>"011101110",
  37660=>"111110111",
  37661=>"001110110",
  37662=>"000100010",
  37663=>"101101110",
  37664=>"110111100",
  37665=>"100010100",
  37666=>"101010100",
  37667=>"110111000",
  37668=>"111110110",
  37669=>"100001000",
  37670=>"001011010",
  37671=>"011101100",
  37672=>"010010101",
  37673=>"101000001",
  37674=>"110010100",
  37675=>"010100111",
  37676=>"000001101",
  37677=>"100101001",
  37678=>"000110001",
  37679=>"100001101",
  37680=>"001100011",
  37681=>"000010000",
  37682=>"010100011",
  37683=>"100010011",
  37684=>"111101100",
  37685=>"001010110",
  37686=>"011000010",
  37687=>"101101110",
  37688=>"110011100",
  37689=>"011101000",
  37690=>"001100100",
  37691=>"011110010",
  37692=>"111010000",
  37693=>"000111100",
  37694=>"101111110",
  37695=>"001000100",
  37696=>"100101010",
  37697=>"101000101",
  37698=>"000101111",
  37699=>"100001011",
  37700=>"111010001",
  37701=>"001011000",
  37702=>"101100100",
  37703=>"000000111",
  37704=>"010100101",
  37705=>"110010000",
  37706=>"000100100",
  37707=>"100101000",
  37708=>"000010011",
  37709=>"011101110",
  37710=>"111010010",
  37711=>"011011110",
  37712=>"100010010",
  37713=>"000101001",
  37714=>"001010100",
  37715=>"100000110",
  37716=>"111000010",
  37717=>"100011011",
  37718=>"101000000",
  37719=>"101111110",
  37720=>"101001001",
  37721=>"000101100",
  37722=>"111001101",
  37723=>"101111110",
  37724=>"111111110",
  37725=>"011110111",
  37726=>"010001001",
  37727=>"001000100",
  37728=>"110101111",
  37729=>"111110001",
  37730=>"101000000",
  37731=>"110000001",
  37732=>"000001111",
  37733=>"101010110",
  37734=>"100110001",
  37735=>"011110010",
  37736=>"100100100",
  37737=>"111000101",
  37738=>"011111110",
  37739=>"110011011",
  37740=>"101111110",
  37741=>"010111111",
  37742=>"011011001",
  37743=>"010010010",
  37744=>"101100110",
  37745=>"111011100",
  37746=>"001011010",
  37747=>"101110110",
  37748=>"100001111",
  37749=>"111111010",
  37750=>"101011000",
  37751=>"000001101",
  37752=>"100010001",
  37753=>"100100101",
  37754=>"111010001",
  37755=>"110000011",
  37756=>"001000100",
  37757=>"001111100",
  37758=>"011111100",
  37759=>"011100111",
  37760=>"101000101",
  37761=>"110100001",
  37762=>"010001000",
  37763=>"111000110",
  37764=>"010100011",
  37765=>"001001011",
  37766=>"111101000",
  37767=>"000101001",
  37768=>"011011100",
  37769=>"001011000",
  37770=>"110001010",
  37771=>"111101111",
  37772=>"000110001",
  37773=>"000001101",
  37774=>"101001000",
  37775=>"001110000",
  37776=>"110011001",
  37777=>"001110001",
  37778=>"001110011",
  37779=>"000011111",
  37780=>"101001001",
  37781=>"101000010",
  37782=>"011001000",
  37783=>"000111100",
  37784=>"101001000",
  37785=>"110100110",
  37786=>"001111001",
  37787=>"100010101",
  37788=>"110011010",
  37789=>"001000000",
  37790=>"000000010",
  37791=>"110000110",
  37792=>"001011000",
  37793=>"111100111",
  37794=>"110100011",
  37795=>"100011101",
  37796=>"110010100",
  37797=>"011000001",
  37798=>"100101100",
  37799=>"000010110",
  37800=>"110001101",
  37801=>"111000011",
  37802=>"111101011",
  37803=>"110100101",
  37804=>"000011010",
  37805=>"001110110",
  37806=>"000100000",
  37807=>"100010010",
  37808=>"010000000",
  37809=>"110100001",
  37810=>"010100111",
  37811=>"000000010",
  37812=>"111100000",
  37813=>"000111100",
  37814=>"001111000",
  37815=>"000101000",
  37816=>"000100000",
  37817=>"001000111",
  37818=>"101000000",
  37819=>"000000010",
  37820=>"101101101",
  37821=>"001011100",
  37822=>"111110110",
  37823=>"100010110",
  37824=>"000011000",
  37825=>"001101110",
  37826=>"011001011",
  37827=>"111100010",
  37828=>"111010101",
  37829=>"111101100",
  37830=>"111101111",
  37831=>"110101001",
  37832=>"100001001",
  37833=>"110011001",
  37834=>"010000000",
  37835=>"010100110",
  37836=>"001100110",
  37837=>"111010101",
  37838=>"110011100",
  37839=>"100000101",
  37840=>"000110101",
  37841=>"001001111",
  37842=>"010011101",
  37843=>"110101101",
  37844=>"000000000",
  37845=>"111111100",
  37846=>"011000010",
  37847=>"001010000",
  37848=>"101000110",
  37849=>"111000111",
  37850=>"010100110",
  37851=>"101010110",
  37852=>"110111011",
  37853=>"010100110",
  37854=>"100000100",
  37855=>"111111111",
  37856=>"111100001",
  37857=>"010110100",
  37858=>"010011000",
  37859=>"000100011",
  37860=>"000000100",
  37861=>"000111110",
  37862=>"011110100",
  37863=>"010000111",
  37864=>"000011100",
  37865=>"101111100",
  37866=>"101101011",
  37867=>"010011001",
  37868=>"111100101",
  37869=>"010110111",
  37870=>"011110000",
  37871=>"000100101",
  37872=>"111101110",
  37873=>"100100000",
  37874=>"100101001",
  37875=>"100001001",
  37876=>"111111000",
  37877=>"111101010",
  37878=>"100010100",
  37879=>"101100001",
  37880=>"000001001",
  37881=>"001001001",
  37882=>"011110001",
  37883=>"011110100",
  37884=>"000010000",
  37885=>"101000100",
  37886=>"100011101",
  37887=>"101011001",
  37888=>"101100111",
  37889=>"001100110",
  37890=>"111110110",
  37891=>"011111100",
  37892=>"100111101",
  37893=>"111010001",
  37894=>"010010110",
  37895=>"110100101",
  37896=>"011001111",
  37897=>"011011100",
  37898=>"000010110",
  37899=>"000011010",
  37900=>"100011011",
  37901=>"110010100",
  37902=>"001010111",
  37903=>"111111101",
  37904=>"000001011",
  37905=>"101110001",
  37906=>"010010111",
  37907=>"110001110",
  37908=>"010000000",
  37909=>"000111011",
  37910=>"011101101",
  37911=>"110101100",
  37912=>"111011100",
  37913=>"001011011",
  37914=>"001000111",
  37915=>"011000000",
  37916=>"100101000",
  37917=>"111001001",
  37918=>"011100111",
  37919=>"011010001",
  37920=>"100100001",
  37921=>"011001111",
  37922=>"001111110",
  37923=>"001011101",
  37924=>"110101000",
  37925=>"101110110",
  37926=>"000110100",
  37927=>"111010100",
  37928=>"111101000",
  37929=>"100011010",
  37930=>"110110001",
  37931=>"100010001",
  37932=>"000100100",
  37933=>"001100110",
  37934=>"011011010",
  37935=>"111100110",
  37936=>"011101010",
  37937=>"111111000",
  37938=>"000010000",
  37939=>"100111001",
  37940=>"011001011",
  37941=>"111001111",
  37942=>"111000001",
  37943=>"010101000",
  37944=>"111111011",
  37945=>"011010011",
  37946=>"000001101",
  37947=>"000111010",
  37948=>"000001111",
  37949=>"000111110",
  37950=>"100111111",
  37951=>"001001101",
  37952=>"101000000",
  37953=>"000010000",
  37954=>"010010110",
  37955=>"111101010",
  37956=>"101101111",
  37957=>"101010110",
  37958=>"101100011",
  37959=>"010000011",
  37960=>"010100011",
  37961=>"111010000",
  37962=>"101000001",
  37963=>"101000000",
  37964=>"101001110",
  37965=>"100110110",
  37966=>"001010111",
  37967=>"011110110",
  37968=>"110110101",
  37969=>"000000100",
  37970=>"011101100",
  37971=>"100011100",
  37972=>"101010101",
  37973=>"001101110",
  37974=>"110000010",
  37975=>"101100101",
  37976=>"101011011",
  37977=>"111111010",
  37978=>"101001001",
  37979=>"011100111",
  37980=>"011011000",
  37981=>"011001110",
  37982=>"010001010",
  37983=>"010101111",
  37984=>"000100011",
  37985=>"011001000",
  37986=>"000011010",
  37987=>"011000010",
  37988=>"101000000",
  37989=>"111101110",
  37990=>"100110110",
  37991=>"110001011",
  37992=>"100100100",
  37993=>"001101110",
  37994=>"111001110",
  37995=>"110000100",
  37996=>"111100010",
  37997=>"000101010",
  37998=>"010001010",
  37999=>"101000001",
  38000=>"000011100",
  38001=>"010110101",
  38002=>"100001100",
  38003=>"010111010",
  38004=>"000010100",
  38005=>"000111000",
  38006=>"010010011",
  38007=>"001100000",
  38008=>"100001001",
  38009=>"001000110",
  38010=>"111101111",
  38011=>"111101000",
  38012=>"000110001",
  38013=>"011111110",
  38014=>"001010000",
  38015=>"000010111",
  38016=>"101101011",
  38017=>"010010000",
  38018=>"000000011",
  38019=>"000000000",
  38020=>"010011001",
  38021=>"111100010",
  38022=>"011110000",
  38023=>"110010000",
  38024=>"000111101",
  38025=>"001000001",
  38026=>"110101000",
  38027=>"000001100",
  38028=>"101110011",
  38029=>"001010010",
  38030=>"010000110",
  38031=>"100000111",
  38032=>"101001110",
  38033=>"100011110",
  38034=>"111000000",
  38035=>"100111011",
  38036=>"100001000",
  38037=>"000011000",
  38038=>"011100011",
  38039=>"011111011",
  38040=>"110010000",
  38041=>"000001010",
  38042=>"011111011",
  38043=>"111110111",
  38044=>"111101000",
  38045=>"000001011",
  38046=>"101100111",
  38047=>"000000000",
  38048=>"101010001",
  38049=>"010111111",
  38050=>"001110001",
  38051=>"101000100",
  38052=>"000111011",
  38053=>"000111001",
  38054=>"001111110",
  38055=>"011011000",
  38056=>"011100111",
  38057=>"001000101",
  38058=>"101101001",
  38059=>"000100101",
  38060=>"001111000",
  38061=>"111111001",
  38062=>"010101000",
  38063=>"010010010",
  38064=>"100010101",
  38065=>"000010010",
  38066=>"011001110",
  38067=>"001001110",
  38068=>"001110000",
  38069=>"010010000",
  38070=>"001101111",
  38071=>"100010100",
  38072=>"001000111",
  38073=>"111011010",
  38074=>"011100110",
  38075=>"001111000",
  38076=>"010110111",
  38077=>"011000011",
  38078=>"010001110",
  38079=>"101110101",
  38080=>"011001111",
  38081=>"000110010",
  38082=>"111000100",
  38083=>"000010100",
  38084=>"010101000",
  38085=>"000000011",
  38086=>"100100010",
  38087=>"000000010",
  38088=>"001111010",
  38089=>"001010111",
  38090=>"010010000",
  38091=>"010100011",
  38092=>"001010100",
  38093=>"010100000",
  38094=>"010000100",
  38095=>"100100111",
  38096=>"110000100",
  38097=>"011010001",
  38098=>"101001000",
  38099=>"011011110",
  38100=>"111110110",
  38101=>"101111000",
  38102=>"000111101",
  38103=>"011010011",
  38104=>"001100010",
  38105=>"000000010",
  38106=>"000010101",
  38107=>"000011001",
  38108=>"010000111",
  38109=>"100100000",
  38110=>"111000111",
  38111=>"000000111",
  38112=>"010110101",
  38113=>"110000010",
  38114=>"011000101",
  38115=>"110001111",
  38116=>"011001110",
  38117=>"011101001",
  38118=>"010111101",
  38119=>"101001011",
  38120=>"000010000",
  38121=>"111110110",
  38122=>"110101010",
  38123=>"101100000",
  38124=>"111100001",
  38125=>"111100010",
  38126=>"100100111",
  38127=>"010001100",
  38128=>"110101100",
  38129=>"101000100",
  38130=>"010110100",
  38131=>"101100111",
  38132=>"111001000",
  38133=>"010111111",
  38134=>"110110110",
  38135=>"000001111",
  38136=>"110100110",
  38137=>"001010011",
  38138=>"000100100",
  38139=>"100110110",
  38140=>"010000100",
  38141=>"101100010",
  38142=>"111001111",
  38143=>"110011011",
  38144=>"110011111",
  38145=>"101011101",
  38146=>"011111000",
  38147=>"110010110",
  38148=>"011001111",
  38149=>"101111101",
  38150=>"101101011",
  38151=>"001000011",
  38152=>"110000000",
  38153=>"110011100",
  38154=>"001010001",
  38155=>"100110000",
  38156=>"100101000",
  38157=>"011000101",
  38158=>"110100000",
  38159=>"101101110",
  38160=>"101001001",
  38161=>"101101110",
  38162=>"111101111",
  38163=>"010101111",
  38164=>"011100000",
  38165=>"011100100",
  38166=>"100001110",
  38167=>"011011101",
  38168=>"000011100",
  38169=>"000110101",
  38170=>"010100000",
  38171=>"001100100",
  38172=>"110101101",
  38173=>"011110011",
  38174=>"001011100",
  38175=>"101110000",
  38176=>"101000000",
  38177=>"001100100",
  38178=>"010111010",
  38179=>"101100111",
  38180=>"010010010",
  38181=>"010101101",
  38182=>"100000000",
  38183=>"000001001",
  38184=>"011000011",
  38185=>"010101010",
  38186=>"111011111",
  38187=>"101001011",
  38188=>"011111010",
  38189=>"111001101",
  38190=>"001100111",
  38191=>"011000010",
  38192=>"001100001",
  38193=>"000001111",
  38194=>"111101111",
  38195=>"101000111",
  38196=>"001010000",
  38197=>"110111110",
  38198=>"101010101",
  38199=>"100001011",
  38200=>"000000101",
  38201=>"110100000",
  38202=>"100000111",
  38203=>"010001111",
  38204=>"010010111",
  38205=>"000100101",
  38206=>"000000111",
  38207=>"011010111",
  38208=>"000100001",
  38209=>"010000101",
  38210=>"101000001",
  38211=>"101110111",
  38212=>"011001001",
  38213=>"010110000",
  38214=>"000010101",
  38215=>"000010110",
  38216=>"110110110",
  38217=>"100011011",
  38218=>"111101000",
  38219=>"001111001",
  38220=>"110111010",
  38221=>"100110100",
  38222=>"000110101",
  38223=>"000111000",
  38224=>"110110000",
  38225=>"010001111",
  38226=>"111100111",
  38227=>"100010011",
  38228=>"010100000",
  38229=>"001000110",
  38230=>"101101011",
  38231=>"111111101",
  38232=>"010000100",
  38233=>"110110111",
  38234=>"101111010",
  38235=>"111110100",
  38236=>"000110010",
  38237=>"010000100",
  38238=>"001000110",
  38239=>"010010100",
  38240=>"000111100",
  38241=>"101101010",
  38242=>"111111011",
  38243=>"001000000",
  38244=>"010110001",
  38245=>"011010010",
  38246=>"111001010",
  38247=>"111000010",
  38248=>"001011101",
  38249=>"010111110",
  38250=>"101000000",
  38251=>"100101101",
  38252=>"001100111",
  38253=>"111110110",
  38254=>"010000000",
  38255=>"010100011",
  38256=>"111101100",
  38257=>"011011111",
  38258=>"110111001",
  38259=>"111010011",
  38260=>"101111010",
  38261=>"011001000",
  38262=>"101101111",
  38263=>"110001100",
  38264=>"010111111",
  38265=>"111000100",
  38266=>"101001101",
  38267=>"100011010",
  38268=>"111100000",
  38269=>"001100110",
  38270=>"011000000",
  38271=>"000111110",
  38272=>"000000111",
  38273=>"000000000",
  38274=>"011010001",
  38275=>"001001110",
  38276=>"011011110",
  38277=>"101001110",
  38278=>"000100101",
  38279=>"111100100",
  38280=>"001000110",
  38281=>"000110100",
  38282=>"111111011",
  38283=>"000111101",
  38284=>"111000011",
  38285=>"111111000",
  38286=>"100110101",
  38287=>"000011100",
  38288=>"111111111",
  38289=>"000101010",
  38290=>"010101001",
  38291=>"001000011",
  38292=>"000001111",
  38293=>"111010010",
  38294=>"010111111",
  38295=>"000010010",
  38296=>"100111100",
  38297=>"011010010",
  38298=>"100010110",
  38299=>"001011011",
  38300=>"000111111",
  38301=>"100010010",
  38302=>"111110010",
  38303=>"001001000",
  38304=>"010010000",
  38305=>"010001011",
  38306=>"000001101",
  38307=>"111001101",
  38308=>"111010100",
  38309=>"000101011",
  38310=>"110101100",
  38311=>"010110011",
  38312=>"100110011",
  38313=>"111110101",
  38314=>"111111100",
  38315=>"000111100",
  38316=>"011001110",
  38317=>"100000010",
  38318=>"001100001",
  38319=>"101010011",
  38320=>"000111001",
  38321=>"111111110",
  38322=>"111111010",
  38323=>"011111111",
  38324=>"110100000",
  38325=>"010010001",
  38326=>"111111000",
  38327=>"001111010",
  38328=>"010100100",
  38329=>"000100011",
  38330=>"110100100",
  38331=>"011011111",
  38332=>"011011101",
  38333=>"101110101",
  38334=>"010001011",
  38335=>"011110001",
  38336=>"110110100",
  38337=>"111110000",
  38338=>"000001101",
  38339=>"101001110",
  38340=>"000000000",
  38341=>"100001010",
  38342=>"001101110",
  38343=>"011100000",
  38344=>"110100010",
  38345=>"011110010",
  38346=>"000000000",
  38347=>"111110111",
  38348=>"100000100",
  38349=>"111011001",
  38350=>"101100011",
  38351=>"000010111",
  38352=>"011110110",
  38353=>"101100110",
  38354=>"111101011",
  38355=>"111101000",
  38356=>"100010110",
  38357=>"001001000",
  38358=>"011000100",
  38359=>"010111101",
  38360=>"100001010",
  38361=>"110111110",
  38362=>"010000010",
  38363=>"110000000",
  38364=>"001000000",
  38365=>"000101110",
  38366=>"100101010",
  38367=>"000000000",
  38368=>"101111101",
  38369=>"110011011",
  38370=>"110110100",
  38371=>"001010000",
  38372=>"110110011",
  38373=>"111110000",
  38374=>"111100000",
  38375=>"011000111",
  38376=>"100100011",
  38377=>"100000111",
  38378=>"001011100",
  38379=>"000010010",
  38380=>"010010010",
  38381=>"011000101",
  38382=>"001110010",
  38383=>"001111110",
  38384=>"010000000",
  38385=>"100011110",
  38386=>"010000110",
  38387=>"110110000",
  38388=>"000010110",
  38389=>"111010011",
  38390=>"111100000",
  38391=>"000111110",
  38392=>"010010011",
  38393=>"111000101",
  38394=>"011101110",
  38395=>"110110000",
  38396=>"001111100",
  38397=>"001100111",
  38398=>"111010111",
  38399=>"101111111",
  38400=>"000110001",
  38401=>"001011100",
  38402=>"100011000",
  38403=>"100110101",
  38404=>"010001000",
  38405=>"001110101",
  38406=>"100000011",
  38407=>"100100001",
  38408=>"101111011",
  38409=>"011001001",
  38410=>"001011010",
  38411=>"101000111",
  38412=>"001000001",
  38413=>"000001000",
  38414=>"100100000",
  38415=>"111110011",
  38416=>"101011111",
  38417=>"001000110",
  38418=>"100000111",
  38419=>"000010011",
  38420=>"111011000",
  38421=>"011110010",
  38422=>"110110000",
  38423=>"110110101",
  38424=>"100110010",
  38425=>"101001001",
  38426=>"010100001",
  38427=>"100110100",
  38428=>"101110100",
  38429=>"100001100",
  38430=>"111111000",
  38431=>"111011001",
  38432=>"001011100",
  38433=>"010000001",
  38434=>"110110111",
  38435=>"001111111",
  38436=>"000001000",
  38437=>"100110111",
  38438=>"101111101",
  38439=>"111001111",
  38440=>"001111001",
  38441=>"100000010",
  38442=>"000000001",
  38443=>"011110011",
  38444=>"000111001",
  38445=>"101101011",
  38446=>"010101111",
  38447=>"001000100",
  38448=>"000001100",
  38449=>"111011010",
  38450=>"110010011",
  38451=>"001010101",
  38452=>"111011010",
  38453=>"000011001",
  38454=>"100011000",
  38455=>"100000000",
  38456=>"001100101",
  38457=>"111000100",
  38458=>"111001101",
  38459=>"011010000",
  38460=>"010110101",
  38461=>"001111000",
  38462=>"010001010",
  38463=>"010010010",
  38464=>"000000010",
  38465=>"000001001",
  38466=>"000010100",
  38467=>"110011001",
  38468=>"001001110",
  38469=>"101111011",
  38470=>"000110010",
  38471=>"110000011",
  38472=>"110100000",
  38473=>"111010011",
  38474=>"111000010",
  38475=>"010111101",
  38476=>"010110000",
  38477=>"001100001",
  38478=>"111011111",
  38479=>"000010000",
  38480=>"110110010",
  38481=>"111100010",
  38482=>"001111010",
  38483=>"000001001",
  38484=>"101011100",
  38485=>"000001000",
  38486=>"100011101",
  38487=>"111100101",
  38488=>"111111111",
  38489=>"011111101",
  38490=>"010100100",
  38491=>"001010000",
  38492=>"011111000",
  38493=>"000110011",
  38494=>"101011010",
  38495=>"010011011",
  38496=>"011101010",
  38497=>"000001001",
  38498=>"101110101",
  38499=>"100010010",
  38500=>"110011001",
  38501=>"010101110",
  38502=>"111110111",
  38503=>"111010011",
  38504=>"001000101",
  38505=>"111001110",
  38506=>"110110011",
  38507=>"001111101",
  38508=>"101110001",
  38509=>"101110110",
  38510=>"100110000",
  38511=>"110011000",
  38512=>"101101111",
  38513=>"010011000",
  38514=>"011010100",
  38515=>"001100111",
  38516=>"100110011",
  38517=>"110010111",
  38518=>"011110010",
  38519=>"010001000",
  38520=>"000011000",
  38521=>"100000000",
  38522=>"000001000",
  38523=>"100011001",
  38524=>"001111010",
  38525=>"010001111",
  38526=>"010111011",
  38527=>"001100011",
  38528=>"011001101",
  38529=>"100110101",
  38530=>"111111110",
  38531=>"110111000",
  38532=>"101010001",
  38533=>"100001001",
  38534=>"001010001",
  38535=>"010100000",
  38536=>"000010001",
  38537=>"010010100",
  38538=>"011101010",
  38539=>"001010100",
  38540=>"111111111",
  38541=>"111101011",
  38542=>"111000110",
  38543=>"000111011",
  38544=>"101010010",
  38545=>"100100000",
  38546=>"100111011",
  38547=>"100010100",
  38548=>"110100011",
  38549=>"100000011",
  38550=>"011100110",
  38551=>"010000001",
  38552=>"111110100",
  38553=>"101111110",
  38554=>"111111011",
  38555=>"101100010",
  38556=>"000101101",
  38557=>"010011010",
  38558=>"000011011",
  38559=>"000111111",
  38560=>"101000110",
  38561=>"101101101",
  38562=>"000111000",
  38563=>"111010101",
  38564=>"010001011",
  38565=>"010011110",
  38566=>"010100101",
  38567=>"000001011",
  38568=>"110101100",
  38569=>"000001101",
  38570=>"100100110",
  38571=>"111111001",
  38572=>"000100110",
  38573=>"111011011",
  38574=>"100010100",
  38575=>"110110111",
  38576=>"101000010",
  38577=>"000010111",
  38578=>"001000011",
  38579=>"110000100",
  38580=>"111110010",
  38581=>"011011010",
  38582=>"101010001",
  38583=>"101111100",
  38584=>"101111110",
  38585=>"110100010",
  38586=>"101111110",
  38587=>"000001000",
  38588=>"101011001",
  38589=>"110010110",
  38590=>"000001010",
  38591=>"110010111",
  38592=>"000001101",
  38593=>"000000001",
  38594=>"100010010",
  38595=>"100110011",
  38596=>"010110100",
  38597=>"111000000",
  38598=>"110001010",
  38599=>"000111011",
  38600=>"011000101",
  38601=>"111011111",
  38602=>"011000100",
  38603=>"101001011",
  38604=>"001000100",
  38605=>"001000011",
  38606=>"001000001",
  38607=>"100001100",
  38608=>"101101010",
  38609=>"011110100",
  38610=>"101110010",
  38611=>"111001000",
  38612=>"001001001",
  38613=>"011011001",
  38614=>"111010001",
  38615=>"101111101",
  38616=>"110010101",
  38617=>"110001000",
  38618=>"000101111",
  38619=>"101000100",
  38620=>"100100010",
  38621=>"101000111",
  38622=>"001111011",
  38623=>"001100010",
  38624=>"000001000",
  38625=>"110010000",
  38626=>"010111111",
  38627=>"101011100",
  38628=>"000111110",
  38629=>"101000110",
  38630=>"000000000",
  38631=>"010000010",
  38632=>"110010011",
  38633=>"100111101",
  38634=>"000000100",
  38635=>"000001100",
  38636=>"010110010",
  38637=>"110110001",
  38638=>"011100010",
  38639=>"000011000",
  38640=>"011000101",
  38641=>"000110011",
  38642=>"000010111",
  38643=>"100110101",
  38644=>"011010001",
  38645=>"111100010",
  38646=>"001000001",
  38647=>"101100100",
  38648=>"101111001",
  38649=>"011010011",
  38650=>"001101101",
  38651=>"110000001",
  38652=>"101001111",
  38653=>"010011110",
  38654=>"110010100",
  38655=>"101101001",
  38656=>"010000101",
  38657=>"101011101",
  38658=>"111001101",
  38659=>"000001110",
  38660=>"010000001",
  38661=>"011000101",
  38662=>"101000010",
  38663=>"010010110",
  38664=>"000110110",
  38665=>"110000011",
  38666=>"001110001",
  38667=>"001100111",
  38668=>"110010101",
  38669=>"100010100",
  38670=>"110110000",
  38671=>"010011111",
  38672=>"101010101",
  38673=>"110010111",
  38674=>"100110101",
  38675=>"110011101",
  38676=>"011010110",
  38677=>"101101111",
  38678=>"101000000",
  38679=>"000101000",
  38680=>"001010001",
  38681=>"000101000",
  38682=>"011010010",
  38683=>"011100010",
  38684=>"101101100",
  38685=>"000000011",
  38686=>"000111100",
  38687=>"111110100",
  38688=>"111110101",
  38689=>"100110000",
  38690=>"010110011",
  38691=>"110011111",
  38692=>"111011111",
  38693=>"010001000",
  38694=>"110010010",
  38695=>"111001000",
  38696=>"101011000",
  38697=>"101111111",
  38698=>"011011001",
  38699=>"110001000",
  38700=>"101111001",
  38701=>"000001011",
  38702=>"111010101",
  38703=>"001010111",
  38704=>"100011100",
  38705=>"000000010",
  38706=>"000100110",
  38707=>"000010000",
  38708=>"010111010",
  38709=>"011000101",
  38710=>"111001011",
  38711=>"101100101",
  38712=>"101110111",
  38713=>"111101001",
  38714=>"100110011",
  38715=>"111100010",
  38716=>"111000010",
  38717=>"010110011",
  38718=>"111010100",
  38719=>"010101010",
  38720=>"000110001",
  38721=>"000010110",
  38722=>"111000011",
  38723=>"001101100",
  38724=>"101100010",
  38725=>"000100101",
  38726=>"001111100",
  38727=>"110011100",
  38728=>"011110010",
  38729=>"001000000",
  38730=>"001111010",
  38731=>"110101101",
  38732=>"100011010",
  38733=>"001101111",
  38734=>"001011000",
  38735=>"100110101",
  38736=>"101001001",
  38737=>"011101111",
  38738=>"010001101",
  38739=>"100111001",
  38740=>"110010011",
  38741=>"000111011",
  38742=>"111111010",
  38743=>"101100110",
  38744=>"001000100",
  38745=>"011100010",
  38746=>"101010011",
  38747=>"100100110",
  38748=>"101010111",
  38749=>"011011101",
  38750=>"000111010",
  38751=>"000000000",
  38752=>"011011100",
  38753=>"000101001",
  38754=>"001000000",
  38755=>"000010010",
  38756=>"100011111",
  38757=>"000100101",
  38758=>"111100011",
  38759=>"101110001",
  38760=>"111000111",
  38761=>"000011111",
  38762=>"110100000",
  38763=>"111110001",
  38764=>"100000100",
  38765=>"000100000",
  38766=>"111001010",
  38767=>"000010101",
  38768=>"000100100",
  38769=>"100010010",
  38770=>"110110010",
  38771=>"101101111",
  38772=>"001101000",
  38773=>"001001100",
  38774=>"000000100",
  38775=>"000010010",
  38776=>"111100111",
  38777=>"110011001",
  38778=>"010000000",
  38779=>"111101000",
  38780=>"010101001",
  38781=>"101000011",
  38782=>"100101011",
  38783=>"000101100",
  38784=>"100011110",
  38785=>"011000010",
  38786=>"110010011",
  38787=>"001011111",
  38788=>"010000001",
  38789=>"001101101",
  38790=>"000001100",
  38791=>"101001111",
  38792=>"100101001",
  38793=>"010011100",
  38794=>"001011101",
  38795=>"010000011",
  38796=>"000011001",
  38797=>"000100000",
  38798=>"100101010",
  38799=>"010010001",
  38800=>"000000000",
  38801=>"001001000",
  38802=>"000110000",
  38803=>"010100001",
  38804=>"011100000",
  38805=>"111101101",
  38806=>"001100000",
  38807=>"011011101",
  38808=>"001111110",
  38809=>"000000100",
  38810=>"000110111",
  38811=>"100010000",
  38812=>"011001110",
  38813=>"100011000",
  38814=>"101000000",
  38815=>"000000011",
  38816=>"000000100",
  38817=>"010110010",
  38818=>"111111000",
  38819=>"001000010",
  38820=>"000000110",
  38821=>"101110110",
  38822=>"010111011",
  38823=>"000101111",
  38824=>"011001001",
  38825=>"111000111",
  38826=>"111110101",
  38827=>"010110101",
  38828=>"001011101",
  38829=>"000100010",
  38830=>"001000101",
  38831=>"100011001",
  38832=>"111111011",
  38833=>"111011101",
  38834=>"011101010",
  38835=>"100000010",
  38836=>"001011111",
  38837=>"011011010",
  38838=>"101010101",
  38839=>"011101001",
  38840=>"101010000",
  38841=>"010110010",
  38842=>"010010110",
  38843=>"101011100",
  38844=>"001101110",
  38845=>"101110010",
  38846=>"010100000",
  38847=>"010010100",
  38848=>"100000011",
  38849=>"100001001",
  38850=>"110111110",
  38851=>"111111111",
  38852=>"010101000",
  38853=>"100110101",
  38854=>"001010110",
  38855=>"101100001",
  38856=>"101101001",
  38857=>"111101000",
  38858=>"010001010",
  38859=>"001100001",
  38860=>"101111001",
  38861=>"010101010",
  38862=>"101010100",
  38863=>"000000011",
  38864=>"100111110",
  38865=>"111101100",
  38866=>"100000001",
  38867=>"101101111",
  38868=>"010011010",
  38869=>"100000001",
  38870=>"011000001",
  38871=>"000000000",
  38872=>"110011010",
  38873=>"100110011",
  38874=>"000100001",
  38875=>"111100111",
  38876=>"111011101",
  38877=>"000010010",
  38878=>"100001100",
  38879=>"011011100",
  38880=>"111111111",
  38881=>"111010000",
  38882=>"110111111",
  38883=>"000111111",
  38884=>"100100001",
  38885=>"000001000",
  38886=>"001100010",
  38887=>"111010000",
  38888=>"111111000",
  38889=>"001110101",
  38890=>"000100010",
  38891=>"111101100",
  38892=>"110111110",
  38893=>"011000000",
  38894=>"010100000",
  38895=>"001010111",
  38896=>"110110001",
  38897=>"010111011",
  38898=>"100100001",
  38899=>"100010111",
  38900=>"000100100",
  38901=>"100000000",
  38902=>"001011100",
  38903=>"000000001",
  38904=>"000111100",
  38905=>"010111011",
  38906=>"011100111",
  38907=>"110111101",
  38908=>"001001010",
  38909=>"010101110",
  38910=>"001100110",
  38911=>"100100001",
  38912=>"010000000",
  38913=>"111100100",
  38914=>"000000101",
  38915=>"011111101",
  38916=>"011011011",
  38917=>"001111100",
  38918=>"111110000",
  38919=>"000111000",
  38920=>"011010100",
  38921=>"110010110",
  38922=>"101100101",
  38923=>"110011100",
  38924=>"011011010",
  38925=>"100110110",
  38926=>"100100100",
  38927=>"100100001",
  38928=>"101111111",
  38929=>"100001100",
  38930=>"101111110",
  38931=>"010111001",
  38932=>"010011000",
  38933=>"011111001",
  38934=>"100110001",
  38935=>"000010110",
  38936=>"100111000",
  38937=>"001100111",
  38938=>"100101010",
  38939=>"111101110",
  38940=>"100001001",
  38941=>"000010010",
  38942=>"000111111",
  38943=>"011000100",
  38944=>"011101000",
  38945=>"110011011",
  38946=>"110111100",
  38947=>"111000010",
  38948=>"000010110",
  38949=>"111010010",
  38950=>"000000100",
  38951=>"110110000",
  38952=>"101001101",
  38953=>"011110100",
  38954=>"011010100",
  38955=>"011110011",
  38956=>"101011000",
  38957=>"000000011",
  38958=>"110010101",
  38959=>"010101111",
  38960=>"010101110",
  38961=>"010001001",
  38962=>"110010110",
  38963=>"100001111",
  38964=>"011010001",
  38965=>"000101000",
  38966=>"011001000",
  38967=>"011000101",
  38968=>"111000100",
  38969=>"101101110",
  38970=>"111111011",
  38971=>"100010000",
  38972=>"010111001",
  38973=>"101010101",
  38974=>"000100010",
  38975=>"101110111",
  38976=>"000001000",
  38977=>"011100101",
  38978=>"101000111",
  38979=>"101010100",
  38980=>"001101001",
  38981=>"011111000",
  38982=>"110101110",
  38983=>"001010011",
  38984=>"111101011",
  38985=>"001101111",
  38986=>"010110001",
  38987=>"111101011",
  38988=>"000001101",
  38989=>"011101101",
  38990=>"011010011",
  38991=>"100000111",
  38992=>"000101100",
  38993=>"010101111",
  38994=>"011101110",
  38995=>"001000001",
  38996=>"110000010",
  38997=>"110000010",
  38998=>"011110110",
  38999=>"110010101",
  39000=>"110010010",
  39001=>"101100110",
  39002=>"100010100",
  39003=>"010001000",
  39004=>"010100000",
  39005=>"100110000",
  39006=>"000011110",
  39007=>"011100101",
  39008=>"011101101",
  39009=>"000011010",
  39010=>"001011100",
  39011=>"000000010",
  39012=>"111111010",
  39013=>"000100011",
  39014=>"010010101",
  39015=>"101000100",
  39016=>"100110101",
  39017=>"000000001",
  39018=>"100100000",
  39019=>"000101110",
  39020=>"110101001",
  39021=>"011011000",
  39022=>"110101011",
  39023=>"101001011",
  39024=>"100100001",
  39025=>"000011110",
  39026=>"001000000",
  39027=>"110110100",
  39028=>"011011101",
  39029=>"011100011",
  39030=>"010101100",
  39031=>"100001101",
  39032=>"101100101",
  39033=>"110111110",
  39034=>"000000101",
  39035=>"101111011",
  39036=>"100011101",
  39037=>"000100001",
  39038=>"101011111",
  39039=>"010110100",
  39040=>"110001100",
  39041=>"000110110",
  39042=>"111011111",
  39043=>"110101010",
  39044=>"011011001",
  39045=>"101000000",
  39046=>"010110000",
  39047=>"110011001",
  39048=>"000011011",
  39049=>"100000010",
  39050=>"100101001",
  39051=>"011000011",
  39052=>"101010011",
  39053=>"100010011",
  39054=>"001101100",
  39055=>"010000101",
  39056=>"111000100",
  39057=>"000110111",
  39058=>"101001001",
  39059=>"100001001",
  39060=>"001000101",
  39061=>"100001001",
  39062=>"100110100",
  39063=>"101011000",
  39064=>"101101001",
  39065=>"110110100",
  39066=>"011001001",
  39067=>"011011100",
  39068=>"111110100",
  39069=>"000100010",
  39070=>"000000100",
  39071=>"111100011",
  39072=>"110100010",
  39073=>"100110011",
  39074=>"110110001",
  39075=>"010000000",
  39076=>"110111100",
  39077=>"000110101",
  39078=>"010101010",
  39079=>"000000000",
  39080=>"100110000",
  39081=>"011010011",
  39082=>"010101011",
  39083=>"011001011",
  39084=>"111100000",
  39085=>"110011011",
  39086=>"111100000",
  39087=>"010101000",
  39088=>"000001001",
  39089=>"000001110",
  39090=>"011010011",
  39091=>"000011101",
  39092=>"100111100",
  39093=>"101100111",
  39094=>"011101110",
  39095=>"111110101",
  39096=>"000010011",
  39097=>"000100000",
  39098=>"000110001",
  39099=>"011011101",
  39100=>"001001000",
  39101=>"000001000",
  39102=>"001110101",
  39103=>"100100001",
  39104=>"111000110",
  39105=>"011100011",
  39106=>"011000000",
  39107=>"001000100",
  39108=>"110110010",
  39109=>"001101111",
  39110=>"111101001",
  39111=>"101011101",
  39112=>"001001100",
  39113=>"111010101",
  39114=>"101001001",
  39115=>"010111101",
  39116=>"011001110",
  39117=>"001100110",
  39118=>"110111110",
  39119=>"001100101",
  39120=>"000101001",
  39121=>"100100111",
  39122=>"000101000",
  39123=>"101111110",
  39124=>"111101101",
  39125=>"111100001",
  39126=>"000010100",
  39127=>"001011001",
  39128=>"101101000",
  39129=>"111010111",
  39130=>"110110101",
  39131=>"000001000",
  39132=>"010000001",
  39133=>"001000000",
  39134=>"011100100",
  39135=>"111110010",
  39136=>"000010100",
  39137=>"000110000",
  39138=>"101010101",
  39139=>"011110111",
  39140=>"110010110",
  39141=>"111101101",
  39142=>"100001101",
  39143=>"100101111",
  39144=>"001110010",
  39145=>"011101100",
  39146=>"101000001",
  39147=>"000001101",
  39148=>"001100100",
  39149=>"100101001",
  39150=>"110000010",
  39151=>"011110011",
  39152=>"000101111",
  39153=>"001011001",
  39154=>"001100101",
  39155=>"000001001",
  39156=>"111011011",
  39157=>"101100001",
  39158=>"111100110",
  39159=>"110010001",
  39160=>"111101000",
  39161=>"110100111",
  39162=>"110000010",
  39163=>"010011001",
  39164=>"100001111",
  39165=>"111111000",
  39166=>"001111111",
  39167=>"010000000",
  39168=>"100101110",
  39169=>"110101111",
  39170=>"011010011",
  39171=>"100101101",
  39172=>"110100010",
  39173=>"101110011",
  39174=>"101110000",
  39175=>"100000101",
  39176=>"110111101",
  39177=>"111111100",
  39178=>"101100101",
  39179=>"010010100",
  39180=>"100011011",
  39181=>"100000001",
  39182=>"111001100",
  39183=>"101101011",
  39184=>"010001010",
  39185=>"100011011",
  39186=>"111111001",
  39187=>"110101001",
  39188=>"000001001",
  39189=>"100100101",
  39190=>"111010111",
  39191=>"001111111",
  39192=>"111110100",
  39193=>"100011000",
  39194=>"100010010",
  39195=>"101001100",
  39196=>"100101011",
  39197=>"000010101",
  39198=>"101011001",
  39199=>"111101001",
  39200=>"011101100",
  39201=>"111110010",
  39202=>"010011000",
  39203=>"011001111",
  39204=>"000010101",
  39205=>"101111010",
  39206=>"100001011",
  39207=>"011000000",
  39208=>"101100111",
  39209=>"101010001",
  39210=>"110110111",
  39211=>"100100010",
  39212=>"110100000",
  39213=>"001000011",
  39214=>"111010010",
  39215=>"100011101",
  39216=>"011001100",
  39217=>"010111101",
  39218=>"111001011",
  39219=>"000100111",
  39220=>"101101100",
  39221=>"001100100",
  39222=>"110110111",
  39223=>"010101100",
  39224=>"011001101",
  39225=>"000101110",
  39226=>"111010000",
  39227=>"111110011",
  39228=>"010111001",
  39229=>"101110111",
  39230=>"000110001",
  39231=>"100001100",
  39232=>"000011110",
  39233=>"010011110",
  39234=>"110101010",
  39235=>"010001111",
  39236=>"011110100",
  39237=>"011000101",
  39238=>"001100001",
  39239=>"000110000",
  39240=>"100001100",
  39241=>"100010101",
  39242=>"001000101",
  39243=>"110010000",
  39244=>"001010111",
  39245=>"110001001",
  39246=>"110110111",
  39247=>"000000001",
  39248=>"101110001",
  39249=>"011101111",
  39250=>"101101101",
  39251=>"010101101",
  39252=>"001110101",
  39253=>"100011110",
  39254=>"100111110",
  39255=>"101100101",
  39256=>"111001111",
  39257=>"010000011",
  39258=>"011101000",
  39259=>"010111110",
  39260=>"100001110",
  39261=>"110000110",
  39262=>"101110111",
  39263=>"101110001",
  39264=>"110100000",
  39265=>"000110000",
  39266=>"001010010",
  39267=>"110001110",
  39268=>"011011101",
  39269=>"100010100",
  39270=>"011011100",
  39271=>"011111000",
  39272=>"011110110",
  39273=>"010010001",
  39274=>"111001011",
  39275=>"111001011",
  39276=>"010100000",
  39277=>"010110110",
  39278=>"011011011",
  39279=>"010100010",
  39280=>"011000101",
  39281=>"110011100",
  39282=>"011110010",
  39283=>"111001100",
  39284=>"000001001",
  39285=>"101011111",
  39286=>"100011111",
  39287=>"110101001",
  39288=>"000101100",
  39289=>"010110111",
  39290=>"011100100",
  39291=>"111011110",
  39292=>"001110100",
  39293=>"010111100",
  39294=>"001110011",
  39295=>"000001100",
  39296=>"001001011",
  39297=>"001011100",
  39298=>"000111010",
  39299=>"100100011",
  39300=>"101100111",
  39301=>"101010101",
  39302=>"111110001",
  39303=>"010010100",
  39304=>"001000001",
  39305=>"110101010",
  39306=>"111011011",
  39307=>"111110111",
  39308=>"001100001",
  39309=>"011101000",
  39310=>"001000011",
  39311=>"011111110",
  39312=>"010110000",
  39313=>"111110110",
  39314=>"110111010",
  39315=>"000011111",
  39316=>"111011100",
  39317=>"001000110",
  39318=>"001100011",
  39319=>"101000000",
  39320=>"001101111",
  39321=>"000010111",
  39322=>"010011110",
  39323=>"101001100",
  39324=>"111010011",
  39325=>"011100001",
  39326=>"011010111",
  39327=>"101101000",
  39328=>"000000100",
  39329=>"000001010",
  39330=>"111000000",
  39331=>"110100000",
  39332=>"001000001",
  39333=>"000100110",
  39334=>"101110111",
  39335=>"111110010",
  39336=>"100011011",
  39337=>"010001000",
  39338=>"111010000",
  39339=>"010101011",
  39340=>"010100011",
  39341=>"101001110",
  39342=>"111111011",
  39343=>"111011101",
  39344=>"001100100",
  39345=>"001010000",
  39346=>"001001000",
  39347=>"111110100",
  39348=>"111111100",
  39349=>"011000001",
  39350=>"100101110",
  39351=>"011101011",
  39352=>"010111100",
  39353=>"000100011",
  39354=>"001000000",
  39355=>"100000101",
  39356=>"011110110",
  39357=>"010011000",
  39358=>"011111100",
  39359=>"011110110",
  39360=>"011111010",
  39361=>"011101011",
  39362=>"111011010",
  39363=>"010110011",
  39364=>"110011011",
  39365=>"100000010",
  39366=>"111001011",
  39367=>"010110010",
  39368=>"011100010",
  39369=>"010010010",
  39370=>"001101010",
  39371=>"010000001",
  39372=>"001111000",
  39373=>"000010011",
  39374=>"000000100",
  39375=>"100101000",
  39376=>"101100011",
  39377=>"010101010",
  39378=>"000000101",
  39379=>"001011001",
  39380=>"011101001",
  39381=>"100011010",
  39382=>"100010001",
  39383=>"100100000",
  39384=>"010101100",
  39385=>"110101010",
  39386=>"011011100",
  39387=>"011110011",
  39388=>"110001000",
  39389=>"110010101",
  39390=>"110010100",
  39391=>"101000111",
  39392=>"011010010",
  39393=>"011000110",
  39394=>"110011000",
  39395=>"100000011",
  39396=>"001100111",
  39397=>"000000101",
  39398=>"001010111",
  39399=>"000011001",
  39400=>"111011101",
  39401=>"111101111",
  39402=>"100011100",
  39403=>"001110000",
  39404=>"110110000",
  39405=>"101000010",
  39406=>"000000001",
  39407=>"001001000",
  39408=>"000000011",
  39409=>"100101110",
  39410=>"011111100",
  39411=>"000011000",
  39412=>"111011010",
  39413=>"011111000",
  39414=>"100011011",
  39415=>"011101001",
  39416=>"111111110",
  39417=>"011010111",
  39418=>"101100011",
  39419=>"001010110",
  39420=>"110011000",
  39421=>"010100001",
  39422=>"110000100",
  39423=>"000101101",
  39424=>"100001000",
  39425=>"011100000",
  39426=>"101001001",
  39427=>"000010001",
  39428=>"111111111",
  39429=>"010010010",
  39430=>"101111111",
  39431=>"001000111",
  39432=>"001001010",
  39433=>"111010111",
  39434=>"101011001",
  39435=>"100100000",
  39436=>"111000010",
  39437=>"011001111",
  39438=>"001011110",
  39439=>"101110011",
  39440=>"010100100",
  39441=>"010101111",
  39442=>"010100010",
  39443=>"000100100",
  39444=>"001111010",
  39445=>"101110100",
  39446=>"010001110",
  39447=>"011100001",
  39448=>"001001110",
  39449=>"001110010",
  39450=>"110111001",
  39451=>"011010100",
  39452=>"001000111",
  39453=>"001011000",
  39454=>"011001000",
  39455=>"001111111",
  39456=>"111101000",
  39457=>"011010010",
  39458=>"111000010",
  39459=>"100100011",
  39460=>"011111101",
  39461=>"100000011",
  39462=>"011111000",
  39463=>"010001110",
  39464=>"000101010",
  39465=>"111101010",
  39466=>"010000010",
  39467=>"000011111",
  39468=>"000000010",
  39469=>"110110001",
  39470=>"010111110",
  39471=>"000000111",
  39472=>"010110010",
  39473=>"111100111",
  39474=>"001111011",
  39475=>"110110111",
  39476=>"001011100",
  39477=>"101010100",
  39478=>"001000000",
  39479=>"010010001",
  39480=>"100110101",
  39481=>"011010110",
  39482=>"001111101",
  39483=>"101100101",
  39484=>"010111101",
  39485=>"000001001",
  39486=>"100001010",
  39487=>"010111101",
  39488=>"101010100",
  39489=>"000011101",
  39490=>"001101100",
  39491=>"101111111",
  39492=>"100000110",
  39493=>"111111001",
  39494=>"110010001",
  39495=>"001010101",
  39496=>"110111000",
  39497=>"110111111",
  39498=>"101100111",
  39499=>"111111010",
  39500=>"111010001",
  39501=>"011111000",
  39502=>"101011010",
  39503=>"010110011",
  39504=>"110110011",
  39505=>"000111000",
  39506=>"110011101",
  39507=>"100100110",
  39508=>"011010100",
  39509=>"111110111",
  39510=>"100001011",
  39511=>"010011011",
  39512=>"010010110",
  39513=>"101100100",
  39514=>"110000000",
  39515=>"000011011",
  39516=>"100101111",
  39517=>"000001101",
  39518=>"010011000",
  39519=>"001110100",
  39520=>"000001011",
  39521=>"100101111",
  39522=>"000001010",
  39523=>"011001110",
  39524=>"010011100",
  39525=>"110100001",
  39526=>"000010000",
  39527=>"111001011",
  39528=>"101011101",
  39529=>"110000111",
  39530=>"110011010",
  39531=>"101001100",
  39532=>"011011001",
  39533=>"100111101",
  39534=>"111101001",
  39535=>"101011011",
  39536=>"111111101",
  39537=>"110001001",
  39538=>"101011011",
  39539=>"000110111",
  39540=>"010111100",
  39541=>"000111110",
  39542=>"100000110",
  39543=>"101100111",
  39544=>"110010111",
  39545=>"111111011",
  39546=>"001100010",
  39547=>"110110110",
  39548=>"100111110",
  39549=>"101100010",
  39550=>"000110101",
  39551=>"100101001",
  39552=>"010010001",
  39553=>"011111110",
  39554=>"101000110",
  39555=>"000000110",
  39556=>"011000111",
  39557=>"010010000",
  39558=>"000010111",
  39559=>"000000100",
  39560=>"001111110",
  39561=>"110010001",
  39562=>"110001100",
  39563=>"011111010",
  39564=>"100101001",
  39565=>"110001110",
  39566=>"110111010",
  39567=>"110010011",
  39568=>"011000011",
  39569=>"011110101",
  39570=>"000000111",
  39571=>"001100111",
  39572=>"011111001",
  39573=>"111010100",
  39574=>"010110000",
  39575=>"101101110",
  39576=>"100010100",
  39577=>"110011011",
  39578=>"001110010",
  39579=>"100100000",
  39580=>"110111110",
  39581=>"101101110",
  39582=>"111000000",
  39583=>"000110001",
  39584=>"111101001",
  39585=>"001000000",
  39586=>"111101110",
  39587=>"100010011",
  39588=>"011000010",
  39589=>"010100010",
  39590=>"100100001",
  39591=>"100000010",
  39592=>"001111100",
  39593=>"001100110",
  39594=>"100110110",
  39595=>"001001010",
  39596=>"000011110",
  39597=>"101100011",
  39598=>"111111000",
  39599=>"010010000",
  39600=>"011010110",
  39601=>"100111101",
  39602=>"010011001",
  39603=>"001101000",
  39604=>"000100101",
  39605=>"110111101",
  39606=>"111000001",
  39607=>"101010000",
  39608=>"011000101",
  39609=>"010101100",
  39610=>"000111111",
  39611=>"110001110",
  39612=>"100100001",
  39613=>"101110001",
  39614=>"111011101",
  39615=>"001001100",
  39616=>"101010011",
  39617=>"001011101",
  39618=>"001000111",
  39619=>"101111101",
  39620=>"111011011",
  39621=>"010110100",
  39622=>"100011111",
  39623=>"101000010",
  39624=>"101000000",
  39625=>"001100010",
  39626=>"111011110",
  39627=>"011011001",
  39628=>"101010011",
  39629=>"000011010",
  39630=>"111101110",
  39631=>"100111001",
  39632=>"101001010",
  39633=>"110000001",
  39634=>"100010010",
  39635=>"000011110",
  39636=>"101001100",
  39637=>"000011001",
  39638=>"100011100",
  39639=>"011111011",
  39640=>"111100000",
  39641=>"100101101",
  39642=>"111001110",
  39643=>"010101100",
  39644=>"100001111",
  39645=>"010101100",
  39646=>"001100100",
  39647=>"111010010",
  39648=>"100101100",
  39649=>"101111001",
  39650=>"001001000",
  39651=>"001101110",
  39652=>"100000110",
  39653=>"101011000",
  39654=>"001110000",
  39655=>"100001100",
  39656=>"001110011",
  39657=>"011110011",
  39658=>"010111010",
  39659=>"010010000",
  39660=>"010110100",
  39661=>"101111010",
  39662=>"110011010",
  39663=>"111010011",
  39664=>"111100000",
  39665=>"101001000",
  39666=>"110011111",
  39667=>"101100101",
  39668=>"011010110",
  39669=>"100100101",
  39670=>"101111011",
  39671=>"101001011",
  39672=>"010000010",
  39673=>"111111101",
  39674=>"000101000",
  39675=>"011111111",
  39676=>"010100111",
  39677=>"100111010",
  39678=>"011100011",
  39679=>"001111011",
  39680=>"010101111",
  39681=>"100100010",
  39682=>"001001001",
  39683=>"100001101",
  39684=>"000010011",
  39685=>"001011000",
  39686=>"111001000",
  39687=>"010101011",
  39688=>"110010100",
  39689=>"111010101",
  39690=>"101101000",
  39691=>"000100000",
  39692=>"101001000",
  39693=>"010000000",
  39694=>"111010110",
  39695=>"011110101",
  39696=>"000000000",
  39697=>"001101000",
  39698=>"110000011",
  39699=>"100001101",
  39700=>"001000000",
  39701=>"110001011",
  39702=>"011011100",
  39703=>"100001011",
  39704=>"000111001",
  39705=>"011101010",
  39706=>"010100000",
  39707=>"110100011",
  39708=>"111111001",
  39709=>"111000101",
  39710=>"000100101",
  39711=>"000110011",
  39712=>"110111010",
  39713=>"110011011",
  39714=>"000011101",
  39715=>"110111111",
  39716=>"101111110",
  39717=>"001010001",
  39718=>"010111100",
  39719=>"000011110",
  39720=>"010001101",
  39721=>"111111000",
  39722=>"111111111",
  39723=>"110101010",
  39724=>"100100101",
  39725=>"000000011",
  39726=>"001111111",
  39727=>"110111010",
  39728=>"100000101",
  39729=>"110011001",
  39730=>"110110110",
  39731=>"001111000",
  39732=>"110010100",
  39733=>"001110000",
  39734=>"101110000",
  39735=>"011000100",
  39736=>"100110000",
  39737=>"111000011",
  39738=>"001100111",
  39739=>"010011111",
  39740=>"111011111",
  39741=>"111110011",
  39742=>"000001000",
  39743=>"101011010",
  39744=>"100101100",
  39745=>"001011010",
  39746=>"001111001",
  39747=>"101110011",
  39748=>"001111110",
  39749=>"000110100",
  39750=>"110100000",
  39751=>"001101011",
  39752=>"000011100",
  39753=>"111100011",
  39754=>"011010110",
  39755=>"100000110",
  39756=>"000101110",
  39757=>"010101111",
  39758=>"110000011",
  39759=>"100111011",
  39760=>"001101101",
  39761=>"000001000",
  39762=>"111111111",
  39763=>"010101010",
  39764=>"000101000",
  39765=>"011110000",
  39766=>"001111011",
  39767=>"101001100",
  39768=>"001111000",
  39769=>"110100111",
  39770=>"000000101",
  39771=>"011100110",
  39772=>"010100110",
  39773=>"100110000",
  39774=>"010010100",
  39775=>"010011110",
  39776=>"100000000",
  39777=>"100010011",
  39778=>"010110100",
  39779=>"110110100",
  39780=>"010000100",
  39781=>"110100101",
  39782=>"100111011",
  39783=>"111110001",
  39784=>"100000010",
  39785=>"001001000",
  39786=>"110000000",
  39787=>"101101101",
  39788=>"111010110",
  39789=>"011100111",
  39790=>"111100111",
  39791=>"110010111",
  39792=>"111000100",
  39793=>"001100101",
  39794=>"001111010",
  39795=>"010011110",
  39796=>"100000001",
  39797=>"110010011",
  39798=>"111010001",
  39799=>"011011000",
  39800=>"000010001",
  39801=>"100000000",
  39802=>"110111011",
  39803=>"111000101",
  39804=>"110100110",
  39805=>"101111101",
  39806=>"101000011",
  39807=>"001011001",
  39808=>"101001000",
  39809=>"001010100",
  39810=>"011100011",
  39811=>"010001111",
  39812=>"111001101",
  39813=>"101100011",
  39814=>"001011110",
  39815=>"011100100",
  39816=>"100010101",
  39817=>"111011100",
  39818=>"110101010",
  39819=>"110101100",
  39820=>"001010110",
  39821=>"010100110",
  39822=>"000111011",
  39823=>"110010110",
  39824=>"011001010",
  39825=>"000000010",
  39826=>"011000011",
  39827=>"101101111",
  39828=>"001001010",
  39829=>"101101100",
  39830=>"010100000",
  39831=>"010110001",
  39832=>"010101010",
  39833=>"000000001",
  39834=>"010101111",
  39835=>"001110001",
  39836=>"100101110",
  39837=>"000101101",
  39838=>"111010010",
  39839=>"100111110",
  39840=>"100100100",
  39841=>"100100110",
  39842=>"100010110",
  39843=>"100000010",
  39844=>"111000100",
  39845=>"011111111",
  39846=>"100001001",
  39847=>"110100100",
  39848=>"000110101",
  39849=>"111011010",
  39850=>"000111010",
  39851=>"001111010",
  39852=>"001010000",
  39853=>"000001100",
  39854=>"010010110",
  39855=>"111000100",
  39856=>"011011100",
  39857=>"000111101",
  39858=>"100110100",
  39859=>"110111101",
  39860=>"111000111",
  39861=>"000010110",
  39862=>"010101001",
  39863=>"111101011",
  39864=>"111101101",
  39865=>"000010110",
  39866=>"011010101",
  39867=>"110000010",
  39868=>"111010010",
  39869=>"001100000",
  39870=>"010000101",
  39871=>"001111100",
  39872=>"010011100",
  39873=>"101111000",
  39874=>"100110010",
  39875=>"100101110",
  39876=>"011001111",
  39877=>"100110101",
  39878=>"010000001",
  39879=>"010100010",
  39880=>"000101111",
  39881=>"010101000",
  39882=>"110000111",
  39883=>"100001001",
  39884=>"011111111",
  39885=>"000000000",
  39886=>"100000001",
  39887=>"010111101",
  39888=>"010001001",
  39889=>"000110101",
  39890=>"010011011",
  39891=>"000110000",
  39892=>"111111111",
  39893=>"110111100",
  39894=>"110010110",
  39895=>"010000010",
  39896=>"100101111",
  39897=>"111101110",
  39898=>"001110101",
  39899=>"111000010",
  39900=>"010001100",
  39901=>"010000111",
  39902=>"010001111",
  39903=>"101000000",
  39904=>"000100100",
  39905=>"000000001",
  39906=>"100000001",
  39907=>"000001100",
  39908=>"011010010",
  39909=>"101010111",
  39910=>"000010100",
  39911=>"100010100",
  39912=>"110010010",
  39913=>"011011011",
  39914=>"001000101",
  39915=>"100001010",
  39916=>"010101100",
  39917=>"110011001",
  39918=>"010110010",
  39919=>"101011010",
  39920=>"101011000",
  39921=>"001101000",
  39922=>"001101101",
  39923=>"100001011",
  39924=>"101101100",
  39925=>"100110100",
  39926=>"001000000",
  39927=>"000010010",
  39928=>"000001010",
  39929=>"101111001",
  39930=>"010000000",
  39931=>"010111001",
  39932=>"010101001",
  39933=>"011100000",
  39934=>"111101011",
  39935=>"011100001",
  39936=>"000101000",
  39937=>"001110010",
  39938=>"010111010",
  39939=>"101001011",
  39940=>"011110001",
  39941=>"010110100",
  39942=>"101011000",
  39943=>"111011010",
  39944=>"010010111",
  39945=>"110000100",
  39946=>"111010100",
  39947=>"100001001",
  39948=>"010010000",
  39949=>"111010111",
  39950=>"011010110",
  39951=>"001111000",
  39952=>"001101010",
  39953=>"001000111",
  39954=>"010011110",
  39955=>"000011000",
  39956=>"111101110",
  39957=>"001001110",
  39958=>"000100110",
  39959=>"101110110",
  39960=>"011101001",
  39961=>"000010000",
  39962=>"101111011",
  39963=>"001101001",
  39964=>"010101000",
  39965=>"111100000",
  39966=>"111001010",
  39967=>"101100100",
  39968=>"101011010",
  39969=>"010001110",
  39970=>"111010000",
  39971=>"100011011",
  39972=>"111101000",
  39973=>"000000001",
  39974=>"010110010",
  39975=>"100001111",
  39976=>"110010000",
  39977=>"001110001",
  39978=>"000010101",
  39979=>"100110111",
  39980=>"000001000",
  39981=>"000111111",
  39982=>"000010110",
  39983=>"010110000",
  39984=>"100011011",
  39985=>"100110010",
  39986=>"110110101",
  39987=>"100010010",
  39988=>"101110110",
  39989=>"000011000",
  39990=>"000000000",
  39991=>"010101001",
  39992=>"111111110",
  39993=>"111101001",
  39994=>"011101011",
  39995=>"101111111",
  39996=>"000010100",
  39997=>"011101000",
  39998=>"001100011",
  39999=>"010101111",
  40000=>"100011101",
  40001=>"001000010",
  40002=>"100000111",
  40003=>"110111111",
  40004=>"110000010",
  40005=>"000010100",
  40006=>"100110011",
  40007=>"111000000",
  40008=>"110111110",
  40009=>"111011111",
  40010=>"101100010",
  40011=>"111000100",
  40012=>"010111010",
  40013=>"100011000",
  40014=>"011011100",
  40015=>"010111100",
  40016=>"100100000",
  40017=>"000000000",
  40018=>"010111110",
  40019=>"101001000",
  40020=>"111100011",
  40021=>"100111100",
  40022=>"101100100",
  40023=>"110100011",
  40024=>"101011011",
  40025=>"100000100",
  40026=>"111001000",
  40027=>"001100111",
  40028=>"001100100",
  40029=>"010110011",
  40030=>"001000001",
  40031=>"011010110",
  40032=>"110010001",
  40033=>"111010100",
  40034=>"001000000",
  40035=>"010010010",
  40036=>"101001000",
  40037=>"011101011",
  40038=>"111111100",
  40039=>"000111100",
  40040=>"001111110",
  40041=>"000010111",
  40042=>"100101001",
  40043=>"111110011",
  40044=>"010001110",
  40045=>"111100101",
  40046=>"001010111",
  40047=>"011011000",
  40048=>"111100100",
  40049=>"010100100",
  40050=>"100101001",
  40051=>"101010111",
  40052=>"110010110",
  40053=>"010101010",
  40054=>"100101100",
  40055=>"011110100",
  40056=>"100001000",
  40057=>"110110000",
  40058=>"011111111",
  40059=>"010110111",
  40060=>"100101001",
  40061=>"000011101",
  40062=>"110010001",
  40063=>"001000000",
  40064=>"100101000",
  40065=>"001101001",
  40066=>"011000110",
  40067=>"100011010",
  40068=>"011010000",
  40069=>"011101110",
  40070=>"101001000",
  40071=>"110100110",
  40072=>"111011100",
  40073=>"001010011",
  40074=>"100000000",
  40075=>"011011011",
  40076=>"110110100",
  40077=>"100000100",
  40078=>"101110101",
  40079=>"001000010",
  40080=>"111100110",
  40081=>"011100011",
  40082=>"001010110",
  40083=>"000000010",
  40084=>"111010000",
  40085=>"011111111",
  40086=>"111110100",
  40087=>"011010000",
  40088=>"111010110",
  40089=>"110100001",
  40090=>"000010001",
  40091=>"110010000",
  40092=>"101011000",
  40093=>"010000010",
  40094=>"011011100",
  40095=>"110110110",
  40096=>"000011100",
  40097=>"111101101",
  40098=>"000111111",
  40099=>"000111111",
  40100=>"111110110",
  40101=>"001011011",
  40102=>"100101011",
  40103=>"111100010",
  40104=>"000111011",
  40105=>"010010001",
  40106=>"101101110",
  40107=>"011100111",
  40108=>"100010111",
  40109=>"111110111",
  40110=>"101101111",
  40111=>"111000111",
  40112=>"100100000",
  40113=>"100001001",
  40114=>"111110000",
  40115=>"010110001",
  40116=>"100111100",
  40117=>"011100000",
  40118=>"111111110",
  40119=>"010111000",
  40120=>"101001101",
  40121=>"011110111",
  40122=>"010010101",
  40123=>"101001110",
  40124=>"101100110",
  40125=>"111010001",
  40126=>"000010111",
  40127=>"100101000",
  40128=>"011011111",
  40129=>"011010000",
  40130=>"101011011",
  40131=>"000001000",
  40132=>"111110010",
  40133=>"010100100",
  40134=>"001100000",
  40135=>"101000010",
  40136=>"000011111",
  40137=>"100010000",
  40138=>"001101111",
  40139=>"111001111",
  40140=>"000101000",
  40141=>"000111110",
  40142=>"100010100",
  40143=>"111000100",
  40144=>"010011111",
  40145=>"110000100",
  40146=>"100011000",
  40147=>"011000110",
  40148=>"010100110",
  40149=>"011001010",
  40150=>"001111101",
  40151=>"111000111",
  40152=>"111100010",
  40153=>"000100100",
  40154=>"110111111",
  40155=>"001000111",
  40156=>"001011010",
  40157=>"110110101",
  40158=>"001101000",
  40159=>"101110010",
  40160=>"001000110",
  40161=>"110000101",
  40162=>"101110100",
  40163=>"000000010",
  40164=>"110010100",
  40165=>"000001010",
  40166=>"011000000",
  40167=>"001111100",
  40168=>"110000100",
  40169=>"111010010",
  40170=>"110110100",
  40171=>"010110011",
  40172=>"111000011",
  40173=>"111010001",
  40174=>"000000101",
  40175=>"001100001",
  40176=>"111111010",
  40177=>"101010001",
  40178=>"010011000",
  40179=>"101101010",
  40180=>"110111100",
  40181=>"110110000",
  40182=>"111010000",
  40183=>"111010000",
  40184=>"011010110",
  40185=>"010101110",
  40186=>"111110100",
  40187=>"111011110",
  40188=>"101110101",
  40189=>"011110100",
  40190=>"010011111",
  40191=>"111100011",
  40192=>"001110111",
  40193=>"100000000",
  40194=>"000101111",
  40195=>"100101101",
  40196=>"110110010",
  40197=>"000000011",
  40198=>"010111000",
  40199=>"011110111",
  40200=>"111101011",
  40201=>"111111110",
  40202=>"111110001",
  40203=>"010010010",
  40204=>"110001010",
  40205=>"011111000",
  40206=>"111101000",
  40207=>"000111110",
  40208=>"011100100",
  40209=>"111000011",
  40210=>"011101111",
  40211=>"100100010",
  40212=>"011000111",
  40213=>"011101011",
  40214=>"011000000",
  40215=>"010111100",
  40216=>"010100110",
  40217=>"100011110",
  40218=>"100001000",
  40219=>"110010111",
  40220=>"110100100",
  40221=>"000000101",
  40222=>"011101011",
  40223=>"000010110",
  40224=>"000101100",
  40225=>"011100101",
  40226=>"110011100",
  40227=>"110100010",
  40228=>"010000100",
  40229=>"110001110",
  40230=>"111001001",
  40231=>"101101011",
  40232=>"001000100",
  40233=>"100001101",
  40234=>"111000010",
  40235=>"100001111",
  40236=>"010101011",
  40237=>"000000000",
  40238=>"000000001",
  40239=>"101000101",
  40240=>"011000001",
  40241=>"100101101",
  40242=>"101100010",
  40243=>"101010000",
  40244=>"010010000",
  40245=>"000111101",
  40246=>"100011101",
  40247=>"100001111",
  40248=>"111110111",
  40249=>"001000011",
  40250=>"000101101",
  40251=>"100011011",
  40252=>"010000111",
  40253=>"010100011",
  40254=>"111111101",
  40255=>"000001100",
  40256=>"100000000",
  40257=>"001010111",
  40258=>"000101101",
  40259=>"100100010",
  40260=>"100101011",
  40261=>"110100111",
  40262=>"011000100",
  40263=>"100010011",
  40264=>"000011000",
  40265=>"001111001",
  40266=>"100010000",
  40267=>"000010000",
  40268=>"001001010",
  40269=>"101111111",
  40270=>"001111111",
  40271=>"001100000",
  40272=>"101001001",
  40273=>"111111100",
  40274=>"000100101",
  40275=>"110001111",
  40276=>"111111011",
  40277=>"001010101",
  40278=>"000000101",
  40279=>"011011100",
  40280=>"111011000",
  40281=>"101001010",
  40282=>"000011111",
  40283=>"010111010",
  40284=>"001101100",
  40285=>"101110101",
  40286=>"111111110",
  40287=>"010100000",
  40288=>"011000000",
  40289=>"000011001",
  40290=>"111101011",
  40291=>"001111111",
  40292=>"101111010",
  40293=>"011001100",
  40294=>"110111100",
  40295=>"010100001",
  40296=>"000111011",
  40297=>"101000000",
  40298=>"101100111",
  40299=>"100000000",
  40300=>"001100110",
  40301=>"001011000",
  40302=>"111011011",
  40303=>"101100100",
  40304=>"100000010",
  40305=>"011001110",
  40306=>"011010011",
  40307=>"111001000",
  40308=>"100010110",
  40309=>"011011010",
  40310=>"110001111",
  40311=>"110011000",
  40312=>"010101001",
  40313=>"111000101",
  40314=>"111100101",
  40315=>"011101001",
  40316=>"011100010",
  40317=>"111101010",
  40318=>"000000001",
  40319=>"001100001",
  40320=>"001110000",
  40321=>"011101010",
  40322=>"100000000",
  40323=>"011110111",
  40324=>"100000010",
  40325=>"100000111",
  40326=>"111001001",
  40327=>"110110111",
  40328=>"011011111",
  40329=>"110101110",
  40330=>"111000110",
  40331=>"110010001",
  40332=>"111101000",
  40333=>"001111010",
  40334=>"001011100",
  40335=>"100000001",
  40336=>"101111000",
  40337=>"000010000",
  40338=>"111100010",
  40339=>"111001101",
  40340=>"110010000",
  40341=>"101000101",
  40342=>"010000000",
  40343=>"001110111",
  40344=>"001111001",
  40345=>"110010111",
  40346=>"000100000",
  40347=>"010100110",
  40348=>"100000110",
  40349=>"010110000",
  40350=>"100000001",
  40351=>"101110001",
  40352=>"000100111",
  40353=>"010110010",
  40354=>"111101101",
  40355=>"000001011",
  40356=>"111000110",
  40357=>"001001010",
  40358=>"000011011",
  40359=>"100110010",
  40360=>"101100110",
  40361=>"011010111",
  40362=>"101000011",
  40363=>"101111110",
  40364=>"000001011",
  40365=>"111100110",
  40366=>"100110001",
  40367=>"011101100",
  40368=>"111111010",
  40369=>"001101110",
  40370=>"000100001",
  40371=>"011100100",
  40372=>"100111001",
  40373=>"011011110",
  40374=>"011000000",
  40375=>"101000001",
  40376=>"001001111",
  40377=>"010101011",
  40378=>"011000010",
  40379=>"000101110",
  40380=>"100100000",
  40381=>"111111001",
  40382=>"111111110",
  40383=>"101110011",
  40384=>"010011000",
  40385=>"100111100",
  40386=>"001011011",
  40387=>"000100011",
  40388=>"100000110",
  40389=>"000011100",
  40390=>"100010101",
  40391=>"000100000",
  40392=>"101000011",
  40393=>"110011110",
  40394=>"111110011",
  40395=>"101111010",
  40396=>"111111111",
  40397=>"001101111",
  40398=>"100110100",
  40399=>"010011001",
  40400=>"110000001",
  40401=>"010101001",
  40402=>"000100011",
  40403=>"111001110",
  40404=>"110011010",
  40405=>"010000001",
  40406=>"000001010",
  40407=>"011111011",
  40408=>"100000100",
  40409=>"010111011",
  40410=>"000000101",
  40411=>"101000101",
  40412=>"110111010",
  40413=>"010110011",
  40414=>"111001011",
  40415=>"001100100",
  40416=>"100001111",
  40417=>"111001101",
  40418=>"111010100",
  40419=>"110011011",
  40420=>"000111011",
  40421=>"110101000",
  40422=>"000111010",
  40423=>"000101110",
  40424=>"000101011",
  40425=>"101100111",
  40426=>"000101010",
  40427=>"000110110",
  40428=>"110011001",
  40429=>"011001100",
  40430=>"100111010",
  40431=>"011101010",
  40432=>"000110110",
  40433=>"011011011",
  40434=>"011111010",
  40435=>"100000100",
  40436=>"110011101",
  40437=>"000001101",
  40438=>"001001100",
  40439=>"000001010",
  40440=>"001111110",
  40441=>"111000101",
  40442=>"110111101",
  40443=>"100000101",
  40444=>"111111110",
  40445=>"010000000",
  40446=>"000010111",
  40447=>"101111110",
  40448=>"000101000",
  40449=>"010001110",
  40450=>"100101001",
  40451=>"010001001",
  40452=>"010011101",
  40453=>"001110001",
  40454=>"111000111",
  40455=>"001011010",
  40456=>"110110010",
  40457=>"110110000",
  40458=>"100100111",
  40459=>"110001101",
  40460=>"011000011",
  40461=>"101001011",
  40462=>"000001000",
  40463=>"000000100",
  40464=>"010001001",
  40465=>"011100101",
  40466=>"111000100",
  40467=>"101010101",
  40468=>"110111011",
  40469=>"000001001",
  40470=>"100101010",
  40471=>"000011011",
  40472=>"101110100",
  40473=>"011001011",
  40474=>"000111011",
  40475=>"010111000",
  40476=>"001110010",
  40477=>"111000101",
  40478=>"000010001",
  40479=>"110110111",
  40480=>"111100111",
  40481=>"101000101",
  40482=>"000011010",
  40483=>"000010101",
  40484=>"111110010",
  40485=>"000001110",
  40486=>"000111110",
  40487=>"111000101",
  40488=>"001010100",
  40489=>"110010011",
  40490=>"100111000",
  40491=>"101001101",
  40492=>"011111110",
  40493=>"111010110",
  40494=>"010101011",
  40495=>"010110100",
  40496=>"110010011",
  40497=>"100110001",
  40498=>"110100110",
  40499=>"100100010",
  40500=>"011100000",
  40501=>"001001111",
  40502=>"110000101",
  40503=>"010110111",
  40504=>"100111110",
  40505=>"001101100",
  40506=>"111010110",
  40507=>"010110001",
  40508=>"100100100",
  40509=>"011110010",
  40510=>"001001110",
  40511=>"110101100",
  40512=>"001011000",
  40513=>"001010000",
  40514=>"011110111",
  40515=>"000010010",
  40516=>"101110100",
  40517=>"111111100",
  40518=>"011100110",
  40519=>"000110011",
  40520=>"111111000",
  40521=>"100101100",
  40522=>"100100101",
  40523=>"001110000",
  40524=>"000101101",
  40525=>"110110101",
  40526=>"101100010",
  40527=>"100100010",
  40528=>"110110101",
  40529=>"000100101",
  40530=>"001000110",
  40531=>"100011110",
  40532=>"100001100",
  40533=>"110110000",
  40534=>"111111100",
  40535=>"111110001",
  40536=>"001011011",
  40537=>"101011101",
  40538=>"001111011",
  40539=>"001000111",
  40540=>"111011100",
  40541=>"101000011",
  40542=>"001110011",
  40543=>"000110001",
  40544=>"100010011",
  40545=>"001001100",
  40546=>"001100000",
  40547=>"000010011",
  40548=>"101110111",
  40549=>"011111110",
  40550=>"100111010",
  40551=>"001011011",
  40552=>"001100101",
  40553=>"010000101",
  40554=>"101111101",
  40555=>"000010111",
  40556=>"101100010",
  40557=>"111011011",
  40558=>"111000011",
  40559=>"101001011",
  40560=>"001110101",
  40561=>"101011001",
  40562=>"011011111",
  40563=>"000011101",
  40564=>"011001101",
  40565=>"001011110",
  40566=>"000010101",
  40567=>"000101000",
  40568=>"001011101",
  40569=>"010001010",
  40570=>"101011000",
  40571=>"000011111",
  40572=>"111000011",
  40573=>"100011100",
  40574=>"010000101",
  40575=>"100010110",
  40576=>"001011101",
  40577=>"010001110",
  40578=>"111101011",
  40579=>"111111110",
  40580=>"101101111",
  40581=>"111111011",
  40582=>"011110011",
  40583=>"111101110",
  40584=>"010111110",
  40585=>"001001111",
  40586=>"110101101",
  40587=>"011011110",
  40588=>"000000010",
  40589=>"010110100",
  40590=>"111111101",
  40591=>"001110111",
  40592=>"110010010",
  40593=>"111100110",
  40594=>"000101100",
  40595=>"110110100",
  40596=>"011000000",
  40597=>"000000101",
  40598=>"110011011",
  40599=>"010111000",
  40600=>"001111101",
  40601=>"001011010",
  40602=>"001000010",
  40603=>"101101001",
  40604=>"010001000",
  40605=>"101101100",
  40606=>"110110101",
  40607=>"101010010",
  40608=>"111111000",
  40609=>"111001011",
  40610=>"001101010",
  40611=>"110011001",
  40612=>"101011011",
  40613=>"111110010",
  40614=>"001110100",
  40615=>"101100111",
  40616=>"000001101",
  40617=>"111111111",
  40618=>"001010101",
  40619=>"000001111",
  40620=>"000011101",
  40621=>"100000010",
  40622=>"011011010",
  40623=>"001111110",
  40624=>"010100111",
  40625=>"010100001",
  40626=>"010010001",
  40627=>"001011001",
  40628=>"100100110",
  40629=>"101100010",
  40630=>"111001011",
  40631=>"101101110",
  40632=>"000100001",
  40633=>"000000000",
  40634=>"101010000",
  40635=>"101010001",
  40636=>"111011111",
  40637=>"001011000",
  40638=>"000010010",
  40639=>"111010111",
  40640=>"101001111",
  40641=>"100011000",
  40642=>"010100001",
  40643=>"100010000",
  40644=>"100110000",
  40645=>"100001101",
  40646=>"100000010",
  40647=>"111011001",
  40648=>"100100011",
  40649=>"100101001",
  40650=>"010110111",
  40651=>"001000111",
  40652=>"000111011",
  40653=>"010000001",
  40654=>"010011001",
  40655=>"111001011",
  40656=>"000000000",
  40657=>"011000111",
  40658=>"100010011",
  40659=>"110010111",
  40660=>"000011110",
  40661=>"101101111",
  40662=>"001110010",
  40663=>"101100100",
  40664=>"100011111",
  40665=>"001001000",
  40666=>"000111001",
  40667=>"000100100",
  40668=>"000000100",
  40669=>"100011111",
  40670=>"001011000",
  40671=>"100100000",
  40672=>"001010101",
  40673=>"111001011",
  40674=>"000010011",
  40675=>"100111000",
  40676=>"011000111",
  40677=>"111111101",
  40678=>"001011000",
  40679=>"000010010",
  40680=>"010110000",
  40681=>"000110010",
  40682=>"100000010",
  40683=>"100100001",
  40684=>"111111000",
  40685=>"100100110",
  40686=>"110110111",
  40687=>"100110001",
  40688=>"100001110",
  40689=>"111001010",
  40690=>"101000111",
  40691=>"101110001",
  40692=>"111100100",
  40693=>"110100101",
  40694=>"100100110",
  40695=>"001100001",
  40696=>"110001000",
  40697=>"111111111",
  40698=>"011110100",
  40699=>"110011110",
  40700=>"110001111",
  40701=>"111111110",
  40702=>"101101010",
  40703=>"001000100",
  40704=>"001011000",
  40705=>"000110000",
  40706=>"110110101",
  40707=>"011110111",
  40708=>"000000110",
  40709=>"111101101",
  40710=>"010100100",
  40711=>"110010001",
  40712=>"001101000",
  40713=>"100011001",
  40714=>"000010100",
  40715=>"011001110",
  40716=>"101110111",
  40717=>"101011111",
  40718=>"010010000",
  40719=>"010000101",
  40720=>"111101110",
  40721=>"011010000",
  40722=>"100000010",
  40723=>"000000001",
  40724=>"011110000",
  40725=>"110110110",
  40726=>"100000111",
  40727=>"011110010",
  40728=>"011101111",
  40729=>"000000111",
  40730=>"010000000",
  40731=>"000101010",
  40732=>"011111111",
  40733=>"001100101",
  40734=>"101000000",
  40735=>"011010001",
  40736=>"101001001",
  40737=>"111010010",
  40738=>"000111100",
  40739=>"101110100",
  40740=>"011000100",
  40741=>"010111100",
  40742=>"000000000",
  40743=>"001100111",
  40744=>"100001010",
  40745=>"111110111",
  40746=>"011100101",
  40747=>"010111111",
  40748=>"111001110",
  40749=>"000010010",
  40750=>"000100100",
  40751=>"001011011",
  40752=>"101000000",
  40753=>"000010101",
  40754=>"001000011",
  40755=>"101110110",
  40756=>"011111000",
  40757=>"101111101",
  40758=>"000000000",
  40759=>"010000010",
  40760=>"001101010",
  40761=>"011101100",
  40762=>"010100010",
  40763=>"110110001",
  40764=>"011100001",
  40765=>"011010101",
  40766=>"000000010",
  40767=>"101000000",
  40768=>"001100101",
  40769=>"010101101",
  40770=>"000000111",
  40771=>"110010111",
  40772=>"110011000",
  40773=>"001110111",
  40774=>"011100100",
  40775=>"100011101",
  40776=>"111110001",
  40777=>"101011101",
  40778=>"110010000",
  40779=>"100011001",
  40780=>"011000110",
  40781=>"100110111",
  40782=>"111110110",
  40783=>"110000100",
  40784=>"000011010",
  40785=>"101011010",
  40786=>"010011000",
  40787=>"000101101",
  40788=>"010111101",
  40789=>"111111111",
  40790=>"000110000",
  40791=>"001111010",
  40792=>"100011101",
  40793=>"111100100",
  40794=>"100000100",
  40795=>"001001010",
  40796=>"011001100",
  40797=>"010011010",
  40798=>"010110010",
  40799=>"000001000",
  40800=>"101100000",
  40801=>"111111101",
  40802=>"100101010",
  40803=>"010011010",
  40804=>"001101100",
  40805=>"011101100",
  40806=>"000100000",
  40807=>"110101101",
  40808=>"000111100",
  40809=>"100111110",
  40810=>"011100110",
  40811=>"011001010",
  40812=>"010100100",
  40813=>"110110011",
  40814=>"101110000",
  40815=>"010001000",
  40816=>"000011000",
  40817=>"110101001",
  40818=>"010101100",
  40819=>"101110110",
  40820=>"101001110",
  40821=>"111101111",
  40822=>"011100011",
  40823=>"110101001",
  40824=>"001111011",
  40825=>"001000100",
  40826=>"100010110",
  40827=>"101001000",
  40828=>"100110010",
  40829=>"110010000",
  40830=>"101111110",
  40831=>"001111000",
  40832=>"000001100",
  40833=>"010001000",
  40834=>"011111010",
  40835=>"100011100",
  40836=>"111011100",
  40837=>"100000001",
  40838=>"100100010",
  40839=>"010001011",
  40840=>"110100000",
  40841=>"011001000",
  40842=>"100100010",
  40843=>"001110101",
  40844=>"000000101",
  40845=>"111011110",
  40846=>"110010011",
  40847=>"110101111",
  40848=>"111110010",
  40849=>"010011101",
  40850=>"101110000",
  40851=>"010001010",
  40852=>"001101110",
  40853=>"000001101",
  40854=>"111101001",
  40855=>"011111000",
  40856=>"111101101",
  40857=>"000010010",
  40858=>"110111011",
  40859=>"011001001",
  40860=>"101110001",
  40861=>"101111101",
  40862=>"010010001",
  40863=>"101011011",
  40864=>"011100101",
  40865=>"010000001",
  40866=>"111000110",
  40867=>"111100111",
  40868=>"001001100",
  40869=>"010111110",
  40870=>"111110100",
  40871=>"110100001",
  40872=>"011101110",
  40873=>"111100001",
  40874=>"111011100",
  40875=>"100000010",
  40876=>"010011010",
  40877=>"011011001",
  40878=>"110010100",
  40879=>"110000101",
  40880=>"111111101",
  40881=>"101001001",
  40882=>"110010100",
  40883=>"110001001",
  40884=>"111100000",
  40885=>"011101110",
  40886=>"001001101",
  40887=>"001011001",
  40888=>"000010111",
  40889=>"100101111",
  40890=>"011110111",
  40891=>"011000111",
  40892=>"100010011",
  40893=>"110010011",
  40894=>"000010001",
  40895=>"010011011",
  40896=>"111110110",
  40897=>"001010111",
  40898=>"010111000",
  40899=>"111111000",
  40900=>"100110001",
  40901=>"000000001",
  40902=>"000100011",
  40903=>"001010101",
  40904=>"000010011",
  40905=>"100000101",
  40906=>"101001010",
  40907=>"001010110",
  40908=>"000000011",
  40909=>"001001110",
  40910=>"100011000",
  40911=>"010000000",
  40912=>"101100000",
  40913=>"011111111",
  40914=>"011001011",
  40915=>"100101111",
  40916=>"010011000",
  40917=>"011111101",
  40918=>"000011010",
  40919=>"101101010",
  40920=>"001000010",
  40921=>"100111001",
  40922=>"110101111",
  40923=>"000110111",
  40924=>"001110111",
  40925=>"000000001",
  40926=>"010001100",
  40927=>"010010110",
  40928=>"011101001",
  40929=>"000100101",
  40930=>"011100100",
  40931=>"000111111",
  40932=>"000010010",
  40933=>"011011000",
  40934=>"000001000",
  40935=>"110010100",
  40936=>"101001010",
  40937=>"010001100",
  40938=>"000000110",
  40939=>"100111101",
  40940=>"100111010",
  40941=>"100101011",
  40942=>"000011011",
  40943=>"001101010",
  40944=>"000001100",
  40945=>"000001110",
  40946=>"111011001",
  40947=>"111111111",
  40948=>"011000011",
  40949=>"111100001",
  40950=>"101111010",
  40951=>"000001010",
  40952=>"011011101",
  40953=>"000101110",
  40954=>"000010011",
  40955=>"001000011",
  40956=>"110111010",
  40957=>"110011100",
  40958=>"111110101",
  40959=>"001100000",
  40960=>"000001111",
  40961=>"010111000",
  40962=>"011000101",
  40963=>"001100111",
  40964=>"111000011",
  40965=>"000100110",
  40966=>"000000001",
  40967=>"101110001",
  40968=>"111011110",
  40969=>"111101110",
  40970=>"011001110",
  40971=>"001011001",
  40972=>"010000001",
  40973=>"100000000",
  40974=>"100010000",
  40975=>"110010100",
  40976=>"100001010",
  40977=>"011110010",
  40978=>"101111101",
  40979=>"111100001",
  40980=>"110011110",
  40981=>"010101001",
  40982=>"011010111",
  40983=>"101001000",
  40984=>"001000110",
  40985=>"011100100",
  40986=>"000100100",
  40987=>"010010101",
  40988=>"100000001",
  40989=>"101000000",
  40990=>"100100011",
  40991=>"100100111",
  40992=>"100010001",
  40993=>"010111101",
  40994=>"010101011",
  40995=>"000000000",
  40996=>"111100101",
  40997=>"011100101",
  40998=>"010110001",
  40999=>"111001101",
  41000=>"000101110",
  41001=>"010100100",
  41002=>"011100111",
  41003=>"000000101",
  41004=>"011110000",
  41005=>"001100000",
  41006=>"110000101",
  41007=>"001110001",
  41008=>"100000111",
  41009=>"100000111",
  41010=>"110110000",
  41011=>"111000100",
  41012=>"100001111",
  41013=>"001000010",
  41014=>"001010101",
  41015=>"110110101",
  41016=>"010011101",
  41017=>"010001100",
  41018=>"011110101",
  41019=>"000110010",
  41020=>"101110010",
  41021=>"010010110",
  41022=>"010011010",
  41023=>"000100011",
  41024=>"000000000",
  41025=>"101010111",
  41026=>"000100111",
  41027=>"000010101",
  41028=>"010110011",
  41029=>"101011110",
  41030=>"000110111",
  41031=>"010010110",
  41032=>"110000010",
  41033=>"011100111",
  41034=>"110101001",
  41035=>"111110011",
  41036=>"101000111",
  41037=>"001110001",
  41038=>"011111010",
  41039=>"110100000",
  41040=>"100001010",
  41041=>"101001110",
  41042=>"100100110",
  41043=>"100011101",
  41044=>"101011011",
  41045=>"111100000",
  41046=>"000100010",
  41047=>"100000001",
  41048=>"011101110",
  41049=>"001011100",
  41050=>"101010100",
  41051=>"111111110",
  41052=>"001100011",
  41053=>"111010000",
  41054=>"010010111",
  41055=>"111110110",
  41056=>"101111101",
  41057=>"101100001",
  41058=>"101010110",
  41059=>"001010000",
  41060=>"111101100",
  41061=>"000101110",
  41062=>"101111111",
  41063=>"100011010",
  41064=>"111111010",
  41065=>"001111011",
  41066=>"000010000",
  41067=>"100001101",
  41068=>"110111100",
  41069=>"010100000",
  41070=>"100001010",
  41071=>"000011101",
  41072=>"000101110",
  41073=>"010001101",
  41074=>"000101101",
  41075=>"101111100",
  41076=>"100110000",
  41077=>"101110011",
  41078=>"000110000",
  41079=>"001110010",
  41080=>"000011011",
  41081=>"010010010",
  41082=>"101100110",
  41083=>"000000110",
  41084=>"001110100",
  41085=>"110000100",
  41086=>"111011101",
  41087=>"111100000",
  41088=>"011100111",
  41089=>"101101101",
  41090=>"011111110",
  41091=>"000001000",
  41092=>"010111101",
  41093=>"111011010",
  41094=>"011010001",
  41095=>"010111001",
  41096=>"100101010",
  41097=>"001000000",
  41098=>"110101110",
  41099=>"111001100",
  41100=>"000000111",
  41101=>"101101011",
  41102=>"100000100",
  41103=>"111111001",
  41104=>"000101111",
  41105=>"100111001",
  41106=>"001111000",
  41107=>"111101010",
  41108=>"110110000",
  41109=>"100100000",
  41110=>"011100000",
  41111=>"000000001",
  41112=>"001100010",
  41113=>"100100000",
  41114=>"111010111",
  41115=>"001101110",
  41116=>"100000111",
  41117=>"100000110",
  41118=>"100100000",
  41119=>"010001001",
  41120=>"111110100",
  41121=>"001100110",
  41122=>"011100001",
  41123=>"111011001",
  41124=>"001111000",
  41125=>"001100110",
  41126=>"001111100",
  41127=>"110111010",
  41128=>"000000111",
  41129=>"001111111",
  41130=>"001010101",
  41131=>"111010000",
  41132=>"100101001",
  41133=>"010110110",
  41134=>"001010010",
  41135=>"010011100",
  41136=>"010100011",
  41137=>"011010101",
  41138=>"000001000",
  41139=>"010001100",
  41140=>"100111101",
  41141=>"001100111",
  41142=>"111101101",
  41143=>"101111110",
  41144=>"000000101",
  41145=>"111111001",
  41146=>"000110110",
  41147=>"111100011",
  41148=>"111011001",
  41149=>"110110010",
  41150=>"011111110",
  41151=>"101111101",
  41152=>"000001001",
  41153=>"000101101",
  41154=>"011001001",
  41155=>"111100101",
  41156=>"101011101",
  41157=>"000111110",
  41158=>"010110100",
  41159=>"000111011",
  41160=>"100100100",
  41161=>"000110010",
  41162=>"101101101",
  41163=>"000101011",
  41164=>"010100011",
  41165=>"111001100",
  41166=>"010011011",
  41167=>"111000100",
  41168=>"101111100",
  41169=>"111110010",
  41170=>"100110010",
  41171=>"011001110",
  41172=>"110100000",
  41173=>"101100001",
  41174=>"001010101",
  41175=>"101010010",
  41176=>"100101110",
  41177=>"100101111",
  41178=>"001100001",
  41179=>"111101001",
  41180=>"001101110",
  41181=>"000110100",
  41182=>"111101000",
  41183=>"011010000",
  41184=>"100011110",
  41185=>"000100111",
  41186=>"101101111",
  41187=>"001010110",
  41188=>"101001000",
  41189=>"100010011",
  41190=>"101001010",
  41191=>"011000101",
  41192=>"111011010",
  41193=>"011100101",
  41194=>"010011101",
  41195=>"000100000",
  41196=>"001101100",
  41197=>"011100000",
  41198=>"010011101",
  41199=>"111101100",
  41200=>"101101101",
  41201=>"110111001",
  41202=>"010110010",
  41203=>"001101001",
  41204=>"110101101",
  41205=>"101110000",
  41206=>"111000101",
  41207=>"101100111",
  41208=>"000000001",
  41209=>"110100111",
  41210=>"001110100",
  41211=>"100110100",
  41212=>"001000101",
  41213=>"000101101",
  41214=>"111000000",
  41215=>"100001100",
  41216=>"000100001",
  41217=>"101000001",
  41218=>"110100111",
  41219=>"100110000",
  41220=>"010010000",
  41221=>"101100111",
  41222=>"010111111",
  41223=>"101010100",
  41224=>"000111000",
  41225=>"101101000",
  41226=>"101010101",
  41227=>"011000011",
  41228=>"010010010",
  41229=>"011010010",
  41230=>"010011000",
  41231=>"110110111",
  41232=>"100000001",
  41233=>"011001011",
  41234=>"011001110",
  41235=>"100010100",
  41236=>"101100111",
  41237=>"110010000",
  41238=>"010000110",
  41239=>"100100111",
  41240=>"110111111",
  41241=>"101000011",
  41242=>"000100010",
  41243=>"100001011",
  41244=>"011101110",
  41245=>"100111111",
  41246=>"011100101",
  41247=>"111010111",
  41248=>"011101110",
  41249=>"000111001",
  41250=>"100011101",
  41251=>"101110101",
  41252=>"010101100",
  41253=>"111110111",
  41254=>"110110001",
  41255=>"010111100",
  41256=>"110000011",
  41257=>"001010001",
  41258=>"000001000",
  41259=>"000111101",
  41260=>"101111011",
  41261=>"101110101",
  41262=>"000111001",
  41263=>"100000110",
  41264=>"001001110",
  41265=>"101010011",
  41266=>"010001011",
  41267=>"011000000",
  41268=>"010000100",
  41269=>"100101010",
  41270=>"010001000",
  41271=>"011111110",
  41272=>"010100000",
  41273=>"011010111",
  41274=>"110100001",
  41275=>"100010111",
  41276=>"110110111",
  41277=>"001001010",
  41278=>"110000101",
  41279=>"000000110",
  41280=>"101001001",
  41281=>"001010110",
  41282=>"111100001",
  41283=>"010000110",
  41284=>"101100110",
  41285=>"101000110",
  41286=>"011101101",
  41287=>"001101010",
  41288=>"011000010",
  41289=>"111010111",
  41290=>"111110001",
  41291=>"010101010",
  41292=>"010111111",
  41293=>"011100111",
  41294=>"010100000",
  41295=>"111001000",
  41296=>"010011011",
  41297=>"111010100",
  41298=>"111011110",
  41299=>"100111011",
  41300=>"101110000",
  41301=>"110010011",
  41302=>"111001101",
  41303=>"000000110",
  41304=>"000000101",
  41305=>"100000100",
  41306=>"111011001",
  41307=>"101100011",
  41308=>"000111101",
  41309=>"100011111",
  41310=>"111111000",
  41311=>"000001001",
  41312=>"111111011",
  41313=>"110100111",
  41314=>"111100010",
  41315=>"111111001",
  41316=>"001100101",
  41317=>"110001000",
  41318=>"011100100",
  41319=>"000011110",
  41320=>"100011000",
  41321=>"001110011",
  41322=>"101110111",
  41323=>"011111111",
  41324=>"101000111",
  41325=>"010000010",
  41326=>"000001110",
  41327=>"010100111",
  41328=>"001010101",
  41329=>"001010101",
  41330=>"101101111",
  41331=>"000110000",
  41332=>"011110100",
  41333=>"010101111",
  41334=>"110111001",
  41335=>"101000000",
  41336=>"010010010",
  41337=>"101100000",
  41338=>"101101000",
  41339=>"000100010",
  41340=>"011000000",
  41341=>"111101111",
  41342=>"010011100",
  41343=>"001001011",
  41344=>"111100101",
  41345=>"111110111",
  41346=>"100111100",
  41347=>"011001010",
  41348=>"011000010",
  41349=>"111100001",
  41350=>"110001001",
  41351=>"100011110",
  41352=>"101100000",
  41353=>"111000000",
  41354=>"111110111",
  41355=>"111111111",
  41356=>"010001110",
  41357=>"010110100",
  41358=>"100111110",
  41359=>"001011000",
  41360=>"011001100",
  41361=>"111011111",
  41362=>"100011011",
  41363=>"101101100",
  41364=>"000000011",
  41365=>"010010101",
  41366=>"000000000",
  41367=>"110010111",
  41368=>"111110100",
  41369=>"010011010",
  41370=>"010010010",
  41371=>"101110000",
  41372=>"101100011",
  41373=>"110000100",
  41374=>"100011111",
  41375=>"011001101",
  41376=>"000000101",
  41377=>"000010000",
  41378=>"011001010",
  41379=>"001010101",
  41380=>"110000110",
  41381=>"000000010",
  41382=>"001110011",
  41383=>"010000011",
  41384=>"010011101",
  41385=>"111010011",
  41386=>"010100001",
  41387=>"000011111",
  41388=>"011001011",
  41389=>"000110010",
  41390=>"111000111",
  41391=>"101010001",
  41392=>"100111101",
  41393=>"110000001",
  41394=>"001010110",
  41395=>"000001011",
  41396=>"011001110",
  41397=>"111101001",
  41398=>"010001101",
  41399=>"001110111",
  41400=>"100100010",
  41401=>"010100000",
  41402=>"101000001",
  41403=>"101011110",
  41404=>"111000110",
  41405=>"011101000",
  41406=>"011001111",
  41407=>"101100000",
  41408=>"110001010",
  41409=>"100011110",
  41410=>"101101001",
  41411=>"010111111",
  41412=>"101101001",
  41413=>"100011000",
  41414=>"000011011",
  41415=>"110101001",
  41416=>"101100001",
  41417=>"010001001",
  41418=>"010101010",
  41419=>"110000001",
  41420=>"101101101",
  41421=>"011100010",
  41422=>"000010011",
  41423=>"111000010",
  41424=>"111001001",
  41425=>"001001101",
  41426=>"110110101",
  41427=>"001100110",
  41428=>"100111100",
  41429=>"000110010",
  41430=>"000000011",
  41431=>"100111010",
  41432=>"011010100",
  41433=>"000010111",
  41434=>"110001101",
  41435=>"000111010",
  41436=>"110101101",
  41437=>"110111001",
  41438=>"100111110",
  41439=>"110011100",
  41440=>"000100111",
  41441=>"000000010",
  41442=>"111011011",
  41443=>"000010000",
  41444=>"100100111",
  41445=>"001101110",
  41446=>"011010000",
  41447=>"010110101",
  41448=>"001010111",
  41449=>"000011011",
  41450=>"010011111",
  41451=>"000010010",
  41452=>"001101001",
  41453=>"100000000",
  41454=>"011011010",
  41455=>"000001000",
  41456=>"001100010",
  41457=>"000011110",
  41458=>"110000111",
  41459=>"000101101",
  41460=>"101001010",
  41461=>"110000011",
  41462=>"100110111",
  41463=>"011010000",
  41464=>"001101001",
  41465=>"001011111",
  41466=>"111000010",
  41467=>"000100001",
  41468=>"000000000",
  41469=>"011010110",
  41470=>"000010000",
  41471=>"111011111",
  41472=>"001101011",
  41473=>"000100100",
  41474=>"100011000",
  41475=>"110011001",
  41476=>"110111111",
  41477=>"110001101",
  41478=>"011101100",
  41479=>"011110110",
  41480=>"010100010",
  41481=>"101000111",
  41482=>"000111110",
  41483=>"110111000",
  41484=>"011101000",
  41485=>"101011010",
  41486=>"101110001",
  41487=>"111000111",
  41488=>"100100100",
  41489=>"001001010",
  41490=>"000000101",
  41491=>"000011011",
  41492=>"100100011",
  41493=>"000011110",
  41494=>"010111101",
  41495=>"110110111",
  41496=>"001101011",
  41497=>"101110001",
  41498=>"000011101",
  41499=>"010110011",
  41500=>"110111000",
  41501=>"111111111",
  41502=>"100000000",
  41503=>"000000011",
  41504=>"100010001",
  41505=>"000111011",
  41506=>"000111111",
  41507=>"100101010",
  41508=>"011111011",
  41509=>"111111101",
  41510=>"001001110",
  41511=>"001001010",
  41512=>"101111010",
  41513=>"001011100",
  41514=>"110110000",
  41515=>"100000010",
  41516=>"101010010",
  41517=>"010001000",
  41518=>"111101001",
  41519=>"001100011",
  41520=>"101100100",
  41521=>"101010010",
  41522=>"111100010",
  41523=>"100010111",
  41524=>"000100011",
  41525=>"011110100",
  41526=>"100010100",
  41527=>"011101111",
  41528=>"010101100",
  41529=>"111011000",
  41530=>"101001101",
  41531=>"010100111",
  41532=>"111101101",
  41533=>"101001100",
  41534=>"000000110",
  41535=>"100011011",
  41536=>"011100100",
  41537=>"010001101",
  41538=>"011010000",
  41539=>"111110110",
  41540=>"101000101",
  41541=>"011011100",
  41542=>"001100111",
  41543=>"000010011",
  41544=>"100110010",
  41545=>"010101001",
  41546=>"011010101",
  41547=>"011000110",
  41548=>"011010101",
  41549=>"001010100",
  41550=>"101100111",
  41551=>"111110111",
  41552=>"001100000",
  41553=>"000100001",
  41554=>"010010111",
  41555=>"100001100",
  41556=>"111101000",
  41557=>"101110110",
  41558=>"010011000",
  41559=>"011000111",
  41560=>"111000110",
  41561=>"010001101",
  41562=>"011000001",
  41563=>"000001000",
  41564=>"100101011",
  41565=>"000111001",
  41566=>"111101110",
  41567=>"111011010",
  41568=>"111111100",
  41569=>"010001000",
  41570=>"000000101",
  41571=>"100101100",
  41572=>"011011100",
  41573=>"101100110",
  41574=>"111110100",
  41575=>"101001110",
  41576=>"010001000",
  41577=>"010111000",
  41578=>"101101101",
  41579=>"000000100",
  41580=>"101011000",
  41581=>"100011011",
  41582=>"111010101",
  41583=>"000010010",
  41584=>"000101001",
  41585=>"000000011",
  41586=>"111101111",
  41587=>"100100011",
  41588=>"110010001",
  41589=>"011101111",
  41590=>"101000000",
  41591=>"000100011",
  41592=>"100001000",
  41593=>"000011101",
  41594=>"111010111",
  41595=>"000000100",
  41596=>"111011001",
  41597=>"110111001",
  41598=>"011101110",
  41599=>"010101110",
  41600=>"001011001",
  41601=>"111001010",
  41602=>"111101010",
  41603=>"110010010",
  41604=>"110010000",
  41605=>"101001101",
  41606=>"101010001",
  41607=>"001100000",
  41608=>"011000010",
  41609=>"010111011",
  41610=>"100011001",
  41611=>"110010101",
  41612=>"101000010",
  41613=>"000110000",
  41614=>"101010111",
  41615=>"010011001",
  41616=>"100001000",
  41617=>"111101010",
  41618=>"010010001",
  41619=>"000100001",
  41620=>"110111111",
  41621=>"010010111",
  41622=>"111100010",
  41623=>"001001000",
  41624=>"111000001",
  41625=>"101001001",
  41626=>"001011001",
  41627=>"011111001",
  41628=>"111101110",
  41629=>"010111011",
  41630=>"011110101",
  41631=>"010011100",
  41632=>"111011101",
  41633=>"010110011",
  41634=>"111101001",
  41635=>"010001011",
  41636=>"001011000",
  41637=>"010000110",
  41638=>"010001000",
  41639=>"010101000",
  41640=>"001110101",
  41641=>"100100100",
  41642=>"001111101",
  41643=>"011100110",
  41644=>"110101111",
  41645=>"110001110",
  41646=>"011001001",
  41647=>"011011101",
  41648=>"001010010",
  41649=>"100000111",
  41650=>"101111001",
  41651=>"000100110",
  41652=>"110001110",
  41653=>"010101100",
  41654=>"111011110",
  41655=>"001000000",
  41656=>"001001100",
  41657=>"000111001",
  41658=>"110110101",
  41659=>"001010011",
  41660=>"101100011",
  41661=>"100110110",
  41662=>"000111010",
  41663=>"010010001",
  41664=>"001001011",
  41665=>"011110100",
  41666=>"101001000",
  41667=>"101100011",
  41668=>"011000011",
  41669=>"111110010",
  41670=>"001100001",
  41671=>"010011100",
  41672=>"101000100",
  41673=>"010101010",
  41674=>"010011011",
  41675=>"101101101",
  41676=>"010100010",
  41677=>"101011010",
  41678=>"111010011",
  41679=>"111101101",
  41680=>"101000100",
  41681=>"101101100",
  41682=>"010011001",
  41683=>"101100000",
  41684=>"001011110",
  41685=>"010100101",
  41686=>"001010011",
  41687=>"001100011",
  41688=>"011011100",
  41689=>"101111101",
  41690=>"110010011",
  41691=>"011000100",
  41692=>"000001110",
  41693=>"101000000",
  41694=>"010111111",
  41695=>"110100000",
  41696=>"001010110",
  41697=>"000101101",
  41698=>"101111101",
  41699=>"001100001",
  41700=>"100010111",
  41701=>"100101010",
  41702=>"011000010",
  41703=>"001110001",
  41704=>"101011101",
  41705=>"001011000",
  41706=>"101111001",
  41707=>"100110000",
  41708=>"110100100",
  41709=>"101111010",
  41710=>"001001011",
  41711=>"111111011",
  41712=>"110000110",
  41713=>"101010010",
  41714=>"110000001",
  41715=>"101010101",
  41716=>"001110000",
  41717=>"100110011",
  41718=>"001001111",
  41719=>"001110111",
  41720=>"100010110",
  41721=>"111000101",
  41722=>"000100101",
  41723=>"111110111",
  41724=>"101011101",
  41725=>"111011010",
  41726=>"010010011",
  41727=>"001000111",
  41728=>"110101011",
  41729=>"011101010",
  41730=>"011000010",
  41731=>"011111100",
  41732=>"111001011",
  41733=>"111000000",
  41734=>"010011100",
  41735=>"111100110",
  41736=>"010001110",
  41737=>"101110110",
  41738=>"110100001",
  41739=>"000101100",
  41740=>"100001110",
  41741=>"000011100",
  41742=>"111000101",
  41743=>"101001100",
  41744=>"011101101",
  41745=>"001111011",
  41746=>"100110011",
  41747=>"011011101",
  41748=>"110010001",
  41749=>"000011000",
  41750=>"110011100",
  41751=>"000001001",
  41752=>"000000010",
  41753=>"011001110",
  41754=>"101111001",
  41755=>"000101111",
  41756=>"001100011",
  41757=>"101010010",
  41758=>"110110011",
  41759=>"111111000",
  41760=>"011010101",
  41761=>"001000000",
  41762=>"000011100",
  41763=>"101110100",
  41764=>"100101010",
  41765=>"110000110",
  41766=>"001100101",
  41767=>"010010010",
  41768=>"011011011",
  41769=>"100101001",
  41770=>"011111001",
  41771=>"010110100",
  41772=>"110010011",
  41773=>"011111111",
  41774=>"111010110",
  41775=>"100101100",
  41776=>"000001100",
  41777=>"100011101",
  41778=>"100010111",
  41779=>"110000001",
  41780=>"101111111",
  41781=>"010010110",
  41782=>"100111010",
  41783=>"110000010",
  41784=>"100111111",
  41785=>"010010000",
  41786=>"110100001",
  41787=>"100001001",
  41788=>"101010111",
  41789=>"101100010",
  41790=>"101100001",
  41791=>"001111110",
  41792=>"101001000",
  41793=>"111110000",
  41794=>"000100100",
  41795=>"111111100",
  41796=>"110000111",
  41797=>"000011000",
  41798=>"000110010",
  41799=>"011010111",
  41800=>"110111100",
  41801=>"101111111",
  41802=>"011111000",
  41803=>"111110101",
  41804=>"100100010",
  41805=>"010100010",
  41806=>"000010000",
  41807=>"101011110",
  41808=>"100010101",
  41809=>"100110010",
  41810=>"011111111",
  41811=>"000101000",
  41812=>"101010011",
  41813=>"111101010",
  41814=>"000000000",
  41815=>"001111010",
  41816=>"100011011",
  41817=>"101111110",
  41818=>"100101001",
  41819=>"101101111",
  41820=>"111111000",
  41821=>"101011111",
  41822=>"000001010",
  41823=>"011000100",
  41824=>"111110110",
  41825=>"111110010",
  41826=>"000001010",
  41827=>"101010111",
  41828=>"011000110",
  41829=>"000001110",
  41830=>"110011101",
  41831=>"001000000",
  41832=>"000000000",
  41833=>"100011100",
  41834=>"010001000",
  41835=>"000110110",
  41836=>"010011110",
  41837=>"000010100",
  41838=>"111110001",
  41839=>"101100010",
  41840=>"110101111",
  41841=>"110001100",
  41842=>"101101000",
  41843=>"100011011",
  41844=>"000111111",
  41845=>"010011001",
  41846=>"011000101",
  41847=>"001010110",
  41848=>"010010100",
  41849=>"000111101",
  41850=>"110100110",
  41851=>"101110100",
  41852=>"010111101",
  41853=>"101101100",
  41854=>"001000000",
  41855=>"010111001",
  41856=>"000111100",
  41857=>"001111011",
  41858=>"001011100",
  41859=>"110001101",
  41860=>"000111000",
  41861=>"110100111",
  41862=>"010101010",
  41863=>"011000001",
  41864=>"101000000",
  41865=>"010001010",
  41866=>"100110000",
  41867=>"000111110",
  41868=>"010100000",
  41869=>"101001000",
  41870=>"011110011",
  41871=>"010000110",
  41872=>"100100100",
  41873=>"111001100",
  41874=>"101111101",
  41875=>"101111011",
  41876=>"010100110",
  41877=>"000011000",
  41878=>"001111011",
  41879=>"011100001",
  41880=>"010001111",
  41881=>"001101011",
  41882=>"100100000",
  41883=>"000010100",
  41884=>"010100110",
  41885=>"010100001",
  41886=>"001010100",
  41887=>"100000000",
  41888=>"011000100",
  41889=>"000111111",
  41890=>"001001110",
  41891=>"101000101",
  41892=>"011010111",
  41893=>"000111100",
  41894=>"010110101",
  41895=>"011000010",
  41896=>"000011101",
  41897=>"010100100",
  41898=>"000101011",
  41899=>"111010111",
  41900=>"000110010",
  41901=>"111010011",
  41902=>"110001011",
  41903=>"001011001",
  41904=>"111111100",
  41905=>"101011000",
  41906=>"010100000",
  41907=>"001010110",
  41908=>"000100010",
  41909=>"001000010",
  41910=>"100001101",
  41911=>"000001100",
  41912=>"101011110",
  41913=>"100000100",
  41914=>"110001100",
  41915=>"000001000",
  41916=>"111111101",
  41917=>"110100110",
  41918=>"001011101",
  41919=>"110110100",
  41920=>"010001101",
  41921=>"110010110",
  41922=>"100101101",
  41923=>"110110000",
  41924=>"001111101",
  41925=>"011111100",
  41926=>"110010001",
  41927=>"101110101",
  41928=>"000101100",
  41929=>"100100101",
  41930=>"110101100",
  41931=>"010000010",
  41932=>"001100010",
  41933=>"000001000",
  41934=>"001000100",
  41935=>"100001100",
  41936=>"101010011",
  41937=>"011100000",
  41938=>"100000101",
  41939=>"101100101",
  41940=>"111110101",
  41941=>"011110110",
  41942=>"001111110",
  41943=>"100101011",
  41944=>"000011110",
  41945=>"011010000",
  41946=>"101011011",
  41947=>"011010010",
  41948=>"101000111",
  41949=>"010010110",
  41950=>"101111111",
  41951=>"010001110",
  41952=>"100011111",
  41953=>"011001010",
  41954=>"011011000",
  41955=>"011011111",
  41956=>"010000111",
  41957=>"010100101",
  41958=>"001101111",
  41959=>"000001000",
  41960=>"001001010",
  41961=>"010010000",
  41962=>"011111010",
  41963=>"110000011",
  41964=>"111000011",
  41965=>"101101101",
  41966=>"100001000",
  41967=>"000100001",
  41968=>"000010010",
  41969=>"111001110",
  41970=>"010100001",
  41971=>"101010111",
  41972=>"001110001",
  41973=>"010011100",
  41974=>"000000000",
  41975=>"000000110",
  41976=>"001111110",
  41977=>"110101100",
  41978=>"000010111",
  41979=>"011010011",
  41980=>"101100101",
  41981=>"011000110",
  41982=>"000010000",
  41983=>"101000000",
  41984=>"000010001",
  41985=>"001010010",
  41986=>"100111101",
  41987=>"101110010",
  41988=>"111000111",
  41989=>"011010101",
  41990=>"010000100",
  41991=>"000101000",
  41992=>"001001000",
  41993=>"001001001",
  41994=>"100001001",
  41995=>"000110101",
  41996=>"000000100",
  41997=>"111110111",
  41998=>"001010101",
  41999=>"101001110",
  42000=>"111000110",
  42001=>"100000000",
  42002=>"010011110",
  42003=>"100000001",
  42004=>"101100010",
  42005=>"100100010",
  42006=>"010110001",
  42007=>"000101101",
  42008=>"001100011",
  42009=>"100000011",
  42010=>"101001101",
  42011=>"010011001",
  42012=>"001001100",
  42013=>"110110101",
  42014=>"110001000",
  42015=>"001111010",
  42016=>"101111000",
  42017=>"001010010",
  42018=>"101001101",
  42019=>"110100000",
  42020=>"101001100",
  42021=>"010100011",
  42022=>"101111111",
  42023=>"101001110",
  42024=>"101000011",
  42025=>"110111001",
  42026=>"110110000",
  42027=>"000100000",
  42028=>"000001001",
  42029=>"101000111",
  42030=>"100011000",
  42031=>"111000101",
  42032=>"011100010",
  42033=>"100001110",
  42034=>"101010000",
  42035=>"011010111",
  42036=>"011100010",
  42037=>"111100000",
  42038=>"100001111",
  42039=>"111010100",
  42040=>"101001000",
  42041=>"011001000",
  42042=>"100101101",
  42043=>"101111110",
  42044=>"100000110",
  42045=>"011011001",
  42046=>"010000100",
  42047=>"100110000",
  42048=>"011100010",
  42049=>"010000001",
  42050=>"100110110",
  42051=>"110000011",
  42052=>"100000110",
  42053=>"001011001",
  42054=>"101001111",
  42055=>"010011010",
  42056=>"011110001",
  42057=>"010000111",
  42058=>"000111010",
  42059=>"001000010",
  42060=>"001000000",
  42061=>"100000000",
  42062=>"001001010",
  42063=>"101010111",
  42064=>"000110111",
  42065=>"001001010",
  42066=>"110011010",
  42067=>"011101111",
  42068=>"001111010",
  42069=>"111111010",
  42070=>"101101111",
  42071=>"101111110",
  42072=>"110111110",
  42073=>"111111001",
  42074=>"111000010",
  42075=>"010000010",
  42076=>"111110111",
  42077=>"110111010",
  42078=>"100011010",
  42079=>"101001100",
  42080=>"001001010",
  42081=>"011001100",
  42082=>"110111110",
  42083=>"101100100",
  42084=>"010000011",
  42085=>"000110111",
  42086=>"001011001",
  42087=>"100110010",
  42088=>"000001000",
  42089=>"010100000",
  42090=>"011001100",
  42091=>"010010101",
  42092=>"001101101",
  42093=>"011101110",
  42094=>"011110100",
  42095=>"010101110",
  42096=>"011000101",
  42097=>"101110111",
  42098=>"010010110",
  42099=>"010011110",
  42100=>"011001100",
  42101=>"000001000",
  42102=>"001000110",
  42103=>"111101010",
  42104=>"000111111",
  42105=>"010100111",
  42106=>"101010001",
  42107=>"110101110",
  42108=>"000101000",
  42109=>"110011110",
  42110=>"010000110",
  42111=>"100101100",
  42112=>"100110001",
  42113=>"001111101",
  42114=>"000111101",
  42115=>"001000100",
  42116=>"111111100",
  42117=>"100000011",
  42118=>"100111110",
  42119=>"111001101",
  42120=>"111101011",
  42121=>"000011110",
  42122=>"110011111",
  42123=>"011011000",
  42124=>"111001100",
  42125=>"100000001",
  42126=>"111111100",
  42127=>"111100010",
  42128=>"001111111",
  42129=>"000001011",
  42130=>"110000101",
  42131=>"111100001",
  42132=>"001001010",
  42133=>"010111111",
  42134=>"001111100",
  42135=>"110100101",
  42136=>"110011000",
  42137=>"000110010",
  42138=>"011001101",
  42139=>"010101010",
  42140=>"100010010",
  42141=>"100100001",
  42142=>"001001001",
  42143=>"001000000",
  42144=>"011010000",
  42145=>"110101100",
  42146=>"011111101",
  42147=>"110110101",
  42148=>"111000001",
  42149=>"111110010",
  42150=>"110100010",
  42151=>"000001110",
  42152=>"011110110",
  42153=>"010011001",
  42154=>"101110011",
  42155=>"100001101",
  42156=>"001001010",
  42157=>"100110010",
  42158=>"111111000",
  42159=>"111111001",
  42160=>"010111000",
  42161=>"000100101",
  42162=>"001101010",
  42163=>"000001101",
  42164=>"010011100",
  42165=>"110100010",
  42166=>"001101110",
  42167=>"101101101",
  42168=>"101101111",
  42169=>"101100100",
  42170=>"101000010",
  42171=>"011001001",
  42172=>"001101000",
  42173=>"011110111",
  42174=>"010110001",
  42175=>"000000011",
  42176=>"011101010",
  42177=>"001111010",
  42178=>"011001000",
  42179=>"110000110",
  42180=>"010000110",
  42181=>"011101101",
  42182=>"100111011",
  42183=>"011110010",
  42184=>"111011011",
  42185=>"110110110",
  42186=>"110111111",
  42187=>"001000000",
  42188=>"000001000",
  42189=>"000100110",
  42190=>"011111101",
  42191=>"010100011",
  42192=>"110000110",
  42193=>"100101111",
  42194=>"101010111",
  42195=>"100110100",
  42196=>"010111111",
  42197=>"101011001",
  42198=>"101000110",
  42199=>"010000111",
  42200=>"111111001",
  42201=>"001110000",
  42202=>"110101010",
  42203=>"101011101",
  42204=>"111110111",
  42205=>"110100000",
  42206=>"001001011",
  42207=>"010111100",
  42208=>"111101100",
  42209=>"100011100",
  42210=>"100100101",
  42211=>"111111111",
  42212=>"110111110",
  42213=>"010111000",
  42214=>"000100100",
  42215=>"000001101",
  42216=>"010110001",
  42217=>"010010100",
  42218=>"001110010",
  42219=>"001111111",
  42220=>"011111100",
  42221=>"010001000",
  42222=>"000101011",
  42223=>"110110111",
  42224=>"000001110",
  42225=>"010001011",
  42226=>"001111010",
  42227=>"011110010",
  42228=>"110101001",
  42229=>"111011010",
  42230=>"110011010",
  42231=>"111111100",
  42232=>"101011111",
  42233=>"100001001",
  42234=>"100000110",
  42235=>"001001101",
  42236=>"000101101",
  42237=>"100101001",
  42238=>"101011110",
  42239=>"101110010",
  42240=>"110000000",
  42241=>"011111011",
  42242=>"011011101",
  42243=>"110001010",
  42244=>"100000000",
  42245=>"000011111",
  42246=>"110011000",
  42247=>"000010111",
  42248=>"000011010",
  42249=>"100111101",
  42250=>"101101111",
  42251=>"101001000",
  42252=>"110100000",
  42253=>"000111010",
  42254=>"001110000",
  42255=>"011110111",
  42256=>"011011111",
  42257=>"000011111",
  42258=>"111000110",
  42259=>"001111011",
  42260=>"000101000",
  42261=>"001101101",
  42262=>"101101100",
  42263=>"110010111",
  42264=>"011111111",
  42265=>"110100011",
  42266=>"101110100",
  42267=>"111001001",
  42268=>"111110100",
  42269=>"101100001",
  42270=>"101111111",
  42271=>"111001100",
  42272=>"010110000",
  42273=>"010000000",
  42274=>"111110111",
  42275=>"011111001",
  42276=>"110000000",
  42277=>"111111010",
  42278=>"011101110",
  42279=>"101011001",
  42280=>"000111000",
  42281=>"001010011",
  42282=>"100011110",
  42283=>"011010011",
  42284=>"111010010",
  42285=>"001100001",
  42286=>"101000100",
  42287=>"111110011",
  42288=>"001000010",
  42289=>"001010100",
  42290=>"011001010",
  42291=>"101100010",
  42292=>"000110110",
  42293=>"000011000",
  42294=>"100100110",
  42295=>"100001011",
  42296=>"000000110",
  42297=>"010111010",
  42298=>"001101100",
  42299=>"011000011",
  42300=>"000111111",
  42301=>"100111111",
  42302=>"110001100",
  42303=>"010100111",
  42304=>"000001110",
  42305=>"011000101",
  42306=>"110011001",
  42307=>"001010000",
  42308=>"110101010",
  42309=>"111000101",
  42310=>"010010001",
  42311=>"101001010",
  42312=>"011011001",
  42313=>"101011001",
  42314=>"111110111",
  42315=>"000000001",
  42316=>"110101001",
  42317=>"111101100",
  42318=>"011111001",
  42319=>"100101110",
  42320=>"001001010",
  42321=>"100010100",
  42322=>"110101110",
  42323=>"100110010",
  42324=>"101100000",
  42325=>"001100111",
  42326=>"100101111",
  42327=>"111000110",
  42328=>"011000010",
  42329=>"110101100",
  42330=>"000001100",
  42331=>"000100000",
  42332=>"100001010",
  42333=>"000001001",
  42334=>"001001010",
  42335=>"100101101",
  42336=>"101110000",
  42337=>"100000011",
  42338=>"001110010",
  42339=>"110101111",
  42340=>"001110100",
  42341=>"010000110",
  42342=>"010011110",
  42343=>"100010001",
  42344=>"000100110",
  42345=>"110111111",
  42346=>"110101101",
  42347=>"010010000",
  42348=>"000101100",
  42349=>"111011111",
  42350=>"000000000",
  42351=>"010100111",
  42352=>"001011000",
  42353=>"111010111",
  42354=>"001001111",
  42355=>"010011101",
  42356=>"111111001",
  42357=>"111001011",
  42358=>"101010110",
  42359=>"110111100",
  42360=>"011000101",
  42361=>"110011000",
  42362=>"101111000",
  42363=>"010101001",
  42364=>"110100011",
  42365=>"101100001",
  42366=>"010010100",
  42367=>"111001001",
  42368=>"001000100",
  42369=>"110111001",
  42370=>"011100000",
  42371=>"000000100",
  42372=>"100011011",
  42373=>"101111001",
  42374=>"111110000",
  42375=>"100101000",
  42376=>"100000011",
  42377=>"110000100",
  42378=>"011011001",
  42379=>"011110001",
  42380=>"001011010",
  42381=>"111010001",
  42382=>"101111111",
  42383=>"110100010",
  42384=>"110111001",
  42385=>"000001011",
  42386=>"000100111",
  42387=>"100000010",
  42388=>"000011001",
  42389=>"101011000",
  42390=>"100000000",
  42391=>"100111011",
  42392=>"010001110",
  42393=>"111101100",
  42394=>"000011010",
  42395=>"100000101",
  42396=>"100111111",
  42397=>"111110110",
  42398=>"110010111",
  42399=>"110000100",
  42400=>"001011011",
  42401=>"001100000",
  42402=>"110001010",
  42403=>"100011110",
  42404=>"110011100",
  42405=>"101001110",
  42406=>"110111001",
  42407=>"011010111",
  42408=>"010111001",
  42409=>"011000000",
  42410=>"000110001",
  42411=>"011000100",
  42412=>"010011100",
  42413=>"001000101",
  42414=>"101111000",
  42415=>"111000001",
  42416=>"011110111",
  42417=>"100101110",
  42418=>"000101000",
  42419=>"111110101",
  42420=>"001100010",
  42421=>"000110100",
  42422=>"100111111",
  42423=>"001001011",
  42424=>"001001001",
  42425=>"100011111",
  42426=>"101011011",
  42427=>"110101001",
  42428=>"101011101",
  42429=>"010100001",
  42430=>"111111110",
  42431=>"101011111",
  42432=>"100110111",
  42433=>"010010100",
  42434=>"110100010",
  42435=>"010101010",
  42436=>"000110111",
  42437=>"110001100",
  42438=>"011110101",
  42439=>"000101101",
  42440=>"101100111",
  42441=>"101000011",
  42442=>"010000011",
  42443=>"110110010",
  42444=>"100000101",
  42445=>"000010000",
  42446=>"001001110",
  42447=>"100011101",
  42448=>"101001101",
  42449=>"110011001",
  42450=>"111001011",
  42451=>"111111010",
  42452=>"011000000",
  42453=>"111100001",
  42454=>"111110010",
  42455=>"000000101",
  42456=>"110001001",
  42457=>"100100010",
  42458=>"000100100",
  42459=>"001010000",
  42460=>"011000110",
  42461=>"010100111",
  42462=>"010010000",
  42463=>"001110110",
  42464=>"110010000",
  42465=>"101000010",
  42466=>"110101001",
  42467=>"010101001",
  42468=>"010100010",
  42469=>"000011000",
  42470=>"010101000",
  42471=>"001101100",
  42472=>"011100111",
  42473=>"110100110",
  42474=>"110010111",
  42475=>"110110110",
  42476=>"000010111",
  42477=>"010000110",
  42478=>"001010000",
  42479=>"011111001",
  42480=>"000010010",
  42481=>"101100110",
  42482=>"010001111",
  42483=>"111000100",
  42484=>"010000100",
  42485=>"010000001",
  42486=>"000010010",
  42487=>"011010011",
  42488=>"111111010",
  42489=>"100000110",
  42490=>"011111010",
  42491=>"001010010",
  42492=>"011011000",
  42493=>"000000011",
  42494=>"111101001",
  42495=>"000110111",
  42496=>"100000000",
  42497=>"001010101",
  42498=>"111000000",
  42499=>"101011000",
  42500=>"100101101",
  42501=>"000111100",
  42502=>"001010000",
  42503=>"010001101",
  42504=>"010001101",
  42505=>"111001111",
  42506=>"010011100",
  42507=>"010010010",
  42508=>"001001101",
  42509=>"101100000",
  42510=>"101110111",
  42511=>"001000111",
  42512=>"111111010",
  42513=>"100011100",
  42514=>"100111110",
  42515=>"010110011",
  42516=>"011001110",
  42517=>"101011111",
  42518=>"101101011",
  42519=>"010000101",
  42520=>"010110110",
  42521=>"001011110",
  42522=>"011001101",
  42523=>"001111110",
  42524=>"001010110",
  42525=>"101111100",
  42526=>"101001011",
  42527=>"011010011",
  42528=>"011100000",
  42529=>"010100111",
  42530=>"101100100",
  42531=>"111011000",
  42532=>"101011001",
  42533=>"101011111",
  42534=>"101100110",
  42535=>"000110011",
  42536=>"101101011",
  42537=>"101001001",
  42538=>"110001001",
  42539=>"111001010",
  42540=>"001111001",
  42541=>"001001110",
  42542=>"100010100",
  42543=>"000010000",
  42544=>"101111101",
  42545=>"111110011",
  42546=>"000111000",
  42547=>"101000001",
  42548=>"111001010",
  42549=>"111110101",
  42550=>"101000011",
  42551=>"011111100",
  42552=>"010100111",
  42553=>"011010001",
  42554=>"101001000",
  42555=>"001010101",
  42556=>"110010010",
  42557=>"101111100",
  42558=>"111001111",
  42559=>"001011000",
  42560=>"111010111",
  42561=>"100011111",
  42562=>"000000100",
  42563=>"010110111",
  42564=>"111101101",
  42565=>"001010010",
  42566=>"101110011",
  42567=>"001110000",
  42568=>"011111011",
  42569=>"100101011",
  42570=>"101001100",
  42571=>"110011101",
  42572=>"111000000",
  42573=>"100000011",
  42574=>"100101000",
  42575=>"001011101",
  42576=>"011111110",
  42577=>"011000001",
  42578=>"110011011",
  42579=>"111010001",
  42580=>"110100101",
  42581=>"010101001",
  42582=>"100000101",
  42583=>"010010010",
  42584=>"101001001",
  42585=>"011101011",
  42586=>"010101001",
  42587=>"010111110",
  42588=>"000000101",
  42589=>"101100000",
  42590=>"001101110",
  42591=>"010000111",
  42592=>"011111100",
  42593=>"111001100",
  42594=>"111110101",
  42595=>"000100001",
  42596=>"011000111",
  42597=>"101111010",
  42598=>"111011101",
  42599=>"110001000",
  42600=>"111010000",
  42601=>"110000010",
  42602=>"100110100",
  42603=>"001010100",
  42604=>"101000011",
  42605=>"110001101",
  42606=>"111000001",
  42607=>"000001100",
  42608=>"011010111",
  42609=>"110001011",
  42610=>"010001001",
  42611=>"000010111",
  42612=>"011000011",
  42613=>"011000100",
  42614=>"011010000",
  42615=>"000001110",
  42616=>"000101000",
  42617=>"010100100",
  42618=>"000010010",
  42619=>"010000101",
  42620=>"111101101",
  42621=>"011000001",
  42622=>"011111000",
  42623=>"001110100",
  42624=>"000100000",
  42625=>"101111111",
  42626=>"111000001",
  42627=>"011110010",
  42628=>"100111110",
  42629=>"000011000",
  42630=>"110000000",
  42631=>"100111001",
  42632=>"100100110",
  42633=>"000100000",
  42634=>"011001101",
  42635=>"100101111",
  42636=>"001111101",
  42637=>"111010100",
  42638=>"101001110",
  42639=>"001111000",
  42640=>"010011101",
  42641=>"111010010",
  42642=>"111010111",
  42643=>"101011011",
  42644=>"001101100",
  42645=>"110101000",
  42646=>"001011000",
  42647=>"000001001",
  42648=>"100011010",
  42649=>"101010101",
  42650=>"110000000",
  42651=>"001101011",
  42652=>"111001001",
  42653=>"010001011",
  42654=>"101000111",
  42655=>"010011000",
  42656=>"111110101",
  42657=>"000000000",
  42658=>"110010011",
  42659=>"110111101",
  42660=>"001100000",
  42661=>"001011010",
  42662=>"101111101",
  42663=>"100010110",
  42664=>"111010101",
  42665=>"111110100",
  42666=>"001000001",
  42667=>"000101011",
  42668=>"111001111",
  42669=>"000010101",
  42670=>"000100001",
  42671=>"000101111",
  42672=>"110111011",
  42673=>"111111110",
  42674=>"110011110",
  42675=>"101111100",
  42676=>"100001111",
  42677=>"100100010",
  42678=>"111101111",
  42679=>"011100101",
  42680=>"101000100",
  42681=>"100001100",
  42682=>"101111001",
  42683=>"100100100",
  42684=>"100000111",
  42685=>"001010001",
  42686=>"000100011",
  42687=>"000101010",
  42688=>"101011101",
  42689=>"100101111",
  42690=>"000100001",
  42691=>"110011100",
  42692=>"110110101",
  42693=>"000011000",
  42694=>"010111001",
  42695=>"111111001",
  42696=>"011010100",
  42697=>"101101110",
  42698=>"010110000",
  42699=>"100000001",
  42700=>"001111000",
  42701=>"111001110",
  42702=>"001011101",
  42703=>"001010100",
  42704=>"100110100",
  42705=>"000110110",
  42706=>"001101111",
  42707=>"111000001",
  42708=>"110001001",
  42709=>"110001010",
  42710=>"101000001",
  42711=>"011011011",
  42712=>"000100000",
  42713=>"111001011",
  42714=>"101000011",
  42715=>"111101101",
  42716=>"101101100",
  42717=>"011000100",
  42718=>"000000110",
  42719=>"000000001",
  42720=>"111000100",
  42721=>"000000100",
  42722=>"110000001",
  42723=>"110110010",
  42724=>"000100000",
  42725=>"011001001",
  42726=>"110111011",
  42727=>"110001010",
  42728=>"010001100",
  42729=>"101110101",
  42730=>"111000011",
  42731=>"111000001",
  42732=>"000010100",
  42733=>"001010111",
  42734=>"100001000",
  42735=>"001101011",
  42736=>"011010111",
  42737=>"011101111",
  42738=>"111000101",
  42739=>"100001010",
  42740=>"000011100",
  42741=>"100110000",
  42742=>"011000000",
  42743=>"110000101",
  42744=>"000000010",
  42745=>"100110010",
  42746=>"100001101",
  42747=>"100001101",
  42748=>"110011000",
  42749=>"110101011",
  42750=>"000000011",
  42751=>"111111111",
  42752=>"000111110",
  42753=>"001100101",
  42754=>"000001011",
  42755=>"000110100",
  42756=>"101100000",
  42757=>"000110001",
  42758=>"011110111",
  42759=>"100100110",
  42760=>"101100000",
  42761=>"011010101",
  42762=>"110001001",
  42763=>"111011010",
  42764=>"111000011",
  42765=>"010011100",
  42766=>"111010000",
  42767=>"111000110",
  42768=>"111100111",
  42769=>"101011111",
  42770=>"010011010",
  42771=>"110000100",
  42772=>"101010010",
  42773=>"001101111",
  42774=>"111100111",
  42775=>"101011101",
  42776=>"001101001",
  42777=>"011000011",
  42778=>"100001010",
  42779=>"101011100",
  42780=>"001001011",
  42781=>"011110011",
  42782=>"110111000",
  42783=>"011111011",
  42784=>"110000001",
  42785=>"101100010",
  42786=>"100100001",
  42787=>"011100011",
  42788=>"101101011",
  42789=>"001101100",
  42790=>"011110010",
  42791=>"010100010",
  42792=>"110011100",
  42793=>"001100101",
  42794=>"100100111",
  42795=>"011011000",
  42796=>"011000001",
  42797=>"001000000",
  42798=>"000111011",
  42799=>"101001110",
  42800=>"101110100",
  42801=>"101011100",
  42802=>"101010001",
  42803=>"000000100",
  42804=>"110010100",
  42805=>"110000000",
  42806=>"100111010",
  42807=>"111100000",
  42808=>"100111101",
  42809=>"000011110",
  42810=>"100000110",
  42811=>"001110111",
  42812=>"100011100",
  42813=>"000011101",
  42814=>"111101110",
  42815=>"111101100",
  42816=>"110101011",
  42817=>"101011111",
  42818=>"101011011",
  42819=>"111111110",
  42820=>"011101110",
  42821=>"011000010",
  42822=>"111101100",
  42823=>"000111011",
  42824=>"010110000",
  42825=>"100101111",
  42826=>"000111100",
  42827=>"100011100",
  42828=>"011100000",
  42829=>"101011111",
  42830=>"111000000",
  42831=>"010111000",
  42832=>"101100011",
  42833=>"010101110",
  42834=>"001001000",
  42835=>"011100111",
  42836=>"011000010",
  42837=>"011010010",
  42838=>"001101101",
  42839=>"011101011",
  42840=>"001100010",
  42841=>"111010001",
  42842=>"001100111",
  42843=>"111001111",
  42844=>"011010000",
  42845=>"000100101",
  42846=>"010000101",
  42847=>"101101001",
  42848=>"101111110",
  42849=>"001101101",
  42850=>"000111011",
  42851=>"010101100",
  42852=>"101001110",
  42853=>"010000010",
  42854=>"000100101",
  42855=>"000110101",
  42856=>"011000101",
  42857=>"001100100",
  42858=>"111100000",
  42859=>"110111100",
  42860=>"100101101",
  42861=>"101101111",
  42862=>"011000000",
  42863=>"001001100",
  42864=>"110110011",
  42865=>"010101000",
  42866=>"000011000",
  42867=>"110101001",
  42868=>"101001001",
  42869=>"011100011",
  42870=>"110111010",
  42871=>"110111001",
  42872=>"100101001",
  42873=>"100000000",
  42874=>"001001111",
  42875=>"001000111",
  42876=>"000111011",
  42877=>"100001111",
  42878=>"111010100",
  42879=>"000010010",
  42880=>"110010010",
  42881=>"000011001",
  42882=>"001100101",
  42883=>"100101001",
  42884=>"100101101",
  42885=>"100010000",
  42886=>"000111011",
  42887=>"100000100",
  42888=>"111000011",
  42889=>"110110110",
  42890=>"011110010",
  42891=>"001010101",
  42892=>"011100110",
  42893=>"000000001",
  42894=>"000101101",
  42895=>"101101000",
  42896=>"000100000",
  42897=>"001110000",
  42898=>"001101101",
  42899=>"010100110",
  42900=>"010010010",
  42901=>"100001110",
  42902=>"011011001",
  42903=>"111101101",
  42904=>"101111000",
  42905=>"010001111",
  42906=>"000111000",
  42907=>"111101001",
  42908=>"001111111",
  42909=>"111101110",
  42910=>"110010101",
  42911=>"010001011",
  42912=>"011001110",
  42913=>"111101000",
  42914=>"111011101",
  42915=>"101000000",
  42916=>"000111111",
  42917=>"110000011",
  42918=>"100000100",
  42919=>"000010100",
  42920=>"011010011",
  42921=>"011110100",
  42922=>"101000010",
  42923=>"101110010",
  42924=>"000010111",
  42925=>"101011100",
  42926=>"101100111",
  42927=>"111001000",
  42928=>"010010110",
  42929=>"100000101",
  42930=>"000100000",
  42931=>"001111010",
  42932=>"011011011",
  42933=>"011110110",
  42934=>"000011010",
  42935=>"111110100",
  42936=>"010011001",
  42937=>"001100001",
  42938=>"110110011",
  42939=>"100111011",
  42940=>"011000111",
  42941=>"100000111",
  42942=>"101111110",
  42943=>"111011011",
  42944=>"000101011",
  42945=>"000000100",
  42946=>"001101001",
  42947=>"110001100",
  42948=>"011111011",
  42949=>"101011110",
  42950=>"101010011",
  42951=>"010011010",
  42952=>"000001101",
  42953=>"101110011",
  42954=>"101010110",
  42955=>"001101001",
  42956=>"011000101",
  42957=>"101100111",
  42958=>"100011100",
  42959=>"001000001",
  42960=>"001000111",
  42961=>"100100001",
  42962=>"110100001",
  42963=>"000000000",
  42964=>"111011101",
  42965=>"100111110",
  42966=>"001111110",
  42967=>"010111010",
  42968=>"100111111",
  42969=>"100101000",
  42970=>"001100001",
  42971=>"111010111",
  42972=>"100010111",
  42973=>"100110001",
  42974=>"000100011",
  42975=>"000001000",
  42976=>"100100101",
  42977=>"000101001",
  42978=>"000001100",
  42979=>"010100101",
  42980=>"001001001",
  42981=>"001100001",
  42982=>"001011100",
  42983=>"000101101",
  42984=>"111110010",
  42985=>"001110001",
  42986=>"011001010",
  42987=>"110111000",
  42988=>"110011010",
  42989=>"000101101",
  42990=>"111111001",
  42991=>"111011001",
  42992=>"000010110",
  42993=>"001000010",
  42994=>"101010010",
  42995=>"111100001",
  42996=>"011100000",
  42997=>"111011101",
  42998=>"010100000",
  42999=>"000011111",
  43000=>"100100100",
  43001=>"100001111",
  43002=>"000001010",
  43003=>"011100000",
  43004=>"111100011",
  43005=>"011101000",
  43006=>"010010011",
  43007=>"011111001",
  43008=>"101000000",
  43009=>"111011011",
  43010=>"100000011",
  43011=>"011010111",
  43012=>"100111100",
  43013=>"010111001",
  43014=>"000010001",
  43015=>"101111101",
  43016=>"110100001",
  43017=>"110111101",
  43018=>"011111100",
  43019=>"101010111",
  43020=>"111100000",
  43021=>"101000111",
  43022=>"100010101",
  43023=>"001110000",
  43024=>"110101010",
  43025=>"111000101",
  43026=>"101101010",
  43027=>"101001001",
  43028=>"001000011",
  43029=>"001010110",
  43030=>"000011011",
  43031=>"000010001",
  43032=>"010101111",
  43033=>"011011110",
  43034=>"010001010",
  43035=>"110001100",
  43036=>"011110000",
  43037=>"011100110",
  43038=>"011001111",
  43039=>"101111001",
  43040=>"111101011",
  43041=>"100001010",
  43042=>"101000010",
  43043=>"011100110",
  43044=>"011001010",
  43045=>"011001011",
  43046=>"101100000",
  43047=>"110101100",
  43048=>"111110110",
  43049=>"000011111",
  43050=>"110111111",
  43051=>"100101000",
  43052=>"010101001",
  43053=>"110111000",
  43054=>"111100010",
  43055=>"110000100",
  43056=>"001101110",
  43057=>"101000000",
  43058=>"101101101",
  43059=>"100001000",
  43060=>"101100111",
  43061=>"111100110",
  43062=>"001001000",
  43063=>"011001100",
  43064=>"001111110",
  43065=>"111000011",
  43066=>"000100011",
  43067=>"010010110",
  43068=>"010001010",
  43069=>"111000011",
  43070=>"100000010",
  43071=>"100000000",
  43072=>"010000010",
  43073=>"000110001",
  43074=>"110110111",
  43075=>"010101010",
  43076=>"010110110",
  43077=>"101010001",
  43078=>"110110110",
  43079=>"011101111",
  43080=>"110100001",
  43081=>"011111100",
  43082=>"001100101",
  43083=>"001100110",
  43084=>"000111011",
  43085=>"111100100",
  43086=>"001100000",
  43087=>"100000001",
  43088=>"000111110",
  43089=>"001011010",
  43090=>"000010001",
  43091=>"000101111",
  43092=>"110111001",
  43093=>"000011011",
  43094=>"111010111",
  43095=>"010110000",
  43096=>"010111111",
  43097=>"101110111",
  43098=>"101011011",
  43099=>"110011111",
  43100=>"000011110",
  43101=>"100110000",
  43102=>"111101011",
  43103=>"000101001",
  43104=>"111001011",
  43105=>"101100101",
  43106=>"000000001",
  43107=>"101101000",
  43108=>"011100101",
  43109=>"100101100",
  43110=>"001100111",
  43111=>"000101100",
  43112=>"111010100",
  43113=>"101100000",
  43114=>"111000011",
  43115=>"000011001",
  43116=>"011001000",
  43117=>"000000001",
  43118=>"110011010",
  43119=>"000100010",
  43120=>"111010000",
  43121=>"001110001",
  43122=>"101111010",
  43123=>"110101101",
  43124=>"100000011",
  43125=>"100011011",
  43126=>"100010101",
  43127=>"010010000",
  43128=>"100111110",
  43129=>"011111100",
  43130=>"111011011",
  43131=>"001111001",
  43132=>"100100101",
  43133=>"111000000",
  43134=>"100000000",
  43135=>"011111010",
  43136=>"011000110",
  43137=>"101100010",
  43138=>"110000011",
  43139=>"010111010",
  43140=>"110101001",
  43141=>"100100010",
  43142=>"011101011",
  43143=>"000010110",
  43144=>"000001000",
  43145=>"101101111",
  43146=>"001000100",
  43147=>"100011111",
  43148=>"001011100",
  43149=>"111110010",
  43150=>"111000000",
  43151=>"000100110",
  43152=>"001100111",
  43153=>"111100001",
  43154=>"110100000",
  43155=>"110101001",
  43156=>"111000000",
  43157=>"001001001",
  43158=>"101011000",
  43159=>"110101000",
  43160=>"011101100",
  43161=>"010001001",
  43162=>"001000011",
  43163=>"000001100",
  43164=>"000101000",
  43165=>"011111100",
  43166=>"110110001",
  43167=>"011011011",
  43168=>"101100010",
  43169=>"100001001",
  43170=>"101001100",
  43171=>"011001010",
  43172=>"100110011",
  43173=>"101100000",
  43174=>"101111111",
  43175=>"101111101",
  43176=>"011011000",
  43177=>"001100101",
  43178=>"011010001",
  43179=>"011101100",
  43180=>"111011010",
  43181=>"100110000",
  43182=>"101000100",
  43183=>"001110101",
  43184=>"101000111",
  43185=>"110000101",
  43186=>"101100110",
  43187=>"000001000",
  43188=>"001001001",
  43189=>"110010011",
  43190=>"000010101",
  43191=>"100110100",
  43192=>"010010010",
  43193=>"001010001",
  43194=>"001000010",
  43195=>"000110011",
  43196=>"001011011",
  43197=>"011000100",
  43198=>"010011101",
  43199=>"100010000",
  43200=>"010101100",
  43201=>"101001001",
  43202=>"001110011",
  43203=>"101011011",
  43204=>"000000111",
  43205=>"100000001",
  43206=>"000101101",
  43207=>"000001000",
  43208=>"101001110",
  43209=>"100001111",
  43210=>"101001110",
  43211=>"011011000",
  43212=>"111100010",
  43213=>"110110011",
  43214=>"001111000",
  43215=>"000011010",
  43216=>"101110101",
  43217=>"011000101",
  43218=>"001100001",
  43219=>"001001101",
  43220=>"110001101",
  43221=>"110100100",
  43222=>"100111000",
  43223=>"000100110",
  43224=>"100101001",
  43225=>"010001100",
  43226=>"110110011",
  43227=>"001101110",
  43228=>"000000011",
  43229=>"000001100",
  43230=>"011010001",
  43231=>"011001110",
  43232=>"011000001",
  43233=>"111011000",
  43234=>"111001011",
  43235=>"010000000",
  43236=>"001011010",
  43237=>"001111100",
  43238=>"001101011",
  43239=>"011100001",
  43240=>"001011000",
  43241=>"001001000",
  43242=>"101111101",
  43243=>"000010001",
  43244=>"010111001",
  43245=>"000000000",
  43246=>"110001001",
  43247=>"110111000",
  43248=>"111110111",
  43249=>"011011000",
  43250=>"010011010",
  43251=>"111010001",
  43252=>"101101100",
  43253=>"111101000",
  43254=>"111011101",
  43255=>"010010001",
  43256=>"101011101",
  43257=>"100101100",
  43258=>"000110001",
  43259=>"000010101",
  43260=>"001110110",
  43261=>"101100001",
  43262=>"001000010",
  43263=>"000101100",
  43264=>"101011110",
  43265=>"011000000",
  43266=>"010010111",
  43267=>"001100010",
  43268=>"001111110",
  43269=>"011100100",
  43270=>"111000110",
  43271=>"001000011",
  43272=>"001000101",
  43273=>"111011101",
  43274=>"101011000",
  43275=>"001000111",
  43276=>"010100001",
  43277=>"010010111",
  43278=>"111100111",
  43279=>"111110101",
  43280=>"110111100",
  43281=>"010100010",
  43282=>"110001100",
  43283=>"011110000",
  43284=>"000000000",
  43285=>"110101010",
  43286=>"010110000",
  43287=>"001110001",
  43288=>"010101000",
  43289=>"100011100",
  43290=>"011100000",
  43291=>"000001000",
  43292=>"000000000",
  43293=>"001000011",
  43294=>"101110000",
  43295=>"011011001",
  43296=>"110110101",
  43297=>"101000000",
  43298=>"011100010",
  43299=>"000010010",
  43300=>"100100010",
  43301=>"000000101",
  43302=>"011011111",
  43303=>"101101010",
  43304=>"000100100",
  43305=>"101100000",
  43306=>"110101001",
  43307=>"010000000",
  43308=>"110010100",
  43309=>"000101010",
  43310=>"111010100",
  43311=>"011000101",
  43312=>"101011001",
  43313=>"101110100",
  43314=>"101000011",
  43315=>"100001010",
  43316=>"110000100",
  43317=>"001001000",
  43318=>"110111100",
  43319=>"011001000",
  43320=>"100000110",
  43321=>"101011000",
  43322=>"011110110",
  43323=>"100101011",
  43324=>"001100000",
  43325=>"001101000",
  43326=>"010001100",
  43327=>"001010001",
  43328=>"011011110",
  43329=>"110010000",
  43330=>"101000010",
  43331=>"111100110",
  43332=>"001100110",
  43333=>"011111110",
  43334=>"011001111",
  43335=>"000001010",
  43336=>"011101010",
  43337=>"000010100",
  43338=>"111100100",
  43339=>"110110110",
  43340=>"001101010",
  43341=>"010100010",
  43342=>"010110000",
  43343=>"001010011",
  43344=>"110001000",
  43345=>"001111010",
  43346=>"011011000",
  43347=>"011101001",
  43348=>"101100100",
  43349=>"011111011",
  43350=>"011100010",
  43351=>"101110011",
  43352=>"000111111",
  43353=>"010010000",
  43354=>"110010000",
  43355=>"110001111",
  43356=>"000101111",
  43357=>"001010011",
  43358=>"100111101",
  43359=>"011110011",
  43360=>"111011011",
  43361=>"001011010",
  43362=>"001110110",
  43363=>"011000101",
  43364=>"001011100",
  43365=>"000110100",
  43366=>"100010101",
  43367=>"011100111",
  43368=>"001100101",
  43369=>"010111010",
  43370=>"010000001",
  43371=>"011010011",
  43372=>"011001100",
  43373=>"000011101",
  43374=>"101000010",
  43375=>"010001101",
  43376=>"101000111",
  43377=>"111010001",
  43378=>"111000000",
  43379=>"001010111",
  43380=>"010000010",
  43381=>"000101000",
  43382=>"110010010",
  43383=>"010101000",
  43384=>"101101100",
  43385=>"110010000",
  43386=>"100110110",
  43387=>"110011100",
  43388=>"000110000",
  43389=>"001001001",
  43390=>"010111110",
  43391=>"000100010",
  43392=>"111001100",
  43393=>"110000010",
  43394=>"011100000",
  43395=>"100100010",
  43396=>"111100110",
  43397=>"000001001",
  43398=>"000000011",
  43399=>"001010101",
  43400=>"000000000",
  43401=>"001011010",
  43402=>"100010111",
  43403=>"010010100",
  43404=>"100010110",
  43405=>"100100111",
  43406=>"010100010",
  43407=>"001100110",
  43408=>"100110001",
  43409=>"001111111",
  43410=>"110111111",
  43411=>"100110110",
  43412=>"001100001",
  43413=>"110110110",
  43414=>"000011111",
  43415=>"011011100",
  43416=>"011011110",
  43417=>"111111001",
  43418=>"111101001",
  43419=>"000011000",
  43420=>"101111111",
  43421=>"101111000",
  43422=>"111010001",
  43423=>"000110010",
  43424=>"011101010",
  43425=>"111011110",
  43426=>"101011001",
  43427=>"110110100",
  43428=>"100001101",
  43429=>"100011101",
  43430=>"011110010",
  43431=>"011100100",
  43432=>"100010110",
  43433=>"001001100",
  43434=>"000111101",
  43435=>"111001001",
  43436=>"011000011",
  43437=>"101010010",
  43438=>"101000101",
  43439=>"111111001",
  43440=>"000101001",
  43441=>"010001111",
  43442=>"011110100",
  43443=>"000011001",
  43444=>"110001110",
  43445=>"000111100",
  43446=>"011111100",
  43447=>"100010101",
  43448=>"111111111",
  43449=>"111010100",
  43450=>"000111001",
  43451=>"011100110",
  43452=>"111110010",
  43453=>"000011101",
  43454=>"110111101",
  43455=>"101110011",
  43456=>"111100011",
  43457=>"000001011",
  43458=>"000110110",
  43459=>"010000100",
  43460=>"000001011",
  43461=>"010110010",
  43462=>"000111110",
  43463=>"110010000",
  43464=>"101101101",
  43465=>"000111011",
  43466=>"111110111",
  43467=>"000101011",
  43468=>"110001011",
  43469=>"000111000",
  43470=>"000010101",
  43471=>"100100100",
  43472=>"111011010",
  43473=>"111000010",
  43474=>"111101101",
  43475=>"000001010",
  43476=>"111111101",
  43477=>"011000111",
  43478=>"000001000",
  43479=>"101011010",
  43480=>"111111110",
  43481=>"101010111",
  43482=>"011011101",
  43483=>"011100001",
  43484=>"011001000",
  43485=>"111011101",
  43486=>"111100001",
  43487=>"001011100",
  43488=>"011010010",
  43489=>"110010001",
  43490=>"101010011",
  43491=>"001010110",
  43492=>"000110001",
  43493=>"111010101",
  43494=>"010111100",
  43495=>"010100110",
  43496=>"101110011",
  43497=>"011000110",
  43498=>"010000110",
  43499=>"110110001",
  43500=>"001011001",
  43501=>"001110001",
  43502=>"011100101",
  43503=>"001010100",
  43504=>"100011111",
  43505=>"011000101",
  43506=>"000000000",
  43507=>"000111000",
  43508=>"110101010",
  43509=>"111100100",
  43510=>"000110100",
  43511=>"100000011",
  43512=>"001010100",
  43513=>"000101110",
  43514=>"101010010",
  43515=>"100011111",
  43516=>"111010100",
  43517=>"001100000",
  43518=>"010100101",
  43519=>"000100110",
  43520=>"101010100",
  43521=>"001000110",
  43522=>"111100001",
  43523=>"100001000",
  43524=>"000100011",
  43525=>"110010111",
  43526=>"111001100",
  43527=>"010011010",
  43528=>"011001000",
  43529=>"101110110",
  43530=>"001000010",
  43531=>"111110110",
  43532=>"100011110",
  43533=>"000100001",
  43534=>"100010110",
  43535=>"011001100",
  43536=>"001101110",
  43537=>"011101000",
  43538=>"100100110",
  43539=>"001110100",
  43540=>"010111010",
  43541=>"101001101",
  43542=>"110101110",
  43543=>"000110010",
  43544=>"010001111",
  43545=>"101111101",
  43546=>"011100001",
  43547=>"111000011",
  43548=>"110100011",
  43549=>"110110011",
  43550=>"000001101",
  43551=>"011111001",
  43552=>"111111001",
  43553=>"111111100",
  43554=>"110100101",
  43555=>"100101010",
  43556=>"011110011",
  43557=>"011011101",
  43558=>"101000010",
  43559=>"010111011",
  43560=>"001001110",
  43561=>"100101111",
  43562=>"101010000",
  43563=>"101111010",
  43564=>"110100000",
  43565=>"011111011",
  43566=>"011111001",
  43567=>"111100101",
  43568=>"010011010",
  43569=>"011001111",
  43570=>"101001101",
  43571=>"010010000",
  43572=>"101010001",
  43573=>"100110111",
  43574=>"101111010",
  43575=>"001001000",
  43576=>"101101111",
  43577=>"001110111",
  43578=>"011100010",
  43579=>"010101010",
  43580=>"111011011",
  43581=>"000000011",
  43582=>"001000110",
  43583=>"111110111",
  43584=>"101111010",
  43585=>"100010000",
  43586=>"001111010",
  43587=>"100100011",
  43588=>"111101110",
  43589=>"001001001",
  43590=>"110001001",
  43591=>"000100001",
  43592=>"000100100",
  43593=>"000100001",
  43594=>"110010011",
  43595=>"001011110",
  43596=>"101110110",
  43597=>"001000001",
  43598=>"011101001",
  43599=>"000011110",
  43600=>"111010111",
  43601=>"111100000",
  43602=>"011110011",
  43603=>"101100100",
  43604=>"000010010",
  43605=>"011100010",
  43606=>"000011111",
  43607=>"000110110",
  43608=>"111011111",
  43609=>"011000001",
  43610=>"010101110",
  43611=>"001001001",
  43612=>"110111110",
  43613=>"100100000",
  43614=>"101101110",
  43615=>"111010111",
  43616=>"011011100",
  43617=>"001010011",
  43618=>"000010100",
  43619=>"101111000",
  43620=>"110000100",
  43621=>"100011101",
  43622=>"001010011",
  43623=>"111111011",
  43624=>"010111101",
  43625=>"010000101",
  43626=>"011100100",
  43627=>"001011010",
  43628=>"000010000",
  43629=>"011000111",
  43630=>"000010011",
  43631=>"101100010",
  43632=>"010000100",
  43633=>"000101010",
  43634=>"111110111",
  43635=>"010111000",
  43636=>"100011011",
  43637=>"101011010",
  43638=>"011101110",
  43639=>"111101100",
  43640=>"011011010",
  43641=>"110111101",
  43642=>"011100001",
  43643=>"010100110",
  43644=>"011100101",
  43645=>"000101000",
  43646=>"111000001",
  43647=>"011000111",
  43648=>"000110001",
  43649=>"111001111",
  43650=>"001001111",
  43651=>"000000100",
  43652=>"101000000",
  43653=>"000010010",
  43654=>"111000101",
  43655=>"000111000",
  43656=>"000111110",
  43657=>"000111000",
  43658=>"110100111",
  43659=>"111101101",
  43660=>"100101011",
  43661=>"100110000",
  43662=>"111001000",
  43663=>"100011111",
  43664=>"111101101",
  43665=>"111101101",
  43666=>"110100011",
  43667=>"100100011",
  43668=>"001100000",
  43669=>"000110110",
  43670=>"010011101",
  43671=>"110011011",
  43672=>"001001101",
  43673=>"100000001",
  43674=>"110010100",
  43675=>"001000110",
  43676=>"100000101",
  43677=>"100100011",
  43678=>"001010010",
  43679=>"011010000",
  43680=>"110111111",
  43681=>"111110101",
  43682=>"101001001",
  43683=>"001010100",
  43684=>"001001001",
  43685=>"011111100",
  43686=>"101001111",
  43687=>"000111001",
  43688=>"001101101",
  43689=>"001110111",
  43690=>"000010111",
  43691=>"111011000",
  43692=>"000101100",
  43693=>"010101011",
  43694=>"011010101",
  43695=>"000000101",
  43696=>"000001000",
  43697=>"010001100",
  43698=>"101010101",
  43699=>"010100101",
  43700=>"110011000",
  43701=>"111110001",
  43702=>"011111111",
  43703=>"010010011",
  43704=>"000001010",
  43705=>"010110110",
  43706=>"001011100",
  43707=>"111110100",
  43708=>"101110010",
  43709=>"011010011",
  43710=>"011101111",
  43711=>"011010110",
  43712=>"011000001",
  43713=>"011100101",
  43714=>"000101111",
  43715=>"101110101",
  43716=>"101100011",
  43717=>"000100101",
  43718=>"111110110",
  43719=>"000100111",
  43720=>"110101110",
  43721=>"010100011",
  43722=>"111101111",
  43723=>"001100010",
  43724=>"111111001",
  43725=>"011011101",
  43726=>"100000000",
  43727=>"010110111",
  43728=>"010101110",
  43729=>"011101100",
  43730=>"101011100",
  43731=>"111111111",
  43732=>"100110100",
  43733=>"010011001",
  43734=>"111101101",
  43735=>"011001101",
  43736=>"011001101",
  43737=>"111001000",
  43738=>"110011100",
  43739=>"111000111",
  43740=>"000111011",
  43741=>"001011001",
  43742=>"111100001",
  43743=>"100000000",
  43744=>"110100101",
  43745=>"000011100",
  43746=>"010101001",
  43747=>"000001001",
  43748=>"110000100",
  43749=>"111111011",
  43750=>"110101010",
  43751=>"000100010",
  43752=>"101011110",
  43753=>"111011011",
  43754=>"111110010",
  43755=>"001011001",
  43756=>"110100110",
  43757=>"011001000",
  43758=>"000000110",
  43759=>"100110011",
  43760=>"110101100",
  43761=>"011111010",
  43762=>"000000110",
  43763=>"011101101",
  43764=>"010101010",
  43765=>"010000101",
  43766=>"111111001",
  43767=>"011000100",
  43768=>"100111100",
  43769=>"111000101",
  43770=>"011111110",
  43771=>"100010010",
  43772=>"010000000",
  43773=>"001000001",
  43774=>"111010110",
  43775=>"001010101",
  43776=>"110010101",
  43777=>"101111100",
  43778=>"011011001",
  43779=>"101111000",
  43780=>"011111111",
  43781=>"001000110",
  43782=>"001001011",
  43783=>"001011111",
  43784=>"001110110",
  43785=>"111001101",
  43786=>"101111111",
  43787=>"001010111",
  43788=>"101000101",
  43789=>"101000110",
  43790=>"101011000",
  43791=>"100010000",
  43792=>"100010000",
  43793=>"000011001",
  43794=>"111011001",
  43795=>"110001111",
  43796=>"101101011",
  43797=>"001000100",
  43798=>"111110011",
  43799=>"101001111",
  43800=>"101011011",
  43801=>"010110111",
  43802=>"100100010",
  43803=>"100100000",
  43804=>"001011010",
  43805=>"001111011",
  43806=>"011110000",
  43807=>"111101100",
  43808=>"000110110",
  43809=>"011111000",
  43810=>"111101001",
  43811=>"100001001",
  43812=>"111110011",
  43813=>"000011011",
  43814=>"100100011",
  43815=>"011101010",
  43816=>"000101101",
  43817=>"100001100",
  43818=>"111111110",
  43819=>"000100010",
  43820=>"110000101",
  43821=>"000111110",
  43822=>"011011011",
  43823=>"101000001",
  43824=>"101111101",
  43825=>"111100001",
  43826=>"010111011",
  43827=>"100011010",
  43828=>"001001110",
  43829=>"111100000",
  43830=>"000000101",
  43831=>"000101100",
  43832=>"101111000",
  43833=>"000111111",
  43834=>"110111011",
  43835=>"000010000",
  43836=>"111001100",
  43837=>"000011010",
  43838=>"000001000",
  43839=>"001001011",
  43840=>"000100110",
  43841=>"001110110",
  43842=>"111111111",
  43843=>"000000000",
  43844=>"111101000",
  43845=>"100001100",
  43846=>"001100010",
  43847=>"111111111",
  43848=>"010110111",
  43849=>"101011000",
  43850=>"010111101",
  43851=>"000010001",
  43852=>"000101110",
  43853=>"001101000",
  43854=>"011100101",
  43855=>"101010010",
  43856=>"100111111",
  43857=>"000000010",
  43858=>"011001010",
  43859=>"001010011",
  43860=>"111111101",
  43861=>"111000101",
  43862=>"010100110",
  43863=>"110100010",
  43864=>"011110111",
  43865=>"101011001",
  43866=>"111110101",
  43867=>"011010111",
  43868=>"001110101",
  43869=>"011111110",
  43870=>"101010000",
  43871=>"010000110",
  43872=>"100000000",
  43873=>"110001111",
  43874=>"010010100",
  43875=>"111110001",
  43876=>"101000001",
  43877=>"100110110",
  43878=>"100101110",
  43879=>"101010000",
  43880=>"111000010",
  43881=>"000100100",
  43882=>"010010111",
  43883=>"101010010",
  43884=>"010101111",
  43885=>"011001100",
  43886=>"000100101",
  43887=>"100000010",
  43888=>"010111111",
  43889=>"111101111",
  43890=>"010111011",
  43891=>"001000100",
  43892=>"011101011",
  43893=>"110110111",
  43894=>"010001010",
  43895=>"100101100",
  43896=>"111000110",
  43897=>"111101000",
  43898=>"111100001",
  43899=>"011000101",
  43900=>"011010000",
  43901=>"011000000",
  43902=>"011100000",
  43903=>"011110000",
  43904=>"100111000",
  43905=>"101010101",
  43906=>"000011000",
  43907=>"010101100",
  43908=>"101101100",
  43909=>"110010101",
  43910=>"000110000",
  43911=>"001010110",
  43912=>"100110000",
  43913=>"111000110",
  43914=>"001001011",
  43915=>"011001101",
  43916=>"111101111",
  43917=>"001111010",
  43918=>"011000101",
  43919=>"110101001",
  43920=>"110001010",
  43921=>"100100100",
  43922=>"000110001",
  43923=>"111000011",
  43924=>"011001100",
  43925=>"101101101",
  43926=>"001110110",
  43927=>"000111000",
  43928=>"111011000",
  43929=>"010100001",
  43930=>"111000011",
  43931=>"011011010",
  43932=>"011111001",
  43933=>"010010010",
  43934=>"101001011",
  43935=>"001000110",
  43936=>"111001110",
  43937=>"011101110",
  43938=>"001001100",
  43939=>"001011101",
  43940=>"010000001",
  43941=>"011001001",
  43942=>"010010000",
  43943=>"010010010",
  43944=>"001000100",
  43945=>"101000110",
  43946=>"010000111",
  43947=>"111001111",
  43948=>"010001101",
  43949=>"011100011",
  43950=>"011011011",
  43951=>"011000001",
  43952=>"101101001",
  43953=>"110001001",
  43954=>"111010010",
  43955=>"101101010",
  43956=>"100000000",
  43957=>"011000110",
  43958=>"101110000",
  43959=>"101110101",
  43960=>"011001100",
  43961=>"000010011",
  43962=>"011000010",
  43963=>"110110100",
  43964=>"111100100",
  43965=>"111101101",
  43966=>"010000100",
  43967=>"000011010",
  43968=>"101100000",
  43969=>"001101011",
  43970=>"000010110",
  43971=>"001011010",
  43972=>"111101101",
  43973=>"101011001",
  43974=>"101110001",
  43975=>"001110111",
  43976=>"110001100",
  43977=>"110111001",
  43978=>"011010000",
  43979=>"001111111",
  43980=>"100010001",
  43981=>"000011001",
  43982=>"100101111",
  43983=>"010000110",
  43984=>"010111011",
  43985=>"000110011",
  43986=>"101110010",
  43987=>"101101000",
  43988=>"010110101",
  43989=>"011111000",
  43990=>"001100101",
  43991=>"100101000",
  43992=>"010011010",
  43993=>"111100100",
  43994=>"011101000",
  43995=>"100010110",
  43996=>"001101101",
  43997=>"111001111",
  43998=>"110110101",
  43999=>"010000111",
  44000=>"101001001",
  44001=>"111101100",
  44002=>"011100000",
  44003=>"010101111",
  44004=>"101010011",
  44005=>"011111011",
  44006=>"100100000",
  44007=>"100010010",
  44008=>"101101100",
  44009=>"111100110",
  44010=>"111011101",
  44011=>"100000101",
  44012=>"011110100",
  44013=>"101001101",
  44014=>"111010010",
  44015=>"110000001",
  44016=>"010010010",
  44017=>"111101000",
  44018=>"000000111",
  44019=>"111110111",
  44020=>"110010100",
  44021=>"111000111",
  44022=>"111110001",
  44023=>"111111000",
  44024=>"101111011",
  44025=>"001101011",
  44026=>"001011001",
  44027=>"111001011",
  44028=>"010001101",
  44029=>"101011110",
  44030=>"111011011",
  44031=>"111001111",
  44032=>"101110101",
  44033=>"111011011",
  44034=>"110100000",
  44035=>"110100110",
  44036=>"100100101",
  44037=>"100010010",
  44038=>"111110011",
  44039=>"010110100",
  44040=>"010111010",
  44041=>"000110010",
  44042=>"111100010",
  44043=>"011111110",
  44044=>"110001011",
  44045=>"001000010",
  44046=>"000010100",
  44047=>"101011011",
  44048=>"011000010",
  44049=>"010101101",
  44050=>"100110111",
  44051=>"011001011",
  44052=>"000010110",
  44053=>"010000011",
  44054=>"000010001",
  44055=>"100111001",
  44056=>"010011100",
  44057=>"000110001",
  44058=>"110101100",
  44059=>"100000100",
  44060=>"110110110",
  44061=>"101100111",
  44062=>"001001110",
  44063=>"100110111",
  44064=>"001101011",
  44065=>"100001101",
  44066=>"111100001",
  44067=>"010101001",
  44068=>"100011100",
  44069=>"000100111",
  44070=>"101111000",
  44071=>"100111011",
  44072=>"101101001",
  44073=>"101001010",
  44074=>"101111001",
  44075=>"111000101",
  44076=>"000010010",
  44077=>"000110010",
  44078=>"011010111",
  44079=>"011010001",
  44080=>"101011111",
  44081=>"000110111",
  44082=>"011110101",
  44083=>"101100000",
  44084=>"001111010",
  44085=>"100101001",
  44086=>"101110100",
  44087=>"111111001",
  44088=>"110000010",
  44089=>"100001010",
  44090=>"101100110",
  44091=>"000100000",
  44092=>"100011100",
  44093=>"110011110",
  44094=>"001001100",
  44095=>"111000011",
  44096=>"100111101",
  44097=>"011001110",
  44098=>"100100001",
  44099=>"010110000",
  44100=>"000010010",
  44101=>"010100101",
  44102=>"001110110",
  44103=>"110001001",
  44104=>"110000001",
  44105=>"101011110",
  44106=>"010001001",
  44107=>"011101011",
  44108=>"110011010",
  44109=>"100011011",
  44110=>"000110111",
  44111=>"101111111",
  44112=>"001111100",
  44113=>"000000100",
  44114=>"100100001",
  44115=>"001010101",
  44116=>"110000011",
  44117=>"000101001",
  44118=>"001011100",
  44119=>"110110011",
  44120=>"111110001",
  44121=>"101111011",
  44122=>"111011110",
  44123=>"001011100",
  44124=>"100001011",
  44125=>"001101100",
  44126=>"001001010",
  44127=>"010001111",
  44128=>"111000000",
  44129=>"111010101",
  44130=>"111110110",
  44131=>"110100110",
  44132=>"110100111",
  44133=>"111010000",
  44134=>"000011001",
  44135=>"000100100",
  44136=>"010111101",
  44137=>"001011010",
  44138=>"000100010",
  44139=>"010110011",
  44140=>"011110111",
  44141=>"101001100",
  44142=>"101011011",
  44143=>"110101011",
  44144=>"010010011",
  44145=>"011011010",
  44146=>"100010100",
  44147=>"111111100",
  44148=>"101011110",
  44149=>"111010101",
  44150=>"111110100",
  44151=>"001011010",
  44152=>"101101000",
  44153=>"110000010",
  44154=>"100011011",
  44155=>"011010100",
  44156=>"011110001",
  44157=>"111111010",
  44158=>"111011100",
  44159=>"101111111",
  44160=>"010110011",
  44161=>"110110100",
  44162=>"100110111",
  44163=>"010000000",
  44164=>"011100100",
  44165=>"111110011",
  44166=>"111111100",
  44167=>"001011000",
  44168=>"111010110",
  44169=>"110101110",
  44170=>"011100001",
  44171=>"101101110",
  44172=>"100000001",
  44173=>"100000001",
  44174=>"000001000",
  44175=>"111011100",
  44176=>"100000110",
  44177=>"110001001",
  44178=>"001001011",
  44179=>"101100010",
  44180=>"101100001",
  44181=>"111010001",
  44182=>"111000000",
  44183=>"000100100",
  44184=>"011101111",
  44185=>"011000000",
  44186=>"011110011",
  44187=>"001100101",
  44188=>"000100101",
  44189=>"000101001",
  44190=>"110011010",
  44191=>"100101001",
  44192=>"000000001",
  44193=>"110101111",
  44194=>"011010100",
  44195=>"000010110",
  44196=>"101100111",
  44197=>"101110010",
  44198=>"000111010",
  44199=>"000100010",
  44200=>"011010100",
  44201=>"010001101",
  44202=>"000111111",
  44203=>"111000110",
  44204=>"001000001",
  44205=>"011111101",
  44206=>"110111011",
  44207=>"110100110",
  44208=>"110000111",
  44209=>"110100101",
  44210=>"101111111",
  44211=>"100011101",
  44212=>"001001010",
  44213=>"110101110",
  44214=>"001000100",
  44215=>"100111001",
  44216=>"110001011",
  44217=>"001111110",
  44218=>"011001111",
  44219=>"101011011",
  44220=>"001010111",
  44221=>"110000111",
  44222=>"100011010",
  44223=>"101111011",
  44224=>"011000100",
  44225=>"001010101",
  44226=>"001100010",
  44227=>"000101110",
  44228=>"010101100",
  44229=>"101100010",
  44230=>"011100001",
  44231=>"011110000",
  44232=>"100000111",
  44233=>"111010111",
  44234=>"011100011",
  44235=>"011000101",
  44236=>"000010111",
  44237=>"011011011",
  44238=>"011110101",
  44239=>"101110110",
  44240=>"110110100",
  44241=>"001100000",
  44242=>"110010111",
  44243=>"001000001",
  44244=>"000000001",
  44245=>"001111010",
  44246=>"011000000",
  44247=>"011001010",
  44248=>"010001001",
  44249=>"101011001",
  44250=>"000111010",
  44251=>"001011100",
  44252=>"100001110",
  44253=>"000111101",
  44254=>"010101011",
  44255=>"001010010",
  44256=>"000010100",
  44257=>"100000000",
  44258=>"110100001",
  44259=>"110111000",
  44260=>"001101010",
  44261=>"111111000",
  44262=>"001011010",
  44263=>"011000110",
  44264=>"111100001",
  44265=>"101010000",
  44266=>"101001000",
  44267=>"101111011",
  44268=>"001000101",
  44269=>"111111101",
  44270=>"110101111",
  44271=>"100111111",
  44272=>"100001100",
  44273=>"111000100",
  44274=>"111001101",
  44275=>"010101110",
  44276=>"101001110",
  44277=>"000101010",
  44278=>"000111000",
  44279=>"001010010",
  44280=>"100100100",
  44281=>"000011100",
  44282=>"110110100",
  44283=>"000101010",
  44284=>"110101010",
  44285=>"101110010",
  44286=>"111101111",
  44287=>"111111011",
  44288=>"100001011",
  44289=>"111100000",
  44290=>"100110110",
  44291=>"111101101",
  44292=>"010000111",
  44293=>"011111011",
  44294=>"010011110",
  44295=>"101010110",
  44296=>"011110101",
  44297=>"100000110",
  44298=>"011101111",
  44299=>"110001110",
  44300=>"000000001",
  44301=>"111000111",
  44302=>"100000110",
  44303=>"111101001",
  44304=>"110000011",
  44305=>"001001110",
  44306=>"001001111",
  44307=>"101011100",
  44308=>"000011110",
  44309=>"110111101",
  44310=>"111000000",
  44311=>"110101101",
  44312=>"101110010",
  44313=>"000000011",
  44314=>"011111000",
  44315=>"000111101",
  44316=>"000001111",
  44317=>"000001100",
  44318=>"100010101",
  44319=>"100101010",
  44320=>"100110110",
  44321=>"111001000",
  44322=>"101111111",
  44323=>"011000001",
  44324=>"000110000",
  44325=>"010110101",
  44326=>"010011100",
  44327=>"100010011",
  44328=>"010111111",
  44329=>"101101101",
  44330=>"001110010",
  44331=>"110100110",
  44332=>"011011100",
  44333=>"101101101",
  44334=>"000000000",
  44335=>"110001000",
  44336=>"101101000",
  44337=>"101110101",
  44338=>"111110100",
  44339=>"101000010",
  44340=>"001100011",
  44341=>"010010110",
  44342=>"110000010",
  44343=>"000101000",
  44344=>"000011010",
  44345=>"111111011",
  44346=>"000011001",
  44347=>"011000010",
  44348=>"001111110",
  44349=>"011000111",
  44350=>"010001000",
  44351=>"101111101",
  44352=>"011001000",
  44353=>"001011011",
  44354=>"000000101",
  44355=>"101001010",
  44356=>"111101000",
  44357=>"101010011",
  44358=>"100000001",
  44359=>"100111000",
  44360=>"010001000",
  44361=>"010011111",
  44362=>"110011111",
  44363=>"111100111",
  44364=>"110001000",
  44365=>"010101011",
  44366=>"000111111",
  44367=>"000100100",
  44368=>"100010001",
  44369=>"010111011",
  44370=>"100101001",
  44371=>"111110011",
  44372=>"100101101",
  44373=>"110011000",
  44374=>"100011011",
  44375=>"100010101",
  44376=>"101111110",
  44377=>"000011001",
  44378=>"100010000",
  44379=>"100001111",
  44380=>"011000110",
  44381=>"111011101",
  44382=>"010011000",
  44383=>"110011000",
  44384=>"101010100",
  44385=>"010011001",
  44386=>"001000100",
  44387=>"110100110",
  44388=>"101110011",
  44389=>"001100010",
  44390=>"111100000",
  44391=>"001001100",
  44392=>"100100101",
  44393=>"111100110",
  44394=>"111111010",
  44395=>"101001110",
  44396=>"110101111",
  44397=>"111010100",
  44398=>"100101000",
  44399=>"000111101",
  44400=>"101000101",
  44401=>"100110111",
  44402=>"100110110",
  44403=>"010000100",
  44404=>"101101110",
  44405=>"010100001",
  44406=>"010000111",
  44407=>"000101100",
  44408=>"000101110",
  44409=>"000110000",
  44410=>"100101111",
  44411=>"101101000",
  44412=>"100001101",
  44413=>"100000010",
  44414=>"111011010",
  44415=>"110111011",
  44416=>"001000110",
  44417=>"100010100",
  44418=>"101100001",
  44419=>"101110001",
  44420=>"110110100",
  44421=>"011011000",
  44422=>"000001001",
  44423=>"110011100",
  44424=>"000010011",
  44425=>"110001000",
  44426=>"110000001",
  44427=>"000000111",
  44428=>"000000000",
  44429=>"000000001",
  44430=>"100000011",
  44431=>"100001110",
  44432=>"001110111",
  44433=>"000010101",
  44434=>"011100110",
  44435=>"000001000",
  44436=>"100010000",
  44437=>"110110001",
  44438=>"100011100",
  44439=>"011001010",
  44440=>"111000111",
  44441=>"000100110",
  44442=>"000001010",
  44443=>"100000100",
  44444=>"100110001",
  44445=>"111111111",
  44446=>"111111010",
  44447=>"110001010",
  44448=>"011010010",
  44449=>"011000101",
  44450=>"101110010",
  44451=>"000100001",
  44452=>"111011101",
  44453=>"011010000",
  44454=>"001111000",
  44455=>"101110100",
  44456=>"011000011",
  44457=>"010000010",
  44458=>"001100011",
  44459=>"011111000",
  44460=>"001100111",
  44461=>"010011111",
  44462=>"011000010",
  44463=>"001101011",
  44464=>"110100010",
  44465=>"101110010",
  44466=>"000101001",
  44467=>"110110101",
  44468=>"100001100",
  44469=>"110100011",
  44470=>"110001110",
  44471=>"011110111",
  44472=>"110011000",
  44473=>"001100010",
  44474=>"000111110",
  44475=>"110111101",
  44476=>"100111111",
  44477=>"010011001",
  44478=>"010110110",
  44479=>"100010010",
  44480=>"101100000",
  44481=>"110010100",
  44482=>"100110000",
  44483=>"001010010",
  44484=>"111101110",
  44485=>"001100100",
  44486=>"001011010",
  44487=>"110100001",
  44488=>"011110100",
  44489=>"111001110",
  44490=>"100010011",
  44491=>"101000001",
  44492=>"010010110",
  44493=>"111000111",
  44494=>"110110101",
  44495=>"101101101",
  44496=>"001010101",
  44497=>"110011000",
  44498=>"111110110",
  44499=>"100100110",
  44500=>"010000011",
  44501=>"000101011",
  44502=>"011001100",
  44503=>"101001010",
  44504=>"011001011",
  44505=>"001111110",
  44506=>"110110111",
  44507=>"010100011",
  44508=>"010001100",
  44509=>"111110010",
  44510=>"100010001",
  44511=>"010110000",
  44512=>"111011010",
  44513=>"111101011",
  44514=>"110000101",
  44515=>"001111011",
  44516=>"110101011",
  44517=>"001011110",
  44518=>"000111000",
  44519=>"101011011",
  44520=>"101111101",
  44521=>"110001010",
  44522=>"001111111",
  44523=>"010111100",
  44524=>"110111000",
  44525=>"111000100",
  44526=>"001000101",
  44527=>"011111011",
  44528=>"101010100",
  44529=>"100110001",
  44530=>"111111111",
  44531=>"011111111",
  44532=>"010111000",
  44533=>"000101011",
  44534=>"101001001",
  44535=>"010100111",
  44536=>"010101010",
  44537=>"111110101",
  44538=>"001001101",
  44539=>"101001100",
  44540=>"000100101",
  44541=>"011100100",
  44542=>"010010001",
  44543=>"101111111",
  44544=>"110001100",
  44545=>"110000110",
  44546=>"010111110",
  44547=>"000011010",
  44548=>"010010111",
  44549=>"011010000",
  44550=>"101011110",
  44551=>"010001100",
  44552=>"010010110",
  44553=>"001001111",
  44554=>"101100110",
  44555=>"111111100",
  44556=>"010011000",
  44557=>"111001000",
  44558=>"001110000",
  44559=>"000110000",
  44560=>"100001110",
  44561=>"111101100",
  44562=>"011011110",
  44563=>"111111111",
  44564=>"110110101",
  44565=>"111100000",
  44566=>"001101000",
  44567=>"001010101",
  44568=>"001111001",
  44569=>"111001000",
  44570=>"110110010",
  44571=>"010110100",
  44572=>"010000111",
  44573=>"111010000",
  44574=>"010011011",
  44575=>"101110000",
  44576=>"111011010",
  44577=>"000111000",
  44578=>"110011010",
  44579=>"100110100",
  44580=>"011000001",
  44581=>"101011100",
  44582=>"001001101",
  44583=>"010001100",
  44584=>"100100101",
  44585=>"010101111",
  44586=>"000000111",
  44587=>"010000000",
  44588=>"101111101",
  44589=>"010011100",
  44590=>"011010001",
  44591=>"110010001",
  44592=>"001001100",
  44593=>"111001100",
  44594=>"110000101",
  44595=>"001010001",
  44596=>"010111111",
  44597=>"010101010",
  44598=>"001010000",
  44599=>"000110111",
  44600=>"101010111",
  44601=>"010001010",
  44602=>"111100011",
  44603=>"010101101",
  44604=>"010000001",
  44605=>"001100011",
  44606=>"001100000",
  44607=>"010101000",
  44608=>"010011000",
  44609=>"100111101",
  44610=>"010110011",
  44611=>"110001101",
  44612=>"000101010",
  44613=>"111000000",
  44614=>"001100101",
  44615=>"111110100",
  44616=>"000100010",
  44617=>"110010011",
  44618=>"110011001",
  44619=>"001010101",
  44620=>"100100001",
  44621=>"001100101",
  44622=>"110010000",
  44623=>"111010101",
  44624=>"011000000",
  44625=>"010010011",
  44626=>"101010011",
  44627=>"000110000",
  44628=>"100110100",
  44629=>"111000000",
  44630=>"100111010",
  44631=>"001100000",
  44632=>"011010010",
  44633=>"101010000",
  44634=>"110010010",
  44635=>"101011100",
  44636=>"010000000",
  44637=>"011110100",
  44638=>"001100010",
  44639=>"111110111",
  44640=>"001000101",
  44641=>"011110011",
  44642=>"110011111",
  44643=>"011111110",
  44644=>"110110110",
  44645=>"111001111",
  44646=>"100001100",
  44647=>"010011001",
  44648=>"010111100",
  44649=>"001100101",
  44650=>"000111111",
  44651=>"000001001",
  44652=>"110100100",
  44653=>"111001111",
  44654=>"100010011",
  44655=>"000011001",
  44656=>"011101111",
  44657=>"110000000",
  44658=>"111101000",
  44659=>"000010110",
  44660=>"000001001",
  44661=>"100100110",
  44662=>"100111011",
  44663=>"101110000",
  44664=>"110101000",
  44665=>"001000101",
  44666=>"110111111",
  44667=>"101010010",
  44668=>"001100110",
  44669=>"110101110",
  44670=>"000000110",
  44671=>"100110000",
  44672=>"010011000",
  44673=>"110001001",
  44674=>"110001010",
  44675=>"110110001",
  44676=>"001101100",
  44677=>"101100110",
  44678=>"011100000",
  44679=>"010111110",
  44680=>"001001110",
  44681=>"010100011",
  44682=>"100001101",
  44683=>"110101001",
  44684=>"100100010",
  44685=>"101111010",
  44686=>"011111001",
  44687=>"100001111",
  44688=>"101101111",
  44689=>"100101000",
  44690=>"011101010",
  44691=>"001000110",
  44692=>"010011111",
  44693=>"110100010",
  44694=>"011010010",
  44695=>"000101110",
  44696=>"011000011",
  44697=>"010100001",
  44698=>"110101000",
  44699=>"101010111",
  44700=>"100000100",
  44701=>"011111010",
  44702=>"000001000",
  44703=>"011111100",
  44704=>"000000001",
  44705=>"000011011",
  44706=>"000011101",
  44707=>"000000110",
  44708=>"011100001",
  44709=>"011011010",
  44710=>"111011001",
  44711=>"000011101",
  44712=>"101111000",
  44713=>"010100010",
  44714=>"000011010",
  44715=>"110011011",
  44716=>"100000110",
  44717=>"001001101",
  44718=>"011000010",
  44719=>"101101111",
  44720=>"101001110",
  44721=>"101110001",
  44722=>"001001011",
  44723=>"100101110",
  44724=>"101101000",
  44725=>"100011101",
  44726=>"100001100",
  44727=>"011010000",
  44728=>"111000111",
  44729=>"110001111",
  44730=>"001011010",
  44731=>"001011100",
  44732=>"011001001",
  44733=>"000100100",
  44734=>"111111111",
  44735=>"011111111",
  44736=>"000001100",
  44737=>"100110011",
  44738=>"001010010",
  44739=>"100110001",
  44740=>"110110110",
  44741=>"001100110",
  44742=>"001010101",
  44743=>"011001011",
  44744=>"010111011",
  44745=>"000010000",
  44746=>"011000001",
  44747=>"000111000",
  44748=>"100010101",
  44749=>"001011001",
  44750=>"100011111",
  44751=>"111010001",
  44752=>"110111001",
  44753=>"001000001",
  44754=>"100001100",
  44755=>"010000010",
  44756=>"001100101",
  44757=>"111100111",
  44758=>"111011110",
  44759=>"001100110",
  44760=>"111000010",
  44761=>"110001110",
  44762=>"000010000",
  44763=>"110110001",
  44764=>"010110111",
  44765=>"010101111",
  44766=>"001011001",
  44767=>"110111111",
  44768=>"101011101",
  44769=>"111010000",
  44770=>"111000010",
  44771=>"101101111",
  44772=>"010000011",
  44773=>"000001011",
  44774=>"111110010",
  44775=>"011100001",
  44776=>"111010100",
  44777=>"001011000",
  44778=>"011111011",
  44779=>"101010000",
  44780=>"000111111",
  44781=>"110111011",
  44782=>"110111001",
  44783=>"101111010",
  44784=>"111011001",
  44785=>"011101011",
  44786=>"001000101",
  44787=>"000001101",
  44788=>"010111110",
  44789=>"110101001",
  44790=>"110010110",
  44791=>"111101100",
  44792=>"001011001",
  44793=>"111100100",
  44794=>"000110100",
  44795=>"011101101",
  44796=>"110001001",
  44797=>"110100110",
  44798=>"101011101",
  44799=>"111111111",
  44800=>"001000011",
  44801=>"111011011",
  44802=>"111101111",
  44803=>"011110101",
  44804=>"111010101",
  44805=>"000000110",
  44806=>"001000010",
  44807=>"001110001",
  44808=>"011010110",
  44809=>"010000110",
  44810=>"111011111",
  44811=>"110110101",
  44812=>"110101110",
  44813=>"011011011",
  44814=>"100101111",
  44815=>"100101100",
  44816=>"101000100",
  44817=>"001000010",
  44818=>"010011011",
  44819=>"000000101",
  44820=>"011000000",
  44821=>"010101101",
  44822=>"010011100",
  44823=>"101100000",
  44824=>"100110100",
  44825=>"100110100",
  44826=>"111111010",
  44827=>"001100000",
  44828=>"001111001",
  44829=>"101011001",
  44830=>"110000110",
  44831=>"001011001",
  44832=>"000100100",
  44833=>"111100001",
  44834=>"000101001",
  44835=>"100100100",
  44836=>"011000011",
  44837=>"011010101",
  44838=>"111101100",
  44839=>"010011110",
  44840=>"111001010",
  44841=>"001111110",
  44842=>"010111111",
  44843=>"111010111",
  44844=>"100011111",
  44845=>"100001101",
  44846=>"000100101",
  44847=>"001011110",
  44848=>"011100111",
  44849=>"100010111",
  44850=>"000010011",
  44851=>"000010001",
  44852=>"000001000",
  44853=>"111000001",
  44854=>"111000011",
  44855=>"110001101",
  44856=>"011110110",
  44857=>"000111100",
  44858=>"110010100",
  44859=>"010101010",
  44860=>"010110010",
  44861=>"000001011",
  44862=>"111010000",
  44863=>"010100101",
  44864=>"000110010",
  44865=>"100111101",
  44866=>"011111110",
  44867=>"101111001",
  44868=>"000010100",
  44869=>"011110000",
  44870=>"001110011",
  44871=>"110001110",
  44872=>"000100000",
  44873=>"010000010",
  44874=>"000101100",
  44875=>"001011000",
  44876=>"010000100",
  44877=>"000111101",
  44878=>"100111000",
  44879=>"101111011",
  44880=>"010111011",
  44881=>"101100101",
  44882=>"111100101",
  44883=>"001101100",
  44884=>"000000111",
  44885=>"101110010",
  44886=>"111100010",
  44887=>"100001101",
  44888=>"010011001",
  44889=>"010110100",
  44890=>"111010111",
  44891=>"111001100",
  44892=>"111001101",
  44893=>"011011001",
  44894=>"111001011",
  44895=>"100100010",
  44896=>"011111101",
  44897=>"100110000",
  44898=>"101000111",
  44899=>"000111001",
  44900=>"001101111",
  44901=>"110000011",
  44902=>"110011011",
  44903=>"010011001",
  44904=>"100000111",
  44905=>"111000100",
  44906=>"110100000",
  44907=>"110101011",
  44908=>"010000011",
  44909=>"101111000",
  44910=>"101100001",
  44911=>"111100011",
  44912=>"010111101",
  44913=>"010101000",
  44914=>"100101110",
  44915=>"101000100",
  44916=>"000001000",
  44917=>"010000000",
  44918=>"010110001",
  44919=>"010000010",
  44920=>"000110111",
  44921=>"001111010",
  44922=>"000000000",
  44923=>"110101100",
  44924=>"111000000",
  44925=>"101000000",
  44926=>"011011110",
  44927=>"100110000",
  44928=>"111100111",
  44929=>"110000110",
  44930=>"010100110",
  44931=>"101000010",
  44932=>"010100000",
  44933=>"100110011",
  44934=>"101110100",
  44935=>"101010111",
  44936=>"110001001",
  44937=>"111000001",
  44938=>"010000110",
  44939=>"000001100",
  44940=>"101011101",
  44941=>"101100101",
  44942=>"111010001",
  44943=>"000111011",
  44944=>"001000011",
  44945=>"010101001",
  44946=>"000010001",
  44947=>"101000000",
  44948=>"011010010",
  44949=>"011100001",
  44950=>"000010111",
  44951=>"001001111",
  44952=>"100001100",
  44953=>"110110010",
  44954=>"010100100",
  44955=>"000000010",
  44956=>"000001101",
  44957=>"001010011",
  44958=>"000110011",
  44959=>"000111100",
  44960=>"000001100",
  44961=>"001110110",
  44962=>"110001100",
  44963=>"000110000",
  44964=>"011111010",
  44965=>"010001110",
  44966=>"000011011",
  44967=>"111101100",
  44968=>"000011000",
  44969=>"001001111",
  44970=>"010110100",
  44971=>"001000100",
  44972=>"111101001",
  44973=>"101001000",
  44974=>"111011100",
  44975=>"001011011",
  44976=>"110101001",
  44977=>"101000000",
  44978=>"001001111",
  44979=>"011100000",
  44980=>"010011100",
  44981=>"000100011",
  44982=>"000010111",
  44983=>"110001001",
  44984=>"011010010",
  44985=>"100111011",
  44986=>"110010111",
  44987=>"000010110",
  44988=>"010110010",
  44989=>"101111100",
  44990=>"010101000",
  44991=>"000000010",
  44992=>"111111101",
  44993=>"001110100",
  44994=>"001101100",
  44995=>"101101100",
  44996=>"111011100",
  44997=>"011110110",
  44998=>"000110011",
  44999=>"101111110",
  45000=>"110001101",
  45001=>"111101111",
  45002=>"111010001",
  45003=>"101111010",
  45004=>"000100010",
  45005=>"110000101",
  45006=>"000100100",
  45007=>"101100100",
  45008=>"101001001",
  45009=>"010000000",
  45010=>"011100111",
  45011=>"001101011",
  45012=>"001011011",
  45013=>"000111010",
  45014=>"001000011",
  45015=>"100110111",
  45016=>"101010011",
  45017=>"000101101",
  45018=>"001101010",
  45019=>"010000011",
  45020=>"001001100",
  45021=>"011111011",
  45022=>"011000111",
  45023=>"010000011",
  45024=>"010101011",
  45025=>"100001010",
  45026=>"101111011",
  45027=>"010011111",
  45028=>"011000101",
  45029=>"111001001",
  45030=>"000111111",
  45031=>"111110111",
  45032=>"000100000",
  45033=>"100000010",
  45034=>"101000010",
  45035=>"001100000",
  45036=>"010111010",
  45037=>"001000010",
  45038=>"110010111",
  45039=>"100001100",
  45040=>"011000000",
  45041=>"101110100",
  45042=>"000011000",
  45043=>"001110010",
  45044=>"001011011",
  45045=>"100010011",
  45046=>"000011001",
  45047=>"000000011",
  45048=>"110011010",
  45049=>"001000001",
  45050=>"100010001",
  45051=>"011101100",
  45052=>"001011111",
  45053=>"000001001",
  45054=>"101001011",
  45055=>"100111100",
  45056=>"000000100",
  45057=>"101010010",
  45058=>"111110101",
  45059=>"001111100",
  45060=>"000111011",
  45061=>"000101010",
  45062=>"000010000",
  45063=>"001001100",
  45064=>"000110000",
  45065=>"010101111",
  45066=>"111011000",
  45067=>"110011011",
  45068=>"101001011",
  45069=>"010111110",
  45070=>"100110011",
  45071=>"111011010",
  45072=>"100001100",
  45073=>"011001101",
  45074=>"101100111",
  45075=>"101100111",
  45076=>"101100111",
  45077=>"111110010",
  45078=>"001000010",
  45079=>"010010100",
  45080=>"000010111",
  45081=>"110101111",
  45082=>"111001001",
  45083=>"000011011",
  45084=>"100011110",
  45085=>"101010110",
  45086=>"001011010",
  45087=>"000110110",
  45088=>"111101001",
  45089=>"011101001",
  45090=>"110011010",
  45091=>"100101011",
  45092=>"000110000",
  45093=>"011100000",
  45094=>"110001111",
  45095=>"101101110",
  45096=>"101000100",
  45097=>"001000011",
  45098=>"100110000",
  45099=>"110010111",
  45100=>"111000100",
  45101=>"010110000",
  45102=>"000100001",
  45103=>"101000011",
  45104=>"011110111",
  45105=>"011000011",
  45106=>"110001011",
  45107=>"010100010",
  45108=>"011000011",
  45109=>"000110001",
  45110=>"111110110",
  45111=>"010100000",
  45112=>"111010111",
  45113=>"010011101",
  45114=>"100010110",
  45115=>"101100110",
  45116=>"100111011",
  45117=>"001101100",
  45118=>"110001001",
  45119=>"000111010",
  45120=>"111100110",
  45121=>"010010111",
  45122=>"101011111",
  45123=>"011010000",
  45124=>"110100011",
  45125=>"111111011",
  45126=>"001110101",
  45127=>"110100110",
  45128=>"100100101",
  45129=>"010001010",
  45130=>"111100010",
  45131=>"011000000",
  45132=>"001000110",
  45133=>"110110110",
  45134=>"010110011",
  45135=>"110110011",
  45136=>"101000111",
  45137=>"100010101",
  45138=>"111100111",
  45139=>"101100000",
  45140=>"000001111",
  45141=>"111101011",
  45142=>"011011000",
  45143=>"001110001",
  45144=>"010110111",
  45145=>"011000100",
  45146=>"101110110",
  45147=>"000000101",
  45148=>"100110100",
  45149=>"011110110",
  45150=>"101010010",
  45151=>"011110110",
  45152=>"010010101",
  45153=>"111011011",
  45154=>"101111100",
  45155=>"101000010",
  45156=>"010010110",
  45157=>"011111011",
  45158=>"011111110",
  45159=>"111000000",
  45160=>"101110100",
  45161=>"110010001",
  45162=>"010010010",
  45163=>"100100110",
  45164=>"011100010",
  45165=>"000000111",
  45166=>"011111101",
  45167=>"001000111",
  45168=>"011110110",
  45169=>"001011100",
  45170=>"111101000",
  45171=>"101001011",
  45172=>"110111010",
  45173=>"010000011",
  45174=>"100110100",
  45175=>"101111111",
  45176=>"011100001",
  45177=>"100000000",
  45178=>"101101110",
  45179=>"111011011",
  45180=>"000101010",
  45181=>"100011110",
  45182=>"010000010",
  45183=>"011001000",
  45184=>"001101101",
  45185=>"101101101",
  45186=>"111100010",
  45187=>"100101111",
  45188=>"110100001",
  45189=>"000111010",
  45190=>"101001100",
  45191=>"111111100",
  45192=>"011011011",
  45193=>"001001001",
  45194=>"001010001",
  45195=>"100010110",
  45196=>"101110000",
  45197=>"101100011",
  45198=>"110100110",
  45199=>"100100110",
  45200=>"100001011",
  45201=>"010000010",
  45202=>"111110100",
  45203=>"000000100",
  45204=>"010011111",
  45205=>"111111101",
  45206=>"000000101",
  45207=>"010101000",
  45208=>"011001100",
  45209=>"000000110",
  45210=>"110010000",
  45211=>"111100101",
  45212=>"000010111",
  45213=>"101110010",
  45214=>"000010110",
  45215=>"001011011",
  45216=>"100101001",
  45217=>"101101001",
  45218=>"001111011",
  45219=>"010100111",
  45220=>"101110010",
  45221=>"010001110",
  45222=>"010101010",
  45223=>"100100100",
  45224=>"111111111",
  45225=>"001110111",
  45226=>"100101110",
  45227=>"000001011",
  45228=>"011110010",
  45229=>"110110111",
  45230=>"001110100",
  45231=>"110110100",
  45232=>"011011100",
  45233=>"001100010",
  45234=>"010001101",
  45235=>"011111001",
  45236=>"110010100",
  45237=>"010011100",
  45238=>"111010111",
  45239=>"110111111",
  45240=>"100010110",
  45241=>"010110010",
  45242=>"011011000",
  45243=>"000001000",
  45244=>"110111101",
  45245=>"011011001",
  45246=>"010010100",
  45247=>"011100110",
  45248=>"111101011",
  45249=>"111011101",
  45250=>"111001111",
  45251=>"111111001",
  45252=>"000100110",
  45253=>"000000111",
  45254=>"011001010",
  45255=>"010111011",
  45256=>"111000101",
  45257=>"001110010",
  45258=>"001001001",
  45259=>"110101101",
  45260=>"101100001",
  45261=>"010010010",
  45262=>"100001000",
  45263=>"111110100",
  45264=>"110110111",
  45265=>"001011100",
  45266=>"100001010",
  45267=>"001101001",
  45268=>"011011101",
  45269=>"100100110",
  45270=>"110101111",
  45271=>"001101001",
  45272=>"010110101",
  45273=>"000110110",
  45274=>"010110101",
  45275=>"001001000",
  45276=>"101111101",
  45277=>"000101101",
  45278=>"011110101",
  45279=>"001011001",
  45280=>"000100011",
  45281=>"111010000",
  45282=>"110101010",
  45283=>"011100110",
  45284=>"000111001",
  45285=>"111011011",
  45286=>"100000000",
  45287=>"000000100",
  45288=>"101101100",
  45289=>"111100110",
  45290=>"011111000",
  45291=>"110101001",
  45292=>"111001000",
  45293=>"011000011",
  45294=>"111001111",
  45295=>"101001000",
  45296=>"000110000",
  45297=>"001001011",
  45298=>"111010000",
  45299=>"111110001",
  45300=>"000110001",
  45301=>"000100110",
  45302=>"111000100",
  45303=>"001001001",
  45304=>"111110110",
  45305=>"110011110",
  45306=>"010110010",
  45307=>"010111111",
  45308=>"010101010",
  45309=>"101011000",
  45310=>"101011010",
  45311=>"000111011",
  45312=>"001000010",
  45313=>"100101100",
  45314=>"101010011",
  45315=>"010111100",
  45316=>"101101001",
  45317=>"111010111",
  45318=>"010101010",
  45319=>"110011101",
  45320=>"001001000",
  45321=>"000010000",
  45322=>"101001000",
  45323=>"001110111",
  45324=>"110001001",
  45325=>"110101100",
  45326=>"011111110",
  45327=>"000000000",
  45328=>"110101100",
  45329=>"111111000",
  45330=>"110001011",
  45331=>"010111100",
  45332=>"100011011",
  45333=>"111010011",
  45334=>"000100011",
  45335=>"111010001",
  45336=>"100011011",
  45337=>"000010111",
  45338=>"111010010",
  45339=>"010110000",
  45340=>"001110100",
  45341=>"011001100",
  45342=>"011111111",
  45343=>"011010000",
  45344=>"110111010",
  45345=>"111100110",
  45346=>"101000010",
  45347=>"010001011",
  45348=>"101110111",
  45349=>"110001110",
  45350=>"011000101",
  45351=>"110010100",
  45352=>"110011100",
  45353=>"010100110",
  45354=>"101011110",
  45355=>"010100110",
  45356=>"110010110",
  45357=>"101000111",
  45358=>"001100001",
  45359=>"101110000",
  45360=>"010100000",
  45361=>"000011001",
  45362=>"110100110",
  45363=>"101000011",
  45364=>"100010111",
  45365=>"100001111",
  45366=>"001001000",
  45367=>"011000011",
  45368=>"000010110",
  45369=>"100111001",
  45370=>"000110111",
  45371=>"110000011",
  45372=>"001100111",
  45373=>"100010101",
  45374=>"110000001",
  45375=>"110010000",
  45376=>"000010001",
  45377=>"011010111",
  45378=>"011111100",
  45379=>"101010010",
  45380=>"000011101",
  45381=>"011111111",
  45382=>"000110110",
  45383=>"110100100",
  45384=>"110111001",
  45385=>"010010010",
  45386=>"101111111",
  45387=>"000001001",
  45388=>"000110010",
  45389=>"001111111",
  45390=>"010010001",
  45391=>"000111000",
  45392=>"010000000",
  45393=>"010001101",
  45394=>"110111011",
  45395=>"011001010",
  45396=>"101100000",
  45397=>"001001011",
  45398=>"101000010",
  45399=>"010001000",
  45400=>"100000011",
  45401=>"011011000",
  45402=>"010110011",
  45403=>"101101000",
  45404=>"010100010",
  45405=>"010101111",
  45406=>"000001111",
  45407=>"100101100",
  45408=>"011011001",
  45409=>"010100000",
  45410=>"000011110",
  45411=>"010111011",
  45412=>"101000101",
  45413=>"011000100",
  45414=>"101110000",
  45415=>"011111100",
  45416=>"110110110",
  45417=>"101111010",
  45418=>"110111111",
  45419=>"011011000",
  45420=>"000011111",
  45421=>"101011010",
  45422=>"011100110",
  45423=>"001111111",
  45424=>"000000110",
  45425=>"110000110",
  45426=>"110100110",
  45427=>"101011101",
  45428=>"000100010",
  45429=>"001110110",
  45430=>"000001111",
  45431=>"011010010",
  45432=>"111000111",
  45433=>"001000110",
  45434=>"110011000",
  45435=>"000000010",
  45436=>"000010000",
  45437=>"111000000",
  45438=>"110011100",
  45439=>"101001000",
  45440=>"100110101",
  45441=>"000000110",
  45442=>"100100001",
  45443=>"001001101",
  45444=>"101000000",
  45445=>"100011001",
  45446=>"010011000",
  45447=>"111110111",
  45448=>"100001000",
  45449=>"111100100",
  45450=>"100101100",
  45451=>"110111111",
  45452=>"000000110",
  45453=>"011001010",
  45454=>"010001000",
  45455=>"111101001",
  45456=>"011110011",
  45457=>"000011111",
  45458=>"101101101",
  45459=>"000001010",
  45460=>"100101101",
  45461=>"001010000",
  45462=>"010101011",
  45463=>"111001010",
  45464=>"110100011",
  45465=>"010111011",
  45466=>"100100100",
  45467=>"000100001",
  45468=>"110110100",
  45469=>"111000100",
  45470=>"110001000",
  45471=>"001111010",
  45472=>"011010011",
  45473=>"001001110",
  45474=>"110000100",
  45475=>"101100111",
  45476=>"101110111",
  45477=>"110100110",
  45478=>"010101111",
  45479=>"000010010",
  45480=>"000011011",
  45481=>"000011110",
  45482=>"001000000",
  45483=>"110100100",
  45484=>"101001010",
  45485=>"011001000",
  45486=>"101100010",
  45487=>"111101100",
  45488=>"010000000",
  45489=>"001010110",
  45490=>"010101100",
  45491=>"001100011",
  45492=>"111110110",
  45493=>"111101101",
  45494=>"110100101",
  45495=>"000000111",
  45496=>"001001000",
  45497=>"100011010",
  45498=>"110001101",
  45499=>"101100111",
  45500=>"111101101",
  45501=>"111110001",
  45502=>"111010011",
  45503=>"010111101",
  45504=>"111110000",
  45505=>"010100111",
  45506=>"110011010",
  45507=>"001000000",
  45508=>"000001111",
  45509=>"001000101",
  45510=>"011101000",
  45511=>"111101001",
  45512=>"001000010",
  45513=>"101101001",
  45514=>"001001001",
  45515=>"110110111",
  45516=>"101001110",
  45517=>"101011010",
  45518=>"010011010",
  45519=>"000001100",
  45520=>"100011110",
  45521=>"111101000",
  45522=>"001111100",
  45523=>"100010001",
  45524=>"011001101",
  45525=>"011110101",
  45526=>"101101100",
  45527=>"001000100",
  45528=>"101010000",
  45529=>"001110111",
  45530=>"001101111",
  45531=>"010000000",
  45532=>"111010011",
  45533=>"100111111",
  45534=>"001100110",
  45535=>"011010011",
  45536=>"000010000",
  45537=>"110100011",
  45538=>"010110001",
  45539=>"001111000",
  45540=>"111101000",
  45541=>"111101110",
  45542=>"010110111",
  45543=>"100001111",
  45544=>"100101111",
  45545=>"110010111",
  45546=>"101101101",
  45547=>"001010110",
  45548=>"011010101",
  45549=>"111110010",
  45550=>"001011001",
  45551=>"010010000",
  45552=>"010011000",
  45553=>"010101011",
  45554=>"011101011",
  45555=>"101101100",
  45556=>"101111011",
  45557=>"100100001",
  45558=>"000110111",
  45559=>"000000111",
  45560=>"011111001",
  45561=>"111010110",
  45562=>"001000010",
  45563=>"010110111",
  45564=>"010111111",
  45565=>"000011011",
  45566=>"011000101",
  45567=>"110010011",
  45568=>"011010101",
  45569=>"100100010",
  45570=>"011100010",
  45571=>"001010110",
  45572=>"010110001",
  45573=>"101010010",
  45574=>"101111010",
  45575=>"110000000",
  45576=>"011110110",
  45577=>"111001010",
  45578=>"111000110",
  45579=>"110001010",
  45580=>"010000010",
  45581=>"010111011",
  45582=>"000110010",
  45583=>"010001110",
  45584=>"000111011",
  45585=>"111111000",
  45586=>"001100011",
  45587=>"111010110",
  45588=>"011111110",
  45589=>"010101010",
  45590=>"110111001",
  45591=>"110110111",
  45592=>"000001101",
  45593=>"011101010",
  45594=>"001100000",
  45595=>"110000110",
  45596=>"010001010",
  45597=>"100000101",
  45598=>"111000011",
  45599=>"000001110",
  45600=>"100110000",
  45601=>"010101011",
  45602=>"010100011",
  45603=>"011001001",
  45604=>"111111010",
  45605=>"001001000",
  45606=>"111111111",
  45607=>"000011111",
  45608=>"010011010",
  45609=>"000001011",
  45610=>"101111111",
  45611=>"110010101",
  45612=>"001010100",
  45613=>"001000111",
  45614=>"011000011",
  45615=>"000001110",
  45616=>"001011001",
  45617=>"011000100",
  45618=>"001100010",
  45619=>"111010110",
  45620=>"110001001",
  45621=>"000000110",
  45622=>"101011010",
  45623=>"000010000",
  45624=>"111111100",
  45625=>"011011011",
  45626=>"110001111",
  45627=>"000111101",
  45628=>"110110100",
  45629=>"101001101",
  45630=>"100011010",
  45631=>"011101000",
  45632=>"101010000",
  45633=>"101110101",
  45634=>"111000111",
  45635=>"000110100",
  45636=>"100111101",
  45637=>"101111010",
  45638=>"111011011",
  45639=>"111101110",
  45640=>"111000100",
  45641=>"001010101",
  45642=>"110101010",
  45643=>"010101111",
  45644=>"111100100",
  45645=>"001110010",
  45646=>"011010001",
  45647=>"100110111",
  45648=>"001011001",
  45649=>"000100101",
  45650=>"010100000",
  45651=>"100000000",
  45652=>"100111000",
  45653=>"011000101",
  45654=>"001101110",
  45655=>"001010110",
  45656=>"111111111",
  45657=>"001110000",
  45658=>"101100011",
  45659=>"100110010",
  45660=>"010000110",
  45661=>"101000111",
  45662=>"000011100",
  45663=>"100000000",
  45664=>"000011011",
  45665=>"111011101",
  45666=>"110111011",
  45667=>"000000010",
  45668=>"001010100",
  45669=>"101110111",
  45670=>"011001110",
  45671=>"111110110",
  45672=>"000001111",
  45673=>"110000110",
  45674=>"100101100",
  45675=>"010011000",
  45676=>"010101011",
  45677=>"110001111",
  45678=>"010011101",
  45679=>"110111100",
  45680=>"010011101",
  45681=>"111110100",
  45682=>"111000011",
  45683=>"010110101",
  45684=>"000111001",
  45685=>"110000010",
  45686=>"010011010",
  45687=>"000001000",
  45688=>"001101110",
  45689=>"110011010",
  45690=>"101011110",
  45691=>"100001110",
  45692=>"011101111",
  45693=>"011111010",
  45694=>"010110111",
  45695=>"100011000",
  45696=>"111000110",
  45697=>"100111001",
  45698=>"000110100",
  45699=>"100110011",
  45700=>"110101100",
  45701=>"100010100",
  45702=>"100010001",
  45703=>"111001110",
  45704=>"011011101",
  45705=>"011001100",
  45706=>"111101110",
  45707=>"000111011",
  45708=>"101000011",
  45709=>"100000001",
  45710=>"010101100",
  45711=>"100010001",
  45712=>"000001000",
  45713=>"110100011",
  45714=>"111001111",
  45715=>"110000101",
  45716=>"011111001",
  45717=>"101001011",
  45718=>"101110111",
  45719=>"001111000",
  45720=>"111100011",
  45721=>"110110001",
  45722=>"101011000",
  45723=>"011110101",
  45724=>"110010110",
  45725=>"110011110",
  45726=>"000001010",
  45727=>"101001101",
  45728=>"010010111",
  45729=>"010011101",
  45730=>"000111101",
  45731=>"100001011",
  45732=>"010101011",
  45733=>"100011110",
  45734=>"011001000",
  45735=>"000110001",
  45736=>"010101110",
  45737=>"000110100",
  45738=>"001011111",
  45739=>"011110000",
  45740=>"100010100",
  45741=>"001100011",
  45742=>"000111011",
  45743=>"110110000",
  45744=>"111100011",
  45745=>"011010100",
  45746=>"111000001",
  45747=>"101001010",
  45748=>"001010100",
  45749=>"000011100",
  45750=>"010001000",
  45751=>"111010101",
  45752=>"010110111",
  45753=>"110101001",
  45754=>"100000000",
  45755=>"010001001",
  45756=>"011010110",
  45757=>"110110011",
  45758=>"010011010",
  45759=>"000110011",
  45760=>"000100011",
  45761=>"100000010",
  45762=>"000100001",
  45763=>"001011101",
  45764=>"001101010",
  45765=>"101110100",
  45766=>"011001110",
  45767=>"111010101",
  45768=>"010100101",
  45769=>"100101001",
  45770=>"001110111",
  45771=>"010101110",
  45772=>"000010111",
  45773=>"000010001",
  45774=>"001101111",
  45775=>"111101101",
  45776=>"000101100",
  45777=>"101100110",
  45778=>"010000110",
  45779=>"111011010",
  45780=>"100000011",
  45781=>"011110001",
  45782=>"010110100",
  45783=>"001001110",
  45784=>"001010111",
  45785=>"011100110",
  45786=>"111011100",
  45787=>"101110110",
  45788=>"010101001",
  45789=>"011011111",
  45790=>"111011001",
  45791=>"001111111",
  45792=>"001000110",
  45793=>"111000001",
  45794=>"100000000",
  45795=>"010001101",
  45796=>"010010010",
  45797=>"101010001",
  45798=>"101010100",
  45799=>"010100110",
  45800=>"110000100",
  45801=>"010110110",
  45802=>"000111010",
  45803=>"100100110",
  45804=>"011000100",
  45805=>"110111110",
  45806=>"111101001",
  45807=>"100000000",
  45808=>"100010010",
  45809=>"001100011",
  45810=>"000100110",
  45811=>"111001110",
  45812=>"011010100",
  45813=>"010011011",
  45814=>"000100101",
  45815=>"000100101",
  45816=>"000101111",
  45817=>"000010001",
  45818=>"101000000",
  45819=>"100101110",
  45820=>"101011111",
  45821=>"011101110",
  45822=>"100110101",
  45823=>"100110011",
  45824=>"000100111",
  45825=>"011101011",
  45826=>"111000011",
  45827=>"000001000",
  45828=>"000011101",
  45829=>"101001001",
  45830=>"001100111",
  45831=>"000110111",
  45832=>"010011011",
  45833=>"100111001",
  45834=>"001101010",
  45835=>"110010001",
  45836=>"001010001",
  45837=>"100100101",
  45838=>"110011101",
  45839=>"110110100",
  45840=>"100000000",
  45841=>"000110001",
  45842=>"010111011",
  45843=>"001110101",
  45844=>"001011111",
  45845=>"111101111",
  45846=>"101101111",
  45847=>"111010101",
  45848=>"111010000",
  45849=>"000110001",
  45850=>"010111111",
  45851=>"101100010",
  45852=>"101001101",
  45853=>"000001100",
  45854=>"110000110",
  45855=>"000100000",
  45856=>"100101101",
  45857=>"001010001",
  45858=>"011001011",
  45859=>"110110001",
  45860=>"110100100",
  45861=>"001111011",
  45862=>"010111010",
  45863=>"010010011",
  45864=>"100000100",
  45865=>"000101100",
  45866=>"110010111",
  45867=>"100101101",
  45868=>"001100001",
  45869=>"100011000",
  45870=>"010000000",
  45871=>"001101100",
  45872=>"101011101",
  45873=>"001010011",
  45874=>"100000101",
  45875=>"100010110",
  45876=>"000001110",
  45877=>"100101100",
  45878=>"001001001",
  45879=>"010100001",
  45880=>"110111001",
  45881=>"100000101",
  45882=>"101011011",
  45883=>"110000101",
  45884=>"010110010",
  45885=>"011000110",
  45886=>"111111101",
  45887=>"111100000",
  45888=>"101011110",
  45889=>"111100111",
  45890=>"001101001",
  45891=>"111001001",
  45892=>"110111111",
  45893=>"000010011",
  45894=>"101101001",
  45895=>"001110110",
  45896=>"000001101",
  45897=>"100000010",
  45898=>"001000100",
  45899=>"111000000",
  45900=>"101010111",
  45901=>"000110111",
  45902=>"111001001",
  45903=>"010100110",
  45904=>"110000101",
  45905=>"001000111",
  45906=>"111110101",
  45907=>"011010001",
  45908=>"010000101",
  45909=>"100111000",
  45910=>"111010010",
  45911=>"000100100",
  45912=>"000100011",
  45913=>"001111001",
  45914=>"100101000",
  45915=>"001100100",
  45916=>"101010011",
  45917=>"010111010",
  45918=>"010000011",
  45919=>"001010010",
  45920=>"001001000",
  45921=>"000011011",
  45922=>"010010000",
  45923=>"001111111",
  45924=>"000101110",
  45925=>"010010111",
  45926=>"100101000",
  45927=>"010011001",
  45928=>"111101100",
  45929=>"010000011",
  45930=>"111000000",
  45931=>"100110011",
  45932=>"111010010",
  45933=>"011010011",
  45934=>"101100011",
  45935=>"101001100",
  45936=>"110100001",
  45937=>"001010110",
  45938=>"110110110",
  45939=>"001110110",
  45940=>"100110110",
  45941=>"110000000",
  45942=>"010101010",
  45943=>"111100000",
  45944=>"001101100",
  45945=>"100010001",
  45946=>"110001000",
  45947=>"011011001",
  45948=>"100111000",
  45949=>"111001111",
  45950=>"110011101",
  45951=>"001101001",
  45952=>"010111100",
  45953=>"001111011",
  45954=>"101000000",
  45955=>"101100101",
  45956=>"111111111",
  45957=>"011110111",
  45958=>"111011111",
  45959=>"101010010",
  45960=>"000010101",
  45961=>"111111011",
  45962=>"000111011",
  45963=>"011111100",
  45964=>"100100011",
  45965=>"000111010",
  45966=>"111100000",
  45967=>"100111001",
  45968=>"011010001",
  45969=>"000100100",
  45970=>"100001100",
  45971=>"000111000",
  45972=>"111110001",
  45973=>"111111000",
  45974=>"100000000",
  45975=>"110011001",
  45976=>"001000100",
  45977=>"101101110",
  45978=>"010010111",
  45979=>"000001100",
  45980=>"100011110",
  45981=>"010010101",
  45982=>"001011010",
  45983=>"011010111",
  45984=>"001000100",
  45985=>"010011110",
  45986=>"100000001",
  45987=>"000010110",
  45988=>"010010111",
  45989=>"011010100",
  45990=>"000110011",
  45991=>"011110110",
  45992=>"100100111",
  45993=>"110011000",
  45994=>"100100011",
  45995=>"111001000",
  45996=>"010011000",
  45997=>"100001111",
  45998=>"100001100",
  45999=>"101110110",
  46000=>"110111001",
  46001=>"111100111",
  46002=>"101011111",
  46003=>"110000001",
  46004=>"110101011",
  46005=>"111101111",
  46006=>"000111010",
  46007=>"000011000",
  46008=>"100111010",
  46009=>"101001101",
  46010=>"101111011",
  46011=>"010000101",
  46012=>"010101010",
  46013=>"011100111",
  46014=>"100101110",
  46015=>"101111000",
  46016=>"000011011",
  46017=>"001110100",
  46018=>"111111000",
  46019=>"001100111",
  46020=>"010101011",
  46021=>"010101010",
  46022=>"001011100",
  46023=>"110100010",
  46024=>"001010001",
  46025=>"000001110",
  46026=>"110010011",
  46027=>"110100101",
  46028=>"010111001",
  46029=>"111010010",
  46030=>"001101001",
  46031=>"000011000",
  46032=>"110110110",
  46033=>"110001001",
  46034=>"101111100",
  46035=>"101000111",
  46036=>"100101100",
  46037=>"000001111",
  46038=>"111110010",
  46039=>"001110010",
  46040=>"000000000",
  46041=>"000110011",
  46042=>"111101110",
  46043=>"101100101",
  46044=>"111000100",
  46045=>"011000110",
  46046=>"100001101",
  46047=>"010110100",
  46048=>"110101100",
  46049=>"110011011",
  46050=>"110100101",
  46051=>"111001011",
  46052=>"010001000",
  46053=>"010000000",
  46054=>"110011110",
  46055=>"001000010",
  46056=>"101010001",
  46057=>"100111101",
  46058=>"111101100",
  46059=>"000101101",
  46060=>"010100111",
  46061=>"110111001",
  46062=>"000010011",
  46063=>"101100111",
  46064=>"111111100",
  46065=>"111110111",
  46066=>"000100010",
  46067=>"110100001",
  46068=>"000010011",
  46069=>"001011001",
  46070=>"111010011",
  46071=>"111101001",
  46072=>"011101111",
  46073=>"101111000",
  46074=>"101101011",
  46075=>"010011110",
  46076=>"011001111",
  46077=>"111110100",
  46078=>"001111011",
  46079=>"000010010",
  46080=>"100000010",
  46081=>"101111100",
  46082=>"101011110",
  46083=>"000011111",
  46084=>"111001101",
  46085=>"111000001",
  46086=>"001101111",
  46087=>"000110011",
  46088=>"011111000",
  46089=>"001100101",
  46090=>"110101100",
  46091=>"010110110",
  46092=>"000001000",
  46093=>"000100010",
  46094=>"110011101",
  46095=>"001000111",
  46096=>"010001111",
  46097=>"101000111",
  46098=>"001001111",
  46099=>"101110100",
  46100=>"010011111",
  46101=>"100110011",
  46102=>"111110101",
  46103=>"000001101",
  46104=>"110011010",
  46105=>"111110011",
  46106=>"110010101",
  46107=>"111001110",
  46108=>"000110101",
  46109=>"000010000",
  46110=>"000010000",
  46111=>"010100000",
  46112=>"011001100",
  46113=>"000011000",
  46114=>"110010010",
  46115=>"110110000",
  46116=>"011010110",
  46117=>"000100001",
  46118=>"001101100",
  46119=>"111110011",
  46120=>"011100000",
  46121=>"001001101",
  46122=>"001100011",
  46123=>"101111001",
  46124=>"100001111",
  46125=>"011000011",
  46126=>"001011100",
  46127=>"000011000",
  46128=>"101111011",
  46129=>"011001111",
  46130=>"101011110",
  46131=>"010001010",
  46132=>"101100010",
  46133=>"000001110",
  46134=>"000101010",
  46135=>"100101110",
  46136=>"001000111",
  46137=>"011111110",
  46138=>"010110011",
  46139=>"101101100",
  46140=>"011000010",
  46141=>"001101100",
  46142=>"000100001",
  46143=>"100000101",
  46144=>"010100011",
  46145=>"111000010",
  46146=>"101001001",
  46147=>"000010000",
  46148=>"100100000",
  46149=>"010100001",
  46150=>"111100001",
  46151=>"011001110",
  46152=>"110011000",
  46153=>"000000000",
  46154=>"001010100",
  46155=>"110110010",
  46156=>"001010111",
  46157=>"100101000",
  46158=>"100000011",
  46159=>"101101100",
  46160=>"110110011",
  46161=>"000011111",
  46162=>"001111110",
  46163=>"000100011",
  46164=>"101101110",
  46165=>"111010011",
  46166=>"110110010",
  46167=>"001111101",
  46168=>"101110100",
  46169=>"101000100",
  46170=>"100010001",
  46171=>"110101001",
  46172=>"111111110",
  46173=>"100101100",
  46174=>"000001110",
  46175=>"010001100",
  46176=>"000110010",
  46177=>"000011001",
  46178=>"000110011",
  46179=>"100001000",
  46180=>"000101011",
  46181=>"111101011",
  46182=>"110111101",
  46183=>"000110011",
  46184=>"111010110",
  46185=>"110110111",
  46186=>"001010110",
  46187=>"111001000",
  46188=>"000100111",
  46189=>"100110100",
  46190=>"101011100",
  46191=>"101001011",
  46192=>"110001011",
  46193=>"000001010",
  46194=>"001011100",
  46195=>"110101010",
  46196=>"000001010",
  46197=>"000001001",
  46198=>"100010100",
  46199=>"010110111",
  46200=>"101101011",
  46201=>"110110111",
  46202=>"000011100",
  46203=>"101000100",
  46204=>"001000110",
  46205=>"101110001",
  46206=>"010011100",
  46207=>"110000111",
  46208=>"000000000",
  46209=>"001010110",
  46210=>"010110110",
  46211=>"010101110",
  46212=>"010100000",
  46213=>"010111101",
  46214=>"111111101",
  46215=>"010000010",
  46216=>"111001000",
  46217=>"010111101",
  46218=>"011001111",
  46219=>"011000001",
  46220=>"011011011",
  46221=>"001111100",
  46222=>"110111001",
  46223=>"110011010",
  46224=>"000111111",
  46225=>"111000000",
  46226=>"101001000",
  46227=>"010011110",
  46228=>"000101001",
  46229=>"110001010",
  46230=>"011111101",
  46231=>"100111110",
  46232=>"001000100",
  46233=>"001011000",
  46234=>"111101100",
  46235=>"100010000",
  46236=>"011110101",
  46237=>"011110100",
  46238=>"001101100",
  46239=>"011010110",
  46240=>"000110111",
  46241=>"111101101",
  46242=>"010101001",
  46243=>"101110101",
  46244=>"110000000",
  46245=>"110110010",
  46246=>"011100000",
  46247=>"011000011",
  46248=>"111111010",
  46249=>"010111010",
  46250=>"001101000",
  46251=>"111000100",
  46252=>"111011001",
  46253=>"010110111",
  46254=>"010000001",
  46255=>"111101101",
  46256=>"001110100",
  46257=>"110101111",
  46258=>"110111001",
  46259=>"011000001",
  46260=>"001000111",
  46261=>"010110001",
  46262=>"010110100",
  46263=>"001110110",
  46264=>"110010110",
  46265=>"000101010",
  46266=>"011011010",
  46267=>"000110000",
  46268=>"111100010",
  46269=>"100001011",
  46270=>"100011111",
  46271=>"111101101",
  46272=>"101101110",
  46273=>"110010100",
  46274=>"011101000",
  46275=>"000110111",
  46276=>"010111001",
  46277=>"011100111",
  46278=>"100001000",
  46279=>"000011000",
  46280=>"011100110",
  46281=>"100100000",
  46282=>"000010011",
  46283=>"001100100",
  46284=>"010001101",
  46285=>"100001101",
  46286=>"100111000",
  46287=>"000101110",
  46288=>"001000101",
  46289=>"001110100",
  46290=>"000100111",
  46291=>"110101001",
  46292=>"100000100",
  46293=>"001000010",
  46294=>"110001100",
  46295=>"111011110",
  46296=>"111101000",
  46297=>"110001010",
  46298=>"010001111",
  46299=>"100010110",
  46300=>"100110111",
  46301=>"101100010",
  46302=>"101000101",
  46303=>"101111010",
  46304=>"001001110",
  46305=>"111010010",
  46306=>"011011101",
  46307=>"000110100",
  46308=>"111111001",
  46309=>"001001000",
  46310=>"000011111",
  46311=>"001111011",
  46312=>"000111011",
  46313=>"100101101",
  46314=>"100010000",
  46315=>"001011001",
  46316=>"111100011",
  46317=>"111000111",
  46318=>"000101010",
  46319=>"011110010",
  46320=>"011110111",
  46321=>"100111000",
  46322=>"100101110",
  46323=>"110101100",
  46324=>"010111001",
  46325=>"000100111",
  46326=>"100000001",
  46327=>"011101110",
  46328=>"101010110",
  46329=>"000101101",
  46330=>"000110100",
  46331=>"000011000",
  46332=>"100101011",
  46333=>"111110111",
  46334=>"111111001",
  46335=>"100010010",
  46336=>"111011100",
  46337=>"010111111",
  46338=>"110110101",
  46339=>"111000111",
  46340=>"111111010",
  46341=>"100001100",
  46342=>"000011100",
  46343=>"101000000",
  46344=>"110011001",
  46345=>"010100000",
  46346=>"111101110",
  46347=>"011001110",
  46348=>"010010010",
  46349=>"001010001",
  46350=>"110100110",
  46351=>"000111101",
  46352=>"011101000",
  46353=>"001111011",
  46354=>"010101101",
  46355=>"111010111",
  46356=>"101010000",
  46357=>"111111011",
  46358=>"000011101",
  46359=>"001001000",
  46360=>"001001010",
  46361=>"000101001",
  46362=>"100110011",
  46363=>"101100110",
  46364=>"000011001",
  46365=>"100100110",
  46366=>"111000000",
  46367=>"000011010",
  46368=>"010111011",
  46369=>"110111100",
  46370=>"110001100",
  46371=>"111111011",
  46372=>"110111111",
  46373=>"110100010",
  46374=>"000100110",
  46375=>"101001010",
  46376=>"010011001",
  46377=>"100101001",
  46378=>"111100010",
  46379=>"010100101",
  46380=>"011100010",
  46381=>"001110101",
  46382=>"100000101",
  46383=>"001000101",
  46384=>"001101001",
  46385=>"101100110",
  46386=>"000110111",
  46387=>"110101000",
  46388=>"001101100",
  46389=>"001010000",
  46390=>"110110100",
  46391=>"111110010",
  46392=>"010001010",
  46393=>"111010100",
  46394=>"100101011",
  46395=>"001110001",
  46396=>"111000011",
  46397=>"100101111",
  46398=>"111100000",
  46399=>"100000111",
  46400=>"010000000",
  46401=>"011101100",
  46402=>"100101010",
  46403=>"011111010",
  46404=>"100000101",
  46405=>"111100111",
  46406=>"000101101",
  46407=>"111111111",
  46408=>"101010001",
  46409=>"001011010",
  46410=>"000011100",
  46411=>"001000000",
  46412=>"111100010",
  46413=>"111100100",
  46414=>"010101111",
  46415=>"110110101",
  46416=>"111101101",
  46417=>"010001110",
  46418=>"011011010",
  46419=>"010111111",
  46420=>"001001001",
  46421=>"001110010",
  46422=>"011001110",
  46423=>"001011010",
  46424=>"100001010",
  46425=>"001101111",
  46426=>"001010001",
  46427=>"101111001",
  46428=>"011111111",
  46429=>"101011011",
  46430=>"100000000",
  46431=>"100111000",
  46432=>"000110001",
  46433=>"011001000",
  46434=>"110101001",
  46435=>"100001110",
  46436=>"001000110",
  46437=>"101010011",
  46438=>"011110000",
  46439=>"101000101",
  46440=>"100001101",
  46441=>"000101001",
  46442=>"111011010",
  46443=>"111111010",
  46444=>"110011010",
  46445=>"001101000",
  46446=>"001000100",
  46447=>"111111010",
  46448=>"010110100",
  46449=>"011111100",
  46450=>"001001101",
  46451=>"111111000",
  46452=>"000111101",
  46453=>"010011011",
  46454=>"110101110",
  46455=>"011101100",
  46456=>"110001010",
  46457=>"100001111",
  46458=>"001111100",
  46459=>"010100010",
  46460=>"100010000",
  46461=>"010111100",
  46462=>"011000101",
  46463=>"101001001",
  46464=>"011111011",
  46465=>"000000000",
  46466=>"110011111",
  46467=>"000001111",
  46468=>"110000111",
  46469=>"010001111",
  46470=>"000010010",
  46471=>"000110100",
  46472=>"011001001",
  46473=>"100010010",
  46474=>"101000010",
  46475=>"111011100",
  46476=>"001011001",
  46477=>"000101111",
  46478=>"101010111",
  46479=>"110100001",
  46480=>"011100011",
  46481=>"100000010",
  46482=>"010100110",
  46483=>"011110110",
  46484=>"000001011",
  46485=>"110110110",
  46486=>"001011011",
  46487=>"100011011",
  46488=>"100111100",
  46489=>"010010101",
  46490=>"000101000",
  46491=>"100010000",
  46492=>"011110110",
  46493=>"000011111",
  46494=>"011100000",
  46495=>"011010011",
  46496=>"100101010",
  46497=>"010111111",
  46498=>"110101001",
  46499=>"010010110",
  46500=>"001100100",
  46501=>"001010011",
  46502=>"000111011",
  46503=>"000100111",
  46504=>"101011101",
  46505=>"001111011",
  46506=>"011001000",
  46507=>"110011001",
  46508=>"001000101",
  46509=>"100110001",
  46510=>"101001001",
  46511=>"011111000",
  46512=>"011010001",
  46513=>"000100000",
  46514=>"011110000",
  46515=>"000000101",
  46516=>"110011111",
  46517=>"000100100",
  46518=>"010110101",
  46519=>"011010010",
  46520=>"101100001",
  46521=>"111010000",
  46522=>"000110111",
  46523=>"110010011",
  46524=>"011110000",
  46525=>"001011101",
  46526=>"011010111",
  46527=>"100100100",
  46528=>"110011000",
  46529=>"010000100",
  46530=>"110010110",
  46531=>"001111110",
  46532=>"000000110",
  46533=>"000010000",
  46534=>"000000110",
  46535=>"000101010",
  46536=>"001111001",
  46537=>"001011010",
  46538=>"010101101",
  46539=>"000001011",
  46540=>"011101011",
  46541=>"011101111",
  46542=>"001000011",
  46543=>"010110001",
  46544=>"000111101",
  46545=>"010101100",
  46546=>"011101111",
  46547=>"110000001",
  46548=>"011011111",
  46549=>"000010100",
  46550=>"101001101",
  46551=>"001000100",
  46552=>"110101100",
  46553=>"101111111",
  46554=>"000010011",
  46555=>"111101010",
  46556=>"100101000",
  46557=>"010110011",
  46558=>"010101100",
  46559=>"111100000",
  46560=>"110010011",
  46561=>"100110111",
  46562=>"100001100",
  46563=>"110100010",
  46564=>"011000111",
  46565=>"011010010",
  46566=>"010001000",
  46567=>"001000011",
  46568=>"001111110",
  46569=>"000001100",
  46570=>"100110100",
  46571=>"110101111",
  46572=>"010111001",
  46573=>"001011010",
  46574=>"101001000",
  46575=>"110010101",
  46576=>"010110110",
  46577=>"010111111",
  46578=>"011100010",
  46579=>"001010010",
  46580=>"000011010",
  46581=>"000110111",
  46582=>"110101100",
  46583=>"011100110",
  46584=>"101100000",
  46585=>"111000101",
  46586=>"110001110",
  46587=>"001010010",
  46588=>"001100011",
  46589=>"101100101",
  46590=>"100101111",
  46591=>"110001110",
  46592=>"011110110",
  46593=>"001101001",
  46594=>"011110010",
  46595=>"001001101",
  46596=>"011110011",
  46597=>"101101010",
  46598=>"000111111",
  46599=>"110011001",
  46600=>"101001011",
  46601=>"000011000",
  46602=>"111111000",
  46603=>"110111010",
  46604=>"100100010",
  46605=>"101100111",
  46606=>"010011110",
  46607=>"110110101",
  46608=>"001001011",
  46609=>"101111110",
  46610=>"010101111",
  46611=>"010111011",
  46612=>"001110001",
  46613=>"001110110",
  46614=>"100111110",
  46615=>"100101000",
  46616=>"011100011",
  46617=>"001100111",
  46618=>"110000011",
  46619=>"110011011",
  46620=>"001000101",
  46621=>"101111000",
  46622=>"101101011",
  46623=>"000011111",
  46624=>"000100011",
  46625=>"001000101",
  46626=>"001000101",
  46627=>"101101110",
  46628=>"011000000",
  46629=>"100011011",
  46630=>"000010010",
  46631=>"010010011",
  46632=>"000000000",
  46633=>"011011111",
  46634=>"101010100",
  46635=>"010000001",
  46636=>"111100100",
  46637=>"110010010",
  46638=>"000000100",
  46639=>"110100100",
  46640=>"001011100",
  46641=>"010001110",
  46642=>"101010101",
  46643=>"000100000",
  46644=>"101000100",
  46645=>"000001100",
  46646=>"000100001",
  46647=>"100000110",
  46648=>"001000010",
  46649=>"101010111",
  46650=>"011110101",
  46651=>"000101011",
  46652=>"011111101",
  46653=>"100111110",
  46654=>"101010010",
  46655=>"101101001",
  46656=>"001101110",
  46657=>"101010001",
  46658=>"001001010",
  46659=>"111001010",
  46660=>"111100101",
  46661=>"101110001",
  46662=>"011111001",
  46663=>"000011010",
  46664=>"000001010",
  46665=>"101000110",
  46666=>"000110001",
  46667=>"100111000",
  46668=>"000100001",
  46669=>"001001000",
  46670=>"101111010",
  46671=>"000110110",
  46672=>"111111101",
  46673=>"000010110",
  46674=>"000100011",
  46675=>"000101011",
  46676=>"101101101",
  46677=>"110101111",
  46678=>"001011000",
  46679=>"001010010",
  46680=>"000110010",
  46681=>"010101000",
  46682=>"000101000",
  46683=>"001101101",
  46684=>"011010110",
  46685=>"000001000",
  46686=>"001100111",
  46687=>"010111001",
  46688=>"011001111",
  46689=>"001010000",
  46690=>"100001001",
  46691=>"001011101",
  46692=>"101010110",
  46693=>"011101000",
  46694=>"110011011",
  46695=>"101110000",
  46696=>"110001000",
  46697=>"000001111",
  46698=>"011100100",
  46699=>"100100000",
  46700=>"001000111",
  46701=>"110111011",
  46702=>"011011001",
  46703=>"010101111",
  46704=>"100011001",
  46705=>"101101111",
  46706=>"010000001",
  46707=>"010110001",
  46708=>"100100000",
  46709=>"100100000",
  46710=>"111001000",
  46711=>"101101110",
  46712=>"110100111",
  46713=>"110111010",
  46714=>"010100001",
  46715=>"111011011",
  46716=>"010000001",
  46717=>"001000111",
  46718=>"001001001",
  46719=>"100111010",
  46720=>"001001000",
  46721=>"000100110",
  46722=>"010001000",
  46723=>"000001101",
  46724=>"000110111",
  46725=>"100010011",
  46726=>"011101111",
  46727=>"010100110",
  46728=>"000100100",
  46729=>"110000100",
  46730=>"111111101",
  46731=>"001101110",
  46732=>"000000101",
  46733=>"111110111",
  46734=>"010000110",
  46735=>"110011000",
  46736=>"001110011",
  46737=>"000010000",
  46738=>"110011101",
  46739=>"010110010",
  46740=>"010000110",
  46741=>"100000001",
  46742=>"011100011",
  46743=>"011101100",
  46744=>"000101111",
  46745=>"110110110",
  46746=>"111101110",
  46747=>"111000010",
  46748=>"000011001",
  46749=>"110110100",
  46750=>"110110110",
  46751=>"110011000",
  46752=>"110100010",
  46753=>"000100011",
  46754=>"001000000",
  46755=>"000001010",
  46756=>"111101000",
  46757=>"111000001",
  46758=>"101111100",
  46759=>"001001000",
  46760=>"010000010",
  46761=>"010001010",
  46762=>"100001101",
  46763=>"101000001",
  46764=>"100010100",
  46765=>"000101000",
  46766=>"100011111",
  46767=>"000010100",
  46768=>"100010110",
  46769=>"010000110",
  46770=>"010010010",
  46771=>"100101001",
  46772=>"010100011",
  46773=>"100111011",
  46774=>"001010110",
  46775=>"111101001",
  46776=>"000100000",
  46777=>"101100011",
  46778=>"010110011",
  46779=>"111001000",
  46780=>"000100110",
  46781=>"010001000",
  46782=>"001001101",
  46783=>"111100110",
  46784=>"101011000",
  46785=>"001010011",
  46786=>"110101010",
  46787=>"111010011",
  46788=>"110011110",
  46789=>"010110001",
  46790=>"111110111",
  46791=>"011011110",
  46792=>"011010000",
  46793=>"010100100",
  46794=>"011000110",
  46795=>"000111000",
  46796=>"111010011",
  46797=>"101101110",
  46798=>"000001111",
  46799=>"001001000",
  46800=>"111000000",
  46801=>"011011100",
  46802=>"110010001",
  46803=>"001101110",
  46804=>"100000001",
  46805=>"011110110",
  46806=>"010100100",
  46807=>"010110001",
  46808=>"001111100",
  46809=>"011011011",
  46810=>"110001111",
  46811=>"111110011",
  46812=>"101101101",
  46813=>"010111100",
  46814=>"101111101",
  46815=>"010111111",
  46816=>"000010001",
  46817=>"000000000",
  46818=>"011111110",
  46819=>"111110001",
  46820=>"001010100",
  46821=>"111010100",
  46822=>"000101101",
  46823=>"001010011",
  46824=>"000101100",
  46825=>"001110100",
  46826=>"011111110",
  46827=>"111101100",
  46828=>"111011011",
  46829=>"001111110",
  46830=>"100111010",
  46831=>"010000110",
  46832=>"011111100",
  46833=>"100010000",
  46834=>"011000111",
  46835=>"100100111",
  46836=>"110000000",
  46837=>"011010001",
  46838=>"110010111",
  46839=>"000110110",
  46840=>"011101010",
  46841=>"011101100",
  46842=>"001011100",
  46843=>"110000010",
  46844=>"111001111",
  46845=>"110101010",
  46846=>"100001100",
  46847=>"111101011",
  46848=>"011100011",
  46849=>"110111111",
  46850=>"110101110",
  46851=>"001101011",
  46852=>"010110001",
  46853=>"101010010",
  46854=>"100101100",
  46855=>"010010111",
  46856=>"111101001",
  46857=>"100100001",
  46858=>"111000000",
  46859=>"010111100",
  46860=>"110001111",
  46861=>"111111010",
  46862=>"100100100",
  46863=>"100111010",
  46864=>"110010001",
  46865=>"000010101",
  46866=>"010100110",
  46867=>"111111100",
  46868=>"111100010",
  46869=>"110111011",
  46870=>"001101001",
  46871=>"101001011",
  46872=>"010100000",
  46873=>"101110110",
  46874=>"011111111",
  46875=>"110010101",
  46876=>"100101011",
  46877=>"000101010",
  46878=>"110000111",
  46879=>"010101011",
  46880=>"001110110",
  46881=>"110010000",
  46882=>"101000100",
  46883=>"000101000",
  46884=>"101001000",
  46885=>"110010010",
  46886=>"110111000",
  46887=>"111010001",
  46888=>"110100101",
  46889=>"001000001",
  46890=>"011101011",
  46891=>"011111101",
  46892=>"100100001",
  46893=>"110010001",
  46894=>"110110101",
  46895=>"000000011",
  46896=>"100110011",
  46897=>"011111111",
  46898=>"000011011",
  46899=>"100111110",
  46900=>"111111000",
  46901=>"111011011",
  46902=>"100011101",
  46903=>"010111111",
  46904=>"011000111",
  46905=>"111001011",
  46906=>"111001110",
  46907=>"001111100",
  46908=>"000010111",
  46909=>"101000110",
  46910=>"000100011",
  46911=>"011011111",
  46912=>"110111010",
  46913=>"000110010",
  46914=>"001100101",
  46915=>"101010101",
  46916=>"100010001",
  46917=>"111111010",
  46918=>"010001000",
  46919=>"111000010",
  46920=>"011000110",
  46921=>"110110001",
  46922=>"101001110",
  46923=>"001011011",
  46924=>"010110001",
  46925=>"010011111",
  46926=>"011111000",
  46927=>"000110011",
  46928=>"110101101",
  46929=>"000011101",
  46930=>"100011011",
  46931=>"010010001",
  46932=>"010101000",
  46933=>"010001011",
  46934=>"000110001",
  46935=>"111011011",
  46936=>"110110011",
  46937=>"101110100",
  46938=>"110111001",
  46939=>"011011010",
  46940=>"010011100",
  46941=>"100111001",
  46942=>"110111010",
  46943=>"010101001",
  46944=>"001000111",
  46945=>"110111100",
  46946=>"110000000",
  46947=>"011111101",
  46948=>"111111101",
  46949=>"100010111",
  46950=>"010001111",
  46951=>"111110110",
  46952=>"011111001",
  46953=>"110000000",
  46954=>"001010101",
  46955=>"011101100",
  46956=>"101110001",
  46957=>"010000000",
  46958=>"100100010",
  46959=>"111001101",
  46960=>"100101110",
  46961=>"001001000",
  46962=>"010100010",
  46963=>"001000001",
  46964=>"011110000",
  46965=>"000110111",
  46966=>"000111010",
  46967=>"110010100",
  46968=>"110001111",
  46969=>"111011101",
  46970=>"101110001",
  46971=>"001000000",
  46972=>"011111000",
  46973=>"011010110",
  46974=>"110111110",
  46975=>"111010110",
  46976=>"100010011",
  46977=>"000001011",
  46978=>"111010011",
  46979=>"001001001",
  46980=>"100010011",
  46981=>"011000001",
  46982=>"110000010",
  46983=>"001110000",
  46984=>"011100001",
  46985=>"110110000",
  46986=>"010100100",
  46987=>"101110010",
  46988=>"001011010",
  46989=>"011100110",
  46990=>"001101000",
  46991=>"100110010",
  46992=>"101011101",
  46993=>"111001010",
  46994=>"000001010",
  46995=>"100011110",
  46996=>"111000011",
  46997=>"110010000",
  46998=>"010110010",
  46999=>"110001000",
  47000=>"100011111",
  47001=>"001011111",
  47002=>"011011110",
  47003=>"100010010",
  47004=>"000111110",
  47005=>"111011011",
  47006=>"110110110",
  47007=>"011011011",
  47008=>"000001000",
  47009=>"010111000",
  47010=>"001101011",
  47011=>"011100010",
  47012=>"011001010",
  47013=>"110001010",
  47014=>"001111001",
  47015=>"010110100",
  47016=>"001001101",
  47017=>"111110011",
  47018=>"010100101",
  47019=>"011011000",
  47020=>"100110110",
  47021=>"001101010",
  47022=>"110011100",
  47023=>"101101001",
  47024=>"100001100",
  47025=>"111111111",
  47026=>"011100000",
  47027=>"011111110",
  47028=>"010000011",
  47029=>"011110111",
  47030=>"110001001",
  47031=>"111001111",
  47032=>"011010110",
  47033=>"101001001",
  47034=>"000001001",
  47035=>"110101101",
  47036=>"010000000",
  47037=>"010001000",
  47038=>"110000001",
  47039=>"000001000",
  47040=>"010000100",
  47041=>"001000010",
  47042=>"000010001",
  47043=>"100010110",
  47044=>"100001111",
  47045=>"110101000",
  47046=>"001000011",
  47047=>"011010111",
  47048=>"000001011",
  47049=>"010001001",
  47050=>"111100111",
  47051=>"001100101",
  47052=>"101100110",
  47053=>"000010010",
  47054=>"001001100",
  47055=>"000010100",
  47056=>"011000110",
  47057=>"111000001",
  47058=>"100010011",
  47059=>"001000001",
  47060=>"100100110",
  47061=>"000001010",
  47062=>"100011000",
  47063=>"111100010",
  47064=>"000001010",
  47065=>"100101110",
  47066=>"111110011",
  47067=>"101111101",
  47068=>"100101010",
  47069=>"111000100",
  47070=>"110000000",
  47071=>"100001110",
  47072=>"100100001",
  47073=>"101011101",
  47074=>"001001110",
  47075=>"001010001",
  47076=>"010010000",
  47077=>"110111011",
  47078=>"000111101",
  47079=>"010110010",
  47080=>"001010101",
  47081=>"011000111",
  47082=>"100011111",
  47083=>"010001110",
  47084=>"011001101",
  47085=>"001001011",
  47086=>"000010000",
  47087=>"100000000",
  47088=>"101010010",
  47089=>"001100010",
  47090=>"010101111",
  47091=>"110001100",
  47092=>"000000110",
  47093=>"000000111",
  47094=>"010001110",
  47095=>"010011100",
  47096=>"100000010",
  47097=>"111010100",
  47098=>"111000110",
  47099=>"000010001",
  47100=>"100101100",
  47101=>"011000010",
  47102=>"100110001",
  47103=>"111010111",
  47104=>"101001010",
  47105=>"011000001",
  47106=>"000000011",
  47107=>"010011010",
  47108=>"111001011",
  47109=>"000011111",
  47110=>"111000110",
  47111=>"011011001",
  47112=>"100110001",
  47113=>"111001000",
  47114=>"001111010",
  47115=>"100111010",
  47116=>"011000111",
  47117=>"000100101",
  47118=>"010101001",
  47119=>"111000001",
  47120=>"001001000",
  47121=>"010010111",
  47122=>"011000001",
  47123=>"000100111",
  47124=>"111100000",
  47125=>"011101100",
  47126=>"000001010",
  47127=>"111101010",
  47128=>"100000010",
  47129=>"101011100",
  47130=>"011001011",
  47131=>"011011111",
  47132=>"111000000",
  47133=>"100111110",
  47134=>"101000101",
  47135=>"110000000",
  47136=>"000100101",
  47137=>"111011101",
  47138=>"110101010",
  47139=>"011100111",
  47140=>"100100010",
  47141=>"100100111",
  47142=>"100100010",
  47143=>"111110101",
  47144=>"010000000",
  47145=>"110000100",
  47146=>"101110001",
  47147=>"110011000",
  47148=>"110011010",
  47149=>"111101111",
  47150=>"001111001",
  47151=>"111001000",
  47152=>"111011111",
  47153=>"010010010",
  47154=>"011110100",
  47155=>"111111110",
  47156=>"000001110",
  47157=>"000111111",
  47158=>"001110110",
  47159=>"001100110",
  47160=>"000001010",
  47161=>"010111101",
  47162=>"000001000",
  47163=>"100110111",
  47164=>"111101000",
  47165=>"111101110",
  47166=>"110101010",
  47167=>"011001111",
  47168=>"001111111",
  47169=>"000111110",
  47170=>"011101001",
  47171=>"001110101",
  47172=>"000010010",
  47173=>"010001010",
  47174=>"101100101",
  47175=>"110101100",
  47176=>"010101101",
  47177=>"001001001",
  47178=>"011101011",
  47179=>"110110000",
  47180=>"111110001",
  47181=>"101100001",
  47182=>"001011111",
  47183=>"100110001",
  47184=>"111101000",
  47185=>"110101101",
  47186=>"010111110",
  47187=>"101100011",
  47188=>"000011111",
  47189=>"110010001",
  47190=>"001010010",
  47191=>"111111101",
  47192=>"110100011",
  47193=>"001101111",
  47194=>"100111111",
  47195=>"001001100",
  47196=>"100000010",
  47197=>"010100000",
  47198=>"110111111",
  47199=>"010100101",
  47200=>"111110100",
  47201=>"111110100",
  47202=>"011000011",
  47203=>"011010000",
  47204=>"111100001",
  47205=>"000010010",
  47206=>"110001001",
  47207=>"110100000",
  47208=>"101100111",
  47209=>"110001011",
  47210=>"010111111",
  47211=>"011111110",
  47212=>"101001101",
  47213=>"100100111",
  47214=>"011101110",
  47215=>"001001000",
  47216=>"110111110",
  47217=>"100000000",
  47218=>"101011100",
  47219=>"101101010",
  47220=>"111001011",
  47221=>"110110001",
  47222=>"110011011",
  47223=>"101101100",
  47224=>"011001011",
  47225=>"111011100",
  47226=>"000000111",
  47227=>"101111111",
  47228=>"101111100",
  47229=>"010101001",
  47230=>"111111001",
  47231=>"010001100",
  47232=>"010101010",
  47233=>"001011101",
  47234=>"110011110",
  47235=>"110101111",
  47236=>"101111101",
  47237=>"110111111",
  47238=>"110100110",
  47239=>"100111111",
  47240=>"011100011",
  47241=>"101011111",
  47242=>"100010001",
  47243=>"110011110",
  47244=>"011010100",
  47245=>"111010010",
  47246=>"011010100",
  47247=>"110010111",
  47248=>"111001000",
  47249=>"000000111",
  47250=>"011111111",
  47251=>"101010001",
  47252=>"101011001",
  47253=>"000100101",
  47254=>"110011101",
  47255=>"001100100",
  47256=>"000001100",
  47257=>"101011110",
  47258=>"010111111",
  47259=>"001010110",
  47260=>"101101111",
  47261=>"100111110",
  47262=>"101000011",
  47263=>"111100000",
  47264=>"000011101",
  47265=>"110101010",
  47266=>"111000011",
  47267=>"001010111",
  47268=>"001011010",
  47269=>"011001011",
  47270=>"011111101",
  47271=>"011111100",
  47272=>"100000011",
  47273=>"111101001",
  47274=>"000110001",
  47275=>"100110111",
  47276=>"100110000",
  47277=>"111011110",
  47278=>"110111100",
  47279=>"100100010",
  47280=>"001110001",
  47281=>"000011100",
  47282=>"011111011",
  47283=>"001111001",
  47284=>"011001001",
  47285=>"000101111",
  47286=>"110001011",
  47287=>"100111011",
  47288=>"000110101",
  47289=>"101000001",
  47290=>"101011100",
  47291=>"000110110",
  47292=>"000101010",
  47293=>"110010000",
  47294=>"000111100",
  47295=>"011000110",
  47296=>"000110010",
  47297=>"001111000",
  47298=>"111010101",
  47299=>"001011001",
  47300=>"000111000",
  47301=>"110100000",
  47302=>"000001100",
  47303=>"101001001",
  47304=>"010101010",
  47305=>"011011110",
  47306=>"000100011",
  47307=>"100100110",
  47308=>"111101000",
  47309=>"100101001",
  47310=>"000001011",
  47311=>"001101111",
  47312=>"010110111",
  47313=>"110100100",
  47314=>"101000000",
  47315=>"110000111",
  47316=>"010010010",
  47317=>"011001000",
  47318=>"111001011",
  47319=>"011010001",
  47320=>"010110001",
  47321=>"000111111",
  47322=>"111000010",
  47323=>"111000110",
  47324=>"000110101",
  47325=>"110100011",
  47326=>"100110111",
  47327=>"010001010",
  47328=>"111100011",
  47329=>"101010111",
  47330=>"101001011",
  47331=>"111100001",
  47332=>"000111100",
  47333=>"111010011",
  47334=>"100010011",
  47335=>"111011111",
  47336=>"011011001",
  47337=>"100000010",
  47338=>"001011000",
  47339=>"010111110",
  47340=>"100111001",
  47341=>"111001011",
  47342=>"011110100",
  47343=>"100110110",
  47344=>"010000000",
  47345=>"011101100",
  47346=>"101011001",
  47347=>"001110001",
  47348=>"010110111",
  47349=>"001111010",
  47350=>"001110110",
  47351=>"011001010",
  47352=>"111010001",
  47353=>"011111111",
  47354=>"001000100",
  47355=>"011110000",
  47356=>"011110110",
  47357=>"101001100",
  47358=>"111110111",
  47359=>"011010111",
  47360=>"100110101",
  47361=>"100111010",
  47362=>"101100100",
  47363=>"110111111",
  47364=>"011000101",
  47365=>"010101011",
  47366=>"101001011",
  47367=>"010101001",
  47368=>"111010101",
  47369=>"000111111",
  47370=>"101000110",
  47371=>"101110100",
  47372=>"000100100",
  47373=>"001000100",
  47374=>"010001110",
  47375=>"011011010",
  47376=>"110111111",
  47377=>"110011001",
  47378=>"101000010",
  47379=>"000001110",
  47380=>"010100100",
  47381=>"111001100",
  47382=>"010111011",
  47383=>"111111111",
  47384=>"011010101",
  47385=>"100011000",
  47386=>"011010110",
  47387=>"001110111",
  47388=>"111101100",
  47389=>"111100101",
  47390=>"101000001",
  47391=>"111010010",
  47392=>"111001111",
  47393=>"111011111",
  47394=>"011111111",
  47395=>"000111001",
  47396=>"100010110",
  47397=>"101000101",
  47398=>"101101011",
  47399=>"011111010",
  47400=>"111010101",
  47401=>"110110000",
  47402=>"011111110",
  47403=>"011111111",
  47404=>"011111100",
  47405=>"110110001",
  47406=>"111010101",
  47407=>"111010111",
  47408=>"101101000",
  47409=>"011111010",
  47410=>"010000101",
  47411=>"111100111",
  47412=>"111001001",
  47413=>"101010000",
  47414=>"000000100",
  47415=>"110001110",
  47416=>"011001110",
  47417=>"110101111",
  47418=>"101001000",
  47419=>"001000111",
  47420=>"000100110",
  47421=>"111001110",
  47422=>"101100100",
  47423=>"100100010",
  47424=>"001110011",
  47425=>"010000001",
  47426=>"010110001",
  47427=>"110111100",
  47428=>"010110100",
  47429=>"011011110",
  47430=>"001111100",
  47431=>"101100100",
  47432=>"000100010",
  47433=>"000110101",
  47434=>"101000111",
  47435=>"010000011",
  47436=>"001010001",
  47437=>"011001010",
  47438=>"010110100",
  47439=>"001000111",
  47440=>"001111110",
  47441=>"011100101",
  47442=>"110100101",
  47443=>"101000011",
  47444=>"111011101",
  47445=>"001101011",
  47446=>"100101011",
  47447=>"111110010",
  47448=>"001110010",
  47449=>"010010001",
  47450=>"110100100",
  47451=>"000111000",
  47452=>"010100101",
  47453=>"011111110",
  47454=>"110011000",
  47455=>"011100110",
  47456=>"010011000",
  47457=>"101100100",
  47458=>"101000101",
  47459=>"100101001",
  47460=>"001000110",
  47461=>"000111110",
  47462=>"100000111",
  47463=>"000100110",
  47464=>"110011110",
  47465=>"111010000",
  47466=>"010101001",
  47467=>"010111001",
  47468=>"110111111",
  47469=>"101001000",
  47470=>"010110010",
  47471=>"110001000",
  47472=>"010000011",
  47473=>"111110000",
  47474=>"001001101",
  47475=>"011111110",
  47476=>"010111110",
  47477=>"000011101",
  47478=>"110011001",
  47479=>"100110100",
  47480=>"000100011",
  47481=>"100110101",
  47482=>"101000111",
  47483=>"010000101",
  47484=>"100101111",
  47485=>"011110100",
  47486=>"110011000",
  47487=>"110000101",
  47488=>"001100100",
  47489=>"110010000",
  47490=>"010010101",
  47491=>"011100111",
  47492=>"111010010",
  47493=>"100100011",
  47494=>"000011000",
  47495=>"011101010",
  47496=>"111000000",
  47497=>"000110110",
  47498=>"111110111",
  47499=>"101111111",
  47500=>"111010011",
  47501=>"111110110",
  47502=>"110110100",
  47503=>"111001011",
  47504=>"011011110",
  47505=>"001110000",
  47506=>"000011001",
  47507=>"010110001",
  47508=>"010000010",
  47509=>"111011001",
  47510=>"100101001",
  47511=>"011111000",
  47512=>"001100000",
  47513=>"000000000",
  47514=>"111010111",
  47515=>"111110000",
  47516=>"010011001",
  47517=>"101101011",
  47518=>"000000011",
  47519=>"011111010",
  47520=>"000001101",
  47521=>"111110000",
  47522=>"100110111",
  47523=>"110011011",
  47524=>"011010110",
  47525=>"100111101",
  47526=>"110111111",
  47527=>"001100100",
  47528=>"000010000",
  47529=>"110110101",
  47530=>"111000000",
  47531=>"001111101",
  47532=>"000001111",
  47533=>"111111001",
  47534=>"011100111",
  47535=>"010111111",
  47536=>"111101101",
  47537=>"000011110",
  47538=>"001010010",
  47539=>"101001001",
  47540=>"001010011",
  47541=>"111111111",
  47542=>"000010011",
  47543=>"100010011",
  47544=>"010010111",
  47545=>"101001111",
  47546=>"101010100",
  47547=>"101000111",
  47548=>"110101110",
  47549=>"000100011",
  47550=>"001110001",
  47551=>"110001110",
  47552=>"111101101",
  47553=>"100011000",
  47554=>"101111100",
  47555=>"101111100",
  47556=>"110110001",
  47557=>"110010110",
  47558=>"110010010",
  47559=>"111011011",
  47560=>"111001000",
  47561=>"110000101",
  47562=>"000001001",
  47563=>"000011000",
  47564=>"110011011",
  47565=>"000100011",
  47566=>"111100100",
  47567=>"110000101",
  47568=>"011010011",
  47569=>"100000010",
  47570=>"001010101",
  47571=>"101000010",
  47572=>"000110101",
  47573=>"000110010",
  47574=>"000001100",
  47575=>"011110001",
  47576=>"100000011",
  47577=>"111000000",
  47578=>"001010011",
  47579=>"111000110",
  47580=>"111111011",
  47581=>"000101111",
  47582=>"000001010",
  47583=>"001010010",
  47584=>"111100000",
  47585=>"100010011",
  47586=>"101001111",
  47587=>"010010001",
  47588=>"101110101",
  47589=>"011110100",
  47590=>"101001110",
  47591=>"111101111",
  47592=>"111100010",
  47593=>"101110110",
  47594=>"111100010",
  47595=>"100000010",
  47596=>"000100100",
  47597=>"111000110",
  47598=>"010111001",
  47599=>"011111111",
  47600=>"010011011",
  47601=>"011111111",
  47602=>"111010110",
  47603=>"100001011",
  47604=>"001001100",
  47605=>"001111001",
  47606=>"100010001",
  47607=>"011110100",
  47608=>"010101000",
  47609=>"010011110",
  47610=>"110110110",
  47611=>"100010101",
  47612=>"111111000",
  47613=>"111110010",
  47614=>"000001010",
  47615=>"111100010",
  47616=>"110000100",
  47617=>"010001000",
  47618=>"100010100",
  47619=>"001111100",
  47620=>"011110111",
  47621=>"100100000",
  47622=>"000000010",
  47623=>"011010100",
  47624=>"010001001",
  47625=>"100100011",
  47626=>"000101010",
  47627=>"110111111",
  47628=>"001110111",
  47629=>"101001110",
  47630=>"110011110",
  47631=>"000000110",
  47632=>"011100110",
  47633=>"100111111",
  47634=>"000101001",
  47635=>"101100101",
  47636=>"111001000",
  47637=>"001110110",
  47638=>"100101100",
  47639=>"111110001",
  47640=>"111011000",
  47641=>"001000011",
  47642=>"101001111",
  47643=>"001110000",
  47644=>"000101001",
  47645=>"111001011",
  47646=>"011101111",
  47647=>"000011101",
  47648=>"110001010",
  47649=>"111101011",
  47650=>"111000110",
  47651=>"011001110",
  47652=>"011011001",
  47653=>"001110111",
  47654=>"100111000",
  47655=>"111111011",
  47656=>"001101001",
  47657=>"011010111",
  47658=>"110101110",
  47659=>"010100111",
  47660=>"001010110",
  47661=>"101111111",
  47662=>"000110111",
  47663=>"000110111",
  47664=>"111010111",
  47665=>"011011001",
  47666=>"101000111",
  47667=>"101100000",
  47668=>"000001101",
  47669=>"110010010",
  47670=>"001001110",
  47671=>"001011101",
  47672=>"110000001",
  47673=>"111111110",
  47674=>"110010100",
  47675=>"110110101",
  47676=>"110100011",
  47677=>"011010010",
  47678=>"111100011",
  47679=>"000101010",
  47680=>"000001111",
  47681=>"101110011",
  47682=>"110001111",
  47683=>"011101100",
  47684=>"101010100",
  47685=>"001101011",
  47686=>"001001011",
  47687=>"001011011",
  47688=>"011010010",
  47689=>"111100110",
  47690=>"000000000",
  47691=>"100011011",
  47692=>"010011010",
  47693=>"001101100",
  47694=>"000111100",
  47695=>"100101000",
  47696=>"101100000",
  47697=>"100111001",
  47698=>"000110111",
  47699=>"001100100",
  47700=>"110000001",
  47701=>"100000101",
  47702=>"000111100",
  47703=>"010000000",
  47704=>"110011100",
  47705=>"010110011",
  47706=>"001001000",
  47707=>"011101010",
  47708=>"111111111",
  47709=>"011010110",
  47710=>"101100101",
  47711=>"010000011",
  47712=>"111110101",
  47713=>"101010001",
  47714=>"101011101",
  47715=>"101110101",
  47716=>"100110110",
  47717=>"111010011",
  47718=>"111111001",
  47719=>"101001111",
  47720=>"011000011",
  47721=>"111000010",
  47722=>"001111001",
  47723=>"111010100",
  47724=>"011100011",
  47725=>"010100110",
  47726=>"000000100",
  47727=>"000000001",
  47728=>"000100010",
  47729=>"101011000",
  47730=>"111100111",
  47731=>"100010111",
  47732=>"011010010",
  47733=>"010010110",
  47734=>"011110101",
  47735=>"101000111",
  47736=>"011011001",
  47737=>"111100000",
  47738=>"100110001",
  47739=>"100101111",
  47740=>"001001001",
  47741=>"110101011",
  47742=>"111101110",
  47743=>"110000011",
  47744=>"110001100",
  47745=>"010100011",
  47746=>"101100101",
  47747=>"100000111",
  47748=>"001100010",
  47749=>"000010110",
  47750=>"101100111",
  47751=>"100010010",
  47752=>"110001001",
  47753=>"110110001",
  47754=>"101000001",
  47755=>"111110010",
  47756=>"101111110",
  47757=>"011101101",
  47758=>"000111011",
  47759=>"111110101",
  47760=>"011111010",
  47761=>"100111101",
  47762=>"001111010",
  47763=>"001000001",
  47764=>"000011001",
  47765=>"011110111",
  47766=>"011101000",
  47767=>"111011110",
  47768=>"101100100",
  47769=>"111111010",
  47770=>"011100011",
  47771=>"001011011",
  47772=>"111101011",
  47773=>"000000110",
  47774=>"001111111",
  47775=>"010011101",
  47776=>"111011101",
  47777=>"111111010",
  47778=>"011110010",
  47779=>"101100010",
  47780=>"001011011",
  47781=>"100101100",
  47782=>"101010101",
  47783=>"010101000",
  47784=>"100100110",
  47785=>"010010010",
  47786=>"111011111",
  47787=>"010111100",
  47788=>"100010101",
  47789=>"100011101",
  47790=>"111001111",
  47791=>"010000101",
  47792=>"110110000",
  47793=>"111101011",
  47794=>"110111000",
  47795=>"000010000",
  47796=>"110010001",
  47797=>"100000110",
  47798=>"000010100",
  47799=>"011111100",
  47800=>"000100001",
  47801=>"000101001",
  47802=>"001000010",
  47803=>"110011101",
  47804=>"110010101",
  47805=>"001100101",
  47806=>"001100000",
  47807=>"100111000",
  47808=>"010000000",
  47809=>"011100010",
  47810=>"101001010",
  47811=>"111001111",
  47812=>"001111001",
  47813=>"111101111",
  47814=>"011111111",
  47815=>"010111010",
  47816=>"001110110",
  47817=>"000011101",
  47818=>"111100010",
  47819=>"101101001",
  47820=>"100101110",
  47821=>"100000011",
  47822=>"010001010",
  47823=>"001111010",
  47824=>"001000011",
  47825=>"101010111",
  47826=>"100100100",
  47827=>"111000010",
  47828=>"010000111",
  47829=>"111000000",
  47830=>"111000111",
  47831=>"110000001",
  47832=>"111010101",
  47833=>"010011110",
  47834=>"111111111",
  47835=>"001101010",
  47836=>"111101100",
  47837=>"110111110",
  47838=>"000100111",
  47839=>"001000110",
  47840=>"000100110",
  47841=>"101000000",
  47842=>"010110110",
  47843=>"111001111",
  47844=>"111101000",
  47845=>"000111111",
  47846=>"100110100",
  47847=>"001000110",
  47848=>"001000011",
  47849=>"010100000",
  47850=>"000011010",
  47851=>"000000010",
  47852=>"000001011",
  47853=>"100000101",
  47854=>"101111010",
  47855=>"001110110",
  47856=>"000000011",
  47857=>"110100000",
  47858=>"000000011",
  47859=>"011110110",
  47860=>"000111101",
  47861=>"110110110",
  47862=>"000101000",
  47863=>"000100101",
  47864=>"110111110",
  47865=>"010010001",
  47866=>"111001010",
  47867=>"111100111",
  47868=>"110111100",
  47869=>"111010010",
  47870=>"110101010",
  47871=>"011101100",
  47872=>"101111000",
  47873=>"010111101",
  47874=>"111111110",
  47875=>"010101110",
  47876=>"011101111",
  47877=>"110101101",
  47878=>"010001001",
  47879=>"111010000",
  47880=>"100010000",
  47881=>"011111011",
  47882=>"001001100",
  47883=>"111111000",
  47884=>"011110011",
  47885=>"110111101",
  47886=>"110110010",
  47887=>"110011110",
  47888=>"110111011",
  47889=>"101101111",
  47890=>"000001001",
  47891=>"100010010",
  47892=>"111000000",
  47893=>"010110101",
  47894=>"101101101",
  47895=>"100111010",
  47896=>"111011001",
  47897=>"001010110",
  47898=>"001111110",
  47899=>"110110111",
  47900=>"110110010",
  47901=>"111110110",
  47902=>"001101100",
  47903=>"010011111",
  47904=>"000011000",
  47905=>"100010100",
  47906=>"000110000",
  47907=>"011111100",
  47908=>"111110111",
  47909=>"110001000",
  47910=>"011010101",
  47911=>"100001110",
  47912=>"000101001",
  47913=>"110111101",
  47914=>"001010010",
  47915=>"111000000",
  47916=>"101111011",
  47917=>"000000110",
  47918=>"110010100",
  47919=>"000100100",
  47920=>"100010111",
  47921=>"010000111",
  47922=>"111110111",
  47923=>"001010111",
  47924=>"101000000",
  47925=>"110000010",
  47926=>"111111001",
  47927=>"111011110",
  47928=>"000110100",
  47929=>"111100111",
  47930=>"111001000",
  47931=>"001010000",
  47932=>"000011000",
  47933=>"111111000",
  47934=>"111011110",
  47935=>"001000000",
  47936=>"010001011",
  47937=>"011010101",
  47938=>"010100111",
  47939=>"111100100",
  47940=>"101001001",
  47941=>"001101110",
  47942=>"000110100",
  47943=>"100010001",
  47944=>"001111000",
  47945=>"100000101",
  47946=>"010110110",
  47947=>"010110001",
  47948=>"000111100",
  47949=>"100101000",
  47950=>"111100111",
  47951=>"100111000",
  47952=>"110100000",
  47953=>"111101110",
  47954=>"101101011",
  47955=>"111100000",
  47956=>"101101000",
  47957=>"111010000",
  47958=>"000111010",
  47959=>"111110101",
  47960=>"110111101",
  47961=>"100000010",
  47962=>"000110111",
  47963=>"111001101",
  47964=>"011010011",
  47965=>"101001111",
  47966=>"100001010",
  47967=>"101010000",
  47968=>"100000000",
  47969=>"010100011",
  47970=>"011000100",
  47971=>"111111101",
  47972=>"000110001",
  47973=>"110110001",
  47974=>"000010010",
  47975=>"000010001",
  47976=>"110101101",
  47977=>"111110111",
  47978=>"010011010",
  47979=>"000001001",
  47980=>"000111111",
  47981=>"101001111",
  47982=>"000111111",
  47983=>"011000111",
  47984=>"100001110",
  47985=>"101010011",
  47986=>"100010010",
  47987=>"010101001",
  47988=>"111101100",
  47989=>"001111100",
  47990=>"000001001",
  47991=>"101100110",
  47992=>"111111001",
  47993=>"001000110",
  47994=>"000010100",
  47995=>"001000111",
  47996=>"100101110",
  47997=>"111011101",
  47998=>"100000110",
  47999=>"110111000",
  48000=>"100001101",
  48001=>"110110111",
  48002=>"110101100",
  48003=>"101100100",
  48004=>"100000011",
  48005=>"100001111",
  48006=>"110101111",
  48007=>"110101011",
  48008=>"011111111",
  48009=>"000111110",
  48010=>"001110000",
  48011=>"110101101",
  48012=>"000011000",
  48013=>"111110011",
  48014=>"010000011",
  48015=>"101101101",
  48016=>"011000010",
  48017=>"001010110",
  48018=>"111000110",
  48019=>"000010100",
  48020=>"000010001",
  48021=>"100010000",
  48022=>"011001101",
  48023=>"001100110",
  48024=>"100011101",
  48025=>"001101100",
  48026=>"110000011",
  48027=>"101101111",
  48028=>"000001100",
  48029=>"101110000",
  48030=>"100011110",
  48031=>"111011001",
  48032=>"001111111",
  48033=>"000100100",
  48034=>"110001000",
  48035=>"011111111",
  48036=>"110011001",
  48037=>"010011001",
  48038=>"100111000",
  48039=>"110011000",
  48040=>"001111000",
  48041=>"111101110",
  48042=>"000101011",
  48043=>"101000000",
  48044=>"110001111",
  48045=>"001111001",
  48046=>"001101110",
  48047=>"111010110",
  48048=>"101110011",
  48049=>"111110111",
  48050=>"000100110",
  48051=>"011111101",
  48052=>"110111010",
  48053=>"101010100",
  48054=>"111110110",
  48055=>"011100111",
  48056=>"100100001",
  48057=>"111000100",
  48058=>"010001110",
  48059=>"110101001",
  48060=>"011011010",
  48061=>"000100011",
  48062=>"100000000",
  48063=>"101111111",
  48064=>"011001100",
  48065=>"000101010",
  48066=>"110010101",
  48067=>"010000101",
  48068=>"011000010",
  48069=>"101001111",
  48070=>"010100101",
  48071=>"111001011",
  48072=>"111011010",
  48073=>"010111011",
  48074=>"100000110",
  48075=>"101011100",
  48076=>"000100100",
  48077=>"111101001",
  48078=>"011001000",
  48079=>"101111100",
  48080=>"000001001",
  48081=>"101101011",
  48082=>"111010011",
  48083=>"101010000",
  48084=>"100110000",
  48085=>"110101011",
  48086=>"110010010",
  48087=>"111010110",
  48088=>"101000011",
  48089=>"000110000",
  48090=>"001111111",
  48091=>"000001001",
  48092=>"010100000",
  48093=>"100111011",
  48094=>"010111001",
  48095=>"100010100",
  48096=>"001000111",
  48097=>"001000100",
  48098=>"000101000",
  48099=>"001100010",
  48100=>"010101000",
  48101=>"110101101",
  48102=>"100110100",
  48103=>"101011101",
  48104=>"111111101",
  48105=>"001010001",
  48106=>"001001001",
  48107=>"110111100",
  48108=>"011101101",
  48109=>"001100010",
  48110=>"001111000",
  48111=>"111101001",
  48112=>"000100111",
  48113=>"110110110",
  48114=>"110000000",
  48115=>"000010010",
  48116=>"110101001",
  48117=>"111011111",
  48118=>"100111010",
  48119=>"110101100",
  48120=>"110100111",
  48121=>"101001000",
  48122=>"000111000",
  48123=>"100111001",
  48124=>"001000100",
  48125=>"010110000",
  48126=>"111001001",
  48127=>"000010110",
  48128=>"000011111",
  48129=>"010011110",
  48130=>"100001000",
  48131=>"110000000",
  48132=>"000001001",
  48133=>"100101011",
  48134=>"101111111",
  48135=>"000000101",
  48136=>"110000101",
  48137=>"011010001",
  48138=>"010110001",
  48139=>"001100000",
  48140=>"101010000",
  48141=>"000000100",
  48142=>"001011001",
  48143=>"010001111",
  48144=>"001010010",
  48145=>"100111010",
  48146=>"001000010",
  48147=>"000100111",
  48148=>"101110000",
  48149=>"101000010",
  48150=>"101000001",
  48151=>"010101101",
  48152=>"111110110",
  48153=>"001011110",
  48154=>"010110001",
  48155=>"001000000",
  48156=>"110000001",
  48157=>"000001001",
  48158=>"111011100",
  48159=>"000110100",
  48160=>"111011010",
  48161=>"011101100",
  48162=>"001010101",
  48163=>"010111011",
  48164=>"111010111",
  48165=>"001110111",
  48166=>"100011100",
  48167=>"101100000",
  48168=>"101111110",
  48169=>"101111111",
  48170=>"101101111",
  48171=>"100110111",
  48172=>"111011111",
  48173=>"101000111",
  48174=>"111000101",
  48175=>"101110011",
  48176=>"000110010",
  48177=>"010111110",
  48178=>"101111010",
  48179=>"000010001",
  48180=>"111011011",
  48181=>"010000001",
  48182=>"111011010",
  48183=>"001011111",
  48184=>"110000110",
  48185=>"011101010",
  48186=>"110010101",
  48187=>"010000010",
  48188=>"110001100",
  48189=>"001100100",
  48190=>"100110011",
  48191=>"111011011",
  48192=>"001110100",
  48193=>"011110100",
  48194=>"110000000",
  48195=>"110001001",
  48196=>"001011011",
  48197=>"100111100",
  48198=>"001101001",
  48199=>"010110100",
  48200=>"111001101",
  48201=>"110001011",
  48202=>"100101100",
  48203=>"111111010",
  48204=>"000111001",
  48205=>"011101000",
  48206=>"110010011",
  48207=>"111100000",
  48208=>"101100100",
  48209=>"111100111",
  48210=>"001111011",
  48211=>"001011010",
  48212=>"001000011",
  48213=>"001111111",
  48214=>"011101011",
  48215=>"011101100",
  48216=>"001010100",
  48217=>"110010101",
  48218=>"111001111",
  48219=>"000111110",
  48220=>"000100110",
  48221=>"001011111",
  48222=>"111100110",
  48223=>"000011110",
  48224=>"111111111",
  48225=>"101000000",
  48226=>"110100110",
  48227=>"110110000",
  48228=>"011010011",
  48229=>"011101001",
  48230=>"010110100",
  48231=>"011101010",
  48232=>"011101111",
  48233=>"000010001",
  48234=>"101111001",
  48235=>"000001001",
  48236=>"001000001",
  48237=>"110001001",
  48238=>"110001000",
  48239=>"111110101",
  48240=>"110101011",
  48241=>"101001011",
  48242=>"110111011",
  48243=>"000000001",
  48244=>"100101111",
  48245=>"111001101",
  48246=>"101010101",
  48247=>"111001000",
  48248=>"100111100",
  48249=>"110010110",
  48250=>"100000000",
  48251=>"011011000",
  48252=>"010010111",
  48253=>"111010000",
  48254=>"101000110",
  48255=>"001101000",
  48256=>"100100001",
  48257=>"110010111",
  48258=>"000001111",
  48259=>"101111101",
  48260=>"110101101",
  48261=>"000111001",
  48262=>"111001101",
  48263=>"111010011",
  48264=>"000110001",
  48265=>"101101111",
  48266=>"110000111",
  48267=>"101011000",
  48268=>"101001101",
  48269=>"010001000",
  48270=>"000011110",
  48271=>"100011100",
  48272=>"110100100",
  48273=>"111101000",
  48274=>"110110010",
  48275=>"010101111",
  48276=>"110001100",
  48277=>"111000111",
  48278=>"110101101",
  48279=>"101001101",
  48280=>"000000001",
  48281=>"000000110",
  48282=>"101110101",
  48283=>"111100110",
  48284=>"001010000",
  48285=>"100011001",
  48286=>"001001111",
  48287=>"010011101",
  48288=>"110010000",
  48289=>"000101001",
  48290=>"010100000",
  48291=>"010110111",
  48292=>"001000110",
  48293=>"111010110",
  48294=>"110100110",
  48295=>"111011100",
  48296=>"110001110",
  48297=>"001111001",
  48298=>"001000000",
  48299=>"111110000",
  48300=>"010010001",
  48301=>"100011110",
  48302=>"100110111",
  48303=>"001100110",
  48304=>"011011111",
  48305=>"010100100",
  48306=>"011000111",
  48307=>"111101100",
  48308=>"110010100",
  48309=>"111011011",
  48310=>"011001101",
  48311=>"111111101",
  48312=>"101010110",
  48313=>"111101001",
  48314=>"000100101",
  48315=>"111001001",
  48316=>"100100111",
  48317=>"101001110",
  48318=>"100000010",
  48319=>"010011101",
  48320=>"011111000",
  48321=>"011100011",
  48322=>"100000010",
  48323=>"111110001",
  48324=>"010001000",
  48325=>"111111101",
  48326=>"111001110",
  48327=>"001111000",
  48328=>"010101011",
  48329=>"011001100",
  48330=>"001101001",
  48331=>"011010101",
  48332=>"000010100",
  48333=>"101110100",
  48334=>"010011111",
  48335=>"101001111",
  48336=>"001100000",
  48337=>"101101010",
  48338=>"001101000",
  48339=>"001110000",
  48340=>"101000111",
  48341=>"010101011",
  48342=>"010010011",
  48343=>"100111110",
  48344=>"110100011",
  48345=>"000001011",
  48346=>"100101000",
  48347=>"000110010",
  48348=>"110011011",
  48349=>"001100111",
  48350=>"000110100",
  48351=>"101001100",
  48352=>"001100101",
  48353=>"101101100",
  48354=>"110000110",
  48355=>"000001100",
  48356=>"111011000",
  48357=>"100000101",
  48358=>"100110000",
  48359=>"100000000",
  48360=>"010101111",
  48361=>"000100100",
  48362=>"110111110",
  48363=>"011101110",
  48364=>"111111111",
  48365=>"100101100",
  48366=>"100101110",
  48367=>"011000000",
  48368=>"101111101",
  48369=>"100010101",
  48370=>"010001000",
  48371=>"110000111",
  48372=>"110010111",
  48373=>"100000000",
  48374=>"010001000",
  48375=>"001111110",
  48376=>"111100000",
  48377=>"111101111",
  48378=>"100110100",
  48379=>"101101100",
  48380=>"101000011",
  48381=>"110110110",
  48382=>"111100000",
  48383=>"001001100",
  48384=>"010111001",
  48385=>"111100101",
  48386=>"001101000",
  48387=>"001000000",
  48388=>"011000101",
  48389=>"111101110",
  48390=>"001001111",
  48391=>"010001001",
  48392=>"011011001",
  48393=>"011001110",
  48394=>"001111101",
  48395=>"000000001",
  48396=>"011111101",
  48397=>"000110101",
  48398=>"000011001",
  48399=>"000011100",
  48400=>"001011111",
  48401=>"101111011",
  48402=>"011100101",
  48403=>"000100100",
  48404=>"001101110",
  48405=>"100100100",
  48406=>"110100111",
  48407=>"111011111",
  48408=>"100000011",
  48409=>"110111001",
  48410=>"111101111",
  48411=>"101110001",
  48412=>"110100111",
  48413=>"010001111",
  48414=>"000000010",
  48415=>"101010011",
  48416=>"111111111",
  48417=>"111100100",
  48418=>"011101011",
  48419=>"000100010",
  48420=>"110100110",
  48421=>"100010100",
  48422=>"000110010",
  48423=>"100101011",
  48424=>"000001110",
  48425=>"011100110",
  48426=>"000110111",
  48427=>"010110101",
  48428=>"100100110",
  48429=>"110010001",
  48430=>"111011110",
  48431=>"110110000",
  48432=>"010011011",
  48433=>"001011011",
  48434=>"010111100",
  48435=>"100101010",
  48436=>"110100111",
  48437=>"010000000",
  48438=>"010011100",
  48439=>"000000111",
  48440=>"111111111",
  48441=>"001000111",
  48442=>"000000110",
  48443=>"001001110",
  48444=>"000111100",
  48445=>"011100000",
  48446=>"100111101",
  48447=>"100111001",
  48448=>"111100100",
  48449=>"101000000",
  48450=>"000000100",
  48451=>"000110010",
  48452=>"111001111",
  48453=>"000000100",
  48454=>"001101001",
  48455=>"111000111",
  48456=>"000011101",
  48457=>"010100001",
  48458=>"110001000",
  48459=>"010001110",
  48460=>"001111001",
  48461=>"100100011",
  48462=>"110101001",
  48463=>"010110011",
  48464=>"100000100",
  48465=>"001001001",
  48466=>"100110000",
  48467=>"100111001",
  48468=>"011100111",
  48469=>"100011110",
  48470=>"110001001",
  48471=>"101011001",
  48472=>"100001101",
  48473=>"010110011",
  48474=>"101011001",
  48475=>"000001100",
  48476=>"010000011",
  48477=>"111011001",
  48478=>"011111011",
  48479=>"100011100",
  48480=>"111101001",
  48481=>"110101000",
  48482=>"100101101",
  48483=>"111100100",
  48484=>"011000010",
  48485=>"111011010",
  48486=>"011000101",
  48487=>"011001000",
  48488=>"011101000",
  48489=>"010111111",
  48490=>"111001111",
  48491=>"011000110",
  48492=>"101010000",
  48493=>"000100100",
  48494=>"111111101",
  48495=>"101010101",
  48496=>"011111100",
  48497=>"101100100",
  48498=>"010011100",
  48499=>"010101111",
  48500=>"101001110",
  48501=>"010110000",
  48502=>"100000000",
  48503=>"101110100",
  48504=>"110001000",
  48505=>"111011010",
  48506=>"100111010",
  48507=>"100110111",
  48508=>"000101100",
  48509=>"011001010",
  48510=>"011100011",
  48511=>"101110110",
  48512=>"101101011",
  48513=>"111010110",
  48514=>"110111110",
  48515=>"011001100",
  48516=>"011010110",
  48517=>"111000001",
  48518=>"001011111",
  48519=>"110100001",
  48520=>"010111000",
  48521=>"111111011",
  48522=>"011000010",
  48523=>"101010011",
  48524=>"010111100",
  48525=>"010000100",
  48526=>"010100101",
  48527=>"010010001",
  48528=>"110000100",
  48529=>"101100011",
  48530=>"010000101",
  48531=>"100100111",
  48532=>"100010111",
  48533=>"111001111",
  48534=>"001100110",
  48535=>"011100110",
  48536=>"000110100",
  48537=>"011110100",
  48538=>"101000000",
  48539=>"010111110",
  48540=>"101011000",
  48541=>"000111000",
  48542=>"100000000",
  48543=>"111010010",
  48544=>"101111001",
  48545=>"111001111",
  48546=>"100000100",
  48547=>"101001111",
  48548=>"001110100",
  48549=>"110011110",
  48550=>"000000111",
  48551=>"011101011",
  48552=>"011101000",
  48553=>"000010101",
  48554=>"011011011",
  48555=>"011100111",
  48556=>"110010000",
  48557=>"010000010",
  48558=>"111010011",
  48559=>"011101101",
  48560=>"001000111",
  48561=>"010010100",
  48562=>"001101100",
  48563=>"001001111",
  48564=>"010110110",
  48565=>"011001000",
  48566=>"100000101",
  48567=>"010110111",
  48568=>"101010011",
  48569=>"001000101",
  48570=>"000000100",
  48571=>"101000011",
  48572=>"101001111",
  48573=>"010100001",
  48574=>"111110010",
  48575=>"101110010",
  48576=>"010011001",
  48577=>"110011010",
  48578=>"100110100",
  48579=>"111101010",
  48580=>"100111101",
  48581=>"100010000",
  48582=>"111100101",
  48583=>"001001001",
  48584=>"101110110",
  48585=>"100111010",
  48586=>"111111011",
  48587=>"101111001",
  48588=>"111100010",
  48589=>"011010000",
  48590=>"000010001",
  48591=>"010101100",
  48592=>"101101100",
  48593=>"111001000",
  48594=>"011011010",
  48595=>"100010011",
  48596=>"010110110",
  48597=>"010010010",
  48598=>"101101001",
  48599=>"000011000",
  48600=>"001000000",
  48601=>"001100100",
  48602=>"001010111",
  48603=>"101100001",
  48604=>"100100101",
  48605=>"110000100",
  48606=>"110110001",
  48607=>"011010011",
  48608=>"100110111",
  48609=>"001011000",
  48610=>"110100111",
  48611=>"101010001",
  48612=>"100000100",
  48613=>"111111110",
  48614=>"100100110",
  48615=>"111111010",
  48616=>"110100010",
  48617=>"010011111",
  48618=>"001011011",
  48619=>"000000000",
  48620=>"000011010",
  48621=>"011011101",
  48622=>"111100101",
  48623=>"111011011",
  48624=>"011000001",
  48625=>"010011101",
  48626=>"100000000",
  48627=>"011000001",
  48628=>"001011010",
  48629=>"010011111",
  48630=>"011010101",
  48631=>"010100110",
  48632=>"000100000",
  48633=>"011111111",
  48634=>"100111011",
  48635=>"100100110",
  48636=>"101111010",
  48637=>"000101100",
  48638=>"110111011",
  48639=>"111011100",
  48640=>"011100110",
  48641=>"010110110",
  48642=>"011101111",
  48643=>"100010010",
  48644=>"000110001",
  48645=>"101110001",
  48646=>"110011011",
  48647=>"110100110",
  48648=>"011101000",
  48649=>"111000111",
  48650=>"101111011",
  48651=>"001000000",
  48652=>"111111111",
  48653=>"111111110",
  48654=>"001011100",
  48655=>"001110011",
  48656=>"001010000",
  48657=>"100000111",
  48658=>"000000111",
  48659=>"011011011",
  48660=>"000111000",
  48661=>"110101100",
  48662=>"111111010",
  48663=>"011101001",
  48664=>"001101101",
  48665=>"110110101",
  48666=>"010111110",
  48667=>"010011000",
  48668=>"000111111",
  48669=>"001001000",
  48670=>"000000100",
  48671=>"111111110",
  48672=>"111001000",
  48673=>"101110100",
  48674=>"000011100",
  48675=>"001101001",
  48676=>"001100100",
  48677=>"111000001",
  48678=>"001011001",
  48679=>"110110001",
  48680=>"001111101",
  48681=>"000011110",
  48682=>"100110101",
  48683=>"101111111",
  48684=>"001010111",
  48685=>"011111110",
  48686=>"111111111",
  48687=>"010100101",
  48688=>"011000101",
  48689=>"001000101",
  48690=>"111111111",
  48691=>"000010110",
  48692=>"000011101",
  48693=>"011110100",
  48694=>"100001110",
  48695=>"111111011",
  48696=>"111011010",
  48697=>"111001010",
  48698=>"101010011",
  48699=>"000100110",
  48700=>"101011101",
  48701=>"101111001",
  48702=>"001110000",
  48703=>"111101110",
  48704=>"011001001",
  48705=>"111010011",
  48706=>"101000111",
  48707=>"111000100",
  48708=>"111000010",
  48709=>"000000000",
  48710=>"000010100",
  48711=>"100010101",
  48712=>"000111101",
  48713=>"111101011",
  48714=>"011111110",
  48715=>"001110000",
  48716=>"100100001",
  48717=>"000000111",
  48718=>"110010010",
  48719=>"001000101",
  48720=>"110110001",
  48721=>"111011101",
  48722=>"100001010",
  48723=>"010011101",
  48724=>"111111001",
  48725=>"011110011",
  48726=>"001000101",
  48727=>"110111001",
  48728=>"111001010",
  48729=>"000100010",
  48730=>"111011000",
  48731=>"000110101",
  48732=>"000111111",
  48733=>"000110001",
  48734=>"010010110",
  48735=>"001110010",
  48736=>"111110001",
  48737=>"011100000",
  48738=>"000101100",
  48739=>"111010001",
  48740=>"000010000",
  48741=>"111011010",
  48742=>"100101011",
  48743=>"000111110",
  48744=>"011110011",
  48745=>"010001010",
  48746=>"101100000",
  48747=>"010110000",
  48748=>"110101010",
  48749=>"110000000",
  48750=>"110101101",
  48751=>"110000110",
  48752=>"111111100",
  48753=>"000010110",
  48754=>"111011000",
  48755=>"111001110",
  48756=>"111110000",
  48757=>"001011111",
  48758=>"100100101",
  48759=>"011000100",
  48760=>"100111110",
  48761=>"111100000",
  48762=>"111111000",
  48763=>"100111010",
  48764=>"110011000",
  48765=>"010110000",
  48766=>"111101011",
  48767=>"101011010",
  48768=>"000010100",
  48769=>"110011100",
  48770=>"100100010",
  48771=>"101100010",
  48772=>"001100100",
  48773=>"100010001",
  48774=>"001001000",
  48775=>"111110100",
  48776=>"101101001",
  48777=>"001011101",
  48778=>"111100000",
  48779=>"111110000",
  48780=>"001101111",
  48781=>"000111101",
  48782=>"001011010",
  48783=>"000011110",
  48784=>"101100101",
  48785=>"101000010",
  48786=>"011110001",
  48787=>"010010011",
  48788=>"000010101",
  48789=>"111110100",
  48790=>"110110101",
  48791=>"000111110",
  48792=>"010101000",
  48793=>"001001110",
  48794=>"110111011",
  48795=>"100110000",
  48796=>"011110000",
  48797=>"111000110",
  48798=>"100111011",
  48799=>"111110100",
  48800=>"111010111",
  48801=>"111011011",
  48802=>"000111111",
  48803=>"000000001",
  48804=>"101110100",
  48805=>"100011010",
  48806=>"011011111",
  48807=>"110111111",
  48808=>"101010001",
  48809=>"000111101",
  48810=>"110100100",
  48811=>"001101001",
  48812=>"011000001",
  48813=>"011011101",
  48814=>"101110001",
  48815=>"000101100",
  48816=>"100110110",
  48817=>"000001001",
  48818=>"111010110",
  48819=>"111110011",
  48820=>"101111010",
  48821=>"000111001",
  48822=>"001110000",
  48823=>"100111000",
  48824=>"010010010",
  48825=>"000000110",
  48826=>"000001111",
  48827=>"000111111",
  48828=>"000011111",
  48829=>"011000110",
  48830=>"011101010",
  48831=>"110101101",
  48832=>"011010010",
  48833=>"100000101",
  48834=>"001101000",
  48835=>"111111110",
  48836=>"010111111",
  48837=>"010111010",
  48838=>"010101010",
  48839=>"110000011",
  48840=>"111010010",
  48841=>"001100111",
  48842=>"101001101",
  48843=>"001001010",
  48844=>"011110000",
  48845=>"000001001",
  48846=>"101110010",
  48847=>"110001000",
  48848=>"011000100",
  48849=>"011001100",
  48850=>"010110010",
  48851=>"001101111",
  48852=>"110110010",
  48853=>"011110011",
  48854=>"001111000",
  48855=>"110100001",
  48856=>"010101011",
  48857=>"101110110",
  48858=>"101101100",
  48859=>"100110110",
  48860=>"111101011",
  48861=>"111111100",
  48862=>"000111110",
  48863=>"111011001",
  48864=>"101110110",
  48865=>"001001010",
  48866=>"101001100",
  48867=>"000001011",
  48868=>"110101000",
  48869=>"011010010",
  48870=>"100011001",
  48871=>"001110000",
  48872=>"101100111",
  48873=>"011010110",
  48874=>"110101011",
  48875=>"110000101",
  48876=>"000001111",
  48877=>"110000010",
  48878=>"111111110",
  48879=>"010100111",
  48880=>"100000000",
  48881=>"110011001",
  48882=>"101100011",
  48883=>"111100011",
  48884=>"000001001",
  48885=>"001101010",
  48886=>"011111100",
  48887=>"000011011",
  48888=>"000110000",
  48889=>"010000001",
  48890=>"100010000",
  48891=>"111101110",
  48892=>"001101100",
  48893=>"111111100",
  48894=>"000000100",
  48895=>"011100110",
  48896=>"001101101",
  48897=>"101101000",
  48898=>"100000000",
  48899=>"011010101",
  48900=>"001111000",
  48901=>"000100001",
  48902=>"100101110",
  48903=>"101101001",
  48904=>"000010000",
  48905=>"101111101",
  48906=>"111111110",
  48907=>"010111110",
  48908=>"000101100",
  48909=>"110010100",
  48910=>"011001110",
  48911=>"110111001",
  48912=>"100110000",
  48913=>"011101011",
  48914=>"111010110",
  48915=>"011000010",
  48916=>"010100111",
  48917=>"000101101",
  48918=>"001000010",
  48919=>"110100011",
  48920=>"101101101",
  48921=>"000000111",
  48922=>"100010111",
  48923=>"000101111",
  48924=>"000010111",
  48925=>"011111011",
  48926=>"110110010",
  48927=>"101010001",
  48928=>"111001110",
  48929=>"001111000",
  48930=>"110001000",
  48931=>"101010010",
  48932=>"110111110",
  48933=>"111101011",
  48934=>"101010100",
  48935=>"001011000",
  48936=>"111001010",
  48937=>"111010011",
  48938=>"010010110",
  48939=>"000000001",
  48940=>"000010011",
  48941=>"000010001",
  48942=>"100010000",
  48943=>"001111011",
  48944=>"001111001",
  48945=>"001000010",
  48946=>"000001101",
  48947=>"100011010",
  48948=>"010001000",
  48949=>"101111010",
  48950=>"011111000",
  48951=>"001001111",
  48952=>"101111101",
  48953=>"111011010",
  48954=>"100100111",
  48955=>"000000110",
  48956=>"111111000",
  48957=>"100101000",
  48958=>"111000111",
  48959=>"010010001",
  48960=>"100000001",
  48961=>"101000101",
  48962=>"000000111",
  48963=>"101100101",
  48964=>"011100001",
  48965=>"000100110",
  48966=>"101111111",
  48967=>"000101100",
  48968=>"111011100",
  48969=>"100000010",
  48970=>"111010111",
  48971=>"011110011",
  48972=>"010001111",
  48973=>"101110111",
  48974=>"110000111",
  48975=>"001100010",
  48976=>"101101101",
  48977=>"111111100",
  48978=>"011100101",
  48979=>"100001111",
  48980=>"000111111",
  48981=>"111111011",
  48982=>"000100011",
  48983=>"100110110",
  48984=>"100000010",
  48985=>"110100100",
  48986=>"001100111",
  48987=>"110001011",
  48988=>"111011001",
  48989=>"011010000",
  48990=>"010000001",
  48991=>"001011100",
  48992=>"101111111",
  48993=>"110001101",
  48994=>"101000111",
  48995=>"000000010",
  48996=>"101001111",
  48997=>"010101111",
  48998=>"100111100",
  48999=>"001010001",
  49000=>"111111111",
  49001=>"100111000",
  49002=>"001001011",
  49003=>"001101111",
  49004=>"100000000",
  49005=>"000010001",
  49006=>"101110000",
  49007=>"100110001",
  49008=>"101100100",
  49009=>"001001010",
  49010=>"001001001",
  49011=>"101011010",
  49012=>"000110000",
  49013=>"011000010",
  49014=>"001111101",
  49015=>"010001001",
  49016=>"100000010",
  49017=>"011111111",
  49018=>"010001111",
  49019=>"001000000",
  49020=>"000111011",
  49021=>"111100100",
  49022=>"111000000",
  49023=>"111101011",
  49024=>"011111001",
  49025=>"000110100",
  49026=>"101110010",
  49027=>"101001010",
  49028=>"001010011",
  49029=>"101110011",
  49030=>"111110101",
  49031=>"111111111",
  49032=>"100101111",
  49033=>"101100000",
  49034=>"111000100",
  49035=>"010110011",
  49036=>"001101011",
  49037=>"111011010",
  49038=>"110100010",
  49039=>"101000110",
  49040=>"100101111",
  49041=>"010111000",
  49042=>"001100100",
  49043=>"110001011",
  49044=>"011111110",
  49045=>"100111111",
  49046=>"100000111",
  49047=>"011000111",
  49048=>"010011101",
  49049=>"100000100",
  49050=>"110101001",
  49051=>"101001111",
  49052=>"000010101",
  49053=>"100000010",
  49054=>"000000100",
  49055=>"110001111",
  49056=>"011010011",
  49057=>"001011111",
  49058=>"011101011",
  49059=>"100011011",
  49060=>"010011100",
  49061=>"101000001",
  49062=>"101001000",
  49063=>"001101001",
  49064=>"101001110",
  49065=>"110111111",
  49066=>"100111111",
  49067=>"010010111",
  49068=>"110100101",
  49069=>"110100110",
  49070=>"001111011",
  49071=>"010000000",
  49072=>"000011000",
  49073=>"111110111",
  49074=>"011101000",
  49075=>"110100110",
  49076=>"111010010",
  49077=>"001011101",
  49078=>"010001100",
  49079=>"001010000",
  49080=>"100100000",
  49081=>"100110101",
  49082=>"011001101",
  49083=>"001110001",
  49084=>"011000001",
  49085=>"010100100",
  49086=>"111011011",
  49087=>"011000110",
  49088=>"010000010",
  49089=>"001110000",
  49090=>"010001000",
  49091=>"000000110",
  49092=>"110001110",
  49093=>"001001011",
  49094=>"000100111",
  49095=>"010101100",
  49096=>"000000001",
  49097=>"111111110",
  49098=>"001110101",
  49099=>"101110110",
  49100=>"011110000",
  49101=>"111111111",
  49102=>"000100110",
  49103=>"111111010",
  49104=>"100100000",
  49105=>"100111100",
  49106=>"100101001",
  49107=>"010001100",
  49108=>"011000111",
  49109=>"110110100",
  49110=>"110111100",
  49111=>"100011110",
  49112=>"100010011",
  49113=>"111000010",
  49114=>"000000111",
  49115=>"000100100",
  49116=>"110011110",
  49117=>"000001010",
  49118=>"001010000",
  49119=>"111011010",
  49120=>"010110111",
  49121=>"110011110",
  49122=>"100110101",
  49123=>"000001110",
  49124=>"000000100",
  49125=>"101110010",
  49126=>"000100011",
  49127=>"000111001",
  49128=>"000100100",
  49129=>"001110110",
  49130=>"010001100",
  49131=>"010001010",
  49132=>"110101110",
  49133=>"010000000",
  49134=>"110000100",
  49135=>"110111101",
  49136=>"111101001",
  49137=>"010001111",
  49138=>"100000001",
  49139=>"101110111",
  49140=>"010001010",
  49141=>"001101100",
  49142=>"111110000",
  49143=>"000000010",
  49144=>"001000000",
  49145=>"001100111",
  49146=>"000100111",
  49147=>"111111100",
  49148=>"011010010",
  49149=>"000111111",
  49150=>"000111011",
  49151=>"010110001",
  49152=>"101001000",
  49153=>"100100000",
  49154=>"101111011",
  49155=>"001000101",
  49156=>"111010000",
  49157=>"111101101",
  49158=>"010111000",
  49159=>"100010101",
  49160=>"110001010",
  49161=>"010010110",
  49162=>"110110000",
  49163=>"011011111",
  49164=>"001000000",
  49165=>"001111100",
  49166=>"001111010",
  49167=>"111110100",
  49168=>"110000110",
  49169=>"110001011",
  49170=>"111010011",
  49171=>"000100000",
  49172=>"000000100",
  49173=>"110011011",
  49174=>"111001110",
  49175=>"010001111",
  49176=>"010000101",
  49177=>"110010101",
  49178=>"110100011",
  49179=>"110111010",
  49180=>"000110011",
  49181=>"001111101",
  49182=>"000001010",
  49183=>"110000011",
  49184=>"011011001",
  49185=>"001100010",
  49186=>"010110000",
  49187=>"100001011",
  49188=>"000101101",
  49189=>"101011001",
  49190=>"111100110",
  49191=>"100110111",
  49192=>"001000000",
  49193=>"100011110",
  49194=>"111000111",
  49195=>"010111100",
  49196=>"100100000",
  49197=>"010011100",
  49198=>"111000110",
  49199=>"101001000",
  49200=>"100000001",
  49201=>"101001111",
  49202=>"111110111",
  49203=>"011110111",
  49204=>"110110111",
  49205=>"110000001",
  49206=>"000010100",
  49207=>"101001010",
  49208=>"000010001",
  49209=>"001010110",
  49210=>"011000110",
  49211=>"100000110",
  49212=>"011101100",
  49213=>"001100001",
  49214=>"100111000",
  49215=>"010001100",
  49216=>"111001111",
  49217=>"000110000",
  49218=>"010000100",
  49219=>"110100010",
  49220=>"000100100",
  49221=>"001010001",
  49222=>"010100101",
  49223=>"110010001",
  49224=>"010010010",
  49225=>"110100011",
  49226=>"000001001",
  49227=>"110110100",
  49228=>"001000110",
  49229=>"010011011",
  49230=>"011011110",
  49231=>"101010101",
  49232=>"010100001",
  49233=>"000010010",
  49234=>"111010011",
  49235=>"111011101",
  49236=>"110101100",
  49237=>"000000110",
  49238=>"111100110",
  49239=>"010000010",
  49240=>"110011011",
  49241=>"100100110",
  49242=>"101010101",
  49243=>"000101101",
  49244=>"100001000",
  49245=>"010010010",
  49246=>"000111100",
  49247=>"101000111",
  49248=>"011010100",
  49249=>"010001111",
  49250=>"010000010",
  49251=>"000001111",
  49252=>"010011111",
  49253=>"000100001",
  49254=>"011000000",
  49255=>"110001111",
  49256=>"000001101",
  49257=>"000011110",
  49258=>"000100110",
  49259=>"001001010",
  49260=>"011011011",
  49261=>"011011101",
  49262=>"110101110",
  49263=>"000111010",
  49264=>"000100101",
  49265=>"010010111",
  49266=>"100011000",
  49267=>"000110110",
  49268=>"100100111",
  49269=>"111001000",
  49270=>"011010000",
  49271=>"101100010",
  49272=>"101100001",
  49273=>"110000011",
  49274=>"100111011",
  49275=>"110100000",
  49276=>"001110001",
  49277=>"000011000",
  49278=>"010101000",
  49279=>"010100010",
  49280=>"111000000",
  49281=>"110001010",
  49282=>"000010100",
  49283=>"010111101",
  49284=>"100001111",
  49285=>"011110000",
  49286=>"100010000",
  49287=>"000011000",
  49288=>"010100101",
  49289=>"000000111",
  49290=>"010001010",
  49291=>"111011010",
  49292=>"010111110",
  49293=>"010000110",
  49294=>"010110010",
  49295=>"000011101",
  49296=>"100100101",
  49297=>"110100111",
  49298=>"001010001",
  49299=>"110000110",
  49300=>"010010100",
  49301=>"100001001",
  49302=>"010010000",
  49303=>"100100011",
  49304=>"110000011",
  49305=>"000111011",
  49306=>"101011001",
  49307=>"111010111",
  49308=>"100000100",
  49309=>"111000101",
  49310=>"111001000",
  49311=>"011110100",
  49312=>"000011010",
  49313=>"110101011",
  49314=>"110010110",
  49315=>"011011000",
  49316=>"010001010",
  49317=>"011111010",
  49318=>"011011101",
  49319=>"001001001",
  49320=>"010010110",
  49321=>"110111100",
  49322=>"101010011",
  49323=>"000111001",
  49324=>"010000000",
  49325=>"001111001",
  49326=>"011011011",
  49327=>"001101001",
  49328=>"011011001",
  49329=>"110001101",
  49330=>"100001101",
  49331=>"000010101",
  49332=>"100001001",
  49333=>"001101000",
  49334=>"000111011",
  49335=>"011000011",
  49336=>"101100000",
  49337=>"010011010",
  49338=>"010111100",
  49339=>"000111110",
  49340=>"010100101",
  49341=>"001001101",
  49342=>"001101001",
  49343=>"010010000",
  49344=>"011111100",
  49345=>"010001100",
  49346=>"100010011",
  49347=>"010110010",
  49348=>"101110011",
  49349=>"000000010",
  49350=>"111001110",
  49351=>"110010111",
  49352=>"001100010",
  49353=>"100111101",
  49354=>"010110110",
  49355=>"111111010",
  49356=>"010100000",
  49357=>"100100010",
  49358=>"110101100",
  49359=>"010101000",
  49360=>"101011010",
  49361=>"101100001",
  49362=>"010001011",
  49363=>"111010111",
  49364=>"001000000",
  49365=>"100111110",
  49366=>"101001100",
  49367=>"011000010",
  49368=>"000111001",
  49369=>"001011100",
  49370=>"010000000",
  49371=>"110000000",
  49372=>"001000101",
  49373=>"101110011",
  49374=>"010100011",
  49375=>"011010010",
  49376=>"010011000",
  49377=>"100011111",
  49378=>"110101111",
  49379=>"011100011",
  49380=>"000001000",
  49381=>"101010101",
  49382=>"000000000",
  49383=>"010010111",
  49384=>"001111000",
  49385=>"110000010",
  49386=>"011100110",
  49387=>"010010100",
  49388=>"011100111",
  49389=>"100000000",
  49390=>"100011100",
  49391=>"010000001",
  49392=>"000110001",
  49393=>"010101110",
  49394=>"111111110",
  49395=>"100000100",
  49396=>"000010101",
  49397=>"000110001",
  49398=>"000000111",
  49399=>"010111010",
  49400=>"100011110",
  49401=>"100100111",
  49402=>"000110010",
  49403=>"101000001",
  49404=>"001111110",
  49405=>"010111111",
  49406=>"010010011",
  49407=>"000000010",
  49408=>"001100101",
  49409=>"000100111",
  49410=>"011101100",
  49411=>"110001110",
  49412=>"111111001",
  49413=>"001110100",
  49414=>"001101001",
  49415=>"111010111",
  49416=>"111111011",
  49417=>"101011111",
  49418=>"011111100",
  49419=>"111101100",
  49420=>"101010111",
  49421=>"100010000",
  49422=>"000111100",
  49423=>"000011000",
  49424=>"001110001",
  49425=>"100100001",
  49426=>"010100000",
  49427=>"010110001",
  49428=>"011000001",
  49429=>"100100100",
  49430=>"101001000",
  49431=>"000010110",
  49432=>"001101011",
  49433=>"011010110",
  49434=>"010101011",
  49435=>"001000100",
  49436=>"110011011",
  49437=>"000111111",
  49438=>"110111001",
  49439=>"010111110",
  49440=>"110000100",
  49441=>"001110100",
  49442=>"100010101",
  49443=>"101101101",
  49444=>"000100010",
  49445=>"101000001",
  49446=>"100110010",
  49447=>"011110011",
  49448=>"010111010",
  49449=>"001010000",
  49450=>"111111110",
  49451=>"111101101",
  49452=>"100010010",
  49453=>"011000000",
  49454=>"000100111",
  49455=>"100001110",
  49456=>"011101010",
  49457=>"111010000",
  49458=>"001100011",
  49459=>"100011001",
  49460=>"111001010",
  49461=>"010001101",
  49462=>"001100011",
  49463=>"010110011",
  49464=>"100000111",
  49465=>"101100000",
  49466=>"001101010",
  49467=>"100100011",
  49468=>"011001110",
  49469=>"010101101",
  49470=>"001000110",
  49471=>"011100000",
  49472=>"101001110",
  49473=>"000001001",
  49474=>"000010011",
  49475=>"110111111",
  49476=>"101110011",
  49477=>"101101010",
  49478=>"100101001",
  49479=>"000010011",
  49480=>"111001000",
  49481=>"111000000",
  49482=>"100010000",
  49483=>"010101100",
  49484=>"110101100",
  49485=>"100000010",
  49486=>"110010010",
  49487=>"000001111",
  49488=>"100101001",
  49489=>"011001110",
  49490=>"110010000",
  49491=>"001110010",
  49492=>"000111100",
  49493=>"111110110",
  49494=>"000000000",
  49495=>"011000000",
  49496=>"010100001",
  49497=>"101110000",
  49498=>"110111000",
  49499=>"111110100",
  49500=>"100111011",
  49501=>"011111000",
  49502=>"010101101",
  49503=>"100001011",
  49504=>"000110001",
  49505=>"010001110",
  49506=>"111001011",
  49507=>"011100001",
  49508=>"111110101",
  49509=>"100011101",
  49510=>"100000001",
  49511=>"111100010",
  49512=>"111001001",
  49513=>"111110011",
  49514=>"010001111",
  49515=>"101010111",
  49516=>"000000010",
  49517=>"111001010",
  49518=>"000100101",
  49519=>"001101111",
  49520=>"111111000",
  49521=>"111101101",
  49522=>"000100001",
  49523=>"001010001",
  49524=>"100000110",
  49525=>"111111110",
  49526=>"001111111",
  49527=>"100011001",
  49528=>"011011101",
  49529=>"100001100",
  49530=>"110000110",
  49531=>"000000101",
  49532=>"110010111",
  49533=>"001000101",
  49534=>"110100100",
  49535=>"101001100",
  49536=>"000000011",
  49537=>"100011000",
  49538=>"111001011",
  49539=>"110010001",
  49540=>"010100000",
  49541=>"110100011",
  49542=>"011110100",
  49543=>"010001101",
  49544=>"000111110",
  49545=>"001000100",
  49546=>"010110000",
  49547=>"000010010",
  49548=>"100100011",
  49549=>"111000011",
  49550=>"110010010",
  49551=>"000101110",
  49552=>"010001110",
  49553=>"100001101",
  49554=>"001100000",
  49555=>"100001010",
  49556=>"111000000",
  49557=>"001111101",
  49558=>"100001000",
  49559=>"110001011",
  49560=>"000110011",
  49561=>"011011111",
  49562=>"010111111",
  49563=>"010000011",
  49564=>"101000001",
  49565=>"000010011",
  49566=>"101101011",
  49567=>"001011101",
  49568=>"000110010",
  49569=>"101100011",
  49570=>"000110000",
  49571=>"110100111",
  49572=>"001010010",
  49573=>"100000101",
  49574=>"011101001",
  49575=>"111100011",
  49576=>"111101110",
  49577=>"100100010",
  49578=>"010000010",
  49579=>"111100111",
  49580=>"000100100",
  49581=>"110100010",
  49582=>"000101001",
  49583=>"111000000",
  49584=>"100100011",
  49585=>"000010101",
  49586=>"110100010",
  49587=>"010001111",
  49588=>"001101000",
  49589=>"101111011",
  49590=>"000111011",
  49591=>"111010111",
  49592=>"111000000",
  49593=>"001101001",
  49594=>"100100111",
  49595=>"100010001",
  49596=>"001101110",
  49597=>"111011111",
  49598=>"100001101",
  49599=>"100011110",
  49600=>"001011011",
  49601=>"100101111",
  49602=>"001100010",
  49603=>"111011001",
  49604=>"100010010",
  49605=>"011100011",
  49606=>"101111011",
  49607=>"011110100",
  49608=>"010110110",
  49609=>"110101010",
  49610=>"000000001",
  49611=>"011011111",
  49612=>"000001010",
  49613=>"010000111",
  49614=>"000101101",
  49615=>"000010010",
  49616=>"000010011",
  49617=>"101101101",
  49618=>"100111011",
  49619=>"101101010",
  49620=>"000000111",
  49621=>"010010000",
  49622=>"010110011",
  49623=>"010110010",
  49624=>"010010011",
  49625=>"000000100",
  49626=>"101000000",
  49627=>"100011000",
  49628=>"011011111",
  49629=>"001000001",
  49630=>"110101111",
  49631=>"111000101",
  49632=>"011110100",
  49633=>"110100101",
  49634=>"010011111",
  49635=>"011110000",
  49636=>"001001111",
  49637=>"111001010",
  49638=>"010011110",
  49639=>"001000010",
  49640=>"110110101",
  49641=>"111010110",
  49642=>"011111101",
  49643=>"000000101",
  49644=>"010101001",
  49645=>"011000000",
  49646=>"001000111",
  49647=>"011111011",
  49648=>"100100011",
  49649=>"100000011",
  49650=>"111010001",
  49651=>"101110001",
  49652=>"000000000",
  49653=>"000011000",
  49654=>"101100011",
  49655=>"110001001",
  49656=>"100011110",
  49657=>"000001001",
  49658=>"110000010",
  49659=>"000111000",
  49660=>"101100010",
  49661=>"101111001",
  49662=>"011011011",
  49663=>"011001100",
  49664=>"001101101",
  49665=>"001000110",
  49666=>"001100001",
  49667=>"000011000",
  49668=>"000111010",
  49669=>"111111100",
  49670=>"011011010",
  49671=>"011110001",
  49672=>"011001110",
  49673=>"101010111",
  49674=>"011100110",
  49675=>"000000010",
  49676=>"100001000",
  49677=>"011001101",
  49678=>"001000110",
  49679=>"101000000",
  49680=>"010010000",
  49681=>"101101111",
  49682=>"110001110",
  49683=>"101000010",
  49684=>"010111000",
  49685=>"000011010",
  49686=>"010010111",
  49687=>"100110001",
  49688=>"101011011",
  49689=>"000100111",
  49690=>"001101000",
  49691=>"000000111",
  49692=>"001101010",
  49693=>"111110011",
  49694=>"101000011",
  49695=>"011011110",
  49696=>"100111101",
  49697=>"101111110",
  49698=>"111010110",
  49699=>"000100000",
  49700=>"110010100",
  49701=>"111101111",
  49702=>"110000010",
  49703=>"100110001",
  49704=>"000111001",
  49705=>"100001101",
  49706=>"111010100",
  49707=>"011001010",
  49708=>"100101101",
  49709=>"100100001",
  49710=>"101110111",
  49711=>"111011101",
  49712=>"000001000",
  49713=>"101010111",
  49714=>"010011110",
  49715=>"000011111",
  49716=>"100101110",
  49717=>"101001010",
  49718=>"111011101",
  49719=>"101011001",
  49720=>"100011000",
  49721=>"101000110",
  49722=>"111101011",
  49723=>"010110111",
  49724=>"011010001",
  49725=>"110010000",
  49726=>"000110110",
  49727=>"011101000",
  49728=>"111011111",
  49729=>"001000101",
  49730=>"001010010",
  49731=>"001110000",
  49732=>"000001010",
  49733=>"011000000",
  49734=>"111011011",
  49735=>"101100000",
  49736=>"010111000",
  49737=>"000100111",
  49738=>"101011001",
  49739=>"001010101",
  49740=>"111100011",
  49741=>"001101001",
  49742=>"100101101",
  49743=>"011100101",
  49744=>"101100100",
  49745=>"110011100",
  49746=>"101000001",
  49747=>"111010010",
  49748=>"001010100",
  49749=>"100110110",
  49750=>"110010000",
  49751=>"011110000",
  49752=>"111101001",
  49753=>"111101011",
  49754=>"111110110",
  49755=>"110001110",
  49756=>"011110100",
  49757=>"011000111",
  49758=>"011000000",
  49759=>"000000101",
  49760=>"101110110",
  49761=>"010110110",
  49762=>"011111100",
  49763=>"111001001",
  49764=>"001111100",
  49765=>"001101011",
  49766=>"111010101",
  49767=>"100110000",
  49768=>"101111101",
  49769=>"000101000",
  49770=>"101111111",
  49771=>"100111110",
  49772=>"000111101",
  49773=>"111001111",
  49774=>"111000110",
  49775=>"010011110",
  49776=>"010101000",
  49777=>"011001110",
  49778=>"001000010",
  49779=>"101101011",
  49780=>"111111101",
  49781=>"100110111",
  49782=>"111010000",
  49783=>"110101001",
  49784=>"111010001",
  49785=>"100100001",
  49786=>"110111001",
  49787=>"010100111",
  49788=>"100100010",
  49789=>"001010111",
  49790=>"000000000",
  49791=>"101010110",
  49792=>"101010100",
  49793=>"010000010",
  49794=>"001101111",
  49795=>"100101001",
  49796=>"001011010",
  49797=>"000100101",
  49798=>"000010010",
  49799=>"101110011",
  49800=>"111111000",
  49801=>"100001010",
  49802=>"100011100",
  49803=>"111101000",
  49804=>"101110101",
  49805=>"000000000",
  49806=>"111010011",
  49807=>"000101001",
  49808=>"001010100",
  49809=>"001101000",
  49810=>"111110101",
  49811=>"001010111",
  49812=>"000001100",
  49813=>"010101101",
  49814=>"011110111",
  49815=>"111111000",
  49816=>"110101000",
  49817=>"111111111",
  49818=>"001010011",
  49819=>"011011100",
  49820=>"110001010",
  49821=>"101111011",
  49822=>"100100001",
  49823=>"000010010",
  49824=>"000001011",
  49825=>"010100010",
  49826=>"010011110",
  49827=>"101100010",
  49828=>"100001001",
  49829=>"010101011",
  49830=>"100001100",
  49831=>"001000000",
  49832=>"111001101",
  49833=>"111001111",
  49834=>"101100100",
  49835=>"110010011",
  49836=>"101011000",
  49837=>"010001011",
  49838=>"110000111",
  49839=>"100010110",
  49840=>"000101010",
  49841=>"110101001",
  49842=>"101011101",
  49843=>"100111011",
  49844=>"110010010",
  49845=>"101111011",
  49846=>"110010010",
  49847=>"000100000",
  49848=>"110001101",
  49849=>"110010001",
  49850=>"100101100",
  49851=>"011000101",
  49852=>"111010010",
  49853=>"010001000",
  49854=>"010010000",
  49855=>"010010000",
  49856=>"111000001",
  49857=>"001100111",
  49858=>"011111110",
  49859=>"001010000",
  49860=>"111011100",
  49861=>"001101010",
  49862=>"110011100",
  49863=>"100000011",
  49864=>"010010000",
  49865=>"110001001",
  49866=>"101111000",
  49867=>"000011010",
  49868=>"111010011",
  49869=>"001111001",
  49870=>"010111110",
  49871=>"001011001",
  49872=>"101000011",
  49873=>"010011000",
  49874=>"000000011",
  49875=>"011001111",
  49876=>"111100001",
  49877=>"010010011",
  49878=>"101101000",
  49879=>"100100110",
  49880=>"101111010",
  49881=>"111001100",
  49882=>"100100010",
  49883=>"100100110",
  49884=>"100101110",
  49885=>"110110011",
  49886=>"111000100",
  49887=>"010010101",
  49888=>"001010110",
  49889=>"110100000",
  49890=>"000100101",
  49891=>"000000110",
  49892=>"011010111",
  49893=>"000010101",
  49894=>"100100010",
  49895=>"101011001",
  49896=>"110001100",
  49897=>"001001001",
  49898=>"000101000",
  49899=>"110100010",
  49900=>"110100000",
  49901=>"000110110",
  49902=>"101000111",
  49903=>"011001101",
  49904=>"110000110",
  49905=>"010011011",
  49906=>"100001000",
  49907=>"110100110",
  49908=>"110010001",
  49909=>"100001111",
  49910=>"111111110",
  49911=>"000001000",
  49912=>"110101101",
  49913=>"110000111",
  49914=>"111010010",
  49915=>"100000000",
  49916=>"100100110",
  49917=>"100110111",
  49918=>"111000110",
  49919=>"011010100",
  49920=>"001101101",
  49921=>"010100000",
  49922=>"110100111",
  49923=>"110011101",
  49924=>"100000110",
  49925=>"100010110",
  49926=>"101110111",
  49927=>"010111010",
  49928=>"001100011",
  49929=>"101101011",
  49930=>"100110001",
  49931=>"000001010",
  49932=>"001010010",
  49933=>"101000111",
  49934=>"101001100",
  49935=>"110110110",
  49936=>"101000000",
  49937=>"000010000",
  49938=>"001011010",
  49939=>"100101101",
  49940=>"100011001",
  49941=>"001001001",
  49942=>"111111000",
  49943=>"111110111",
  49944=>"010010010",
  49945=>"111001110",
  49946=>"000110000",
  49947=>"001001111",
  49948=>"001100111",
  49949=>"010100000",
  49950=>"000000001",
  49951=>"110001001",
  49952=>"011100011",
  49953=>"101110010",
  49954=>"011010111",
  49955=>"011001101",
  49956=>"001111001",
  49957=>"100111000",
  49958=>"100000101",
  49959=>"101000001",
  49960=>"010101001",
  49961=>"110010110",
  49962=>"010000111",
  49963=>"101100001",
  49964=>"000101111",
  49965=>"110010111",
  49966=>"010110011",
  49967=>"101000111",
  49968=>"010010010",
  49969=>"110110001",
  49970=>"110000010",
  49971=>"111010111",
  49972=>"101010011",
  49973=>"011000101",
  49974=>"001000101",
  49975=>"011010111",
  49976=>"100000000",
  49977=>"000110010",
  49978=>"000010010",
  49979=>"010000011",
  49980=>"010100100",
  49981=>"111000100",
  49982=>"100101100",
  49983=>"010010001",
  49984=>"110111110",
  49985=>"111101010",
  49986=>"010100101",
  49987=>"100001001",
  49988=>"010000100",
  49989=>"101100100",
  49990=>"011000010",
  49991=>"000100100",
  49992=>"101101101",
  49993=>"010101000",
  49994=>"111011110",
  49995=>"101001110",
  49996=>"110111001",
  49997=>"010011011",
  49998=>"010011011",
  49999=>"111110011",
  50000=>"010100010",
  50001=>"111101110",
  50002=>"110010011",
  50003=>"010010110",
  50004=>"011010001",
  50005=>"101101010",
  50006=>"011101100",
  50007=>"101010111",
  50008=>"010011011",
  50009=>"010110110",
  50010=>"111001010",
  50011=>"101101111",
  50012=>"100011011",
  50013=>"110101100",
  50014=>"011001001",
  50015=>"010100000",
  50016=>"111000101",
  50017=>"011101010",
  50018=>"010100000",
  50019=>"100011100",
  50020=>"011100100",
  50021=>"110110010",
  50022=>"101001001",
  50023=>"001101010",
  50024=>"000111011",
  50025=>"001110011",
  50026=>"111001111",
  50027=>"111110011",
  50028=>"101101000",
  50029=>"000010010",
  50030=>"011000100",
  50031=>"100110111",
  50032=>"000110010",
  50033=>"100101000",
  50034=>"100101010",
  50035=>"000010011",
  50036=>"110000010",
  50037=>"001000100",
  50038=>"000100110",
  50039=>"100110111",
  50040=>"101001011",
  50041=>"111110101",
  50042=>"000010110",
  50043=>"101100000",
  50044=>"000000000",
  50045=>"101001110",
  50046=>"000100010",
  50047=>"111111111",
  50048=>"011001010",
  50049=>"101011011",
  50050=>"100111111",
  50051=>"000011000",
  50052=>"010000010",
  50053=>"111101000",
  50054=>"001100000",
  50055=>"011000001",
  50056=>"110111000",
  50057=>"111001011",
  50058=>"101000110",
  50059=>"011101111",
  50060=>"100000110",
  50061=>"110000001",
  50062=>"000111100",
  50063=>"100010001",
  50064=>"010011100",
  50065=>"101010111",
  50066=>"111010000",
  50067=>"100011110",
  50068=>"000001011",
  50069=>"010001000",
  50070=>"010001010",
  50071=>"000111100",
  50072=>"011000001",
  50073=>"000100000",
  50074=>"011111001",
  50075=>"011011011",
  50076=>"101000111",
  50077=>"100000110",
  50078=>"011111100",
  50079=>"110010101",
  50080=>"011111100",
  50081=>"110001001",
  50082=>"110001000",
  50083=>"101011100",
  50084=>"000001000",
  50085=>"000000000",
  50086=>"101010000",
  50087=>"111010000",
  50088=>"111100100",
  50089=>"100101111",
  50090=>"101001000",
  50091=>"011100010",
  50092=>"000101001",
  50093=>"111101110",
  50094=>"010100011",
  50095=>"011110010",
  50096=>"110101000",
  50097=>"011011101",
  50098=>"000011101",
  50099=>"100101101",
  50100=>"101001111",
  50101=>"011110001",
  50102=>"111110100",
  50103=>"100001100",
  50104=>"001100110",
  50105=>"100101010",
  50106=>"111110000",
  50107=>"111101011",
  50108=>"110001000",
  50109=>"011101100",
  50110=>"100010100",
  50111=>"010010110",
  50112=>"010001010",
  50113=>"000100000",
  50114=>"011101100",
  50115=>"011010110",
  50116=>"000100001",
  50117=>"110000110",
  50118=>"110111001",
  50119=>"001001101",
  50120=>"011100011",
  50121=>"000111101",
  50122=>"100110001",
  50123=>"011110010",
  50124=>"010100010",
  50125=>"011000011",
  50126=>"100000001",
  50127=>"111001000",
  50128=>"100011111",
  50129=>"010011100",
  50130=>"010110100",
  50131=>"010001000",
  50132=>"000000111",
  50133=>"111000101",
  50134=>"001110001",
  50135=>"010101111",
  50136=>"100111100",
  50137=>"000101101",
  50138=>"010110001",
  50139=>"110110111",
  50140=>"110010111",
  50141=>"011000111",
  50142=>"110110111",
  50143=>"010011011",
  50144=>"011101111",
  50145=>"001101010",
  50146=>"000011110",
  50147=>"010101100",
  50148=>"000010110",
  50149=>"011100111",
  50150=>"100010010",
  50151=>"000000001",
  50152=>"000110100",
  50153=>"100100000",
  50154=>"110110000",
  50155=>"010001111",
  50156=>"011110100",
  50157=>"010000101",
  50158=>"110000001",
  50159=>"011110011",
  50160=>"010111000",
  50161=>"001010101",
  50162=>"100011001",
  50163=>"010100100",
  50164=>"111001100",
  50165=>"100011000",
  50166=>"001111000",
  50167=>"000000010",
  50168=>"110011101",
  50169=>"011010011",
  50170=>"100101000",
  50171=>"001100100",
  50172=>"000100100",
  50173=>"011001100",
  50174=>"100111101",
  50175=>"001101001",
  50176=>"000001001",
  50177=>"111000101",
  50178=>"000000011",
  50179=>"101100010",
  50180=>"011011010",
  50181=>"000011111",
  50182=>"101001010",
  50183=>"000001000",
  50184=>"110110010",
  50185=>"101110100",
  50186=>"101110100",
  50187=>"111100101",
  50188=>"010001001",
  50189=>"000011010",
  50190=>"011101101",
  50191=>"100000111",
  50192=>"110101100",
  50193=>"010101101",
  50194=>"011001000",
  50195=>"101111101",
  50196=>"010001010",
  50197=>"100000001",
  50198=>"010010111",
  50199=>"010001011",
  50200=>"011001010",
  50201=>"101001000",
  50202=>"100011010",
  50203=>"001000101",
  50204=>"101010000",
  50205=>"111100111",
  50206=>"101000110",
  50207=>"000001111",
  50208=>"111000001",
  50209=>"001011010",
  50210=>"011010001",
  50211=>"011010000",
  50212=>"101101011",
  50213=>"111011001",
  50214=>"111111001",
  50215=>"111101111",
  50216=>"100001001",
  50217=>"101000111",
  50218=>"011100110",
  50219=>"000111101",
  50220=>"100111111",
  50221=>"110110110",
  50222=>"101010110",
  50223=>"110000101",
  50224=>"111010000",
  50225=>"011000011",
  50226=>"110100001",
  50227=>"100111010",
  50228=>"110100111",
  50229=>"111000010",
  50230=>"100100100",
  50231=>"111001100",
  50232=>"111111010",
  50233=>"100011110",
  50234=>"100000100",
  50235=>"010010000",
  50236=>"100010000",
  50237=>"111010011",
  50238=>"100100001",
  50239=>"010011011",
  50240=>"111010110",
  50241=>"001010010",
  50242=>"001000110",
  50243=>"100011001",
  50244=>"100101011",
  50245=>"110101100",
  50246=>"011000110",
  50247=>"000100011",
  50248=>"000010100",
  50249=>"001101010",
  50250=>"010100100",
  50251=>"000110000",
  50252=>"011001001",
  50253=>"110110001",
  50254=>"101000010",
  50255=>"111100100",
  50256=>"101001100",
  50257=>"010111001",
  50258=>"011010110",
  50259=>"001010011",
  50260=>"110010100",
  50261=>"100001111",
  50262=>"010010001",
  50263=>"111010110",
  50264=>"101010010",
  50265=>"000101111",
  50266=>"001100111",
  50267=>"000101110",
  50268=>"100001000",
  50269=>"010110111",
  50270=>"010001110",
  50271=>"001101100",
  50272=>"010110101",
  50273=>"001011111",
  50274=>"001000000",
  50275=>"100100000",
  50276=>"001010011",
  50277=>"100000111",
  50278=>"111011111",
  50279=>"010101011",
  50280=>"000000111",
  50281=>"011011010",
  50282=>"110110100",
  50283=>"111110001",
  50284=>"110111010",
  50285=>"110011011",
  50286=>"010011011",
  50287=>"000111101",
  50288=>"010110010",
  50289=>"110101011",
  50290=>"110101110",
  50291=>"101011110",
  50292=>"011111100",
  50293=>"111111001",
  50294=>"100011001",
  50295=>"111100000",
  50296=>"010001010",
  50297=>"101111001",
  50298=>"001101010",
  50299=>"000111011",
  50300=>"001011101",
  50301=>"110010000",
  50302=>"110011001",
  50303=>"011011110",
  50304=>"110001000",
  50305=>"011111010",
  50306=>"011110011",
  50307=>"001100011",
  50308=>"110001100",
  50309=>"111111111",
  50310=>"101100101",
  50311=>"001110111",
  50312=>"110011111",
  50313=>"110010110",
  50314=>"100000000",
  50315=>"010100001",
  50316=>"100010001",
  50317=>"011110111",
  50318=>"010111010",
  50319=>"110001101",
  50320=>"101011001",
  50321=>"000011000",
  50322=>"011000011",
  50323=>"000111000",
  50324=>"001101100",
  50325=>"011110111",
  50326=>"000101000",
  50327=>"100000101",
  50328=>"010001110",
  50329=>"011101001",
  50330=>"101000101",
  50331=>"011101111",
  50332=>"001010111",
  50333=>"100001100",
  50334=>"010010011",
  50335=>"110011011",
  50336=>"010001111",
  50337=>"010010100",
  50338=>"100101100",
  50339=>"010001000",
  50340=>"010001101",
  50341=>"101000011",
  50342=>"101011011",
  50343=>"000010100",
  50344=>"011111110",
  50345=>"011110111",
  50346=>"101000000",
  50347=>"110101101",
  50348=>"010101001",
  50349=>"000011111",
  50350=>"011010000",
  50351=>"010100111",
  50352=>"110000100",
  50353=>"000100000",
  50354=>"111010101",
  50355=>"000101110",
  50356=>"110110101",
  50357=>"110011110",
  50358=>"001100100",
  50359=>"101101000",
  50360=>"101110111",
  50361=>"100111111",
  50362=>"101100100",
  50363=>"111101100",
  50364=>"100111100",
  50365=>"010001001",
  50366=>"000011100",
  50367=>"011001000",
  50368=>"010100101",
  50369=>"101011110",
  50370=>"001110101",
  50371=>"011011110",
  50372=>"011100010",
  50373=>"000111000",
  50374=>"101100110",
  50375=>"000111001",
  50376=>"111001111",
  50377=>"000100101",
  50378=>"011100100",
  50379=>"110100100",
  50380=>"111010111",
  50381=>"111101010",
  50382=>"110111100",
  50383=>"100011110",
  50384=>"001010010",
  50385=>"110100001",
  50386=>"001001001",
  50387=>"110111001",
  50388=>"110000001",
  50389=>"001001011",
  50390=>"111111001",
  50391=>"110100101",
  50392=>"011100000",
  50393=>"000101100",
  50394=>"000001010",
  50395=>"011110000",
  50396=>"110001000",
  50397=>"110100101",
  50398=>"111100100",
  50399=>"111011011",
  50400=>"111001001",
  50401=>"000111010",
  50402=>"110111110",
  50403=>"001000100",
  50404=>"111011111",
  50405=>"100110111",
  50406=>"000001001",
  50407=>"011011001",
  50408=>"101111001",
  50409=>"011101111",
  50410=>"000101111",
  50411=>"010010101",
  50412=>"100010100",
  50413=>"100001100",
  50414=>"100011011",
  50415=>"110110101",
  50416=>"001111100",
  50417=>"010111100",
  50418=>"110001001",
  50419=>"001001110",
  50420=>"110110011",
  50421=>"101010011",
  50422=>"010110001",
  50423=>"010001011",
  50424=>"100101101",
  50425=>"100101101",
  50426=>"011110111",
  50427=>"000011101",
  50428=>"011110100",
  50429=>"100001111",
  50430=>"010100000",
  50431=>"101111110",
  50432=>"001110000",
  50433=>"010111111",
  50434=>"010110001",
  50435=>"110000000",
  50436=>"001001001",
  50437=>"000001111",
  50438=>"100100000",
  50439=>"101010101",
  50440=>"001011110",
  50441=>"000100100",
  50442=>"001110000",
  50443=>"000111100",
  50444=>"110101000",
  50445=>"010111101",
  50446=>"011001011",
  50447=>"011000000",
  50448=>"100110001",
  50449=>"100100010",
  50450=>"010001110",
  50451=>"011100000",
  50452=>"111001110",
  50453=>"101111110",
  50454=>"110111100",
  50455=>"011000111",
  50456=>"011101000",
  50457=>"110011011",
  50458=>"100000001",
  50459=>"100011100",
  50460=>"100010011",
  50461=>"101011110",
  50462=>"011101111",
  50463=>"100101011",
  50464=>"001010100",
  50465=>"010111001",
  50466=>"000011011",
  50467=>"010100111",
  50468=>"101011100",
  50469=>"011011111",
  50470=>"011101111",
  50471=>"010110111",
  50472=>"000100010",
  50473=>"000000101",
  50474=>"001001100",
  50475=>"000100011",
  50476=>"111011110",
  50477=>"110001000",
  50478=>"001001100",
  50479=>"101100001",
  50480=>"001010100",
  50481=>"111011101",
  50482=>"011011000",
  50483=>"000000010",
  50484=>"111111111",
  50485=>"011011100",
  50486=>"110101010",
  50487=>"100110000",
  50488=>"110001101",
  50489=>"000001100",
  50490=>"110100111",
  50491=>"100101010",
  50492=>"001111111",
  50493=>"110101110",
  50494=>"111110100",
  50495=>"110110011",
  50496=>"111101101",
  50497=>"010011011",
  50498=>"100111001",
  50499=>"110111100",
  50500=>"000110110",
  50501=>"111010010",
  50502=>"011000000",
  50503=>"000001100",
  50504=>"000011111",
  50505=>"000010111",
  50506=>"001011101",
  50507=>"010011100",
  50508=>"010000100",
  50509=>"011100101",
  50510=>"001011110",
  50511=>"010110010",
  50512=>"110110101",
  50513=>"101000100",
  50514=>"010001000",
  50515=>"000100001",
  50516=>"000011101",
  50517=>"110010100",
  50518=>"100000110",
  50519=>"111101001",
  50520=>"101001110",
  50521=>"010111010",
  50522=>"111111110",
  50523=>"101000001",
  50524=>"101011110",
  50525=>"100111011",
  50526=>"011000011",
  50527=>"111101001",
  50528=>"011000110",
  50529=>"000101111",
  50530=>"000111101",
  50531=>"101001111",
  50532=>"010101010",
  50533=>"100110011",
  50534=>"110000011",
  50535=>"010010100",
  50536=>"100010011",
  50537=>"010000001",
  50538=>"011101011",
  50539=>"010100100",
  50540=>"001111010",
  50541=>"111011001",
  50542=>"110111110",
  50543=>"101011101",
  50544=>"010101001",
  50545=>"000100010",
  50546=>"011010111",
  50547=>"110001101",
  50548=>"100010100",
  50549=>"111101000",
  50550=>"110001011",
  50551=>"111101110",
  50552=>"000101000",
  50553=>"010000011",
  50554=>"011111111",
  50555=>"001100100",
  50556=>"101100011",
  50557=>"101110000",
  50558=>"101001000",
  50559=>"011101000",
  50560=>"100011001",
  50561=>"010110101",
  50562=>"001111001",
  50563=>"010101111",
  50564=>"001011000",
  50565=>"110001001",
  50566=>"111110111",
  50567=>"001111110",
  50568=>"000000110",
  50569=>"000110110",
  50570=>"011110001",
  50571=>"101100001",
  50572=>"000100000",
  50573=>"001000000",
  50574=>"011000100",
  50575=>"011101010",
  50576=>"101101011",
  50577=>"101000100",
  50578=>"111010010",
  50579=>"111010101",
  50580=>"111111010",
  50581=>"011110010",
  50582=>"010010010",
  50583=>"110000010",
  50584=>"010101010",
  50585=>"100100011",
  50586=>"001111110",
  50587=>"011001100",
  50588=>"000110111",
  50589=>"101101101",
  50590=>"001110000",
  50591=>"011001011",
  50592=>"100010011",
  50593=>"000111000",
  50594=>"111110010",
  50595=>"001000111",
  50596=>"100101110",
  50597=>"000011100",
  50598=>"100000101",
  50599=>"000000111",
  50600=>"001001110",
  50601=>"000110100",
  50602=>"011101111",
  50603=>"101111010",
  50604=>"101011001",
  50605=>"101001100",
  50606=>"111110101",
  50607=>"101101100",
  50608=>"011000011",
  50609=>"011001110",
  50610=>"100011111",
  50611=>"000110100",
  50612=>"111111100",
  50613=>"001001100",
  50614=>"000011000",
  50615=>"010001001",
  50616=>"011110001",
  50617=>"110000101",
  50618=>"110011001",
  50619=>"011011100",
  50620=>"010110000",
  50621=>"111011010",
  50622=>"001010001",
  50623=>"100000001",
  50624=>"011001000",
  50625=>"011101000",
  50626=>"011000001",
  50627=>"111010001",
  50628=>"100100110",
  50629=>"111001000",
  50630=>"110100110",
  50631=>"011101101",
  50632=>"101001101",
  50633=>"101111001",
  50634=>"000000000",
  50635=>"101100000",
  50636=>"101011011",
  50637=>"110100010",
  50638=>"000101110",
  50639=>"111011110",
  50640=>"010010000",
  50641=>"001110000",
  50642=>"001001100",
  50643=>"110111000",
  50644=>"101000110",
  50645=>"101100010",
  50646=>"110111011",
  50647=>"100010001",
  50648=>"001001000",
  50649=>"111101100",
  50650=>"100100100",
  50651=>"000110011",
  50652=>"010101001",
  50653=>"111010000",
  50654=>"100101001",
  50655=>"010000011",
  50656=>"001110100",
  50657=>"001010110",
  50658=>"111000100",
  50659=>"001101011",
  50660=>"011110100",
  50661=>"111101110",
  50662=>"101000010",
  50663=>"000101101",
  50664=>"111001001",
  50665=>"110000011",
  50666=>"010011011",
  50667=>"001001101",
  50668=>"110011111",
  50669=>"110011001",
  50670=>"000111100",
  50671=>"001010100",
  50672=>"101001001",
  50673=>"111110101",
  50674=>"100011011",
  50675=>"101010100",
  50676=>"001001111",
  50677=>"000110011",
  50678=>"101100100",
  50679=>"110010111",
  50680=>"110110101",
  50681=>"011001001",
  50682=>"010110011",
  50683=>"111011101",
  50684=>"100111110",
  50685=>"000010001",
  50686=>"011001000",
  50687=>"110011000",
  50688=>"111110011",
  50689=>"000111010",
  50690=>"000010110",
  50691=>"010011011",
  50692=>"000000000",
  50693=>"001000101",
  50694=>"010000001",
  50695=>"010001100",
  50696=>"010000011",
  50697=>"001011111",
  50698=>"000101011",
  50699=>"110010000",
  50700=>"011000010",
  50701=>"101000000",
  50702=>"010100011",
  50703=>"000010011",
  50704=>"110111110",
  50705=>"100000000",
  50706=>"000101110",
  50707=>"001101111",
  50708=>"010000000",
  50709=>"010110111",
  50710=>"011011000",
  50711=>"011101111",
  50712=>"101100010",
  50713=>"011010111",
  50714=>"101101110",
  50715=>"000000100",
  50716=>"000011010",
  50717=>"010010011",
  50718=>"111011110",
  50719=>"100100010",
  50720=>"110000001",
  50721=>"111101011",
  50722=>"010001100",
  50723=>"000001000",
  50724=>"111010101",
  50725=>"101101010",
  50726=>"100101101",
  50727=>"110001110",
  50728=>"110001000",
  50729=>"001011010",
  50730=>"011000001",
  50731=>"001000011",
  50732=>"101101101",
  50733=>"100101110",
  50734=>"011101010",
  50735=>"101000001",
  50736=>"000110111",
  50737=>"100110100",
  50738=>"011011000",
  50739=>"000001011",
  50740=>"010001000",
  50741=>"011001010",
  50742=>"111111010",
  50743=>"100010111",
  50744=>"110111000",
  50745=>"101001100",
  50746=>"100110101",
  50747=>"111100110",
  50748=>"101110000",
  50749=>"110100000",
  50750=>"001000001",
  50751=>"001011101",
  50752=>"111011111",
  50753=>"010011011",
  50754=>"110011111",
  50755=>"110111000",
  50756=>"011010110",
  50757=>"110011110",
  50758=>"010000011",
  50759=>"001010000",
  50760=>"101111100",
  50761=>"110100000",
  50762=>"010011100",
  50763=>"001011010",
  50764=>"000100101",
  50765=>"001001010",
  50766=>"100011100",
  50767=>"010011101",
  50768=>"000110111",
  50769=>"000101101",
  50770=>"011100110",
  50771=>"001010001",
  50772=>"100100111",
  50773=>"001010001",
  50774=>"100011000",
  50775=>"001100101",
  50776=>"100011101",
  50777=>"010001010",
  50778=>"011000001",
  50779=>"000110000",
  50780=>"011000001",
  50781=>"011011010",
  50782=>"000000000",
  50783=>"111110111",
  50784=>"101000010",
  50785=>"011001110",
  50786=>"011100000",
  50787=>"010100101",
  50788=>"011101010",
  50789=>"001000001",
  50790=>"111001110",
  50791=>"010011100",
  50792=>"111101111",
  50793=>"111010000",
  50794=>"110011011",
  50795=>"010000100",
  50796=>"111011111",
  50797=>"001000101",
  50798=>"001001110",
  50799=>"001000000",
  50800=>"001000110",
  50801=>"000011000",
  50802=>"101000111",
  50803=>"001111111",
  50804=>"011111111",
  50805=>"001110010",
  50806=>"111011000",
  50807=>"101110100",
  50808=>"110000011",
  50809=>"111101100",
  50810=>"111100111",
  50811=>"000000000",
  50812=>"010001111",
  50813=>"011101101",
  50814=>"110101101",
  50815=>"110010100",
  50816=>"010101101",
  50817=>"010011100",
  50818=>"011001111",
  50819=>"001101100",
  50820=>"110100101",
  50821=>"101100011",
  50822=>"100101001",
  50823=>"000010100",
  50824=>"101011010",
  50825=>"100000101",
  50826=>"011010001",
  50827=>"010111100",
  50828=>"101010001",
  50829=>"010101111",
  50830=>"111110011",
  50831=>"101000101",
  50832=>"001011001",
  50833=>"000111011",
  50834=>"010001001",
  50835=>"111010011",
  50836=>"000100110",
  50837=>"011000011",
  50838=>"010001000",
  50839=>"010010010",
  50840=>"010010101",
  50841=>"110011010",
  50842=>"111100000",
  50843=>"001111111",
  50844=>"110001001",
  50845=>"001000100",
  50846=>"000011000",
  50847=>"010101011",
  50848=>"001110000",
  50849=>"110001111",
  50850=>"000110011",
  50851=>"001000111",
  50852=>"011011111",
  50853=>"100111011",
  50854=>"000000101",
  50855=>"000111110",
  50856=>"110111001",
  50857=>"001110111",
  50858=>"010011010",
  50859=>"010100001",
  50860=>"111010010",
  50861=>"010010000",
  50862=>"000011110",
  50863=>"111100111",
  50864=>"111010011",
  50865=>"000011010",
  50866=>"001100010",
  50867=>"001000100",
  50868=>"110111100",
  50869=>"010000111",
  50870=>"111011000",
  50871=>"010111111",
  50872=>"100101110",
  50873=>"111011111",
  50874=>"111111000",
  50875=>"000101000",
  50876=>"000011011",
  50877=>"100010011",
  50878=>"111111011",
  50879=>"010110111",
  50880=>"110011001",
  50881=>"000100100",
  50882=>"110011001",
  50883=>"101011110",
  50884=>"000001100",
  50885=>"100011000",
  50886=>"101000001",
  50887=>"101010101",
  50888=>"110100100",
  50889=>"011101110",
  50890=>"100101101",
  50891=>"101100011",
  50892=>"110101011",
  50893=>"011001001",
  50894=>"010101101",
  50895=>"000100010",
  50896=>"100011000",
  50897=>"000000001",
  50898=>"011110010",
  50899=>"010001100",
  50900=>"100010011",
  50901=>"001001101",
  50902=>"000101010",
  50903=>"111001101",
  50904=>"101001000",
  50905=>"000110101",
  50906=>"110000100",
  50907=>"110010100",
  50908=>"111100011",
  50909=>"110011000",
  50910=>"101010111",
  50911=>"100010010",
  50912=>"000111001",
  50913=>"101001101",
  50914=>"100100100",
  50915=>"000011111",
  50916=>"011011110",
  50917=>"101101101",
  50918=>"000001110",
  50919=>"010000001",
  50920=>"000011010",
  50921=>"001100011",
  50922=>"101101010",
  50923=>"111111011",
  50924=>"010011001",
  50925=>"110000001",
  50926=>"010111011",
  50927=>"110001100",
  50928=>"011110001",
  50929=>"110111011",
  50930=>"000100000",
  50931=>"101010110",
  50932=>"000100101",
  50933=>"100000100",
  50934=>"111110111",
  50935=>"100001000",
  50936=>"100000000",
  50937=>"111010010",
  50938=>"100000101",
  50939=>"110000011",
  50940=>"100001011",
  50941=>"010100110",
  50942=>"000000111",
  50943=>"001000010",
  50944=>"010101100",
  50945=>"111000010",
  50946=>"110101000",
  50947=>"001101110",
  50948=>"110110111",
  50949=>"000000110",
  50950=>"011101010",
  50951=>"010001010",
  50952=>"110011101",
  50953=>"111000111",
  50954=>"101110110",
  50955=>"100111110",
  50956=>"000000100",
  50957=>"000000111",
  50958=>"010101110",
  50959=>"010100010",
  50960=>"011100110",
  50961=>"001110000",
  50962=>"100000000",
  50963=>"110111000",
  50964=>"101111100",
  50965=>"001101010",
  50966=>"011100001",
  50967=>"110001000",
  50968=>"110101110",
  50969=>"011010011",
  50970=>"010010010",
  50971=>"001001001",
  50972=>"010000110",
  50973=>"101101100",
  50974=>"110010111",
  50975=>"100110110",
  50976=>"010011011",
  50977=>"100001001",
  50978=>"101110111",
  50979=>"001010011",
  50980=>"001010000",
  50981=>"111001111",
  50982=>"110111010",
  50983=>"100100000",
  50984=>"110101000",
  50985=>"000111001",
  50986=>"110001111",
  50987=>"100011100",
  50988=>"111111011",
  50989=>"110010101",
  50990=>"100111110",
  50991=>"110100001",
  50992=>"000110110",
  50993=>"000001100",
  50994=>"010001001",
  50995=>"111100010",
  50996=>"111111111",
  50997=>"111111110",
  50998=>"110000010",
  50999=>"100110001",
  51000=>"000011000",
  51001=>"000001011",
  51002=>"000110001",
  51003=>"100010101",
  51004=>"100111001",
  51005=>"000011010",
  51006=>"010000100",
  51007=>"110100001",
  51008=>"110110001",
  51009=>"111111101",
  51010=>"011011000",
  51011=>"110100101",
  51012=>"000101000",
  51013=>"110010001",
  51014=>"100101110",
  51015=>"111111111",
  51016=>"011001111",
  51017=>"000111111",
  51018=>"001110100",
  51019=>"000001000",
  51020=>"000000010",
  51021=>"111100010",
  51022=>"001111001",
  51023=>"111010010",
  51024=>"010010000",
  51025=>"100110110",
  51026=>"110000001",
  51027=>"011010100",
  51028=>"000000000",
  51029=>"111010101",
  51030=>"100010000",
  51031=>"000101111",
  51032=>"000011000",
  51033=>"110001111",
  51034=>"011000000",
  51035=>"110010100",
  51036=>"101111100",
  51037=>"101001000",
  51038=>"010111111",
  51039=>"110000110",
  51040=>"111111010",
  51041=>"111000011",
  51042=>"001101011",
  51043=>"101110001",
  51044=>"001000010",
  51045=>"010000001",
  51046=>"100110011",
  51047=>"101000011",
  51048=>"110101100",
  51049=>"011110010",
  51050=>"101010100",
  51051=>"001111111",
  51052=>"110100001",
  51053=>"100110110",
  51054=>"110111111",
  51055=>"111001011",
  51056=>"001010111",
  51057=>"011101100",
  51058=>"110101111",
  51059=>"011100110",
  51060=>"101110100",
  51061=>"100000010",
  51062=>"010010011",
  51063=>"010011101",
  51064=>"111011001",
  51065=>"001001011",
  51066=>"000010011",
  51067=>"010111111",
  51068=>"000010010",
  51069=>"011100001",
  51070=>"010100010",
  51071=>"011100011",
  51072=>"000110001",
  51073=>"000101001",
  51074=>"101111101",
  51075=>"100111000",
  51076=>"110001100",
  51077=>"010001001",
  51078=>"001010110",
  51079=>"011000110",
  51080=>"111110111",
  51081=>"101111011",
  51082=>"000001110",
  51083=>"111100011",
  51084=>"001101110",
  51085=>"011000000",
  51086=>"010011001",
  51087=>"010101110",
  51088=>"111111111",
  51089=>"101100101",
  51090=>"000000111",
  51091=>"101110011",
  51092=>"001101110",
  51093=>"100111010",
  51094=>"011110001",
  51095=>"010011010",
  51096=>"001010111",
  51097=>"101000101",
  51098=>"110101100",
  51099=>"100100011",
  51100=>"100111110",
  51101=>"011011001",
  51102=>"001010100",
  51103=>"110100000",
  51104=>"111011010",
  51105=>"101101010",
  51106=>"111010001",
  51107=>"000000011",
  51108=>"000000111",
  51109=>"111000101",
  51110=>"010001010",
  51111=>"100000100",
  51112=>"000111011",
  51113=>"010000000",
  51114=>"110000101",
  51115=>"000101000",
  51116=>"110100000",
  51117=>"000101101",
  51118=>"110111111",
  51119=>"010101001",
  51120=>"001011111",
  51121=>"110110101",
  51122=>"011001010",
  51123=>"110001000",
  51124=>"100111100",
  51125=>"001110010",
  51126=>"010110001",
  51127=>"101000001",
  51128=>"000101010",
  51129=>"100010111",
  51130=>"110010011",
  51131=>"001001011",
  51132=>"011000001",
  51133=>"000001000",
  51134=>"000010000",
  51135=>"100100011",
  51136=>"100010110",
  51137=>"001100100",
  51138=>"110011100",
  51139=>"100011000",
  51140=>"010101001",
  51141=>"110110101",
  51142=>"111101000",
  51143=>"011101100",
  51144=>"000000000",
  51145=>"010100001",
  51146=>"100010010",
  51147=>"110101011",
  51148=>"001111111",
  51149=>"011110010",
  51150=>"011010111",
  51151=>"110000010",
  51152=>"011100111",
  51153=>"000110111",
  51154=>"010000000",
  51155=>"110000110",
  51156=>"010100010",
  51157=>"000010110",
  51158=>"101000001",
  51159=>"001101100",
  51160=>"001000100",
  51161=>"110101001",
  51162=>"010100000",
  51163=>"111111110",
  51164=>"100010010",
  51165=>"000101111",
  51166=>"010100011",
  51167=>"101111001",
  51168=>"010111110",
  51169=>"100100010",
  51170=>"001000100",
  51171=>"000110111",
  51172=>"010001100",
  51173=>"100001001",
  51174=>"101010100",
  51175=>"110101010",
  51176=>"011010010",
  51177=>"100010001",
  51178=>"011101101",
  51179=>"101010110",
  51180=>"010100110",
  51181=>"000111010",
  51182=>"101110011",
  51183=>"111110111",
  51184=>"001011101",
  51185=>"000101001",
  51186=>"010000001",
  51187=>"101000110",
  51188=>"101000111",
  51189=>"010100010",
  51190=>"010001100",
  51191=>"111001110",
  51192=>"011111010",
  51193=>"011110001",
  51194=>"011010111",
  51195=>"111100110",
  51196=>"011100000",
  51197=>"111010010",
  51198=>"010010010",
  51199=>"001001110",
  51200=>"000101000",
  51201=>"101111100",
  51202=>"101100111",
  51203=>"111011101",
  51204=>"110001101",
  51205=>"101110111",
  51206=>"100011101",
  51207=>"000010101",
  51208=>"001111001",
  51209=>"100011101",
  51210=>"011001111",
  51211=>"100000111",
  51212=>"110000011",
  51213=>"101011000",
  51214=>"011011010",
  51215=>"111101001",
  51216=>"010010000",
  51217=>"000010010",
  51218=>"010001100",
  51219=>"001000010",
  51220=>"100001110",
  51221=>"001001011",
  51222=>"001110010",
  51223=>"100010001",
  51224=>"110111100",
  51225=>"100011000",
  51226=>"011111011",
  51227=>"101111110",
  51228=>"110001000",
  51229=>"101011101",
  51230=>"111100110",
  51231=>"011011111",
  51232=>"110011010",
  51233=>"011100111",
  51234=>"100100111",
  51235=>"010100101",
  51236=>"001110111",
  51237=>"101001101",
  51238=>"111000001",
  51239=>"101010101",
  51240=>"110111111",
  51241=>"000001000",
  51242=>"110011110",
  51243=>"000010101",
  51244=>"011001011",
  51245=>"010000111",
  51246=>"111111110",
  51247=>"100110011",
  51248=>"011010001",
  51249=>"100110010",
  51250=>"111110011",
  51251=>"111011111",
  51252=>"101010111",
  51253=>"110110110",
  51254=>"111100100",
  51255=>"101110100",
  51256=>"101101000",
  51257=>"011011010",
  51258=>"001011111",
  51259=>"001101011",
  51260=>"011011000",
  51261=>"110111110",
  51262=>"011100000",
  51263=>"011110110",
  51264=>"111010110",
  51265=>"010100011",
  51266=>"011010010",
  51267=>"111101110",
  51268=>"001101101",
  51269=>"011100110",
  51270=>"011000001",
  51271=>"100000011",
  51272=>"110100101",
  51273=>"010001000",
  51274=>"111100011",
  51275=>"110010110",
  51276=>"010110100",
  51277=>"111010101",
  51278=>"101000000",
  51279=>"100101101",
  51280=>"101010110",
  51281=>"110110011",
  51282=>"101000011",
  51283=>"110010011",
  51284=>"100110101",
  51285=>"111100100",
  51286=>"000100010",
  51287=>"000011010",
  51288=>"010101110",
  51289=>"111010010",
  51290=>"110110001",
  51291=>"010110110",
  51292=>"000101001",
  51293=>"000001111",
  51294=>"001110010",
  51295=>"001010000",
  51296=>"010001000",
  51297=>"001100100",
  51298=>"101101010",
  51299=>"010110100",
  51300=>"111100101",
  51301=>"111011100",
  51302=>"011101110",
  51303=>"011011001",
  51304=>"010100110",
  51305=>"100110000",
  51306=>"001000110",
  51307=>"001100101",
  51308=>"011010101",
  51309=>"110110111",
  51310=>"100010101",
  51311=>"110001100",
  51312=>"110110110",
  51313=>"100001000",
  51314=>"100110110",
  51315=>"111100010",
  51316=>"101010000",
  51317=>"010111110",
  51318=>"001010110",
  51319=>"011010111",
  51320=>"100011000",
  51321=>"000000111",
  51322=>"010010001",
  51323=>"000011111",
  51324=>"000010011",
  51325=>"000011001",
  51326=>"111011101",
  51327=>"111000001",
  51328=>"110001101",
  51329=>"101011111",
  51330=>"101000000",
  51331=>"010101010",
  51332=>"100111110",
  51333=>"010000011",
  51334=>"011101100",
  51335=>"101100110",
  51336=>"000110100",
  51337=>"010110101",
  51338=>"011011101",
  51339=>"110001000",
  51340=>"001100010",
  51341=>"110111001",
  51342=>"011011011",
  51343=>"010101100",
  51344=>"101001111",
  51345=>"111111111",
  51346=>"111111011",
  51347=>"111101000",
  51348=>"011110110",
  51349=>"100111101",
  51350=>"000100011",
  51351=>"011011111",
  51352=>"000010100",
  51353=>"001000100",
  51354=>"110111111",
  51355=>"001100110",
  51356=>"110000101",
  51357=>"111000010",
  51358=>"010111100",
  51359=>"101001001",
  51360=>"101101101",
  51361=>"001111011",
  51362=>"100100100",
  51363=>"010011011",
  51364=>"101011000",
  51365=>"110001000",
  51366=>"001110010",
  51367=>"101111010",
  51368=>"011111111",
  51369=>"101011100",
  51370=>"000100110",
  51371=>"001001000",
  51372=>"010010111",
  51373=>"111010100",
  51374=>"111111100",
  51375=>"000011011",
  51376=>"100101001",
  51377=>"000011011",
  51378=>"110100001",
  51379=>"111100011",
  51380=>"000110100",
  51381=>"101000110",
  51382=>"100101000",
  51383=>"001000001",
  51384=>"111100010",
  51385=>"001101000",
  51386=>"010001011",
  51387=>"011111100",
  51388=>"110101011",
  51389=>"100101000",
  51390=>"111111110",
  51391=>"000101111",
  51392=>"001000010",
  51393=>"011010000",
  51394=>"011100010",
  51395=>"110111101",
  51396=>"101010000",
  51397=>"001000000",
  51398=>"101111111",
  51399=>"001000110",
  51400=>"010101111",
  51401=>"001011101",
  51402=>"100110011",
  51403=>"100010101",
  51404=>"101011010",
  51405=>"011001110",
  51406=>"000000001",
  51407=>"101011110",
  51408=>"001101000",
  51409=>"001001111",
  51410=>"000101100",
  51411=>"110011001",
  51412=>"110011000",
  51413=>"111111111",
  51414=>"010011001",
  51415=>"101100010",
  51416=>"000100010",
  51417=>"010110011",
  51418=>"010010011",
  51419=>"110011101",
  51420=>"111011000",
  51421=>"111010000",
  51422=>"110000101",
  51423=>"101100101",
  51424=>"010000100",
  51425=>"001101010",
  51426=>"011111100",
  51427=>"110110000",
  51428=>"100001001",
  51429=>"001111000",
  51430=>"111110110",
  51431=>"110010101",
  51432=>"110110101",
  51433=>"011001110",
  51434=>"011010110",
  51435=>"000110110",
  51436=>"011111101",
  51437=>"001000111",
  51438=>"100000101",
  51439=>"001100100",
  51440=>"010110100",
  51441=>"011010110",
  51442=>"110100001",
  51443=>"110110010",
  51444=>"000100101",
  51445=>"101001111",
  51446=>"110100000",
  51447=>"000111000",
  51448=>"101101101",
  51449=>"011011111",
  51450=>"111111001",
  51451=>"110000001",
  51452=>"011100101",
  51453=>"011000001",
  51454=>"100100111",
  51455=>"000101000",
  51456=>"011100111",
  51457=>"110110100",
  51458=>"010110110",
  51459=>"111000100",
  51460=>"000100101",
  51461=>"010010110",
  51462=>"001000000",
  51463=>"101100101",
  51464=>"101111110",
  51465=>"010001100",
  51466=>"011001000",
  51467=>"010111000",
  51468=>"100000001",
  51469=>"100100011",
  51470=>"011001110",
  51471=>"001100100",
  51472=>"001010111",
  51473=>"101001111",
  51474=>"111101110",
  51475=>"011111101",
  51476=>"000010111",
  51477=>"011011111",
  51478=>"101111010",
  51479=>"011111011",
  51480=>"001011010",
  51481=>"110110111",
  51482=>"010111011",
  51483=>"010001011",
  51484=>"101001010",
  51485=>"110000100",
  51486=>"101111001",
  51487=>"000100111",
  51488=>"001010101",
  51489=>"011010000",
  51490=>"010110110",
  51491=>"001001111",
  51492=>"011111100",
  51493=>"100110001",
  51494=>"000011010",
  51495=>"010111111",
  51496=>"111010110",
  51497=>"011101110",
  51498=>"110111111",
  51499=>"101010001",
  51500=>"110110111",
  51501=>"111110111",
  51502=>"001000111",
  51503=>"001111001",
  51504=>"110110111",
  51505=>"101011000",
  51506=>"011010011",
  51507=>"100101101",
  51508=>"011010110",
  51509=>"000001001",
  51510=>"011011101",
  51511=>"011010011",
  51512=>"111101010",
  51513=>"011000001",
  51514=>"011110000",
  51515=>"101100000",
  51516=>"101101001",
  51517=>"101011011",
  51518=>"100000101",
  51519=>"111001110",
  51520=>"010101111",
  51521=>"011101110",
  51522=>"000111001",
  51523=>"010000101",
  51524=>"110100011",
  51525=>"010100110",
  51526=>"100000111",
  51527=>"111111010",
  51528=>"101000010",
  51529=>"110101000",
  51530=>"000000110",
  51531=>"100110111",
  51532=>"101010110",
  51533=>"000110010",
  51534=>"100011010",
  51535=>"000100000",
  51536=>"110000001",
  51537=>"010111011",
  51538=>"111010010",
  51539=>"010000011",
  51540=>"010101010",
  51541=>"101010110",
  51542=>"001011110",
  51543=>"101001101",
  51544=>"001111111",
  51545=>"000010010",
  51546=>"010000001",
  51547=>"111100011",
  51548=>"000110011",
  51549=>"101000010",
  51550=>"100000110",
  51551=>"100100000",
  51552=>"001010111",
  51553=>"100001110",
  51554=>"010111101",
  51555=>"000010010",
  51556=>"000101010",
  51557=>"000111101",
  51558=>"111111100",
  51559=>"000100001",
  51560=>"111000110",
  51561=>"000101101",
  51562=>"101011001",
  51563=>"001011000",
  51564=>"110111111",
  51565=>"111101110",
  51566=>"010101100",
  51567=>"101110100",
  51568=>"000010101",
  51569=>"000010100",
  51570=>"011100001",
  51571=>"000111110",
  51572=>"001000001",
  51573=>"111111110",
  51574=>"010001110",
  51575=>"000101000",
  51576=>"110110011",
  51577=>"011101111",
  51578=>"101011111",
  51579=>"000000101",
  51580=>"111110001",
  51581=>"111100000",
  51582=>"010111100",
  51583=>"111011001",
  51584=>"111100111",
  51585=>"101001011",
  51586=>"111001010",
  51587=>"111011010",
  51588=>"001100110",
  51589=>"010111111",
  51590=>"101111110",
  51591=>"111100000",
  51592=>"011010011",
  51593=>"011011110",
  51594=>"110101110",
  51595=>"100100000",
  51596=>"011010100",
  51597=>"100001010",
  51598=>"001001000",
  51599=>"000000001",
  51600=>"110100111",
  51601=>"110110100",
  51602=>"011100001",
  51603=>"010001001",
  51604=>"101000000",
  51605=>"111101011",
  51606=>"111010011",
  51607=>"001011100",
  51608=>"100100011",
  51609=>"110100101",
  51610=>"101101010",
  51611=>"000001000",
  51612=>"001001110",
  51613=>"111011100",
  51614=>"101010100",
  51615=>"000011011",
  51616=>"010100010",
  51617=>"010000000",
  51618=>"000011100",
  51619=>"110001111",
  51620=>"000001010",
  51621=>"001110001",
  51622=>"001110111",
  51623=>"001110101",
  51624=>"110010010",
  51625=>"010010111",
  51626=>"000111111",
  51627=>"111111110",
  51628=>"011001001",
  51629=>"101101101",
  51630=>"110111010",
  51631=>"111111111",
  51632=>"101001110",
  51633=>"110110100",
  51634=>"111100011",
  51635=>"001110000",
  51636=>"010101011",
  51637=>"111100110",
  51638=>"100111000",
  51639=>"101111111",
  51640=>"011000011",
  51641=>"100001100",
  51642=>"111010000",
  51643=>"101001001",
  51644=>"110000010",
  51645=>"001101011",
  51646=>"110101111",
  51647=>"011111111",
  51648=>"001100101",
  51649=>"000001000",
  51650=>"011011100",
  51651=>"011000001",
  51652=>"111110111",
  51653=>"000001000",
  51654=>"000001010",
  51655=>"010101101",
  51656=>"111010000",
  51657=>"011100100",
  51658=>"111011111",
  51659=>"111001110",
  51660=>"010000011",
  51661=>"010111011",
  51662=>"101110000",
  51663=>"111001011",
  51664=>"000100101",
  51665=>"111110101",
  51666=>"111001100",
  51667=>"011111000",
  51668=>"111001110",
  51669=>"010101101",
  51670=>"100001101",
  51671=>"100010001",
  51672=>"001100000",
  51673=>"001110110",
  51674=>"111010001",
  51675=>"100110011",
  51676=>"001101001",
  51677=>"101011111",
  51678=>"101111101",
  51679=>"001101100",
  51680=>"000001011",
  51681=>"100111011",
  51682=>"011110101",
  51683=>"011100011",
  51684=>"110010110",
  51685=>"011111010",
  51686=>"011101111",
  51687=>"101110101",
  51688=>"100010100",
  51689=>"000111001",
  51690=>"101101001",
  51691=>"011000111",
  51692=>"011000011",
  51693=>"001001111",
  51694=>"100000011",
  51695=>"010001110",
  51696=>"001100000",
  51697=>"010000011",
  51698=>"010100000",
  51699=>"001001000",
  51700=>"111110101",
  51701=>"101000111",
  51702=>"111001100",
  51703=>"100010000",
  51704=>"000110000",
  51705=>"101110100",
  51706=>"000110001",
  51707=>"100110110",
  51708=>"010010000",
  51709=>"111101010",
  51710=>"011001110",
  51711=>"111001011",
  51712=>"001101101",
  51713=>"011101011",
  51714=>"111000111",
  51715=>"101001000",
  51716=>"111100011",
  51717=>"001001000",
  51718=>"010100101",
  51719=>"010100000",
  51720=>"101110001",
  51721=>"010011011",
  51722=>"100111100",
  51723=>"010110001",
  51724=>"101111101",
  51725=>"010000011",
  51726=>"100100011",
  51727=>"110001011",
  51728=>"101010011",
  51729=>"011010000",
  51730=>"110111110",
  51731=>"111000101",
  51732=>"011000101",
  51733=>"111010101",
  51734=>"000000010",
  51735=>"111111110",
  51736=>"010010111",
  51737=>"100100101",
  51738=>"010001101",
  51739=>"000000101",
  51740=>"001011000",
  51741=>"101011000",
  51742=>"010000011",
  51743=>"101111101",
  51744=>"110101101",
  51745=>"010101101",
  51746=>"010001011",
  51747=>"111110111",
  51748=>"101101101",
  51749=>"110001110",
  51750=>"100010001",
  51751=>"100110111",
  51752=>"001111001",
  51753=>"011110111",
  51754=>"111100100",
  51755=>"101001000",
  51756=>"011011100",
  51757=>"110100110",
  51758=>"100111100",
  51759=>"011010111",
  51760=>"110111011",
  51761=>"000001100",
  51762=>"111100100",
  51763=>"000010011",
  51764=>"001010100",
  51765=>"101010111",
  51766=>"011111111",
  51767=>"011010000",
  51768=>"101011110",
  51769=>"111100011",
  51770=>"011110110",
  51771=>"011001011",
  51772=>"100010110",
  51773=>"110001111",
  51774=>"001000101",
  51775=>"100010100",
  51776=>"101101011",
  51777=>"000111110",
  51778=>"110100100",
  51779=>"100110010",
  51780=>"110011100",
  51781=>"001001010",
  51782=>"001111110",
  51783=>"111110111",
  51784=>"000000000",
  51785=>"011000111",
  51786=>"011000101",
  51787=>"111000011",
  51788=>"000100001",
  51789=>"010000101",
  51790=>"000000000",
  51791=>"000110011",
  51792=>"111111111",
  51793=>"110001111",
  51794=>"111011011",
  51795=>"110000100",
  51796=>"110100010",
  51797=>"000010100",
  51798=>"001001001",
  51799=>"011010001",
  51800=>"111100000",
  51801=>"100011000",
  51802=>"101111110",
  51803=>"001110000",
  51804=>"111100111",
  51805=>"000010110",
  51806=>"000110100",
  51807=>"111110111",
  51808=>"100101101",
  51809=>"010001000",
  51810=>"100000000",
  51811=>"111110010",
  51812=>"111011001",
  51813=>"011010110",
  51814=>"101011111",
  51815=>"000111000",
  51816=>"101111111",
  51817=>"010011110",
  51818=>"101000101",
  51819=>"001100110",
  51820=>"000100101",
  51821=>"100101111",
  51822=>"111100011",
  51823=>"100110101",
  51824=>"000011101",
  51825=>"100010100",
  51826=>"100101100",
  51827=>"100100010",
  51828=>"111101100",
  51829=>"000001010",
  51830=>"000000011",
  51831=>"011011100",
  51832=>"001101110",
  51833=>"101110010",
  51834=>"100100111",
  51835=>"000010101",
  51836=>"111110111",
  51837=>"110011101",
  51838=>"110111101",
  51839=>"000010010",
  51840=>"011101110",
  51841=>"011000000",
  51842=>"111101111",
  51843=>"010010111",
  51844=>"101101010",
  51845=>"100110011",
  51846=>"110110100",
  51847=>"100001100",
  51848=>"111011110",
  51849=>"010010001",
  51850=>"100100011",
  51851=>"011010100",
  51852=>"001101001",
  51853=>"000001000",
  51854=>"010011111",
  51855=>"001100001",
  51856=>"000011011",
  51857=>"001000010",
  51858=>"011011100",
  51859=>"111000011",
  51860=>"001100101",
  51861=>"011010001",
  51862=>"100000111",
  51863=>"101101110",
  51864=>"011110000",
  51865=>"100100101",
  51866=>"101010011",
  51867=>"011010110",
  51868=>"010000111",
  51869=>"110110000",
  51870=>"001011110",
  51871=>"011011110",
  51872=>"110110101",
  51873=>"100110110",
  51874=>"011001001",
  51875=>"111010101",
  51876=>"110010000",
  51877=>"110101001",
  51878=>"110110001",
  51879=>"011011100",
  51880=>"000100000",
  51881=>"111111011",
  51882=>"001000010",
  51883=>"111100000",
  51884=>"001101100",
  51885=>"001011110",
  51886=>"101010011",
  51887=>"101110100",
  51888=>"001010111",
  51889=>"101101001",
  51890=>"111001000",
  51891=>"100100111",
  51892=>"111101101",
  51893=>"100010001",
  51894=>"100111111",
  51895=>"100101101",
  51896=>"100110000",
  51897=>"101100111",
  51898=>"001100011",
  51899=>"110100101",
  51900=>"010101011",
  51901=>"111010011",
  51902=>"110011111",
  51903=>"101101110",
  51904=>"001001011",
  51905=>"000100010",
  51906=>"011111101",
  51907=>"011000010",
  51908=>"110001110",
  51909=>"001001011",
  51910=>"110010001",
  51911=>"010101010",
  51912=>"111111100",
  51913=>"000001111",
  51914=>"111000011",
  51915=>"010011000",
  51916=>"001010001",
  51917=>"010100000",
  51918=>"001111100",
  51919=>"101011011",
  51920=>"001100110",
  51921=>"101000100",
  51922=>"100111101",
  51923=>"001101100",
  51924=>"101001111",
  51925=>"000011011",
  51926=>"001110110",
  51927=>"100101100",
  51928=>"101001001",
  51929=>"001101101",
  51930=>"010001101",
  51931=>"001001100",
  51932=>"111101000",
  51933=>"010110001",
  51934=>"000010001",
  51935=>"011111011",
  51936=>"011011001",
  51937=>"111110000",
  51938=>"111010001",
  51939=>"101101111",
  51940=>"100000000",
  51941=>"000111110",
  51942=>"011011011",
  51943=>"101100010",
  51944=>"011101110",
  51945=>"010111000",
  51946=>"001011011",
  51947=>"011110011",
  51948=>"110001011",
  51949=>"001101101",
  51950=>"111010010",
  51951=>"010010011",
  51952=>"001000101",
  51953=>"110101000",
  51954=>"001001101",
  51955=>"010111000",
  51956=>"110011111",
  51957=>"000111101",
  51958=>"010101001",
  51959=>"001001111",
  51960=>"101101110",
  51961=>"000000000",
  51962=>"010011001",
  51963=>"110100001",
  51964=>"101001000",
  51965=>"111000111",
  51966=>"001111000",
  51967=>"011011010",
  51968=>"011001001",
  51969=>"010001100",
  51970=>"001100011",
  51971=>"010010000",
  51972=>"110100000",
  51973=>"110011000",
  51974=>"001111001",
  51975=>"001000000",
  51976=>"001101010",
  51977=>"010011010",
  51978=>"111000001",
  51979=>"011100000",
  51980=>"111110000",
  51981=>"101001010",
  51982=>"011111111",
  51983=>"101010110",
  51984=>"010011000",
  51985=>"111110010",
  51986=>"101001011",
  51987=>"101101010",
  51988=>"101101010",
  51989=>"110101011",
  51990=>"100111011",
  51991=>"111111011",
  51992=>"001000001",
  51993=>"001011001",
  51994=>"100110010",
  51995=>"001000110",
  51996=>"110010100",
  51997=>"110010101",
  51998=>"111101101",
  51999=>"101101001",
  52000=>"111100011",
  52001=>"010001101",
  52002=>"110111010",
  52003=>"111010111",
  52004=>"011101101",
  52005=>"100110100",
  52006=>"011101111",
  52007=>"010010110",
  52008=>"111010011",
  52009=>"000101110",
  52010=>"100000001",
  52011=>"101110111",
  52012=>"100110110",
  52013=>"111011100",
  52014=>"011000001",
  52015=>"101111000",
  52016=>"000000000",
  52017=>"000010110",
  52018=>"110100010",
  52019=>"010101110",
  52020=>"000000000",
  52021=>"110111110",
  52022=>"100110110",
  52023=>"001011111",
  52024=>"010011001",
  52025=>"010100101",
  52026=>"110001100",
  52027=>"000011011",
  52028=>"101001010",
  52029=>"110100100",
  52030=>"101110100",
  52031=>"101001000",
  52032=>"110101000",
  52033=>"101111111",
  52034=>"001010000",
  52035=>"100000001",
  52036=>"001000111",
  52037=>"110010001",
  52038=>"101100110",
  52039=>"110111001",
  52040=>"001011001",
  52041=>"011101100",
  52042=>"010100000",
  52043=>"000100100",
  52044=>"101010011",
  52045=>"011000100",
  52046=>"100111001",
  52047=>"100011110",
  52048=>"010100101",
  52049=>"010000000",
  52050=>"101011010",
  52051=>"010000000",
  52052=>"010000001",
  52053=>"011110100",
  52054=>"001001001",
  52055=>"101000101",
  52056=>"111110111",
  52057=>"100111101",
  52058=>"110110000",
  52059=>"011100010",
  52060=>"011010000",
  52061=>"100101010",
  52062=>"001001100",
  52063=>"001001010",
  52064=>"011010010",
  52065=>"010110001",
  52066=>"101001110",
  52067=>"011101101",
  52068=>"010001001",
  52069=>"101011000",
  52070=>"110001100",
  52071=>"111011101",
  52072=>"011010110",
  52073=>"110011001",
  52074=>"001011100",
  52075=>"111001000",
  52076=>"000110100",
  52077=>"001001110",
  52078=>"100000000",
  52079=>"100110000",
  52080=>"010011100",
  52081=>"001110011",
  52082=>"010000101",
  52083=>"111010100",
  52084=>"000001100",
  52085=>"110111000",
  52086=>"100001100",
  52087=>"010111000",
  52088=>"100011011",
  52089=>"010100100",
  52090=>"000111101",
  52091=>"110110010",
  52092=>"111111111",
  52093=>"100100011",
  52094=>"000111111",
  52095=>"100101111",
  52096=>"110101100",
  52097=>"101101100",
  52098=>"001100000",
  52099=>"100111010",
  52100=>"100001111",
  52101=>"110011100",
  52102=>"101111111",
  52103=>"000100001",
  52104=>"101100101",
  52105=>"100100001",
  52106=>"110101111",
  52107=>"000000100",
  52108=>"100000111",
  52109=>"001100111",
  52110=>"010001010",
  52111=>"000000110",
  52112=>"000010110",
  52113=>"110101000",
  52114=>"010100100",
  52115=>"000000111",
  52116=>"101010010",
  52117=>"011111001",
  52118=>"000100111",
  52119=>"000101101",
  52120=>"111000010",
  52121=>"101101001",
  52122=>"000001101",
  52123=>"110100010",
  52124=>"100101010",
  52125=>"000110001",
  52126=>"101110111",
  52127=>"111011001",
  52128=>"101001001",
  52129=>"001001111",
  52130=>"000101100",
  52131=>"110111010",
  52132=>"000111110",
  52133=>"110111011",
  52134=>"100001111",
  52135=>"001001001",
  52136=>"010010011",
  52137=>"110111100",
  52138=>"111111001",
  52139=>"010011101",
  52140=>"110110000",
  52141=>"010111101",
  52142=>"000011001",
  52143=>"011110010",
  52144=>"001100111",
  52145=>"111110011",
  52146=>"001101111",
  52147=>"011101111",
  52148=>"101011100",
  52149=>"011001100",
  52150=>"111101000",
  52151=>"111001101",
  52152=>"100110110",
  52153=>"000100000",
  52154=>"011010010",
  52155=>"011100011",
  52156=>"010011100",
  52157=>"100000111",
  52158=>"111010111",
  52159=>"111110101",
  52160=>"101110111",
  52161=>"011011110",
  52162=>"000100000",
  52163=>"010000100",
  52164=>"010001100",
  52165=>"100001011",
  52166=>"101101010",
  52167=>"111110010",
  52168=>"010000011",
  52169=>"001011000",
  52170=>"101010110",
  52171=>"111111011",
  52172=>"100000011",
  52173=>"111010010",
  52174=>"011001001",
  52175=>"000101111",
  52176=>"111111110",
  52177=>"110101111",
  52178=>"101000101",
  52179=>"110111110",
  52180=>"100010000",
  52181=>"111110111",
  52182=>"101001010",
  52183=>"001101001",
  52184=>"100000010",
  52185=>"101000110",
  52186=>"010101011",
  52187=>"000011111",
  52188=>"010001001",
  52189=>"000001110",
  52190=>"101000101",
  52191=>"000110001",
  52192=>"000110101",
  52193=>"110000100",
  52194=>"010110011",
  52195=>"000101111",
  52196=>"011110011",
  52197=>"001011010",
  52198=>"010000100",
  52199=>"000100110",
  52200=>"000001001",
  52201=>"111001011",
  52202=>"011101010",
  52203=>"010010110",
  52204=>"111100011",
  52205=>"111000100",
  52206=>"101110111",
  52207=>"101001111",
  52208=>"000001110",
  52209=>"000101001",
  52210=>"010011111",
  52211=>"110011001",
  52212=>"010000101",
  52213=>"111111101",
  52214=>"011110010",
  52215=>"110011001",
  52216=>"101010001",
  52217=>"110000100",
  52218=>"001000000",
  52219=>"000010100",
  52220=>"001111001",
  52221=>"001100000",
  52222=>"000011001",
  52223=>"111000111",
  52224=>"000000010",
  52225=>"101110110",
  52226=>"000000000",
  52227=>"000001010",
  52228=>"100010100",
  52229=>"001011111",
  52230=>"010000101",
  52231=>"001001001",
  52232=>"000000001",
  52233=>"101011111",
  52234=>"011000000",
  52235=>"111101111",
  52236=>"110110000",
  52237=>"111000001",
  52238=>"110010100",
  52239=>"011001110",
  52240=>"010010000",
  52241=>"001001000",
  52242=>"100111110",
  52243=>"010011101",
  52244=>"101010111",
  52245=>"001010111",
  52246=>"001100100",
  52247=>"100011010",
  52248=>"011010100",
  52249=>"001111010",
  52250=>"001101111",
  52251=>"111100100",
  52252=>"111101000",
  52253=>"001010100",
  52254=>"100011100",
  52255=>"011010001",
  52256=>"001001001",
  52257=>"110000011",
  52258=>"000100001",
  52259=>"101011101",
  52260=>"100100100",
  52261=>"111100011",
  52262=>"000000100",
  52263=>"000000111",
  52264=>"111101111",
  52265=>"011110000",
  52266=>"111100111",
  52267=>"001010011",
  52268=>"110111000",
  52269=>"110010101",
  52270=>"100010010",
  52271=>"001111010",
  52272=>"100111010",
  52273=>"110011000",
  52274=>"101101101",
  52275=>"001110111",
  52276=>"011000001",
  52277=>"111101010",
  52278=>"100011001",
  52279=>"001111111",
  52280=>"100100010",
  52281=>"010011110",
  52282=>"111000101",
  52283=>"001101000",
  52284=>"010100111",
  52285=>"001111101",
  52286=>"101101000",
  52287=>"001111101",
  52288=>"100100000",
  52289=>"000010101",
  52290=>"101000100",
  52291=>"011011000",
  52292=>"011111010",
  52293=>"110000010",
  52294=>"111000101",
  52295=>"100111001",
  52296=>"010110101",
  52297=>"101000010",
  52298=>"000001010",
  52299=>"001101000",
  52300=>"110101000",
  52301=>"100011111",
  52302=>"101011101",
  52303=>"110110101",
  52304=>"101001000",
  52305=>"011101010",
  52306=>"011101110",
  52307=>"110110000",
  52308=>"110110101",
  52309=>"111010100",
  52310=>"110110011",
  52311=>"111110101",
  52312=>"000001100",
  52313=>"100010110",
  52314=>"111101010",
  52315=>"101010010",
  52316=>"101001110",
  52317=>"001100010",
  52318=>"111100110",
  52319=>"001100001",
  52320=>"000100010",
  52321=>"110010111",
  52322=>"010011010",
  52323=>"000000000",
  52324=>"010110011",
  52325=>"010101011",
  52326=>"010001100",
  52327=>"000000101",
  52328=>"000010110",
  52329=>"101111101",
  52330=>"101001011",
  52331=>"000011100",
  52332=>"010111000",
  52333=>"000010100",
  52334=>"010000000",
  52335=>"000110101",
  52336=>"010000100",
  52337=>"111000011",
  52338=>"110111100",
  52339=>"000100010",
  52340=>"101111001",
  52341=>"101110101",
  52342=>"000100001",
  52343=>"100111111",
  52344=>"011111011",
  52345=>"011011111",
  52346=>"110100101",
  52347=>"110111010",
  52348=>"010111000",
  52349=>"011011001",
  52350=>"010001000",
  52351=>"010000010",
  52352=>"100001000",
  52353=>"100110111",
  52354=>"000000110",
  52355=>"101000110",
  52356=>"010001010",
  52357=>"100010111",
  52358=>"100001001",
  52359=>"000010100",
  52360=>"010011000",
  52361=>"100101001",
  52362=>"100101011",
  52363=>"010101001",
  52364=>"000000110",
  52365=>"111110111",
  52366=>"101100111",
  52367=>"110011111",
  52368=>"101011111",
  52369=>"100101010",
  52370=>"111001011",
  52371=>"000110111",
  52372=>"000000011",
  52373=>"001010001",
  52374=>"110010110",
  52375=>"101010010",
  52376=>"110110000",
  52377=>"100111100",
  52378=>"011001011",
  52379=>"000000111",
  52380=>"001011001",
  52381=>"001111011",
  52382=>"011001111",
  52383=>"101111011",
  52384=>"010100111",
  52385=>"001001100",
  52386=>"110110011",
  52387=>"000000010",
  52388=>"010000101",
  52389=>"000110111",
  52390=>"011101101",
  52391=>"001110111",
  52392=>"011111110",
  52393=>"100011000",
  52394=>"110110000",
  52395=>"000101011",
  52396=>"011101111",
  52397=>"101110101",
  52398=>"001110100",
  52399=>"011010111",
  52400=>"001010001",
  52401=>"000010011",
  52402=>"000000010",
  52403=>"101111001",
  52404=>"100011010",
  52405=>"111001100",
  52406=>"011000111",
  52407=>"100010111",
  52408=>"111001111",
  52409=>"110111110",
  52410=>"100100100",
  52411=>"011100110",
  52412=>"010000111",
  52413=>"011100110",
  52414=>"011010111",
  52415=>"100011011",
  52416=>"001011001",
  52417=>"011110100",
  52418=>"011010011",
  52419=>"000110111",
  52420=>"011001001",
  52421=>"110110111",
  52422=>"101001001",
  52423=>"111000111",
  52424=>"111000110",
  52425=>"111101100",
  52426=>"010010000",
  52427=>"111010100",
  52428=>"011010001",
  52429=>"001011001",
  52430=>"000010010",
  52431=>"111110001",
  52432=>"001101100",
  52433=>"101011100",
  52434=>"011111011",
  52435=>"011001001",
  52436=>"010000110",
  52437=>"000111100",
  52438=>"000010110",
  52439=>"010010001",
  52440=>"100111000",
  52441=>"111011000",
  52442=>"000110000",
  52443=>"111111011",
  52444=>"010000000",
  52445=>"111010011",
  52446=>"100101110",
  52447=>"101000101",
  52448=>"111011010",
  52449=>"001010011",
  52450=>"110100111",
  52451=>"100110111",
  52452=>"001001001",
  52453=>"001110110",
  52454=>"011111001",
  52455=>"111110001",
  52456=>"001110101",
  52457=>"101011100",
  52458=>"111010100",
  52459=>"010111010",
  52460=>"001100001",
  52461=>"101011100",
  52462=>"111000110",
  52463=>"000000111",
  52464=>"101110001",
  52465=>"010010010",
  52466=>"100000011",
  52467=>"100110000",
  52468=>"010011101",
  52469=>"110100010",
  52470=>"101010000",
  52471=>"110101010",
  52472=>"001101100",
  52473=>"101011111",
  52474=>"000100100",
  52475=>"000100101",
  52476=>"011011110",
  52477=>"110100110",
  52478=>"000101000",
  52479=>"010000101",
  52480=>"001100111",
  52481=>"000010111",
  52482=>"110101000",
  52483=>"011100110",
  52484=>"101101111",
  52485=>"010111100",
  52486=>"110010110",
  52487=>"101000110",
  52488=>"100001100",
  52489=>"100011000",
  52490=>"011101100",
  52491=>"111111100",
  52492=>"011011101",
  52493=>"101110110",
  52494=>"101100011",
  52495=>"000100010",
  52496=>"110001001",
  52497=>"110111000",
  52498=>"000110011",
  52499=>"111010100",
  52500=>"000010101",
  52501=>"110001011",
  52502=>"000100000",
  52503=>"001111001",
  52504=>"100011011",
  52505=>"001100100",
  52506=>"011100000",
  52507=>"000101000",
  52508=>"110101111",
  52509=>"110011001",
  52510=>"011110011",
  52511=>"110110010",
  52512=>"110101111",
  52513=>"100111101",
  52514=>"001101110",
  52515=>"000111111",
  52516=>"000000011",
  52517=>"001100011",
  52518=>"011001111",
  52519=>"100010011",
  52520=>"100000001",
  52521=>"111110001",
  52522=>"110111110",
  52523=>"100010101",
  52524=>"111000111",
  52525=>"011010100",
  52526=>"000000110",
  52527=>"101110010",
  52528=>"000010001",
  52529=>"111001001",
  52530=>"111011100",
  52531=>"110001000",
  52532=>"011001001",
  52533=>"110001001",
  52534=>"110111011",
  52535=>"000101001",
  52536=>"010101011",
  52537=>"010100101",
  52538=>"010011010",
  52539=>"001000001",
  52540=>"000000001",
  52541=>"010101000",
  52542=>"111011100",
  52543=>"000111011",
  52544=>"011001001",
  52545=>"100001001",
  52546=>"011010101",
  52547=>"000000001",
  52548=>"101110111",
  52549=>"101101100",
  52550=>"110100000",
  52551=>"001000111",
  52552=>"011011111",
  52553=>"001001111",
  52554=>"110000000",
  52555=>"000000011",
  52556=>"100100101",
  52557=>"011011011",
  52558=>"001010110",
  52559=>"000111111",
  52560=>"101011010",
  52561=>"100110111",
  52562=>"100000000",
  52563=>"010010001",
  52564=>"000000000",
  52565=>"011010101",
  52566=>"010001101",
  52567=>"111100001",
  52568=>"101001011",
  52569=>"001001110",
  52570=>"111000100",
  52571=>"000101100",
  52572=>"001111100",
  52573=>"111100001",
  52574=>"001000100",
  52575=>"111101100",
  52576=>"110100010",
  52577=>"100101011",
  52578=>"010001001",
  52579=>"101011110",
  52580=>"110100001",
  52581=>"111101010",
  52582=>"101111100",
  52583=>"000100100",
  52584=>"100100000",
  52585=>"010110000",
  52586=>"000010100",
  52587=>"000000111",
  52588=>"110111000",
  52589=>"010111000",
  52590=>"011100101",
  52591=>"110000001",
  52592=>"100001100",
  52593=>"011010010",
  52594=>"101110011",
  52595=>"001001000",
  52596=>"100011101",
  52597=>"000010010",
  52598=>"000100000",
  52599=>"001000110",
  52600=>"000001011",
  52601=>"011001000",
  52602=>"111111001",
  52603=>"101101010",
  52604=>"100101010",
  52605=>"110011001",
  52606=>"110100001",
  52607=>"000000100",
  52608=>"110101111",
  52609=>"110110100",
  52610=>"111100110",
  52611=>"001100101",
  52612=>"111101010",
  52613=>"011100010",
  52614=>"110001111",
  52615=>"010011000",
  52616=>"011101011",
  52617=>"101001001",
  52618=>"011101001",
  52619=>"000000000",
  52620=>"101100110",
  52621=>"001001001",
  52622=>"110010110",
  52623=>"001010001",
  52624=>"100001110",
  52625=>"011010000",
  52626=>"100000010",
  52627=>"001001000",
  52628=>"000011011",
  52629=>"000100101",
  52630=>"010001000",
  52631=>"110010000",
  52632=>"000000011",
  52633=>"011011001",
  52634=>"000001101",
  52635=>"110001101",
  52636=>"111011001",
  52637=>"111110101",
  52638=>"011011001",
  52639=>"101100000",
  52640=>"000111111",
  52641=>"001000010",
  52642=>"111010011",
  52643=>"010110110",
  52644=>"101001010",
  52645=>"001111001",
  52646=>"000011001",
  52647=>"100010001",
  52648=>"100010000",
  52649=>"000110001",
  52650=>"110000010",
  52651=>"111010000",
  52652=>"100101101",
  52653=>"101001110",
  52654=>"000001011",
  52655=>"110000001",
  52656=>"111100110",
  52657=>"000001001",
  52658=>"101010010",
  52659=>"110110011",
  52660=>"100111110",
  52661=>"000001111",
  52662=>"110001110",
  52663=>"100010111",
  52664=>"010001111",
  52665=>"000101101",
  52666=>"010011001",
  52667=>"110001010",
  52668=>"001101001",
  52669=>"111111011",
  52670=>"011111010",
  52671=>"001000101",
  52672=>"101101010",
  52673=>"001101100",
  52674=>"100100111",
  52675=>"101011101",
  52676=>"011011010",
  52677=>"111010000",
  52678=>"100111001",
  52679=>"011011110",
  52680=>"110011101",
  52681=>"111010011",
  52682=>"010110110",
  52683=>"011001100",
  52684=>"101000101",
  52685=>"111111100",
  52686=>"100001010",
  52687=>"101110010",
  52688=>"011110011",
  52689=>"011011001",
  52690=>"000101011",
  52691=>"010000110",
  52692=>"000001000",
  52693=>"001101101",
  52694=>"011101011",
  52695=>"111011010",
  52696=>"101001110",
  52697=>"110000000",
  52698=>"111101110",
  52699=>"010010101",
  52700=>"111010101",
  52701=>"111010001",
  52702=>"111111010",
  52703=>"110010111",
  52704=>"001100101",
  52705=>"100001000",
  52706=>"101100011",
  52707=>"001101100",
  52708=>"010000000",
  52709=>"010101000",
  52710=>"001000101",
  52711=>"100001101",
  52712=>"110111001",
  52713=>"011111110",
  52714=>"100100101",
  52715=>"110101101",
  52716=>"101010010",
  52717=>"000011110",
  52718=>"010100011",
  52719=>"111000011",
  52720=>"000100010",
  52721=>"000011110",
  52722=>"110111111",
  52723=>"110000011",
  52724=>"101000010",
  52725=>"001000010",
  52726=>"001111000",
  52727=>"101110010",
  52728=>"001101011",
  52729=>"111101110",
  52730=>"011111100",
  52731=>"110100001",
  52732=>"110111011",
  52733=>"101011100",
  52734=>"101101001",
  52735=>"100110111",
  52736=>"000011001",
  52737=>"110000011",
  52738=>"100000100",
  52739=>"100000000",
  52740=>"100110110",
  52741=>"100011101",
  52742=>"010010101",
  52743=>"001000110",
  52744=>"010001010",
  52745=>"101011000",
  52746=>"111110101",
  52747=>"000000110",
  52748=>"100001011",
  52749=>"011000010",
  52750=>"000111000",
  52751=>"000110000",
  52752=>"101011010",
  52753=>"101110100",
  52754=>"010101111",
  52755=>"111010101",
  52756=>"001011000",
  52757=>"111100010",
  52758=>"001101100",
  52759=>"100111010",
  52760=>"001101011",
  52761=>"000000011",
  52762=>"111101100",
  52763=>"110001011",
  52764=>"111011101",
  52765=>"001100111",
  52766=>"001101001",
  52767=>"001100110",
  52768=>"000011011",
  52769=>"000011011",
  52770=>"100100000",
  52771=>"111000111",
  52772=>"111101101",
  52773=>"011110101",
  52774=>"011110011",
  52775=>"000001100",
  52776=>"110010010",
  52777=>"011101010",
  52778=>"100111101",
  52779=>"110110000",
  52780=>"001101100",
  52781=>"011100111",
  52782=>"001101101",
  52783=>"001110111",
  52784=>"101100010",
  52785=>"010001101",
  52786=>"101010001",
  52787=>"010100010",
  52788=>"000111111",
  52789=>"011100110",
  52790=>"111111101",
  52791=>"001110001",
  52792=>"100001000",
  52793=>"000111011",
  52794=>"101111111",
  52795=>"111101110",
  52796=>"101011011",
  52797=>"010111110",
  52798=>"011111101",
  52799=>"001101001",
  52800=>"110110110",
  52801=>"011110111",
  52802=>"000010111",
  52803=>"111011101",
  52804=>"110101111",
  52805=>"000101011",
  52806=>"000110101",
  52807=>"000110110",
  52808=>"001000101",
  52809=>"101010010",
  52810=>"101001101",
  52811=>"110110100",
  52812=>"110001011",
  52813=>"000111100",
  52814=>"010110010",
  52815=>"100101011",
  52816=>"000110010",
  52817=>"000010111",
  52818=>"011011010",
  52819=>"011111111",
  52820=>"011010001",
  52821=>"000000110",
  52822=>"010010011",
  52823=>"001000110",
  52824=>"110000001",
  52825=>"000010001",
  52826=>"001011110",
  52827=>"001011100",
  52828=>"001000000",
  52829=>"011011111",
  52830=>"010110100",
  52831=>"111100100",
  52832=>"111010011",
  52833=>"011101100",
  52834=>"110101100",
  52835=>"110001110",
  52836=>"010011100",
  52837=>"011110111",
  52838=>"110101110",
  52839=>"001101110",
  52840=>"101011101",
  52841=>"001110001",
  52842=>"101110101",
  52843=>"010001011",
  52844=>"100110011",
  52845=>"010101100",
  52846=>"001000101",
  52847=>"111000001",
  52848=>"110011010",
  52849=>"100000011",
  52850=>"100101000",
  52851=>"011100101",
  52852=>"111110011",
  52853=>"100011101",
  52854=>"100111100",
  52855=>"000110111",
  52856=>"111100100",
  52857=>"010101110",
  52858=>"100110010",
  52859=>"011110001",
  52860=>"001001101",
  52861=>"101111010",
  52862=>"110001111",
  52863=>"110110011",
  52864=>"001100001",
  52865=>"011000010",
  52866=>"000011000",
  52867=>"001001010",
  52868=>"000011110",
  52869=>"001110110",
  52870=>"001111111",
  52871=>"101000111",
  52872=>"101100101",
  52873=>"011001100",
  52874=>"010011001",
  52875=>"110011100",
  52876=>"100100010",
  52877=>"000110000",
  52878=>"100110101",
  52879=>"101100010",
  52880=>"001100010",
  52881=>"110101011",
  52882=>"011101100",
  52883=>"001111011",
  52884=>"101111101",
  52885=>"101010011",
  52886=>"011010100",
  52887=>"111101100",
  52888=>"100111000",
  52889=>"100001111",
  52890=>"011011000",
  52891=>"010100100",
  52892=>"001101100",
  52893=>"100011010",
  52894=>"101000101",
  52895=>"111001101",
  52896=>"111000011",
  52897=>"010111011",
  52898=>"000011000",
  52899=>"010000110",
  52900=>"000111011",
  52901=>"010000000",
  52902=>"000010100",
  52903=>"110001011",
  52904=>"100100000",
  52905=>"111110010",
  52906=>"110000010",
  52907=>"100010111",
  52908=>"010101100",
  52909=>"100001000",
  52910=>"110100000",
  52911=>"111001011",
  52912=>"101101011",
  52913=>"110011010",
  52914=>"100110110",
  52915=>"011010010",
  52916=>"011011010",
  52917=>"101111011",
  52918=>"001011110",
  52919=>"011001100",
  52920=>"110000100",
  52921=>"100110011",
  52922=>"011110000",
  52923=>"100011001",
  52924=>"111010011",
  52925=>"100000010",
  52926=>"011000111",
  52927=>"111011110",
  52928=>"010101111",
  52929=>"111010001",
  52930=>"000110001",
  52931=>"110011110",
  52932=>"011001011",
  52933=>"001110000",
  52934=>"010100110",
  52935=>"111011110",
  52936=>"001100111",
  52937=>"100101100",
  52938=>"101100100",
  52939=>"100110011",
  52940=>"000001010",
  52941=>"100101101",
  52942=>"000010111",
  52943=>"010101001",
  52944=>"111000101",
  52945=>"010010000",
  52946=>"011011111",
  52947=>"010111110",
  52948=>"000011011",
  52949=>"111101111",
  52950=>"100110111",
  52951=>"101011110",
  52952=>"000110111",
  52953=>"010101010",
  52954=>"000010001",
  52955=>"011101101",
  52956=>"100001110",
  52957=>"011100010",
  52958=>"101101001",
  52959=>"000110101",
  52960=>"111001110",
  52961=>"000010100",
  52962=>"010111001",
  52963=>"011101110",
  52964=>"000101101",
  52965=>"100101001",
  52966=>"000001000",
  52967=>"010001000",
  52968=>"011101100",
  52969=>"111011100",
  52970=>"011011111",
  52971=>"000101000",
  52972=>"000110001",
  52973=>"011010100",
  52974=>"110101110",
  52975=>"000100101",
  52976=>"111000010",
  52977=>"110000010",
  52978=>"000011000",
  52979=>"111001110",
  52980=>"111110111",
  52981=>"100000000",
  52982=>"111010010",
  52983=>"000011000",
  52984=>"100010110",
  52985=>"001001100",
  52986=>"011010100",
  52987=>"000110100",
  52988=>"010111011",
  52989=>"101001001",
  52990=>"011001101",
  52991=>"001100100",
  52992=>"101001110",
  52993=>"010010010",
  52994=>"011111000",
  52995=>"101101110",
  52996=>"011010101",
  52997=>"101010010",
  52998=>"010110010",
  52999=>"000010100",
  53000=>"001100010",
  53001=>"111101011",
  53002=>"010011101",
  53003=>"000100010",
  53004=>"101011101",
  53005=>"101011111",
  53006=>"111010110",
  53007=>"100011000",
  53008=>"011011110",
  53009=>"000111111",
  53010=>"100000110",
  53011=>"011111010",
  53012=>"111001001",
  53013=>"010111000",
  53014=>"001010100",
  53015=>"010010011",
  53016=>"000001100",
  53017=>"100010101",
  53018=>"000000111",
  53019=>"111010000",
  53020=>"100001101",
  53021=>"111111111",
  53022=>"100110101",
  53023=>"100100000",
  53024=>"110010011",
  53025=>"100110110",
  53026=>"111101101",
  53027=>"000001111",
  53028=>"010011000",
  53029=>"110110011",
  53030=>"010010001",
  53031=>"001011110",
  53032=>"010110100",
  53033=>"101010100",
  53034=>"000011111",
  53035=>"000110111",
  53036=>"001001110",
  53037=>"000011011",
  53038=>"011101011",
  53039=>"010111110",
  53040=>"010111110",
  53041=>"101101001",
  53042=>"000011000",
  53043=>"001010000",
  53044=>"101110101",
  53045=>"111010010",
  53046=>"001101111",
  53047=>"110100100",
  53048=>"101010011",
  53049=>"111100011",
  53050=>"000000110",
  53051=>"001101001",
  53052=>"000000010",
  53053=>"100100111",
  53054=>"110011101",
  53055=>"100001011",
  53056=>"101011000",
  53057=>"000111001",
  53058=>"001110100",
  53059=>"110110011",
  53060=>"000100100",
  53061=>"001101101",
  53062=>"101011010",
  53063=>"010100111",
  53064=>"101010101",
  53065=>"001010000",
  53066=>"111010000",
  53067=>"011010111",
  53068=>"100010000",
  53069=>"101100001",
  53070=>"100111111",
  53071=>"011000011",
  53072=>"001010010",
  53073=>"011111011",
  53074=>"011100011",
  53075=>"100100110",
  53076=>"111110011",
  53077=>"000001100",
  53078=>"010100001",
  53079=>"011100101",
  53080=>"110100101",
  53081=>"001101111",
  53082=>"000011110",
  53083=>"000101010",
  53084=>"110000101",
  53085=>"101001110",
  53086=>"001010001",
  53087=>"000010100",
  53088=>"001111010",
  53089=>"101101000",
  53090=>"011100011",
  53091=>"100110101",
  53092=>"000011011",
  53093=>"000011010",
  53094=>"001000011",
  53095=>"001101111",
  53096=>"110011100",
  53097=>"110110101",
  53098=>"110011111",
  53099=>"101010010",
  53100=>"101000010",
  53101=>"110001111",
  53102=>"001001111",
  53103=>"010011101",
  53104=>"011010101",
  53105=>"100011011",
  53106=>"110111001",
  53107=>"101100110",
  53108=>"000011000",
  53109=>"100101111",
  53110=>"011010110",
  53111=>"011001100",
  53112=>"011111101",
  53113=>"111100110",
  53114=>"101100011",
  53115=>"011111110",
  53116=>"000000101",
  53117=>"010001000",
  53118=>"111011000",
  53119=>"101011101",
  53120=>"111011101",
  53121=>"000111100",
  53122=>"000000001",
  53123=>"111111101",
  53124=>"001011001",
  53125=>"110100001",
  53126=>"110010001",
  53127=>"110000000",
  53128=>"011011011",
  53129=>"110101111",
  53130=>"111111000",
  53131=>"101110010",
  53132=>"111011101",
  53133=>"011010010",
  53134=>"110011111",
  53135=>"010010001",
  53136=>"000011011",
  53137=>"010011110",
  53138=>"111111011",
  53139=>"010000001",
  53140=>"000000110",
  53141=>"011010011",
  53142=>"110000001",
  53143=>"111001100",
  53144=>"000001011",
  53145=>"111010010",
  53146=>"000000111",
  53147=>"100010001",
  53148=>"011101011",
  53149=>"111000000",
  53150=>"011110111",
  53151=>"011110010",
  53152=>"110101101",
  53153=>"010110111",
  53154=>"110110010",
  53155=>"111010001",
  53156=>"010010000",
  53157=>"010101011",
  53158=>"000010011",
  53159=>"001001001",
  53160=>"100001100",
  53161=>"000000000",
  53162=>"110101101",
  53163=>"011111100",
  53164=>"110000110",
  53165=>"000000110",
  53166=>"110100111",
  53167=>"010111110",
  53168=>"111010110",
  53169=>"001101010",
  53170=>"111111100",
  53171=>"100101100",
  53172=>"010110000",
  53173=>"010001011",
  53174=>"101010111",
  53175=>"011101111",
  53176=>"000101111",
  53177=>"100100000",
  53178=>"111100111",
  53179=>"110101110",
  53180=>"011001010",
  53181=>"100010011",
  53182=>"101001101",
  53183=>"000001010",
  53184=>"010010100",
  53185=>"001100101",
  53186=>"111101100",
  53187=>"101101111",
  53188=>"000000010",
  53189=>"100000010",
  53190=>"111001100",
  53191=>"101001101",
  53192=>"111101010",
  53193=>"001110001",
  53194=>"001111110",
  53195=>"111011010",
  53196=>"010010000",
  53197=>"010000000",
  53198=>"101110001",
  53199=>"011010111",
  53200=>"111111000",
  53201=>"111001011",
  53202=>"101100011",
  53203=>"010100101",
  53204=>"111100111",
  53205=>"100011011",
  53206=>"010100011",
  53207=>"010010010",
  53208=>"001010101",
  53209=>"001010011",
  53210=>"010000001",
  53211=>"010100110",
  53212=>"000010011",
  53213=>"010100111",
  53214=>"000111110",
  53215=>"100011000",
  53216=>"100010101",
  53217=>"000000010",
  53218=>"001001111",
  53219=>"110001010",
  53220=>"101010110",
  53221=>"111000011",
  53222=>"100111100",
  53223=>"101010101",
  53224=>"010110001",
  53225=>"000101111",
  53226=>"111000110",
  53227=>"100100001",
  53228=>"100100010",
  53229=>"110100000",
  53230=>"001000111",
  53231=>"101100010",
  53232=>"010111000",
  53233=>"011100110",
  53234=>"100000001",
  53235=>"000110010",
  53236=>"111011011",
  53237=>"011111100",
  53238=>"110010110",
  53239=>"010010100",
  53240=>"001101111",
  53241=>"101100111",
  53242=>"011010001",
  53243=>"010100111",
  53244=>"010000101",
  53245=>"101111101",
  53246=>"111101111",
  53247=>"100100111",
  53248=>"010100000",
  53249=>"010101001",
  53250=>"111011111",
  53251=>"110011010",
  53252=>"101100011",
  53253=>"001010111",
  53254=>"001010100",
  53255=>"010000100",
  53256=>"100000001",
  53257=>"001010000",
  53258=>"101010011",
  53259=>"111100101",
  53260=>"000010000",
  53261=>"000000100",
  53262=>"111000000",
  53263=>"000100110",
  53264=>"010011001",
  53265=>"110110001",
  53266=>"011001000",
  53267=>"111100100",
  53268=>"110000110",
  53269=>"101011011",
  53270=>"111001001",
  53271=>"111000111",
  53272=>"000101011",
  53273=>"101001010",
  53274=>"110000001",
  53275=>"110001100",
  53276=>"111100101",
  53277=>"101101000",
  53278=>"000100000",
  53279=>"010001001",
  53280=>"000011011",
  53281=>"110111111",
  53282=>"111101010",
  53283=>"010000011",
  53284=>"011111111",
  53285=>"000100100",
  53286=>"110110011",
  53287=>"000000110",
  53288=>"111000000",
  53289=>"010010100",
  53290=>"100010101",
  53291=>"011100110",
  53292=>"110110101",
  53293=>"100111110",
  53294=>"000110011",
  53295=>"100001011",
  53296=>"110100100",
  53297=>"110101010",
  53298=>"101001000",
  53299=>"111011110",
  53300=>"000010110",
  53301=>"000011101",
  53302=>"111101100",
  53303=>"001100110",
  53304=>"001001101",
  53305=>"101110110",
  53306=>"001001000",
  53307=>"111110101",
  53308=>"011100100",
  53309=>"111111011",
  53310=>"111011111",
  53311=>"011011111",
  53312=>"111101010",
  53313=>"001010110",
  53314=>"011011101",
  53315=>"110110111",
  53316=>"111100100",
  53317=>"000110010",
  53318=>"011100001",
  53319=>"111010111",
  53320=>"001100011",
  53321=>"000011111",
  53322=>"010100000",
  53323=>"001000100",
  53324=>"000011110",
  53325=>"011010011",
  53326=>"001110110",
  53327=>"010011100",
  53328=>"010101001",
  53329=>"111001000",
  53330=>"000101010",
  53331=>"101111001",
  53332=>"010100110",
  53333=>"001111110",
  53334=>"011101101",
  53335=>"001000101",
  53336=>"111000011",
  53337=>"111110110",
  53338=>"001010001",
  53339=>"011011001",
  53340=>"101110010",
  53341=>"000101101",
  53342=>"000111111",
  53343=>"011101000",
  53344=>"100001010",
  53345=>"100111111",
  53346=>"111001111",
  53347=>"001101100",
  53348=>"000000101",
  53349=>"111111010",
  53350=>"101010010",
  53351=>"101110000",
  53352=>"000010011",
  53353=>"000011011",
  53354=>"111010111",
  53355=>"111001101",
  53356=>"100110010",
  53357=>"000010111",
  53358=>"111000010",
  53359=>"101101111",
  53360=>"100111001",
  53361=>"000011100",
  53362=>"011110000",
  53363=>"000100001",
  53364=>"101110010",
  53365=>"100111101",
  53366=>"111110010",
  53367=>"010011010",
  53368=>"011000001",
  53369=>"110011111",
  53370=>"110000000",
  53371=>"001000101",
  53372=>"111101110",
  53373=>"000001111",
  53374=>"001001110",
  53375=>"110111100",
  53376=>"011100110",
  53377=>"100001011",
  53378=>"111001110",
  53379=>"000010111",
  53380=>"011101111",
  53381=>"001000001",
  53382=>"100101011",
  53383=>"110111000",
  53384=>"001110111",
  53385=>"110001000",
  53386=>"001000110",
  53387=>"001101001",
  53388=>"110011110",
  53389=>"011011000",
  53390=>"110000111",
  53391=>"000111101",
  53392=>"110001111",
  53393=>"111110011",
  53394=>"001011011",
  53395=>"011011101",
  53396=>"110100001",
  53397=>"110011101",
  53398=>"000010100",
  53399=>"010111000",
  53400=>"011110010",
  53401=>"010101000",
  53402=>"100101100",
  53403=>"101011111",
  53404=>"001000100",
  53405=>"000000101",
  53406=>"000000001",
  53407=>"000000011",
  53408=>"000001010",
  53409=>"111110100",
  53410=>"101110000",
  53411=>"110110100",
  53412=>"101010000",
  53413=>"010101001",
  53414=>"111010101",
  53415=>"100001101",
  53416=>"010101100",
  53417=>"001100110",
  53418=>"101100000",
  53419=>"001101111",
  53420=>"111000010",
  53421=>"111110110",
  53422=>"110010011",
  53423=>"000000010",
  53424=>"010101010",
  53425=>"110001001",
  53426=>"011100011",
  53427=>"110111101",
  53428=>"111110111",
  53429=>"101100001",
  53430=>"010101111",
  53431=>"100011101",
  53432=>"000000011",
  53433=>"100111100",
  53434=>"111000101",
  53435=>"100001111",
  53436=>"101000111",
  53437=>"010111000",
  53438=>"110001111",
  53439=>"101110000",
  53440=>"000010101",
  53441=>"110110111",
  53442=>"111001011",
  53443=>"001110101",
  53444=>"000010000",
  53445=>"001100011",
  53446=>"100011001",
  53447=>"001010010",
  53448=>"010100001",
  53449=>"010001011",
  53450=>"011100000",
  53451=>"110110110",
  53452=>"011110001",
  53453=>"111000011",
  53454=>"111100011",
  53455=>"000110001",
  53456=>"110110010",
  53457=>"000011001",
  53458=>"110111111",
  53459=>"001000101",
  53460=>"111001100",
  53461=>"001010000",
  53462=>"000101110",
  53463=>"001000110",
  53464=>"001110111",
  53465=>"100110011",
  53466=>"011011110",
  53467=>"010000000",
  53468=>"010010010",
  53469=>"001100001",
  53470=>"001101110",
  53471=>"110000000",
  53472=>"110010110",
  53473=>"101101000",
  53474=>"011011101",
  53475=>"101101100",
  53476=>"100000100",
  53477=>"111101001",
  53478=>"001110111",
  53479=>"000001101",
  53480=>"110001000",
  53481=>"111110100",
  53482=>"000001000",
  53483=>"000010111",
  53484=>"001010110",
  53485=>"001011111",
  53486=>"110111100",
  53487=>"011101101",
  53488=>"000001100",
  53489=>"110001001",
  53490=>"100001011",
  53491=>"010110100",
  53492=>"011111000",
  53493=>"100111001",
  53494=>"011100010",
  53495=>"110000011",
  53496=>"011110111",
  53497=>"010011110",
  53498=>"011011011",
  53499=>"101101111",
  53500=>"101100101",
  53501=>"100100110",
  53502=>"110001001",
  53503=>"010111001",
  53504=>"011010110",
  53505=>"100111000",
  53506=>"100000001",
  53507=>"101111000",
  53508=>"001010000",
  53509=>"110001101",
  53510=>"001000011",
  53511=>"001111110",
  53512=>"111111011",
  53513=>"001010100",
  53514=>"101111100",
  53515=>"010111111",
  53516=>"011001101",
  53517=>"100001110",
  53518=>"011101011",
  53519=>"111000001",
  53520=>"001010010",
  53521=>"010101111",
  53522=>"111111111",
  53523=>"011111111",
  53524=>"100100000",
  53525=>"110100010",
  53526=>"101011000",
  53527=>"001111010",
  53528=>"100111000",
  53529=>"001110000",
  53530=>"011001101",
  53531=>"001001101",
  53532=>"000110111",
  53533=>"110000110",
  53534=>"100011001",
  53535=>"010111000",
  53536=>"011110111",
  53537=>"110001010",
  53538=>"011010011",
  53539=>"000100011",
  53540=>"011110110",
  53541=>"001100100",
  53542=>"101111100",
  53543=>"010111111",
  53544=>"110010111",
  53545=>"001001111",
  53546=>"110111111",
  53547=>"100101001",
  53548=>"101001111",
  53549=>"001001010",
  53550=>"111011110",
  53551=>"001111010",
  53552=>"001000110",
  53553=>"100011111",
  53554=>"000110001",
  53555=>"001010010",
  53556=>"101110001",
  53557=>"011111000",
  53558=>"110111010",
  53559=>"001111111",
  53560=>"011000000",
  53561=>"011100110",
  53562=>"100110000",
  53563=>"110100011",
  53564=>"100001010",
  53565=>"110100011",
  53566=>"111110001",
  53567=>"101011100",
  53568=>"011101011",
  53569=>"011001101",
  53570=>"000100100",
  53571=>"000010011",
  53572=>"001010110",
  53573=>"111010110",
  53574=>"101011100",
  53575=>"011110110",
  53576=>"111001110",
  53577=>"100100001",
  53578=>"000001111",
  53579=>"010001000",
  53580=>"100100001",
  53581=>"010010000",
  53582=>"010100111",
  53583=>"110011001",
  53584=>"101011110",
  53585=>"000000110",
  53586=>"101100110",
  53587=>"010010011",
  53588=>"111111000",
  53589=>"101001110",
  53590=>"011100001",
  53591=>"001010110",
  53592=>"101111110",
  53593=>"111101011",
  53594=>"110101001",
  53595=>"100011110",
  53596=>"101110100",
  53597=>"001001010",
  53598=>"110011110",
  53599=>"011000100",
  53600=>"010001000",
  53601=>"001011110",
  53602=>"001101101",
  53603=>"101001101",
  53604=>"000111000",
  53605=>"100101110",
  53606=>"001100101",
  53607=>"011100000",
  53608=>"000110111",
  53609=>"001111110",
  53610=>"000010011",
  53611=>"000000110",
  53612=>"010101001",
  53613=>"011100010",
  53614=>"110000111",
  53615=>"100100001",
  53616=>"101010000",
  53617=>"010100111",
  53618=>"100101000",
  53619=>"001111101",
  53620=>"101010101",
  53621=>"111011101",
  53622=>"101011111",
  53623=>"001110101",
  53624=>"010010100",
  53625=>"010010011",
  53626=>"110000010",
  53627=>"110110111",
  53628=>"011011100",
  53629=>"100000110",
  53630=>"000000110",
  53631=>"100100110",
  53632=>"000111001",
  53633=>"001000000",
  53634=>"111010110",
  53635=>"101110000",
  53636=>"111111000",
  53637=>"010100010",
  53638=>"111111111",
  53639=>"110111000",
  53640=>"111010100",
  53641=>"110101101",
  53642=>"110000001",
  53643=>"101000010",
  53644=>"001001100",
  53645=>"010000011",
  53646=>"111010001",
  53647=>"100011011",
  53648=>"111101110",
  53649=>"001111000",
  53650=>"101010101",
  53651=>"101010001",
  53652=>"000000101",
  53653=>"001011101",
  53654=>"000011100",
  53655=>"010111000",
  53656=>"100011010",
  53657=>"110001001",
  53658=>"111001000",
  53659=>"001011000",
  53660=>"000010100",
  53661=>"000100000",
  53662=>"110000100",
  53663=>"100010100",
  53664=>"111001110",
  53665=>"000011001",
  53666=>"100010110",
  53667=>"000100110",
  53668=>"001000000",
  53669=>"111010111",
  53670=>"111110101",
  53671=>"111000001",
  53672=>"011001000",
  53673=>"110100111",
  53674=>"110111011",
  53675=>"010000000",
  53676=>"011110111",
  53677=>"100001010",
  53678=>"000110000",
  53679=>"010100000",
  53680=>"100010100",
  53681=>"100000000",
  53682=>"011101001",
  53683=>"010110010",
  53684=>"111001110",
  53685=>"001111000",
  53686=>"110000111",
  53687=>"001110001",
  53688=>"001111101",
  53689=>"001001111",
  53690=>"111001011",
  53691=>"000100011",
  53692=>"001100100",
  53693=>"010101001",
  53694=>"111001001",
  53695=>"110010100",
  53696=>"101001011",
  53697=>"111101111",
  53698=>"111100010",
  53699=>"101101001",
  53700=>"111111011",
  53701=>"110110001",
  53702=>"110111001",
  53703=>"010101100",
  53704=>"101011100",
  53705=>"011110000",
  53706=>"110100111",
  53707=>"111001011",
  53708=>"111010101",
  53709=>"010000110",
  53710=>"110001000",
  53711=>"111100011",
  53712=>"000111001",
  53713=>"011110101",
  53714=>"001100111",
  53715=>"111101111",
  53716=>"111101111",
  53717=>"000111101",
  53718=>"000110010",
  53719=>"010000110",
  53720=>"001110011",
  53721=>"101001101",
  53722=>"010011000",
  53723=>"000111111",
  53724=>"110110001",
  53725=>"011100110",
  53726=>"110000000",
  53727=>"001101100",
  53728=>"011111101",
  53729=>"000111011",
  53730=>"101101001",
  53731=>"010111100",
  53732=>"000100110",
  53733=>"110010100",
  53734=>"110001100",
  53735=>"010011111",
  53736=>"011100101",
  53737=>"101011101",
  53738=>"011010100",
  53739=>"011000101",
  53740=>"000000001",
  53741=>"111111101",
  53742=>"011101111",
  53743=>"110010101",
  53744=>"111001101",
  53745=>"011110001",
  53746=>"100111101",
  53747=>"011100000",
  53748=>"000100001",
  53749=>"100010100",
  53750=>"001100110",
  53751=>"100000101",
  53752=>"010010000",
  53753=>"111101100",
  53754=>"110010100",
  53755=>"001000010",
  53756=>"110010100",
  53757=>"111110110",
  53758=>"010011000",
  53759=>"001100001",
  53760=>"000111010",
  53761=>"010111001",
  53762=>"101011111",
  53763=>"110000010",
  53764=>"010101010",
  53765=>"111101111",
  53766=>"010001010",
  53767=>"111111111",
  53768=>"010110001",
  53769=>"001100000",
  53770=>"011000100",
  53771=>"000001000",
  53772=>"110100001",
  53773=>"000101100",
  53774=>"000110101",
  53775=>"100010111",
  53776=>"111101110",
  53777=>"101111000",
  53778=>"100000110",
  53779=>"101000111",
  53780=>"110010111",
  53781=>"000111101",
  53782=>"110011001",
  53783=>"100010111",
  53784=>"110111010",
  53785=>"101001110",
  53786=>"000100000",
  53787=>"100101111",
  53788=>"010101011",
  53789=>"100100100",
  53790=>"011010010",
  53791=>"100110101",
  53792=>"000011011",
  53793=>"110110010",
  53794=>"011010100",
  53795=>"101001111",
  53796=>"000010111",
  53797=>"110000100",
  53798=>"111001110",
  53799=>"110110010",
  53800=>"001001100",
  53801=>"110010101",
  53802=>"101110011",
  53803=>"011000000",
  53804=>"110110010",
  53805=>"010100110",
  53806=>"101001011",
  53807=>"000110011",
  53808=>"001011001",
  53809=>"100111100",
  53810=>"010000111",
  53811=>"111101011",
  53812=>"100110010",
  53813=>"111110001",
  53814=>"010000101",
  53815=>"100001100",
  53816=>"110101001",
  53817=>"101011100",
  53818=>"100111000",
  53819=>"010111010",
  53820=>"101011011",
  53821=>"001001101",
  53822=>"001001100",
  53823=>"100101111",
  53824=>"110011101",
  53825=>"110110001",
  53826=>"111000100",
  53827=>"001111011",
  53828=>"110110100",
  53829=>"100000011",
  53830=>"111000001",
  53831=>"101001110",
  53832=>"101100010",
  53833=>"111110011",
  53834=>"011000100",
  53835=>"001100101",
  53836=>"110000101",
  53837=>"110000000",
  53838=>"000111111",
  53839=>"101010111",
  53840=>"101101001",
  53841=>"010000010",
  53842=>"100100110",
  53843=>"000101101",
  53844=>"001010011",
  53845=>"100001010",
  53846=>"101100011",
  53847=>"000011110",
  53848=>"010110010",
  53849=>"110100101",
  53850=>"010001110",
  53851=>"111101110",
  53852=>"011111011",
  53853=>"000110011",
  53854=>"100001111",
  53855=>"111101100",
  53856=>"001000100",
  53857=>"111100000",
  53858=>"100100010",
  53859=>"111101110",
  53860=>"001000101",
  53861=>"010111001",
  53862=>"011100011",
  53863=>"100000000",
  53864=>"101000001",
  53865=>"000100001",
  53866=>"010111111",
  53867=>"000001100",
  53868=>"010011010",
  53869=>"001010101",
  53870=>"000011011",
  53871=>"100010011",
  53872=>"010101011",
  53873=>"101010111",
  53874=>"011010111",
  53875=>"100000001",
  53876=>"100110001",
  53877=>"111110010",
  53878=>"001010111",
  53879=>"111110110",
  53880=>"000110111",
  53881=>"111001101",
  53882=>"110110001",
  53883=>"010001111",
  53884=>"000101111",
  53885=>"000001010",
  53886=>"001111001",
  53887=>"011100111",
  53888=>"110101110",
  53889=>"110011100",
  53890=>"010010101",
  53891=>"100001000",
  53892=>"110000101",
  53893=>"000011010",
  53894=>"001100000",
  53895=>"001000011",
  53896=>"001101110",
  53897=>"010000100",
  53898=>"010101111",
  53899=>"010110011",
  53900=>"101001001",
  53901=>"100000011",
  53902=>"110110110",
  53903=>"111100001",
  53904=>"111110110",
  53905=>"111010101",
  53906=>"110110111",
  53907=>"011100110",
  53908=>"111100110",
  53909=>"101101000",
  53910=>"010111100",
  53911=>"010001000",
  53912=>"110111101",
  53913=>"001101100",
  53914=>"111100011",
  53915=>"111000001",
  53916=>"011100000",
  53917=>"001010111",
  53918=>"010010000",
  53919=>"110110000",
  53920=>"011100001",
  53921=>"101000110",
  53922=>"110000111",
  53923=>"000110010",
  53924=>"100011000",
  53925=>"100111111",
  53926=>"110111101",
  53927=>"110000110",
  53928=>"001101100",
  53929=>"111101000",
  53930=>"110010010",
  53931=>"111100011",
  53932=>"011101100",
  53933=>"000101000",
  53934=>"011100010",
  53935=>"100010001",
  53936=>"111100100",
  53937=>"100010100",
  53938=>"010001000",
  53939=>"001100111",
  53940=>"111000110",
  53941=>"111011100",
  53942=>"000000101",
  53943=>"010110110",
  53944=>"010111111",
  53945=>"011011000",
  53946=>"011101001",
  53947=>"110000001",
  53948=>"001110011",
  53949=>"000101000",
  53950=>"000100010",
  53951=>"100001100",
  53952=>"010001001",
  53953=>"010001000",
  53954=>"101111010",
  53955=>"010101000",
  53956=>"100100100",
  53957=>"110101100",
  53958=>"110010010",
  53959=>"001011000",
  53960=>"101100011",
  53961=>"001000100",
  53962=>"000000011",
  53963=>"000111011",
  53964=>"111001111",
  53965=>"001111111",
  53966=>"100100011",
  53967=>"111001101",
  53968=>"000100000",
  53969=>"110110111",
  53970=>"111100010",
  53971=>"100001000",
  53972=>"000010100",
  53973=>"011011101",
  53974=>"110100011",
  53975=>"101000100",
  53976=>"000001010",
  53977=>"101111110",
  53978=>"010111011",
  53979=>"001011100",
  53980=>"101101101",
  53981=>"010000011",
  53982=>"110011000",
  53983=>"000011000",
  53984=>"100000100",
  53985=>"110111011",
  53986=>"001000111",
  53987=>"110110001",
  53988=>"000001011",
  53989=>"010111100",
  53990=>"011111010",
  53991=>"011001001",
  53992=>"100000111",
  53993=>"111110111",
  53994=>"111000000",
  53995=>"001101011",
  53996=>"111001000",
  53997=>"000001100",
  53998=>"000101000",
  53999=>"011111001",
  54000=>"101110111",
  54001=>"110110011",
  54002=>"101101111",
  54003=>"101010011",
  54004=>"111101111",
  54005=>"010010010",
  54006=>"110010101",
  54007=>"010101101",
  54008=>"001011011",
  54009=>"110001011",
  54010=>"110101100",
  54011=>"101010011",
  54012=>"101010101",
  54013=>"100001010",
  54014=>"011110101",
  54015=>"101101011",
  54016=>"101010100",
  54017=>"100010011",
  54018=>"011000100",
  54019=>"100000010",
  54020=>"111010010",
  54021=>"001000101",
  54022=>"100011000",
  54023=>"000111011",
  54024=>"001111011",
  54025=>"110010111",
  54026=>"001100110",
  54027=>"110010010",
  54028=>"101010100",
  54029=>"101110101",
  54030=>"110010001",
  54031=>"101111101",
  54032=>"010010001",
  54033=>"010011101",
  54034=>"001111001",
  54035=>"000111111",
  54036=>"110110110",
  54037=>"100111110",
  54038=>"010010001",
  54039=>"000101101",
  54040=>"000011000",
  54041=>"000111111",
  54042=>"010111010",
  54043=>"010110111",
  54044=>"100011010",
  54045=>"110110011",
  54046=>"110000010",
  54047=>"011001000",
  54048=>"110011101",
  54049=>"110000010",
  54050=>"010001110",
  54051=>"101000001",
  54052=>"111000111",
  54053=>"100000001",
  54054=>"000010011",
  54055=>"011101110",
  54056=>"000000111",
  54057=>"111011111",
  54058=>"001111110",
  54059=>"110110111",
  54060=>"000111001",
  54061=>"000001000",
  54062=>"000000001",
  54063=>"101001000",
  54064=>"001011000",
  54065=>"011101100",
  54066=>"001010111",
  54067=>"000111100",
  54068=>"111001101",
  54069=>"111001001",
  54070=>"000000000",
  54071=>"000111010",
  54072=>"110100010",
  54073=>"010100110",
  54074=>"000001010",
  54075=>"101100111",
  54076=>"100100001",
  54077=>"101110011",
  54078=>"100000100",
  54079=>"111011110",
  54080=>"110010001",
  54081=>"010111000",
  54082=>"111011100",
  54083=>"001111100",
  54084=>"101100011",
  54085=>"100010100",
  54086=>"010000010",
  54087=>"101001110",
  54088=>"000010010",
  54089=>"000011110",
  54090=>"011111010",
  54091=>"000000111",
  54092=>"111000011",
  54093=>"000010001",
  54094=>"100000010",
  54095=>"011011011",
  54096=>"011101010",
  54097=>"000101010",
  54098=>"110101000",
  54099=>"010111010",
  54100=>"001000101",
  54101=>"100000111",
  54102=>"000101111",
  54103=>"111111000",
  54104=>"101101011",
  54105=>"111001100",
  54106=>"111111001",
  54107=>"010101101",
  54108=>"000010101",
  54109=>"101011010",
  54110=>"110000101",
  54111=>"001100001",
  54112=>"000010100",
  54113=>"101111001",
  54114=>"111001001",
  54115=>"001010110",
  54116=>"000010101",
  54117=>"010111101",
  54118=>"110000011",
  54119=>"001000011",
  54120=>"000001001",
  54121=>"000001001",
  54122=>"001011110",
  54123=>"000101000",
  54124=>"010110111",
  54125=>"111100001",
  54126=>"111001100",
  54127=>"111110010",
  54128=>"100000000",
  54129=>"000001010",
  54130=>"001001011",
  54131=>"010110101",
  54132=>"010001110",
  54133=>"010111101",
  54134=>"100010001",
  54135=>"100100101",
  54136=>"111000010",
  54137=>"110011100",
  54138=>"101100101",
  54139=>"011011101",
  54140=>"010001101",
  54141=>"000111101",
  54142=>"001001000",
  54143=>"111010101",
  54144=>"100010010",
  54145=>"111110100",
  54146=>"000111101",
  54147=>"111101010",
  54148=>"000100100",
  54149=>"010001000",
  54150=>"011110111",
  54151=>"000000000",
  54152=>"110000101",
  54153=>"000110010",
  54154=>"001010110",
  54155=>"001010110",
  54156=>"001011000",
  54157=>"000000000",
  54158=>"110110000",
  54159=>"100001010",
  54160=>"110000001",
  54161=>"111101000",
  54162=>"100101000",
  54163=>"011010101",
  54164=>"100101011",
  54165=>"001010111",
  54166=>"110100111",
  54167=>"011010000",
  54168=>"010011001",
  54169=>"000001001",
  54170=>"100110101",
  54171=>"100000010",
  54172=>"100000001",
  54173=>"011100110",
  54174=>"000101000",
  54175=>"001000101",
  54176=>"010111110",
  54177=>"000011011",
  54178=>"110101110",
  54179=>"000100100",
  54180=>"101001000",
  54181=>"101101101",
  54182=>"100111000",
  54183=>"100100101",
  54184=>"001101001",
  54185=>"101111101",
  54186=>"010000101",
  54187=>"001110100",
  54188=>"000000110",
  54189=>"010000000",
  54190=>"001101001",
  54191=>"011100101",
  54192=>"010000100",
  54193=>"011111110",
  54194=>"010100110",
  54195=>"110010000",
  54196=>"101100110",
  54197=>"100100010",
  54198=>"011000110",
  54199=>"001011111",
  54200=>"000000110",
  54201=>"101100110",
  54202=>"011010111",
  54203=>"011000110",
  54204=>"000000101",
  54205=>"010110001",
  54206=>"010001101",
  54207=>"000010111",
  54208=>"001110110",
  54209=>"110101101",
  54210=>"100101110",
  54211=>"001110010",
  54212=>"001110111",
  54213=>"111111100",
  54214=>"001110000",
  54215=>"111001111",
  54216=>"000100011",
  54217=>"010111110",
  54218=>"011010001",
  54219=>"111110001",
  54220=>"011000100",
  54221=>"101101011",
  54222=>"011011100",
  54223=>"000110111",
  54224=>"101011000",
  54225=>"110101101",
  54226=>"011000111",
  54227=>"100001000",
  54228=>"101000000",
  54229=>"010000010",
  54230=>"000100011",
  54231=>"111010111",
  54232=>"101001111",
  54233=>"101001001",
  54234=>"100000101",
  54235=>"111110111",
  54236=>"000001111",
  54237=>"110111001",
  54238=>"000010011",
  54239=>"001101100",
  54240=>"011001101",
  54241=>"010000001",
  54242=>"010010101",
  54243=>"101110000",
  54244=>"011110101",
  54245=>"100101000",
  54246=>"001010010",
  54247=>"100100010",
  54248=>"100100101",
  54249=>"010100100",
  54250=>"001001101",
  54251=>"101000010",
  54252=>"101000000",
  54253=>"100011100",
  54254=>"110011010",
  54255=>"011111000",
  54256=>"011110111",
  54257=>"111100000",
  54258=>"111111101",
  54259=>"011001011",
  54260=>"011100000",
  54261=>"000001010",
  54262=>"111110010",
  54263=>"001000101",
  54264=>"010100110",
  54265=>"110111100",
  54266=>"000110011",
  54267=>"111111101",
  54268=>"000110101",
  54269=>"011100110",
  54270=>"001000010",
  54271=>"001110101",
  54272=>"110111100",
  54273=>"100101101",
  54274=>"111111100",
  54275=>"100001011",
  54276=>"000001000",
  54277=>"110101110",
  54278=>"100011001",
  54279=>"010010011",
  54280=>"001111101",
  54281=>"111110011",
  54282=>"001000111",
  54283=>"100111111",
  54284=>"001011110",
  54285=>"010100111",
  54286=>"010110000",
  54287=>"111111001",
  54288=>"100001000",
  54289=>"110010011",
  54290=>"101100000",
  54291=>"111101001",
  54292=>"111111011",
  54293=>"000100111",
  54294=>"001100010",
  54295=>"111010001",
  54296=>"111011111",
  54297=>"000100101",
  54298=>"101010101",
  54299=>"000111001",
  54300=>"110111010",
  54301=>"100000000",
  54302=>"100000110",
  54303=>"110011001",
  54304=>"111111001",
  54305=>"110000000",
  54306=>"110000001",
  54307=>"010111010",
  54308=>"111101100",
  54309=>"010010111",
  54310=>"111111010",
  54311=>"111110101",
  54312=>"000100111",
  54313=>"111010110",
  54314=>"010001001",
  54315=>"110100111",
  54316=>"111010000",
  54317=>"001011101",
  54318=>"101001111",
  54319=>"101100101",
  54320=>"000010001",
  54321=>"111100110",
  54322=>"000001110",
  54323=>"111111011",
  54324=>"111011111",
  54325=>"001110010",
  54326=>"110101000",
  54327=>"001101000",
  54328=>"000010111",
  54329=>"101001110",
  54330=>"000000011",
  54331=>"101000101",
  54332=>"111111010",
  54333=>"000010010",
  54334=>"101110010",
  54335=>"010010111",
  54336=>"010101000",
  54337=>"010110000",
  54338=>"000110000",
  54339=>"111101011",
  54340=>"110001000",
  54341=>"111110010",
  54342=>"101110100",
  54343=>"001111100",
  54344=>"100011100",
  54345=>"001011110",
  54346=>"100000110",
  54347=>"110101100",
  54348=>"101001111",
  54349=>"110111011",
  54350=>"010100001",
  54351=>"101011000",
  54352=>"001110100",
  54353=>"011000101",
  54354=>"100001100",
  54355=>"010011000",
  54356=>"111111110",
  54357=>"000001001",
  54358=>"010001111",
  54359=>"011010010",
  54360=>"011010000",
  54361=>"110110110",
  54362=>"011111101",
  54363=>"010011001",
  54364=>"001100111",
  54365=>"001000010",
  54366=>"010111101",
  54367=>"101110001",
  54368=>"001001001",
  54369=>"101011000",
  54370=>"011001000",
  54371=>"001101010",
  54372=>"011010101",
  54373=>"110001101",
  54374=>"100011001",
  54375=>"010010110",
  54376=>"111100001",
  54377=>"111000010",
  54378=>"011010111",
  54379=>"011010100",
  54380=>"010100111",
  54381=>"010001000",
  54382=>"100101001",
  54383=>"000101001",
  54384=>"010101011",
  54385=>"010100010",
  54386=>"010101111",
  54387=>"010001101",
  54388=>"000100100",
  54389=>"101111000",
  54390=>"111101111",
  54391=>"100101000",
  54392=>"001100111",
  54393=>"001001001",
  54394=>"101111011",
  54395=>"111001001",
  54396=>"101000111",
  54397=>"111011010",
  54398=>"111100000",
  54399=>"000010001",
  54400=>"111000100",
  54401=>"110010011",
  54402=>"000111101",
  54403=>"011100000",
  54404=>"100010110",
  54405=>"101011110",
  54406=>"011011110",
  54407=>"000011000",
  54408=>"011001010",
  54409=>"101010010",
  54410=>"101011011",
  54411=>"111001101",
  54412=>"100101110",
  54413=>"110111110",
  54414=>"100000000",
  54415=>"101111111",
  54416=>"000000101",
  54417=>"101001010",
  54418=>"111111101",
  54419=>"000000010",
  54420=>"010110110",
  54421=>"101111000",
  54422=>"111111010",
  54423=>"110011110",
  54424=>"000001000",
  54425=>"111110111",
  54426=>"001000000",
  54427=>"000101011",
  54428=>"010111101",
  54429=>"111100000",
  54430=>"010111100",
  54431=>"101111100",
  54432=>"111011101",
  54433=>"010001110",
  54434=>"111101111",
  54435=>"011101010",
  54436=>"100100110",
  54437=>"111010010",
  54438=>"111111000",
  54439=>"110101000",
  54440=>"111000100",
  54441=>"110001100",
  54442=>"101101000",
  54443=>"010010010",
  54444=>"110011101",
  54445=>"111100001",
  54446=>"100111101",
  54447=>"110110111",
  54448=>"011011001",
  54449=>"110010011",
  54450=>"010011100",
  54451=>"111101101",
  54452=>"100111111",
  54453=>"000000010",
  54454=>"111111101",
  54455=>"011111111",
  54456=>"001011110",
  54457=>"000001000",
  54458=>"111010011",
  54459=>"010111010",
  54460=>"000110101",
  54461=>"101011101",
  54462=>"001100011",
  54463=>"101010100",
  54464=>"100110001",
  54465=>"101100110",
  54466=>"100111010",
  54467=>"000000110",
  54468=>"111111100",
  54469=>"010000000",
  54470=>"110111001",
  54471=>"001011110",
  54472=>"000100001",
  54473=>"010111011",
  54474=>"111110001",
  54475=>"001010100",
  54476=>"111101101",
  54477=>"100111111",
  54478=>"111110101",
  54479=>"110111100",
  54480=>"100011011",
  54481=>"110010000",
  54482=>"010001000",
  54483=>"010010110",
  54484=>"000011100",
  54485=>"101110111",
  54486=>"101000010",
  54487=>"101011011",
  54488=>"101110110",
  54489=>"000100011",
  54490=>"101111101",
  54491=>"111001001",
  54492=>"111110111",
  54493=>"010110010",
  54494=>"010110010",
  54495=>"000000110",
  54496=>"111111110",
  54497=>"100111001",
  54498=>"010000100",
  54499=>"000111111",
  54500=>"011110001",
  54501=>"100101101",
  54502=>"000110110",
  54503=>"101110000",
  54504=>"111011001",
  54505=>"111101010",
  54506=>"010001011",
  54507=>"101010010",
  54508=>"010010000",
  54509=>"011100011",
  54510=>"000101100",
  54511=>"011011111",
  54512=>"110111111",
  54513=>"000101011",
  54514=>"110111011",
  54515=>"101100010",
  54516=>"110110000",
  54517=>"111101001",
  54518=>"010101101",
  54519=>"001010100",
  54520=>"001010101",
  54521=>"100000100",
  54522=>"101011101",
  54523=>"000101010",
  54524=>"111001110",
  54525=>"010111001",
  54526=>"101111101",
  54527=>"100001010",
  54528=>"001110000",
  54529=>"000111100",
  54530=>"000001100",
  54531=>"100000111",
  54532=>"010001010",
  54533=>"001001011",
  54534=>"010011111",
  54535=>"110110100",
  54536=>"111111010",
  54537=>"101001000",
  54538=>"011111000",
  54539=>"100010100",
  54540=>"001101111",
  54541=>"010011110",
  54542=>"000111010",
  54543=>"101111110",
  54544=>"001000001",
  54545=>"000010011",
  54546=>"101110100",
  54547=>"011000110",
  54548=>"011110101",
  54549=>"001011010",
  54550=>"001101111",
  54551=>"100000100",
  54552=>"001101111",
  54553=>"000110111",
  54554=>"000001100",
  54555=>"100100100",
  54556=>"011101011",
  54557=>"110110111",
  54558=>"111111111",
  54559=>"110011011",
  54560=>"111000011",
  54561=>"001101011",
  54562=>"000110000",
  54563=>"111101101",
  54564=>"101110110",
  54565=>"111111011",
  54566=>"111110100",
  54567=>"001010100",
  54568=>"111011110",
  54569=>"000010010",
  54570=>"111011001",
  54571=>"111110101",
  54572=>"010100000",
  54573=>"001000000",
  54574=>"000000000",
  54575=>"110100010",
  54576=>"101110101",
  54577=>"010101000",
  54578=>"111110000",
  54579=>"000110111",
  54580=>"000110110",
  54581=>"000000100",
  54582=>"000110010",
  54583=>"110001101",
  54584=>"111101111",
  54585=>"011000010",
  54586=>"101100100",
  54587=>"010000010",
  54588=>"100000110",
  54589=>"010010001",
  54590=>"101111110",
  54591=>"101011110",
  54592=>"111010101",
  54593=>"100010000",
  54594=>"000110001",
  54595=>"111000010",
  54596=>"101001111",
  54597=>"101101011",
  54598=>"010111111",
  54599=>"101000101",
  54600=>"110111111",
  54601=>"111110111",
  54602=>"000001111",
  54603=>"000001010",
  54604=>"101100001",
  54605=>"011101000",
  54606=>"111111110",
  54607=>"110111101",
  54608=>"000010100",
  54609=>"111111001",
  54610=>"110000000",
  54611=>"111101110",
  54612=>"101010001",
  54613=>"001101100",
  54614=>"001100110",
  54615=>"111111111",
  54616=>"010001010",
  54617=>"001011011",
  54618=>"000001000",
  54619=>"000011001",
  54620=>"101001111",
  54621=>"110001111",
  54622=>"101110010",
  54623=>"001101100",
  54624=>"000000111",
  54625=>"010001000",
  54626=>"100011001",
  54627=>"010000001",
  54628=>"010101001",
  54629=>"110100011",
  54630=>"101110111",
  54631=>"011101001",
  54632=>"000010011",
  54633=>"100010101",
  54634=>"101101100",
  54635=>"000011000",
  54636=>"110001000",
  54637=>"100111010",
  54638=>"100101001",
  54639=>"110101100",
  54640=>"010001000",
  54641=>"110001101",
  54642=>"101101110",
  54643=>"111100011",
  54644=>"110111110",
  54645=>"000111100",
  54646=>"110111101",
  54647=>"100000011",
  54648=>"000001000",
  54649=>"011011000",
  54650=>"110001111",
  54651=>"000001100",
  54652=>"010100001",
  54653=>"001000011",
  54654=>"101010001",
  54655=>"110100110",
  54656=>"001101110",
  54657=>"001100010",
  54658=>"010110000",
  54659=>"000000001",
  54660=>"011011110",
  54661=>"101001001",
  54662=>"101111110",
  54663=>"100100001",
  54664=>"011011001",
  54665=>"011100110",
  54666=>"000100101",
  54667=>"100110001",
  54668=>"100111101",
  54669=>"110001111",
  54670=>"011101110",
  54671=>"000101110",
  54672=>"111000101",
  54673=>"000000111",
  54674=>"111111111",
  54675=>"001000000",
  54676=>"001101100",
  54677=>"011101000",
  54678=>"000111101",
  54679=>"000110101",
  54680=>"100100101",
  54681=>"010011011",
  54682=>"010100000",
  54683=>"000000101",
  54684=>"111110101",
  54685=>"110110010",
  54686=>"011101111",
  54687=>"101001110",
  54688=>"001100100",
  54689=>"011011000",
  54690=>"011110101",
  54691=>"111011110",
  54692=>"111010100",
  54693=>"111101111",
  54694=>"000100100",
  54695=>"111111000",
  54696=>"101000100",
  54697=>"000101111",
  54698=>"011000001",
  54699=>"001110111",
  54700=>"111111101",
  54701=>"001100001",
  54702=>"110110000",
  54703=>"110111001",
  54704=>"011111010",
  54705=>"111110101",
  54706=>"101111000",
  54707=>"000000110",
  54708=>"001001010",
  54709=>"011010101",
  54710=>"111001111",
  54711=>"100010000",
  54712=>"000101000",
  54713=>"001010110",
  54714=>"100100010",
  54715=>"011010100",
  54716=>"111111011",
  54717=>"101100111",
  54718=>"110110100",
  54719=>"111010101",
  54720=>"100111010",
  54721=>"001011111",
  54722=>"011000101",
  54723=>"100110101",
  54724=>"000101001",
  54725=>"100011101",
  54726=>"010111011",
  54727=>"111011111",
  54728=>"001010011",
  54729=>"011111011",
  54730=>"111101101",
  54731=>"011110111",
  54732=>"001000000",
  54733=>"001011111",
  54734=>"011111011",
  54735=>"110110001",
  54736=>"111110011",
  54737=>"110011110",
  54738=>"011101011",
  54739=>"001110000",
  54740=>"000111101",
  54741=>"010100101",
  54742=>"101111110",
  54743=>"010101101",
  54744=>"101011101",
  54745=>"110001110",
  54746=>"111100011",
  54747=>"101000011",
  54748=>"111101111",
  54749=>"000000010",
  54750=>"111011111",
  54751=>"101000000",
  54752=>"000011001",
  54753=>"000000000",
  54754=>"111110000",
  54755=>"001010011",
  54756=>"000110001",
  54757=>"010001000",
  54758=>"000011001",
  54759=>"001011011",
  54760=>"101000011",
  54761=>"000000100",
  54762=>"110011111",
  54763=>"010000111",
  54764=>"001011000",
  54765=>"111100101",
  54766=>"101011011",
  54767=>"111010101",
  54768=>"111111011",
  54769=>"000011100",
  54770=>"000011111",
  54771=>"011011110",
  54772=>"110101011",
  54773=>"001001000",
  54774=>"110110111",
  54775=>"010100101",
  54776=>"000110011",
  54777=>"000111101",
  54778=>"110101010",
  54779=>"110010010",
  54780=>"110110100",
  54781=>"101001011",
  54782=>"001110111",
  54783=>"000110110",
  54784=>"000011011",
  54785=>"100100010",
  54786=>"011011001",
  54787=>"001001001",
  54788=>"111001110",
  54789=>"100111001",
  54790=>"010110111",
  54791=>"110001110",
  54792=>"110000010",
  54793=>"111111110",
  54794=>"101111110",
  54795=>"110110110",
  54796=>"011001110",
  54797=>"110110000",
  54798=>"010001000",
  54799=>"110110111",
  54800=>"111001010",
  54801=>"100100111",
  54802=>"101001101",
  54803=>"110010010",
  54804=>"100010110",
  54805=>"010001011",
  54806=>"101001110",
  54807=>"100000000",
  54808=>"011110011",
  54809=>"011010011",
  54810=>"011010000",
  54811=>"000001011",
  54812=>"111111011",
  54813=>"110010011",
  54814=>"000010000",
  54815=>"001001011",
  54816=>"010100011",
  54817=>"000011001",
  54818=>"110001111",
  54819=>"010000100",
  54820=>"010101000",
  54821=>"010011010",
  54822=>"111111111",
  54823=>"110010110",
  54824=>"101100101",
  54825=>"111010101",
  54826=>"111101011",
  54827=>"100110000",
  54828=>"101111100",
  54829=>"011010111",
  54830=>"110101100",
  54831=>"011101111",
  54832=>"011011010",
  54833=>"110001110",
  54834=>"010111010",
  54835=>"011010000",
  54836=>"111100100",
  54837=>"100100100",
  54838=>"101111001",
  54839=>"101101111",
  54840=>"010110000",
  54841=>"000001010",
  54842=>"001000101",
  54843=>"110111101",
  54844=>"000011111",
  54845=>"101001011",
  54846=>"001101010",
  54847=>"001110000",
  54848=>"010010111",
  54849=>"000001111",
  54850=>"000101010",
  54851=>"100000111",
  54852=>"001011011",
  54853=>"111111101",
  54854=>"111011010",
  54855=>"000011110",
  54856=>"000010000",
  54857=>"110100100",
  54858=>"110101110",
  54859=>"000110101",
  54860=>"001000101",
  54861=>"110010111",
  54862=>"100101110",
  54863=>"010110100",
  54864=>"011110001",
  54865=>"000110011",
  54866=>"010110111",
  54867=>"000100000",
  54868=>"101111111",
  54869=>"010101011",
  54870=>"110111111",
  54871=>"110100111",
  54872=>"000001101",
  54873=>"101000000",
  54874=>"111111110",
  54875=>"110101011",
  54876=>"101011010",
  54877=>"001001010",
  54878=>"111110101",
  54879=>"000101110",
  54880=>"000101001",
  54881=>"011100111",
  54882=>"100000101",
  54883=>"011101000",
  54884=>"111100010",
  54885=>"100000001",
  54886=>"000000101",
  54887=>"101001111",
  54888=>"011101111",
  54889=>"101101000",
  54890=>"001010100",
  54891=>"100000111",
  54892=>"101000010",
  54893=>"001100000",
  54894=>"111100001",
  54895=>"110011011",
  54896=>"001101110",
  54897=>"101100000",
  54898=>"011010100",
  54899=>"100000001",
  54900=>"010000001",
  54901=>"110101101",
  54902=>"001011000",
  54903=>"000000011",
  54904=>"101111111",
  54905=>"100000110",
  54906=>"101111010",
  54907=>"001101111",
  54908=>"010101111",
  54909=>"001011001",
  54910=>"001011011",
  54911=>"001000101",
  54912=>"000001110",
  54913=>"001000110",
  54914=>"101101000",
  54915=>"111010110",
  54916=>"000111100",
  54917=>"000110000",
  54918=>"001100011",
  54919=>"000111011",
  54920=>"101111100",
  54921=>"000010000",
  54922=>"011010011",
  54923=>"110011100",
  54924=>"000001010",
  54925=>"010001001",
  54926=>"000101101",
  54927=>"101011000",
  54928=>"000000111",
  54929=>"001000000",
  54930=>"011110011",
  54931=>"101101010",
  54932=>"000110011",
  54933=>"001101110",
  54934=>"010010110",
  54935=>"100000010",
  54936=>"100111001",
  54937=>"011001101",
  54938=>"101111100",
  54939=>"110000111",
  54940=>"000001010",
  54941=>"011011111",
  54942=>"011000111",
  54943=>"101111110",
  54944=>"110111010",
  54945=>"100001010",
  54946=>"111110010",
  54947=>"011001111",
  54948=>"101111000",
  54949=>"010011010",
  54950=>"010101010",
  54951=>"000010110",
  54952=>"111011001",
  54953=>"111111110",
  54954=>"101100100",
  54955=>"000000101",
  54956=>"110111101",
  54957=>"100010011",
  54958=>"010111000",
  54959=>"110101101",
  54960=>"100000110",
  54961=>"001011100",
  54962=>"101111100",
  54963=>"100011000",
  54964=>"111111101",
  54965=>"010100001",
  54966=>"010011111",
  54967=>"111100000",
  54968=>"010100101",
  54969=>"101011110",
  54970=>"001111011",
  54971=>"001111000",
  54972=>"000011101",
  54973=>"010101011",
  54974=>"010011100",
  54975=>"110101100",
  54976=>"110000000",
  54977=>"000101000",
  54978=>"010010000",
  54979=>"000110001",
  54980=>"111000001",
  54981=>"101000110",
  54982=>"010100100",
  54983=>"000100100",
  54984=>"001101000",
  54985=>"111111111",
  54986=>"010011111",
  54987=>"111011101",
  54988=>"001010000",
  54989=>"101100010",
  54990=>"111010111",
  54991=>"101100111",
  54992=>"111001000",
  54993=>"100111110",
  54994=>"011100100",
  54995=>"010011011",
  54996=>"000010011",
  54997=>"111111110",
  54998=>"010111110",
  54999=>"001000001",
  55000=>"011000101",
  55001=>"011100101",
  55002=>"111111010",
  55003=>"011000100",
  55004=>"011001110",
  55005=>"000011110",
  55006=>"010110100",
  55007=>"100000011",
  55008=>"100000001",
  55009=>"000110110",
  55010=>"010000101",
  55011=>"000101011",
  55012=>"110101011",
  55013=>"011011001",
  55014=>"110001010",
  55015=>"011111001",
  55016=>"001011010",
  55017=>"111001101",
  55018=>"000000011",
  55019=>"100111010",
  55020=>"010011110",
  55021=>"010110000",
  55022=>"100111100",
  55023=>"010100011",
  55024=>"101101001",
  55025=>"101001101",
  55026=>"001010111",
  55027=>"110010101",
  55028=>"110111011",
  55029=>"100111100",
  55030=>"110111100",
  55031=>"000000010",
  55032=>"110110101",
  55033=>"010010011",
  55034=>"010111011",
  55035=>"000000010",
  55036=>"101101111",
  55037=>"110101001",
  55038=>"100011111",
  55039=>"010101001",
  55040=>"010110110",
  55041=>"000011100",
  55042=>"011111111",
  55043=>"110011101",
  55044=>"101011110",
  55045=>"000000000",
  55046=>"001100100",
  55047=>"100010010",
  55048=>"101010100",
  55049=>"001100010",
  55050=>"111101000",
  55051=>"110101111",
  55052=>"110001111",
  55053=>"001000100",
  55054=>"111101001",
  55055=>"000100100",
  55056=>"000001111",
  55057=>"100011110",
  55058=>"111001101",
  55059=>"000110111",
  55060=>"000000000",
  55061=>"001011100",
  55062=>"110000000",
  55063=>"000111110",
  55064=>"011001001",
  55065=>"101011101",
  55066=>"101001010",
  55067=>"011001111",
  55068=>"110011101",
  55069=>"111100010",
  55070=>"100001001",
  55071=>"101110111",
  55072=>"010101111",
  55073=>"010010110",
  55074=>"100010001",
  55075=>"000000011",
  55076=>"000110110",
  55077=>"000100111",
  55078=>"110000000",
  55079=>"100010100",
  55080=>"110111111",
  55081=>"100100100",
  55082=>"100001000",
  55083=>"100010010",
  55084=>"011100000",
  55085=>"000000101",
  55086=>"101111110",
  55087=>"110001100",
  55088=>"100010101",
  55089=>"001011100",
  55090=>"000001101",
  55091=>"001000000",
  55092=>"110001010",
  55093=>"101010001",
  55094=>"011100110",
  55095=>"110101011",
  55096=>"111011011",
  55097=>"101000110",
  55098=>"011001010",
  55099=>"111011100",
  55100=>"101000100",
  55101=>"101001011",
  55102=>"101011011",
  55103=>"001100100",
  55104=>"101011000",
  55105=>"000110110",
  55106=>"111000010",
  55107=>"111011111",
  55108=>"100010010",
  55109=>"110100011",
  55110=>"111000101",
  55111=>"011111011",
  55112=>"100011010",
  55113=>"101011111",
  55114=>"111000010",
  55115=>"110010101",
  55116=>"110101110",
  55117=>"101001011",
  55118=>"111010001",
  55119=>"110000110",
  55120=>"001000111",
  55121=>"111110011",
  55122=>"001011001",
  55123=>"011111001",
  55124=>"101000111",
  55125=>"001101101",
  55126=>"001010110",
  55127=>"100110001",
  55128=>"101001110",
  55129=>"111100000",
  55130=>"001101111",
  55131=>"010000000",
  55132=>"001001011",
  55133=>"000011011",
  55134=>"000110100",
  55135=>"111010101",
  55136=>"110001010",
  55137=>"111001000",
  55138=>"011110110",
  55139=>"010100110",
  55140=>"001001101",
  55141=>"010100010",
  55142=>"011111000",
  55143=>"001010101",
  55144=>"111111111",
  55145=>"111101010",
  55146=>"110111111",
  55147=>"110100001",
  55148=>"011010010",
  55149=>"011111000",
  55150=>"010111100",
  55151=>"010101000",
  55152=>"101110111",
  55153=>"011011111",
  55154=>"101111101",
  55155=>"001100010",
  55156=>"101001010",
  55157=>"000100010",
  55158=>"110001000",
  55159=>"111110101",
  55160=>"011010011",
  55161=>"111110100",
  55162=>"100100111",
  55163=>"001110010",
  55164=>"110001100",
  55165=>"011011111",
  55166=>"101100001",
  55167=>"110000011",
  55168=>"011011001",
  55169=>"101101000",
  55170=>"111010111",
  55171=>"010010111",
  55172=>"101000100",
  55173=>"111111111",
  55174=>"110000100",
  55175=>"101100110",
  55176=>"111100001",
  55177=>"101101101",
  55178=>"000101001",
  55179=>"010011101",
  55180=>"111110111",
  55181=>"110101110",
  55182=>"000100011",
  55183=>"100100101",
  55184=>"010100101",
  55185=>"111101100",
  55186=>"111100010",
  55187=>"010110001",
  55188=>"001011110",
  55189=>"010111110",
  55190=>"110110001",
  55191=>"011100001",
  55192=>"000000001",
  55193=>"010110110",
  55194=>"100101111",
  55195=>"100100001",
  55196=>"010001011",
  55197=>"100110010",
  55198=>"111110001",
  55199=>"101011011",
  55200=>"000011000",
  55201=>"110111001",
  55202=>"110000101",
  55203=>"101011001",
  55204=>"111101110",
  55205=>"011001001",
  55206=>"100011011",
  55207=>"111110010",
  55208=>"100101111",
  55209=>"111101011",
  55210=>"110001010",
  55211=>"000010011",
  55212=>"100111110",
  55213=>"111000011",
  55214=>"011101111",
  55215=>"100000100",
  55216=>"101101001",
  55217=>"111110101",
  55218=>"010100010",
  55219=>"001100010",
  55220=>"101100010",
  55221=>"000110110",
  55222=>"010001011",
  55223=>"001101000",
  55224=>"111011110",
  55225=>"101011111",
  55226=>"110101010",
  55227=>"000001000",
  55228=>"111101100",
  55229=>"111010101",
  55230=>"111000010",
  55231=>"101010100",
  55232=>"111111110",
  55233=>"010000101",
  55234=>"110111010",
  55235=>"010111000",
  55236=>"101111011",
  55237=>"100001100",
  55238=>"000100000",
  55239=>"111010111",
  55240=>"101101111",
  55241=>"111100001",
  55242=>"100100100",
  55243=>"111000110",
  55244=>"000011111",
  55245=>"001100000",
  55246=>"110010001",
  55247=>"010100100",
  55248=>"100101111",
  55249=>"101101111",
  55250=>"111000010",
  55251=>"110111101",
  55252=>"011001001",
  55253=>"101000000",
  55254=>"010110001",
  55255=>"110110111",
  55256=>"011011110",
  55257=>"110000100",
  55258=>"001011101",
  55259=>"000011110",
  55260=>"111101010",
  55261=>"100111011",
  55262=>"101100101",
  55263=>"001100100",
  55264=>"110111110",
  55265=>"101001010",
  55266=>"011000010",
  55267=>"010101111",
  55268=>"111111111",
  55269=>"000000110",
  55270=>"010000010",
  55271=>"111111011",
  55272=>"001101101",
  55273=>"000101001",
  55274=>"001100001",
  55275=>"011110110",
  55276=>"111111001",
  55277=>"100010000",
  55278=>"011001101",
  55279=>"010011111",
  55280=>"001000010",
  55281=>"101101101",
  55282=>"111001110",
  55283=>"110001101",
  55284=>"011001101",
  55285=>"000011010",
  55286=>"100001101",
  55287=>"000100111",
  55288=>"001110001",
  55289=>"101000000",
  55290=>"000001111",
  55291=>"111111001",
  55292=>"111110000",
  55293=>"111001110",
  55294=>"000010110",
  55295=>"111101011",
  55296=>"001101001",
  55297=>"000000111",
  55298=>"100101110",
  55299=>"011101111",
  55300=>"000000111",
  55301=>"101000100",
  55302=>"111100101",
  55303=>"000001110",
  55304=>"111101011",
  55305=>"110100000",
  55306=>"111001000",
  55307=>"111110011",
  55308=>"000011000",
  55309=>"000110000",
  55310=>"100000100",
  55311=>"000010011",
  55312=>"011110000",
  55313=>"000001000",
  55314=>"100010011",
  55315=>"000000001",
  55316=>"000000100",
  55317=>"101100101",
  55318=>"010001110",
  55319=>"110100001",
  55320=>"000000010",
  55321=>"011000000",
  55322=>"000011101",
  55323=>"000001111",
  55324=>"101001001",
  55325=>"000110111",
  55326=>"110010001",
  55327=>"111111010",
  55328=>"111001100",
  55329=>"010001011",
  55330=>"101100111",
  55331=>"011010101",
  55332=>"101101010",
  55333=>"111011111",
  55334=>"101101110",
  55335=>"010000001",
  55336=>"101101110",
  55337=>"010010111",
  55338=>"000111111",
  55339=>"011111101",
  55340=>"110000010",
  55341=>"010100011",
  55342=>"011000101",
  55343=>"100110011",
  55344=>"101010011",
  55345=>"110010000",
  55346=>"100100110",
  55347=>"000010101",
  55348=>"111111111",
  55349=>"100000000",
  55350=>"100010010",
  55351=>"111101111",
  55352=>"000111111",
  55353=>"000001101",
  55354=>"001011000",
  55355=>"100110111",
  55356=>"101100011",
  55357=>"001110000",
  55358=>"001101011",
  55359=>"010111001",
  55360=>"101001001",
  55361=>"001111011",
  55362=>"111111010",
  55363=>"110010001",
  55364=>"010101011",
  55365=>"011000001",
  55366=>"111101110",
  55367=>"011110101",
  55368=>"111001000",
  55369=>"101111000",
  55370=>"101000000",
  55371=>"000110110",
  55372=>"000011101",
  55373=>"111001110",
  55374=>"010000100",
  55375=>"011000111",
  55376=>"010111110",
  55377=>"100111101",
  55378=>"011000001",
  55379=>"011000100",
  55380=>"011010110",
  55381=>"010101010",
  55382=>"100100011",
  55383=>"001101111",
  55384=>"101111111",
  55385=>"011011100",
  55386=>"101101010",
  55387=>"001110110",
  55388=>"001001100",
  55389=>"000000110",
  55390=>"100100111",
  55391=>"100111001",
  55392=>"010010101",
  55393=>"000010010",
  55394=>"000001101",
  55395=>"011010100",
  55396=>"001101111",
  55397=>"110010001",
  55398=>"011101010",
  55399=>"000101011",
  55400=>"000000001",
  55401=>"111011111",
  55402=>"011101000",
  55403=>"100011101",
  55404=>"000010101",
  55405=>"110100010",
  55406=>"101011001",
  55407=>"101001011",
  55408=>"011001010",
  55409=>"110110010",
  55410=>"110111010",
  55411=>"111110110",
  55412=>"101101111",
  55413=>"101101010",
  55414=>"101111001",
  55415=>"000111001",
  55416=>"011010010",
  55417=>"110011101",
  55418=>"110001111",
  55419=>"000110111",
  55420=>"101110011",
  55421=>"010001111",
  55422=>"100111000",
  55423=>"010000111",
  55424=>"011110000",
  55425=>"011010111",
  55426=>"010000101",
  55427=>"110111010",
  55428=>"001000000",
  55429=>"001101111",
  55430=>"100110111",
  55431=>"001100000",
  55432=>"101111100",
  55433=>"001011001",
  55434=>"010000101",
  55435=>"011101011",
  55436=>"001001100",
  55437=>"111110011",
  55438=>"111010100",
  55439=>"111010111",
  55440=>"011010000",
  55441=>"110001111",
  55442=>"110001110",
  55443=>"011000101",
  55444=>"100011001",
  55445=>"001110011",
  55446=>"110001101",
  55447=>"110111111",
  55448=>"001001101",
  55449=>"001101001",
  55450=>"001101011",
  55451=>"010100000",
  55452=>"000000100",
  55453=>"010010000",
  55454=>"010111011",
  55455=>"000000010",
  55456=>"011100111",
  55457=>"101000000",
  55458=>"000010111",
  55459=>"101100001",
  55460=>"010011100",
  55461=>"000110111",
  55462=>"001101000",
  55463=>"100111001",
  55464=>"011010000",
  55465=>"000001001",
  55466=>"111111001",
  55467=>"011111011",
  55468=>"010001011",
  55469=>"110011101",
  55470=>"110111111",
  55471=>"000000001",
  55472=>"110110110",
  55473=>"111000000",
  55474=>"011001100",
  55475=>"101000101",
  55476=>"001011100",
  55477=>"000000011",
  55478=>"011000111",
  55479=>"010000001",
  55480=>"101110001",
  55481=>"101000110",
  55482=>"000010000",
  55483=>"001011010",
  55484=>"010101000",
  55485=>"101111010",
  55486=>"101111011",
  55487=>"011111111",
  55488=>"100110111",
  55489=>"001001100",
  55490=>"011111000",
  55491=>"011101101",
  55492=>"010011010",
  55493=>"100000011",
  55494=>"111111100",
  55495=>"110011101",
  55496=>"001000100",
  55497=>"010011000",
  55498=>"101010010",
  55499=>"000110011",
  55500=>"010101001",
  55501=>"101101100",
  55502=>"000011010",
  55503=>"110111101",
  55504=>"000010110",
  55505=>"000111011",
  55506=>"100000000",
  55507=>"101101101",
  55508=>"001010111",
  55509=>"101010010",
  55510=>"011111011",
  55511=>"011010110",
  55512=>"101111101",
  55513=>"111001110",
  55514=>"100010011",
  55515=>"001000000",
  55516=>"010011011",
  55517=>"111110110",
  55518=>"000111000",
  55519=>"110101011",
  55520=>"100101111",
  55521=>"110011010",
  55522=>"101110011",
  55523=>"000101100",
  55524=>"110111111",
  55525=>"111101001",
  55526=>"110111100",
  55527=>"000011000",
  55528=>"001011010",
  55529=>"001101011",
  55530=>"110010110",
  55531=>"011101111",
  55532=>"110111100",
  55533=>"010011010",
  55534=>"101111110",
  55535=>"011001100",
  55536=>"111001000",
  55537=>"111000000",
  55538=>"010001010",
  55539=>"100000111",
  55540=>"011000011",
  55541=>"111001001",
  55542=>"011010110",
  55543=>"001010001",
  55544=>"100000000",
  55545=>"011010101",
  55546=>"100001011",
  55547=>"100011100",
  55548=>"111100000",
  55549=>"011010010",
  55550=>"111110111",
  55551=>"111100000",
  55552=>"011100101",
  55553=>"101100100",
  55554=>"110100001",
  55555=>"110001111",
  55556=>"001000101",
  55557=>"011011010",
  55558=>"110110010",
  55559=>"100111111",
  55560=>"101111011",
  55561=>"000000111",
  55562=>"111010101",
  55563=>"110111110",
  55564=>"010110000",
  55565=>"010010011",
  55566=>"010000001",
  55567=>"010100011",
  55568=>"100011101",
  55569=>"100110010",
  55570=>"000100100",
  55571=>"000110001",
  55572=>"110000101",
  55573=>"100100001",
  55574=>"101100000",
  55575=>"000001000",
  55576=>"001001010",
  55577=>"100011011",
  55578=>"001011000",
  55579=>"011101111",
  55580=>"101110001",
  55581=>"110011001",
  55582=>"010011101",
  55583=>"101001001",
  55584=>"001010000",
  55585=>"000000000",
  55586=>"101010000",
  55587=>"100011011",
  55588=>"101000100",
  55589=>"101010101",
  55590=>"010001110",
  55591=>"110010100",
  55592=>"111011011",
  55593=>"010001100",
  55594=>"001111111",
  55595=>"111010100",
  55596=>"101011100",
  55597=>"110101111",
  55598=>"001001100",
  55599=>"100011001",
  55600=>"101101111",
  55601=>"011000000",
  55602=>"011111010",
  55603=>"111000000",
  55604=>"100101011",
  55605=>"011111100",
  55606=>"010101111",
  55607=>"110110101",
  55608=>"000010011",
  55609=>"100011000",
  55610=>"000110001",
  55611=>"100101001",
  55612=>"111101100",
  55613=>"101001101",
  55614=>"100100100",
  55615=>"001000001",
  55616=>"010100011",
  55617=>"010101101",
  55618=>"010101111",
  55619=>"000101101",
  55620=>"110101110",
  55621=>"111010011",
  55622=>"100010111",
  55623=>"101001111",
  55624=>"111010110",
  55625=>"011110100",
  55626=>"001101110",
  55627=>"011011010",
  55628=>"111101001",
  55629=>"100101100",
  55630=>"100111110",
  55631=>"100111000",
  55632=>"011111111",
  55633=>"100100111",
  55634=>"101011001",
  55635=>"110001011",
  55636=>"110000100",
  55637=>"010111011",
  55638=>"000000000",
  55639=>"101101110",
  55640=>"110010011",
  55641=>"101111111",
  55642=>"111110101",
  55643=>"011000110",
  55644=>"111110001",
  55645=>"001110101",
  55646=>"100001010",
  55647=>"001101000",
  55648=>"101001100",
  55649=>"000001011",
  55650=>"011000110",
  55651=>"001110001",
  55652=>"000100010",
  55653=>"111001001",
  55654=>"001101001",
  55655=>"011110011",
  55656=>"010001010",
  55657=>"000000000",
  55658=>"001010111",
  55659=>"010000011",
  55660=>"000000101",
  55661=>"010101010",
  55662=>"000001001",
  55663=>"011001111",
  55664=>"000000001",
  55665=>"110101110",
  55666=>"111100011",
  55667=>"100011110",
  55668=>"110001100",
  55669=>"001001110",
  55670=>"011000111",
  55671=>"010000111",
  55672=>"001111111",
  55673=>"010010001",
  55674=>"011100110",
  55675=>"101010000",
  55676=>"100011110",
  55677=>"101001011",
  55678=>"011111101",
  55679=>"101000011",
  55680=>"000000111",
  55681=>"001000111",
  55682=>"101000101",
  55683=>"100001111",
  55684=>"101011101",
  55685=>"011000000",
  55686=>"001011000",
  55687=>"101110000",
  55688=>"110110101",
  55689=>"101010010",
  55690=>"110111100",
  55691=>"010010100",
  55692=>"000111100",
  55693=>"111101001",
  55694=>"101001010",
  55695=>"111010001",
  55696=>"111101001",
  55697=>"001110110",
  55698=>"000101000",
  55699=>"001001000",
  55700=>"010110111",
  55701=>"101011001",
  55702=>"000110001",
  55703=>"111111001",
  55704=>"000000101",
  55705=>"101110101",
  55706=>"000001100",
  55707=>"101101111",
  55708=>"000101010",
  55709=>"110011011",
  55710=>"110011110",
  55711=>"111010101",
  55712=>"011001001",
  55713=>"011011111",
  55714=>"010001001",
  55715=>"010101000",
  55716=>"011001100",
  55717=>"010011111",
  55718=>"010000000",
  55719=>"101111010",
  55720=>"100011101",
  55721=>"011010101",
  55722=>"001110111",
  55723=>"010000111",
  55724=>"001011011",
  55725=>"101110100",
  55726=>"111000001",
  55727=>"110101110",
  55728=>"011110010",
  55729=>"100101001",
  55730=>"000010001",
  55731=>"010010010",
  55732=>"111111001",
  55733=>"000110000",
  55734=>"110010110",
  55735=>"101011000",
  55736=>"111011101",
  55737=>"110101011",
  55738=>"101101010",
  55739=>"011110000",
  55740=>"000001001",
  55741=>"000111011",
  55742=>"100110100",
  55743=>"000010000",
  55744=>"001101101",
  55745=>"100001010",
  55746=>"001110100",
  55747=>"010111101",
  55748=>"011010000",
  55749=>"010011010",
  55750=>"011011100",
  55751=>"000000010",
  55752=>"000001111",
  55753=>"010101011",
  55754=>"001111000",
  55755=>"101100010",
  55756=>"110010010",
  55757=>"000110101",
  55758=>"011100100",
  55759=>"100001101",
  55760=>"111001110",
  55761=>"101111110",
  55762=>"100011100",
  55763=>"011000000",
  55764=>"000110001",
  55765=>"001011111",
  55766=>"001010100",
  55767=>"101001111",
  55768=>"000100101",
  55769=>"001110010",
  55770=>"010111111",
  55771=>"000000001",
  55772=>"001010010",
  55773=>"011000110",
  55774=>"011011001",
  55775=>"000111100",
  55776=>"101011111",
  55777=>"101110010",
  55778=>"001011001",
  55779=>"111101100",
  55780=>"011101110",
  55781=>"101000100",
  55782=>"111000101",
  55783=>"110100110",
  55784=>"011000111",
  55785=>"101010100",
  55786=>"010100001",
  55787=>"111111100",
  55788=>"010111100",
  55789=>"001101000",
  55790=>"111011110",
  55791=>"101111010",
  55792=>"011111101",
  55793=>"001010110",
  55794=>"011100001",
  55795=>"000100001",
  55796=>"100110010",
  55797=>"110101110",
  55798=>"110111001",
  55799=>"010100010",
  55800=>"000111011",
  55801=>"011001110",
  55802=>"001000001",
  55803=>"101111101",
  55804=>"111111011",
  55805=>"101001111",
  55806=>"110000011",
  55807=>"010001000",
  55808=>"011000101",
  55809=>"100001010",
  55810=>"110001111",
  55811=>"000011100",
  55812=>"010111101",
  55813=>"000100000",
  55814=>"011101100",
  55815=>"100100010",
  55816=>"110001111",
  55817=>"000111100",
  55818=>"100011111",
  55819=>"001000000",
  55820=>"100100111",
  55821=>"000000100",
  55822=>"000001011",
  55823=>"100011010",
  55824=>"011000000",
  55825=>"111101010",
  55826=>"001110011",
  55827=>"111010011",
  55828=>"001011110",
  55829=>"011110111",
  55830=>"101100010",
  55831=>"111010000",
  55832=>"111011111",
  55833=>"000111010",
  55834=>"110100110",
  55835=>"110110111",
  55836=>"010110000",
  55837=>"111001001",
  55838=>"101100101",
  55839=>"010101110",
  55840=>"001000011",
  55841=>"110100000",
  55842=>"011100010",
  55843=>"010110100",
  55844=>"101101010",
  55845=>"110000100",
  55846=>"000101101",
  55847=>"010111001",
  55848=>"001100101",
  55849=>"001011101",
  55850=>"011000011",
  55851=>"100011001",
  55852=>"000001110",
  55853=>"100000110",
  55854=>"010011100",
  55855=>"001011010",
  55856=>"001011010",
  55857=>"111001000",
  55858=>"111011100",
  55859=>"110111010",
  55860=>"000110110",
  55861=>"101110100",
  55862=>"010111100",
  55863=>"101011011",
  55864=>"001111000",
  55865=>"011011000",
  55866=>"101100100",
  55867=>"111100011",
  55868=>"100100010",
  55869=>"110011111",
  55870=>"101000111",
  55871=>"101100110",
  55872=>"010011101",
  55873=>"011010111",
  55874=>"010111011",
  55875=>"011100100",
  55876=>"100111010",
  55877=>"111001110",
  55878=>"101110111",
  55879=>"010011000",
  55880=>"010100000",
  55881=>"000010000",
  55882=>"100101011",
  55883=>"100001100",
  55884=>"111011000",
  55885=>"100001010",
  55886=>"011011000",
  55887=>"010110011",
  55888=>"110011111",
  55889=>"001011010",
  55890=>"110100001",
  55891=>"110100111",
  55892=>"000000110",
  55893=>"010110110",
  55894=>"011100011",
  55895=>"000111011",
  55896=>"001001100",
  55897=>"110000010",
  55898=>"100100001",
  55899=>"101001000",
  55900=>"110110011",
  55901=>"010100001",
  55902=>"000010000",
  55903=>"110001111",
  55904=>"001101100",
  55905=>"010001010",
  55906=>"110011010",
  55907=>"001111001",
  55908=>"101100100",
  55909=>"010001110",
  55910=>"110101100",
  55911=>"101000111",
  55912=>"011100101",
  55913=>"101011111",
  55914=>"111100000",
  55915=>"110100110",
  55916=>"011001111",
  55917=>"001010110",
  55918=>"010000100",
  55919=>"110101110",
  55920=>"100011010",
  55921=>"011000000",
  55922=>"010100100",
  55923=>"011100111",
  55924=>"011000000",
  55925=>"010001000",
  55926=>"100010100",
  55927=>"100111000",
  55928=>"011111100",
  55929=>"110100001",
  55930=>"000001110",
  55931=>"000001001",
  55932=>"101110011",
  55933=>"100110100",
  55934=>"110100010",
  55935=>"100101101",
  55936=>"001011000",
  55937=>"010101011",
  55938=>"011110110",
  55939=>"000100010",
  55940=>"101101011",
  55941=>"100100000",
  55942=>"111110011",
  55943=>"110111111",
  55944=>"011011000",
  55945=>"110000000",
  55946=>"010101111",
  55947=>"010001001",
  55948=>"111011010",
  55949=>"111000110",
  55950=>"110000010",
  55951=>"010010111",
  55952=>"101101111",
  55953=>"101001001",
  55954=>"111100001",
  55955=>"001110000",
  55956=>"001010000",
  55957=>"101011111",
  55958=>"000010101",
  55959=>"110100100",
  55960=>"000101111",
  55961=>"111011010",
  55962=>"000000001",
  55963=>"101100100",
  55964=>"010101000",
  55965=>"101010100",
  55966=>"001110001",
  55967=>"100000000",
  55968=>"111100101",
  55969=>"001000110",
  55970=>"001011010",
  55971=>"100110010",
  55972=>"001001011",
  55973=>"011001100",
  55974=>"110100010",
  55975=>"001100000",
  55976=>"000011100",
  55977=>"010100000",
  55978=>"100100101",
  55979=>"110001101",
  55980=>"101111011",
  55981=>"000100101",
  55982=>"010111001",
  55983=>"101011111",
  55984=>"011000010",
  55985=>"110110111",
  55986=>"101101001",
  55987=>"101111111",
  55988=>"101100010",
  55989=>"010110100",
  55990=>"101101001",
  55991=>"111100000",
  55992=>"110011011",
  55993=>"011111010",
  55994=>"010101000",
  55995=>"111101101",
  55996=>"110010101",
  55997=>"110011011",
  55998=>"011101101",
  55999=>"010111110",
  56000=>"000101000",
  56001=>"011111111",
  56002=>"001101010",
  56003=>"011110101",
  56004=>"010111001",
  56005=>"110100101",
  56006=>"101100101",
  56007=>"111100111",
  56008=>"000010010",
  56009=>"000111110",
  56010=>"110110010",
  56011=>"000010100",
  56012=>"111010110",
  56013=>"000110110",
  56014=>"110000010",
  56015=>"101100101",
  56016=>"010000110",
  56017=>"000100100",
  56018=>"010010100",
  56019=>"101100100",
  56020=>"000111101",
  56021=>"110011001",
  56022=>"001111110",
  56023=>"001110101",
  56024=>"010110111",
  56025=>"110000010",
  56026=>"011000111",
  56027=>"101001100",
  56028=>"010010000",
  56029=>"100100100",
  56030=>"111001010",
  56031=>"010100101",
  56032=>"110000101",
  56033=>"110111100",
  56034=>"110110010",
  56035=>"001010001",
  56036=>"110100001",
  56037=>"100011011",
  56038=>"000000110",
  56039=>"001100101",
  56040=>"100101100",
  56041=>"110000010",
  56042=>"100001100",
  56043=>"001001111",
  56044=>"000000001",
  56045=>"000111100",
  56046=>"001110010",
  56047=>"100111010",
  56048=>"111101101",
  56049=>"111000010",
  56050=>"111110101",
  56051=>"111111101",
  56052=>"001101101",
  56053=>"111001110",
  56054=>"100101001",
  56055=>"101010000",
  56056=>"111111110",
  56057=>"011000000",
  56058=>"111101111",
  56059=>"111011001",
  56060=>"011000111",
  56061=>"011111001",
  56062=>"001100100",
  56063=>"111010000",
  56064=>"010101110",
  56065=>"001000100",
  56066=>"011011101",
  56067=>"000010001",
  56068=>"000110111",
  56069=>"110010110",
  56070=>"111101000",
  56071=>"111011000",
  56072=>"100001100",
  56073=>"000110000",
  56074=>"010101010",
  56075=>"011000110",
  56076=>"011101110",
  56077=>"111011010",
  56078=>"101011010",
  56079=>"111101001",
  56080=>"001100100",
  56081=>"000101010",
  56082=>"001011011",
  56083=>"100111010",
  56084=>"111100011",
  56085=>"101101010",
  56086=>"011110101",
  56087=>"011100000",
  56088=>"001011001",
  56089=>"100000111",
  56090=>"110100111",
  56091=>"110011111",
  56092=>"110110011",
  56093=>"011110000",
  56094=>"011001110",
  56095=>"001011110",
  56096=>"111111010",
  56097=>"011000001",
  56098=>"000101110",
  56099=>"011010001",
  56100=>"101001111",
  56101=>"010110001",
  56102=>"100100011",
  56103=>"100100101",
  56104=>"110110010",
  56105=>"101111110",
  56106=>"010101001",
  56107=>"110011011",
  56108=>"011111001",
  56109=>"001100001",
  56110=>"101110111",
  56111=>"100110001",
  56112=>"010110101",
  56113=>"100000110",
  56114=>"101000111",
  56115=>"100000101",
  56116=>"110100000",
  56117=>"000101100",
  56118=>"111100010",
  56119=>"001000001",
  56120=>"100011011",
  56121=>"000000001",
  56122=>"001100000",
  56123=>"110101100",
  56124=>"100000011",
  56125=>"011101110",
  56126=>"111100000",
  56127=>"010101110",
  56128=>"000100001",
  56129=>"010011100",
  56130=>"111010111",
  56131=>"000101000",
  56132=>"001000011",
  56133=>"110011111",
  56134=>"000110011",
  56135=>"011100001",
  56136=>"111010111",
  56137=>"001010000",
  56138=>"011111100",
  56139=>"101000111",
  56140=>"111111011",
  56141=>"000001000",
  56142=>"011000000",
  56143=>"000011000",
  56144=>"010100111",
  56145=>"000101100",
  56146=>"101001010",
  56147=>"111110111",
  56148=>"001011010",
  56149=>"101100000",
  56150=>"010110001",
  56151=>"000001101",
  56152=>"111111001",
  56153=>"110010001",
  56154=>"010000111",
  56155=>"110101110",
  56156=>"110110110",
  56157=>"100110110",
  56158=>"011111111",
  56159=>"100110111",
  56160=>"000000010",
  56161=>"110111101",
  56162=>"110100110",
  56163=>"011111011",
  56164=>"101010010",
  56165=>"011100110",
  56166=>"010011111",
  56167=>"110011011",
  56168=>"000100010",
  56169=>"001100010",
  56170=>"011101011",
  56171=>"100111111",
  56172=>"000001010",
  56173=>"100011000",
  56174=>"110010011",
  56175=>"111011100",
  56176=>"111100000",
  56177=>"011101110",
  56178=>"110100010",
  56179=>"000011110",
  56180=>"010011000",
  56181=>"000001110",
  56182=>"101100001",
  56183=>"001000100",
  56184=>"111110100",
  56185=>"101011110",
  56186=>"000000101",
  56187=>"110111101",
  56188=>"100100100",
  56189=>"101100000",
  56190=>"100100101",
  56191=>"101000100",
  56192=>"110110100",
  56193=>"101010101",
  56194=>"010000111",
  56195=>"101011010",
  56196=>"000011011",
  56197=>"001101110",
  56198=>"011011111",
  56199=>"101110000",
  56200=>"000100101",
  56201=>"001010010",
  56202=>"011100111",
  56203=>"010000001",
  56204=>"111110111",
  56205=>"101100101",
  56206=>"111101111",
  56207=>"101101110",
  56208=>"100100010",
  56209=>"111001111",
  56210=>"100111000",
  56211=>"010001111",
  56212=>"111000000",
  56213=>"100111111",
  56214=>"110000101",
  56215=>"010000110",
  56216=>"111000000",
  56217=>"010110001",
  56218=>"110001000",
  56219=>"111011000",
  56220=>"010000111",
  56221=>"001111111",
  56222=>"101001011",
  56223=>"111110111",
  56224=>"101111010",
  56225=>"011100000",
  56226=>"001000110",
  56227=>"001100110",
  56228=>"101000001",
  56229=>"110111111",
  56230=>"111100101",
  56231=>"010011010",
  56232=>"010001001",
  56233=>"010110001",
  56234=>"101011110",
  56235=>"100101110",
  56236=>"000000001",
  56237=>"110000010",
  56238=>"011011000",
  56239=>"000110011",
  56240=>"001000110",
  56241=>"001010011",
  56242=>"100010001",
  56243=>"111000111",
  56244=>"001110010",
  56245=>"110111100",
  56246=>"111110100",
  56247=>"111001111",
  56248=>"100100111",
  56249=>"111110010",
  56250=>"000100000",
  56251=>"000101010",
  56252=>"010101001",
  56253=>"100110010",
  56254=>"101100001",
  56255=>"000011000",
  56256=>"110001001",
  56257=>"110000011",
  56258=>"001100001",
  56259=>"000001110",
  56260=>"000111011",
  56261=>"111000000",
  56262=>"001000000",
  56263=>"010000111",
  56264=>"000000011",
  56265=>"011100000",
  56266=>"001111110",
  56267=>"000100001",
  56268=>"110010010",
  56269=>"011010111",
  56270=>"000001001",
  56271=>"000111001",
  56272=>"000100111",
  56273=>"000000010",
  56274=>"000011011",
  56275=>"010000111",
  56276=>"101111111",
  56277=>"000110001",
  56278=>"000000010",
  56279=>"111000101",
  56280=>"001101000",
  56281=>"011010101",
  56282=>"101110111",
  56283=>"111101000",
  56284=>"000111111",
  56285=>"101010111",
  56286=>"001100101",
  56287=>"110110010",
  56288=>"001110110",
  56289=>"111110010",
  56290=>"010000000",
  56291=>"101111111",
  56292=>"101101111",
  56293=>"000010110",
  56294=>"111010101",
  56295=>"100010011",
  56296=>"101010000",
  56297=>"110011100",
  56298=>"011101111",
  56299=>"011011111",
  56300=>"101111000",
  56301=>"101101110",
  56302=>"111001010",
  56303=>"110110010",
  56304=>"001111111",
  56305=>"101111110",
  56306=>"101000111",
  56307=>"101000110",
  56308=>"001000100",
  56309=>"000110000",
  56310=>"111101001",
  56311=>"111100101",
  56312=>"100110000",
  56313=>"110010000",
  56314=>"010000101",
  56315=>"010110011",
  56316=>"010100001",
  56317=>"000000001",
  56318=>"101001000",
  56319=>"101111101",
  56320=>"100110000",
  56321=>"000101011",
  56322=>"000111110",
  56323=>"101001001",
  56324=>"001100010",
  56325=>"001001001",
  56326=>"010000101",
  56327=>"101011000",
  56328=>"101110000",
  56329=>"011110101",
  56330=>"011000111",
  56331=>"101000101",
  56332=>"001001001",
  56333=>"101011010",
  56334=>"010010011",
  56335=>"011010001",
  56336=>"100110000",
  56337=>"001011000",
  56338=>"001110111",
  56339=>"000010000",
  56340=>"010111101",
  56341=>"001111101",
  56342=>"111111011",
  56343=>"000111011",
  56344=>"101010100",
  56345=>"101001111",
  56346=>"000010010",
  56347=>"011010111",
  56348=>"010100100",
  56349=>"000110010",
  56350=>"111100001",
  56351=>"001001111",
  56352=>"001011111",
  56353=>"100110010",
  56354=>"000000010",
  56355=>"110111001",
  56356=>"000111100",
  56357=>"100010001",
  56358=>"101001100",
  56359=>"000101110",
  56360=>"010010010",
  56361=>"010000011",
  56362=>"101000101",
  56363=>"001000111",
  56364=>"010010101",
  56365=>"100001000",
  56366=>"111001010",
  56367=>"101001100",
  56368=>"110011101",
  56369=>"010110011",
  56370=>"000010011",
  56371=>"111001000",
  56372=>"001001010",
  56373=>"100000000",
  56374=>"110001011",
  56375=>"011111100",
  56376=>"000100010",
  56377=>"001110100",
  56378=>"001001100",
  56379=>"111100001",
  56380=>"000110000",
  56381=>"011101010",
  56382=>"010100001",
  56383=>"101011111",
  56384=>"111010111",
  56385=>"101000101",
  56386=>"011000100",
  56387=>"110001111",
  56388=>"011001110",
  56389=>"000010110",
  56390=>"111000010",
  56391=>"010001000",
  56392=>"100101001",
  56393=>"010011000",
  56394=>"101101101",
  56395=>"101011100",
  56396=>"000001110",
  56397=>"110000100",
  56398=>"101011100",
  56399=>"011010000",
  56400=>"000100110",
  56401=>"011101001",
  56402=>"011100110",
  56403=>"101111011",
  56404=>"011110001",
  56405=>"111011110",
  56406=>"011100101",
  56407=>"010010101",
  56408=>"010101100",
  56409=>"001111001",
  56410=>"000011110",
  56411=>"001000110",
  56412=>"011011000",
  56413=>"111100001",
  56414=>"110010100",
  56415=>"010010100",
  56416=>"011110110",
  56417=>"111011100",
  56418=>"000001101",
  56419=>"000111011",
  56420=>"110000100",
  56421=>"110110001",
  56422=>"100100110",
  56423=>"101100101",
  56424=>"101010010",
  56425=>"111110101",
  56426=>"100100000",
  56427=>"100010001",
  56428=>"101100011",
  56429=>"100101011",
  56430=>"111100011",
  56431=>"010010100",
  56432=>"011011001",
  56433=>"111000001",
  56434=>"000010001",
  56435=>"100000100",
  56436=>"010111110",
  56437=>"100001111",
  56438=>"111100011",
  56439=>"000001100",
  56440=>"110110011",
  56441=>"100001010",
  56442=>"110000111",
  56443=>"110100001",
  56444=>"101010000",
  56445=>"110101010",
  56446=>"001010010",
  56447=>"100011100",
  56448=>"011011010",
  56449=>"011000000",
  56450=>"011001100",
  56451=>"000000011",
  56452=>"110010000",
  56453=>"001000000",
  56454=>"000111111",
  56455=>"110100111",
  56456=>"010010101",
  56457=>"011011110",
  56458=>"011011100",
  56459=>"101100010",
  56460=>"111110110",
  56461=>"011001010",
  56462=>"100000101",
  56463=>"010011100",
  56464=>"000111111",
  56465=>"100101000",
  56466=>"101100111",
  56467=>"100011001",
  56468=>"101101000",
  56469=>"010111011",
  56470=>"010011110",
  56471=>"011111101",
  56472=>"111110001",
  56473=>"100010011",
  56474=>"000001001",
  56475=>"101111111",
  56476=>"101000101",
  56477=>"011000111",
  56478=>"010000101",
  56479=>"000011001",
  56480=>"110110010",
  56481=>"101011010",
  56482=>"001011111",
  56483=>"011000011",
  56484=>"011101101",
  56485=>"010101010",
  56486=>"010110110",
  56487=>"100000000",
  56488=>"011101000",
  56489=>"110111110",
  56490=>"101101110",
  56491=>"101000101",
  56492=>"000101111",
  56493=>"010000000",
  56494=>"010100011",
  56495=>"100110101",
  56496=>"101000111",
  56497=>"011100010",
  56498=>"011111101",
  56499=>"011111100",
  56500=>"111001001",
  56501=>"000111000",
  56502=>"111101110",
  56503=>"110110111",
  56504=>"010000010",
  56505=>"011111000",
  56506=>"010101100",
  56507=>"011101001",
  56508=>"100010110",
  56509=>"011100111",
  56510=>"110011010",
  56511=>"110001100",
  56512=>"011000000",
  56513=>"100000110",
  56514=>"011000101",
  56515=>"100100110",
  56516=>"111000001",
  56517=>"001100110",
  56518=>"010000001",
  56519=>"100000011",
  56520=>"001001001",
  56521=>"111101001",
  56522=>"111111111",
  56523=>"111100111",
  56524=>"001001100",
  56525=>"100000001",
  56526=>"110101110",
  56527=>"111010010",
  56528=>"111111011",
  56529=>"100101010",
  56530=>"010001111",
  56531=>"010110111",
  56532=>"011001001",
  56533=>"001001000",
  56534=>"101001110",
  56535=>"111001111",
  56536=>"100100001",
  56537=>"110001001",
  56538=>"001111111",
  56539=>"011001001",
  56540=>"110001000",
  56541=>"011001100",
  56542=>"110001111",
  56543=>"000010001",
  56544=>"111100001",
  56545=>"001010001",
  56546=>"001000001",
  56547=>"000000010",
  56548=>"000100010",
  56549=>"100000101",
  56550=>"100100011",
  56551=>"010001000",
  56552=>"110110111",
  56553=>"111110110",
  56554=>"010111010",
  56555=>"101010011",
  56556=>"111111110",
  56557=>"011110101",
  56558=>"001101001",
  56559=>"000011010",
  56560=>"110111000",
  56561=>"101011101",
  56562=>"110001110",
  56563=>"100111111",
  56564=>"010100011",
  56565=>"100101110",
  56566=>"010100111",
  56567=>"110000011",
  56568=>"010011001",
  56569=>"011000011",
  56570=>"000010000",
  56571=>"000010011",
  56572=>"111111101",
  56573=>"001110000",
  56574=>"110001000",
  56575=>"110011001",
  56576=>"100101111",
  56577=>"111000101",
  56578=>"011000011",
  56579=>"010011101",
  56580=>"001111001",
  56581=>"000111101",
  56582=>"011000011",
  56583=>"111011111",
  56584=>"111111110",
  56585=>"100101011",
  56586=>"010100010",
  56587=>"011011000",
  56588=>"101001111",
  56589=>"010111010",
  56590=>"010001000",
  56591=>"111001100",
  56592=>"001000000",
  56593=>"001101110",
  56594=>"000000000",
  56595=>"011011111",
  56596=>"001110000",
  56597=>"011001111",
  56598=>"000001011",
  56599=>"101111111",
  56600=>"101001010",
  56601=>"110110100",
  56602=>"100001101",
  56603=>"111010000",
  56604=>"010111111",
  56605=>"001100000",
  56606=>"001101110",
  56607=>"001000010",
  56608=>"001110100",
  56609=>"111010100",
  56610=>"000110110",
  56611=>"010000110",
  56612=>"011000010",
  56613=>"101110000",
  56614=>"001101011",
  56615=>"111111001",
  56616=>"000111011",
  56617=>"110110111",
  56618=>"010001111",
  56619=>"101110001",
  56620=>"001100110",
  56621=>"111011001",
  56622=>"001101100",
  56623=>"111110010",
  56624=>"111010000",
  56625=>"111110011",
  56626=>"010101101",
  56627=>"010000000",
  56628=>"101000110",
  56629=>"100101100",
  56630=>"000011000",
  56631=>"101000100",
  56632=>"010010001",
  56633=>"001000111",
  56634=>"100111101",
  56635=>"100111111",
  56636=>"001001100",
  56637=>"000010010",
  56638=>"111111100",
  56639=>"111011001",
  56640=>"011101101",
  56641=>"111110111",
  56642=>"011100010",
  56643=>"110110000",
  56644=>"111111011",
  56645=>"011100111",
  56646=>"010001100",
  56647=>"011111000",
  56648=>"101101111",
  56649=>"100101111",
  56650=>"111010000",
  56651=>"000111101",
  56652=>"010110100",
  56653=>"001110110",
  56654=>"011010000",
  56655=>"111001000",
  56656=>"101110111",
  56657=>"001011010",
  56658=>"000110100",
  56659=>"010111111",
  56660=>"110111000",
  56661=>"110110110",
  56662=>"000100101",
  56663=>"011110111",
  56664=>"100101110",
  56665=>"011001000",
  56666=>"110000011",
  56667=>"011001000",
  56668=>"110111000",
  56669=>"010000010",
  56670=>"110100100",
  56671=>"100101111",
  56672=>"101110010",
  56673=>"000110000",
  56674=>"000111001",
  56675=>"011110110",
  56676=>"101110011",
  56677=>"000000101",
  56678=>"001001000",
  56679=>"000001011",
  56680=>"110101100",
  56681=>"101011011",
  56682=>"101110000",
  56683=>"110100010",
  56684=>"100110000",
  56685=>"101100011",
  56686=>"011111111",
  56687=>"111111001",
  56688=>"110101101",
  56689=>"101011010",
  56690=>"101100001",
  56691=>"001001101",
  56692=>"011110100",
  56693=>"111010100",
  56694=>"010100100",
  56695=>"010000001",
  56696=>"111100001",
  56697=>"100011010",
  56698=>"000010101",
  56699=>"111000000",
  56700=>"011010101",
  56701=>"101100010",
  56702=>"101010101",
  56703=>"101011010",
  56704=>"000000111",
  56705=>"010010100",
  56706=>"010101101",
  56707=>"000010111",
  56708=>"010100001",
  56709=>"000100000",
  56710=>"101101111",
  56711=>"010010010",
  56712=>"111110000",
  56713=>"001100011",
  56714=>"011100001",
  56715=>"101001000",
  56716=>"000111000",
  56717=>"011111010",
  56718=>"011000110",
  56719=>"110101011",
  56720=>"000000000",
  56721=>"101001110",
  56722=>"110001000",
  56723=>"001111010",
  56724=>"010111110",
  56725=>"111100110",
  56726=>"101100101",
  56727=>"111000101",
  56728=>"001010011",
  56729=>"011010100",
  56730=>"101110011",
  56731=>"110110011",
  56732=>"100010010",
  56733=>"011100001",
  56734=>"001100000",
  56735=>"010000110",
  56736=>"100001000",
  56737=>"000010110",
  56738=>"011001000",
  56739=>"110000111",
  56740=>"111110010",
  56741=>"010101000",
  56742=>"110110111",
  56743=>"101101001",
  56744=>"111000010",
  56745=>"011001111",
  56746=>"000001101",
  56747=>"011111010",
  56748=>"100001111",
  56749=>"101110011",
  56750=>"001100100",
  56751=>"011100000",
  56752=>"110101111",
  56753=>"110010011",
  56754=>"000111110",
  56755=>"111011110",
  56756=>"001010000",
  56757=>"101111010",
  56758=>"100100111",
  56759=>"000001000",
  56760=>"000101101",
  56761=>"000010110",
  56762=>"100110000",
  56763=>"101011100",
  56764=>"110001100",
  56765=>"001001001",
  56766=>"011100011",
  56767=>"010100110",
  56768=>"001110010",
  56769=>"011001010",
  56770=>"011000000",
  56771=>"101100101",
  56772=>"010000000",
  56773=>"000010110",
  56774=>"111011000",
  56775=>"001101011",
  56776=>"000100101",
  56777=>"000000101",
  56778=>"000110011",
  56779=>"101010110",
  56780=>"000101100",
  56781=>"000111011",
  56782=>"100110010",
  56783=>"101011100",
  56784=>"101100001",
  56785=>"100101010",
  56786=>"000100000",
  56787=>"000010001",
  56788=>"000101101",
  56789=>"001110001",
  56790=>"011011111",
  56791=>"011110111",
  56792=>"101111011",
  56793=>"100111100",
  56794=>"010011111",
  56795=>"011000010",
  56796=>"101100110",
  56797=>"000100100",
  56798=>"110111010",
  56799=>"111110010",
  56800=>"001101010",
  56801=>"111010011",
  56802=>"001011011",
  56803=>"100111101",
  56804=>"010100010",
  56805=>"011001011",
  56806=>"100010101",
  56807=>"000000101",
  56808=>"010010100",
  56809=>"001100011",
  56810=>"000011110",
  56811=>"100001111",
  56812=>"101010010",
  56813=>"011001100",
  56814=>"000010001",
  56815=>"000011000",
  56816=>"110110100",
  56817=>"111011001",
  56818=>"110110000",
  56819=>"110001101",
  56820=>"101011110",
  56821=>"101010001",
  56822=>"110111000",
  56823=>"011111111",
  56824=>"011011001",
  56825=>"010100100",
  56826=>"100001100",
  56827=>"110111000",
  56828=>"001100001",
  56829=>"110111100",
  56830=>"100001001",
  56831=>"001101100",
  56832=>"110100111",
  56833=>"000001101",
  56834=>"011000111",
  56835=>"101000011",
  56836=>"010111101",
  56837=>"010001011",
  56838=>"111000010",
  56839=>"010101000",
  56840=>"110100111",
  56841=>"000011110",
  56842=>"111001001",
  56843=>"111001110",
  56844=>"010110011",
  56845=>"101001001",
  56846=>"001100110",
  56847=>"100000000",
  56848=>"011001111",
  56849=>"001100101",
  56850=>"011110011",
  56851=>"000011110",
  56852=>"100100000",
  56853=>"110100000",
  56854=>"101110011",
  56855=>"110011000",
  56856=>"111110011",
  56857=>"001011010",
  56858=>"010010011",
  56859=>"111011100",
  56860=>"001000010",
  56861=>"001111110",
  56862=>"111111000",
  56863=>"010010011",
  56864=>"011010001",
  56865=>"100100110",
  56866=>"000001101",
  56867=>"000111101",
  56868=>"101000110",
  56869=>"100110101",
  56870=>"111110111",
  56871=>"001000010",
  56872=>"000101110",
  56873=>"010110001",
  56874=>"101110000",
  56875=>"100111001",
  56876=>"101011000",
  56877=>"111110000",
  56878=>"010001000",
  56879=>"101100000",
  56880=>"110000111",
  56881=>"101110010",
  56882=>"001000000",
  56883=>"011010111",
  56884=>"111000000",
  56885=>"010000110",
  56886=>"010101101",
  56887=>"000001010",
  56888=>"011000001",
  56889=>"100000000",
  56890=>"011111001",
  56891=>"100000110",
  56892=>"001010111",
  56893=>"100101101",
  56894=>"101001100",
  56895=>"001010101",
  56896=>"011101000",
  56897=>"110000011",
  56898=>"010010000",
  56899=>"010111010",
  56900=>"011111110",
  56901=>"010001011",
  56902=>"000111001",
  56903=>"011101010",
  56904=>"011111101",
  56905=>"100010111",
  56906=>"010101111",
  56907=>"000001101",
  56908=>"011000001",
  56909=>"010000000",
  56910=>"011101000",
  56911=>"000010011",
  56912=>"001111011",
  56913=>"001111101",
  56914=>"110100000",
  56915=>"001000101",
  56916=>"001111000",
  56917=>"101111101",
  56918=>"001011010",
  56919=>"010101010",
  56920=>"111110101",
  56921=>"001101011",
  56922=>"011000100",
  56923=>"010011110",
  56924=>"100101011",
  56925=>"000100001",
  56926=>"101111100",
  56927=>"111110000",
  56928=>"001011110",
  56929=>"101001010",
  56930=>"100100110",
  56931=>"110101101",
  56932=>"100000110",
  56933=>"100111011",
  56934=>"100010010",
  56935=>"110011111",
  56936=>"110000001",
  56937=>"110010000",
  56938=>"110100100",
  56939=>"000001100",
  56940=>"101101001",
  56941=>"011100010",
  56942=>"011011000",
  56943=>"001100011",
  56944=>"011101101",
  56945=>"100000000",
  56946=>"011111001",
  56947=>"011110111",
  56948=>"001011001",
  56949=>"011100010",
  56950=>"110111011",
  56951=>"100000110",
  56952=>"010001111",
  56953=>"010000010",
  56954=>"101111011",
  56955=>"011111100",
  56956=>"001001101",
  56957=>"011010111",
  56958=>"110101011",
  56959=>"101111100",
  56960=>"010011001",
  56961=>"001010000",
  56962=>"000110111",
  56963=>"111101111",
  56964=>"100000101",
  56965=>"011100111",
  56966=>"010000000",
  56967=>"010110111",
  56968=>"100111101",
  56969=>"101000011",
  56970=>"111111010",
  56971=>"011110001",
  56972=>"010111101",
  56973=>"011000101",
  56974=>"111110001",
  56975=>"111111011",
  56976=>"101110011",
  56977=>"010001100",
  56978=>"010111111",
  56979=>"100111011",
  56980=>"111101110",
  56981=>"110011011",
  56982=>"111001110",
  56983=>"100001010",
  56984=>"111101100",
  56985=>"110001000",
  56986=>"111001011",
  56987=>"010110000",
  56988=>"000000000",
  56989=>"110001110",
  56990=>"010110011",
  56991=>"011110110",
  56992=>"001100001",
  56993=>"010000100",
  56994=>"101010010",
  56995=>"011000010",
  56996=>"110100001",
  56997=>"000011100",
  56998=>"001110100",
  56999=>"111010000",
  57000=>"101000111",
  57001=>"110001011",
  57002=>"011110011",
  57003=>"000010000",
  57004=>"010001011",
  57005=>"111101100",
  57006=>"010010010",
  57007=>"000101000",
  57008=>"100111111",
  57009=>"001000010",
  57010=>"010010110",
  57011=>"010011010",
  57012=>"100111100",
  57013=>"101011001",
  57014=>"000000101",
  57015=>"100001011",
  57016=>"011011010",
  57017=>"110010100",
  57018=>"110101001",
  57019=>"111011011",
  57020=>"001010010",
  57021=>"001000000",
  57022=>"001010101",
  57023=>"001001111",
  57024=>"000001010",
  57025=>"100010010",
  57026=>"000001110",
  57027=>"100110000",
  57028=>"111100110",
  57029=>"001010011",
  57030=>"011110101",
  57031=>"101000010",
  57032=>"011010000",
  57033=>"001001000",
  57034=>"011110010",
  57035=>"110100110",
  57036=>"110100111",
  57037=>"100001000",
  57038=>"000100010",
  57039=>"011001101",
  57040=>"011011010",
  57041=>"010101110",
  57042=>"111000001",
  57043=>"001001010",
  57044=>"010011100",
  57045=>"001001001",
  57046=>"110100101",
  57047=>"001000011",
  57048=>"000110000",
  57049=>"011011111",
  57050=>"100101100",
  57051=>"111100101",
  57052=>"010110101",
  57053=>"001110000",
  57054=>"111010100",
  57055=>"101100000",
  57056=>"010011111",
  57057=>"010010110",
  57058=>"011101000",
  57059=>"110111000",
  57060=>"001101000",
  57061=>"000111100",
  57062=>"011101101",
  57063=>"001111101",
  57064=>"000011000",
  57065=>"011011000",
  57066=>"100001100",
  57067=>"111111100",
  57068=>"111110100",
  57069=>"011001100",
  57070=>"100111101",
  57071=>"000111011",
  57072=>"001000001",
  57073=>"111101101",
  57074=>"101010010",
  57075=>"011000011",
  57076=>"101011000",
  57077=>"001111101",
  57078=>"010011010",
  57079=>"010110100",
  57080=>"100110110",
  57081=>"110011001",
  57082=>"000110101",
  57083=>"000011100",
  57084=>"011001000",
  57085=>"010101010",
  57086=>"011000001",
  57087=>"111001111",
  57088=>"111110111",
  57089=>"010100110",
  57090=>"100001001",
  57091=>"101100011",
  57092=>"000000100",
  57093=>"100011100",
  57094=>"000111110",
  57095=>"011111110",
  57096=>"001101000",
  57097=>"010011010",
  57098=>"101010101",
  57099=>"100001111",
  57100=>"000101001",
  57101=>"111110111",
  57102=>"011001100",
  57103=>"100110101",
  57104=>"110001001",
  57105=>"011100111",
  57106=>"101101110",
  57107=>"011100111",
  57108=>"101001000",
  57109=>"011110110",
  57110=>"100010001",
  57111=>"101001000",
  57112=>"010001000",
  57113=>"010100000",
  57114=>"001011101",
  57115=>"100100000",
  57116=>"001110101",
  57117=>"010011001",
  57118=>"101101010",
  57119=>"011110011",
  57120=>"100001111",
  57121=>"111010010",
  57122=>"010001111",
  57123=>"100111101",
  57124=>"001010001",
  57125=>"000100100",
  57126=>"001001100",
  57127=>"000000101",
  57128=>"011100010",
  57129=>"011001010",
  57130=>"111000110",
  57131=>"111111101",
  57132=>"101000111",
  57133=>"010100101",
  57134=>"100001010",
  57135=>"101100001",
  57136=>"100011111",
  57137=>"101000100",
  57138=>"001100010",
  57139=>"111011111",
  57140=>"100010101",
  57141=>"111100110",
  57142=>"000010001",
  57143=>"110000000",
  57144=>"111000100",
  57145=>"010111111",
  57146=>"111001111",
  57147=>"000010011",
  57148=>"011111001",
  57149=>"100011000",
  57150=>"111011101",
  57151=>"100010011",
  57152=>"110000100",
  57153=>"000110100",
  57154=>"100011010",
  57155=>"111011100",
  57156=>"000100000",
  57157=>"011101011",
  57158=>"101011000",
  57159=>"111011010",
  57160=>"110000111",
  57161=>"110010001",
  57162=>"101001000",
  57163=>"011000100",
  57164=>"000100010",
  57165=>"000011000",
  57166=>"110111100",
  57167=>"101000010",
  57168=>"110101010",
  57169=>"110110000",
  57170=>"010000010",
  57171=>"101010111",
  57172=>"010111011",
  57173=>"011100111",
  57174=>"011111001",
  57175=>"111010010",
  57176=>"100010000",
  57177=>"100111010",
  57178=>"011101011",
  57179=>"110111101",
  57180=>"001101011",
  57181=>"011001010",
  57182=>"101001010",
  57183=>"111011111",
  57184=>"111011001",
  57185=>"001011001",
  57186=>"001000110",
  57187=>"100100011",
  57188=>"011110000",
  57189=>"010011000",
  57190=>"101010001",
  57191=>"011010010",
  57192=>"000000111",
  57193=>"110100100",
  57194=>"010100000",
  57195=>"001011100",
  57196=>"101010111",
  57197=>"011010110",
  57198=>"101010101",
  57199=>"110000011",
  57200=>"111010011",
  57201=>"100001000",
  57202=>"111000011",
  57203=>"111110010",
  57204=>"100100110",
  57205=>"100000010",
  57206=>"100010000",
  57207=>"010010001",
  57208=>"001010100",
  57209=>"101001111",
  57210=>"010100110",
  57211=>"000101011",
  57212=>"000101111",
  57213=>"100000100",
  57214=>"000001111",
  57215=>"001101100",
  57216=>"011110010",
  57217=>"011111100",
  57218=>"011000000",
  57219=>"110010101",
  57220=>"001110100",
  57221=>"000110010",
  57222=>"010010111",
  57223=>"110010111",
  57224=>"001011100",
  57225=>"011101100",
  57226=>"010010010",
  57227=>"000001010",
  57228=>"110011101",
  57229=>"100101010",
  57230=>"001010101",
  57231=>"000001000",
  57232=>"000011010",
  57233=>"001110111",
  57234=>"000000000",
  57235=>"011110000",
  57236=>"111110101",
  57237=>"010101000",
  57238=>"010110111",
  57239=>"111110001",
  57240=>"001000000",
  57241=>"001101001",
  57242=>"000001000",
  57243=>"001010000",
  57244=>"111010001",
  57245=>"111010111",
  57246=>"101000110",
  57247=>"110000001",
  57248=>"000000101",
  57249=>"001011010",
  57250=>"001100011",
  57251=>"001010110",
  57252=>"101111001",
  57253=>"100101100",
  57254=>"000110011",
  57255=>"000001001",
  57256=>"111001000",
  57257=>"100001100",
  57258=>"110110011",
  57259=>"011110111",
  57260=>"010110001",
  57261=>"011011111",
  57262=>"111111011",
  57263=>"100110100",
  57264=>"010111101",
  57265=>"010000000",
  57266=>"001100110",
  57267=>"111110000",
  57268=>"001100011",
  57269=>"011011000",
  57270=>"101101000",
  57271=>"001111110",
  57272=>"011001110",
  57273=>"101101101",
  57274=>"000110111",
  57275=>"000110010",
  57276=>"011001000",
  57277=>"001011000",
  57278=>"010000101",
  57279=>"111111101",
  57280=>"010110000",
  57281=>"110010011",
  57282=>"110101100",
  57283=>"111100001",
  57284=>"111110001",
  57285=>"111101111",
  57286=>"001101000",
  57287=>"001110111",
  57288=>"110100011",
  57289=>"010110100",
  57290=>"000100110",
  57291=>"111110101",
  57292=>"000101101",
  57293=>"011111111",
  57294=>"011111010",
  57295=>"111011110",
  57296=>"100001010",
  57297=>"010010111",
  57298=>"010001010",
  57299=>"100110101",
  57300=>"101011111",
  57301=>"101000110",
  57302=>"010011000",
  57303=>"001101010",
  57304=>"010100011",
  57305=>"001010001",
  57306=>"100001111",
  57307=>"110010011",
  57308=>"100111010",
  57309=>"110100010",
  57310=>"111001111",
  57311=>"011110101",
  57312=>"111101111",
  57313=>"010011010",
  57314=>"111111100",
  57315=>"101010010",
  57316=>"010101010",
  57317=>"100010111",
  57318=>"110001100",
  57319=>"110000001",
  57320=>"000101001",
  57321=>"000011011",
  57322=>"000000010",
  57323=>"101010110",
  57324=>"111011111",
  57325=>"111010101",
  57326=>"111000011",
  57327=>"011000010",
  57328=>"101011000",
  57329=>"111000011",
  57330=>"011110111",
  57331=>"000000010",
  57332=>"010111101",
  57333=>"100110011",
  57334=>"010101111",
  57335=>"010010111",
  57336=>"001100011",
  57337=>"001001001",
  57338=>"100101111",
  57339=>"101101001",
  57340=>"001101000",
  57341=>"111001110",
  57342=>"010011010",
  57343=>"100101010",
  57344=>"011111011",
  57345=>"111111100",
  57346=>"001010100",
  57347=>"010001011",
  57348=>"010010011",
  57349=>"101101101",
  57350=>"110001010",
  57351=>"011101010",
  57352=>"011101001",
  57353=>"100000010",
  57354=>"010001001",
  57355=>"100001111",
  57356=>"111100111",
  57357=>"010110100",
  57358=>"000001001",
  57359=>"100110011",
  57360=>"000001001",
  57361=>"110101111",
  57362=>"110110000",
  57363=>"010101100",
  57364=>"110111110",
  57365=>"001001011",
  57366=>"101101011",
  57367=>"111110110",
  57368=>"100010011",
  57369=>"100010001",
  57370=>"111100001",
  57371=>"100101101",
  57372=>"101001111",
  57373=>"010110001",
  57374=>"111000110",
  57375=>"101000010",
  57376=>"111111111",
  57377=>"011101111",
  57378=>"101110101",
  57379=>"011100010",
  57380=>"010110111",
  57381=>"010000000",
  57382=>"101000011",
  57383=>"100110110",
  57384=>"111001010",
  57385=>"111001100",
  57386=>"100011100",
  57387=>"001010110",
  57388=>"101111010",
  57389=>"110100011",
  57390=>"100100111",
  57391=>"111001101",
  57392=>"100101100",
  57393=>"001110011",
  57394=>"000001100",
  57395=>"110001111",
  57396=>"111010111",
  57397=>"010110000",
  57398=>"010010011",
  57399=>"010001011",
  57400=>"000011111",
  57401=>"111011001",
  57402=>"110100111",
  57403=>"010101111",
  57404=>"101101111",
  57405=>"001101101",
  57406=>"100111111",
  57407=>"010101010",
  57408=>"111110010",
  57409=>"101010101",
  57410=>"000001110",
  57411=>"110110110",
  57412=>"111010110",
  57413=>"000110011",
  57414=>"010011000",
  57415=>"111111101",
  57416=>"101001111",
  57417=>"000100001",
  57418=>"110000000",
  57419=>"000000100",
  57420=>"110110110",
  57421=>"100111100",
  57422=>"101111110",
  57423=>"010000010",
  57424=>"001001111",
  57425=>"100001101",
  57426=>"100101011",
  57427=>"011000011",
  57428=>"111100001",
  57429=>"000010111",
  57430=>"010000001",
  57431=>"111000111",
  57432=>"010110000",
  57433=>"011001111",
  57434=>"111000111",
  57435=>"110110110",
  57436=>"010000000",
  57437=>"100001000",
  57438=>"111010100",
  57439=>"101001011",
  57440=>"100111001",
  57441=>"001011101",
  57442=>"111100101",
  57443=>"000011000",
  57444=>"111011111",
  57445=>"110001000",
  57446=>"010100001",
  57447=>"100011010",
  57448=>"110110110",
  57449=>"011001101",
  57450=>"100100100",
  57451=>"110010101",
  57452=>"110100111",
  57453=>"001010000",
  57454=>"110100010",
  57455=>"001110111",
  57456=>"010100010",
  57457=>"101110011",
  57458=>"110010000",
  57459=>"100001001",
  57460=>"011001010",
  57461=>"001100000",
  57462=>"110110111",
  57463=>"110001111",
  57464=>"011110010",
  57465=>"101110011",
  57466=>"100010001",
  57467=>"000101101",
  57468=>"101001111",
  57469=>"010100011",
  57470=>"101100101",
  57471=>"011000000",
  57472=>"001101101",
  57473=>"001001010",
  57474=>"000000101",
  57475=>"100001101",
  57476=>"000011111",
  57477=>"111000000",
  57478=>"100101000",
  57479=>"101111110",
  57480=>"010010110",
  57481=>"101111010",
  57482=>"010010111",
  57483=>"100110111",
  57484=>"110000100",
  57485=>"111111000",
  57486=>"111011101",
  57487=>"000100001",
  57488=>"101000000",
  57489=>"100010101",
  57490=>"011010110",
  57491=>"101111010",
  57492=>"110000011",
  57493=>"000111101",
  57494=>"111011100",
  57495=>"110100111",
  57496=>"010010000",
  57497=>"100110001",
  57498=>"111111100",
  57499=>"111001000",
  57500=>"101011001",
  57501=>"011011000",
  57502=>"110000010",
  57503=>"100011010",
  57504=>"001111100",
  57505=>"001101111",
  57506=>"011101000",
  57507=>"011111110",
  57508=>"111111100",
  57509=>"100100001",
  57510=>"000111011",
  57511=>"000111011",
  57512=>"001000101",
  57513=>"111010011",
  57514=>"001100111",
  57515=>"101000010",
  57516=>"101000000",
  57517=>"011011001",
  57518=>"001001110",
  57519=>"111010010",
  57520=>"001011001",
  57521=>"100110011",
  57522=>"000101010",
  57523=>"111100110",
  57524=>"011110011",
  57525=>"111101010",
  57526=>"100110110",
  57527=>"100011110",
  57528=>"011010101",
  57529=>"011100011",
  57530=>"101100000",
  57531=>"101011110",
  57532=>"011000100",
  57533=>"100111011",
  57534=>"111110010",
  57535=>"011110011",
  57536=>"111110001",
  57537=>"111101000",
  57538=>"111110001",
  57539=>"111000000",
  57540=>"010000010",
  57541=>"101010000",
  57542=>"110010001",
  57543=>"011010000",
  57544=>"100010100",
  57545=>"111001111",
  57546=>"111010000",
  57547=>"010100000",
  57548=>"110111111",
  57549=>"000110000",
  57550=>"100111101",
  57551=>"000001000",
  57552=>"110110110",
  57553=>"010001100",
  57554=>"110100100",
  57555=>"110100001",
  57556=>"000100010",
  57557=>"100100011",
  57558=>"001110011",
  57559=>"011001100",
  57560=>"101010110",
  57561=>"011100000",
  57562=>"100001010",
  57563=>"000010010",
  57564=>"001111100",
  57565=>"110010001",
  57566=>"000100110",
  57567=>"010000110",
  57568=>"001000101",
  57569=>"101110001",
  57570=>"010010000",
  57571=>"010000001",
  57572=>"100001011",
  57573=>"011101011",
  57574=>"101000001",
  57575=>"100111001",
  57576=>"000110111",
  57577=>"010101100",
  57578=>"111111111",
  57579=>"011110011",
  57580=>"100000101",
  57581=>"110110100",
  57582=>"001001010",
  57583=>"001000010",
  57584=>"111001100",
  57585=>"101111111",
  57586=>"000101000",
  57587=>"110001110",
  57588=>"000111010",
  57589=>"110110010",
  57590=>"101010011",
  57591=>"011010001",
  57592=>"001000100",
  57593=>"111010101",
  57594=>"001110110",
  57595=>"101111010",
  57596=>"101000000",
  57597=>"000001110",
  57598=>"011100011",
  57599=>"101110101",
  57600=>"101100100",
  57601=>"100111101",
  57602=>"001001101",
  57603=>"011100000",
  57604=>"101000011",
  57605=>"111110110",
  57606=>"110010011",
  57607=>"001110011",
  57608=>"101100101",
  57609=>"110001111",
  57610=>"111011011",
  57611=>"101111100",
  57612=>"110110110",
  57613=>"101100010",
  57614=>"111111011",
  57615=>"011000111",
  57616=>"111111110",
  57617=>"111001010",
  57618=>"000101100",
  57619=>"110111001",
  57620=>"000011010",
  57621=>"101001010",
  57622=>"100110001",
  57623=>"100101110",
  57624=>"000100101",
  57625=>"100100000",
  57626=>"001000001",
  57627=>"010001101",
  57628=>"011100111",
  57629=>"010001101",
  57630=>"111011100",
  57631=>"100001011",
  57632=>"111000011",
  57633=>"110101101",
  57634=>"000110110",
  57635=>"101100011",
  57636=>"101011000",
  57637=>"011001000",
  57638=>"010110111",
  57639=>"011111101",
  57640=>"111111001",
  57641=>"111001111",
  57642=>"100100001",
  57643=>"111001111",
  57644=>"111110110",
  57645=>"001010111",
  57646=>"001101111",
  57647=>"011111000",
  57648=>"111101111",
  57649=>"000110110",
  57650=>"101111000",
  57651=>"110110010",
  57652=>"010010110",
  57653=>"110101110",
  57654=>"100100011",
  57655=>"010111101",
  57656=>"010011110",
  57657=>"110000011",
  57658=>"001100011",
  57659=>"001001100",
  57660=>"111100000",
  57661=>"111101001",
  57662=>"001001010",
  57663=>"001101000",
  57664=>"001000111",
  57665=>"001001110",
  57666=>"111001101",
  57667=>"101100111",
  57668=>"001100001",
  57669=>"000011000",
  57670=>"010011001",
  57671=>"110001111",
  57672=>"011100001",
  57673=>"101011000",
  57674=>"101011001",
  57675=>"100110110",
  57676=>"111110110",
  57677=>"100110110",
  57678=>"000000111",
  57679=>"011100010",
  57680=>"001001110",
  57681=>"001111010",
  57682=>"111110001",
  57683=>"010101001",
  57684=>"010101000",
  57685=>"010001011",
  57686=>"110001110",
  57687=>"010100001",
  57688=>"101010001",
  57689=>"100000000",
  57690=>"011101111",
  57691=>"001110110",
  57692=>"000011011",
  57693=>"100111110",
  57694=>"010010011",
  57695=>"000101010",
  57696=>"100111101",
  57697=>"111111100",
  57698=>"101010111",
  57699=>"100000000",
  57700=>"110101101",
  57701=>"011001001",
  57702=>"100111110",
  57703=>"001100111",
  57704=>"101101010",
  57705=>"000010100",
  57706=>"000110001",
  57707=>"100101110",
  57708=>"001110001",
  57709=>"111010011",
  57710=>"110010101",
  57711=>"101101101",
  57712=>"101110110",
  57713=>"101101101",
  57714=>"000100011",
  57715=>"011001001",
  57716=>"101011000",
  57717=>"001100000",
  57718=>"011111000",
  57719=>"000101000",
  57720=>"001001000",
  57721=>"001000000",
  57722=>"100111111",
  57723=>"011100011",
  57724=>"010011101",
  57725=>"010001000",
  57726=>"011111100",
  57727=>"101001100",
  57728=>"000101100",
  57729=>"000111100",
  57730=>"101101000",
  57731=>"011100011",
  57732=>"001010001",
  57733=>"110001101",
  57734=>"100101001",
  57735=>"100000001",
  57736=>"011001110",
  57737=>"110001010",
  57738=>"100100101",
  57739=>"100111101",
  57740=>"100101011",
  57741=>"100101011",
  57742=>"100001101",
  57743=>"111010001",
  57744=>"100111011",
  57745=>"011010000",
  57746=>"011000111",
  57747=>"110010100",
  57748=>"011011100",
  57749=>"100000101",
  57750=>"010011001",
  57751=>"000011011",
  57752=>"011111011",
  57753=>"011101100",
  57754=>"101101100",
  57755=>"110111100",
  57756=>"000110100",
  57757=>"111001101",
  57758=>"101010011",
  57759=>"000111010",
  57760=>"011100101",
  57761=>"101001111",
  57762=>"111000110",
  57763=>"110101100",
  57764=>"010001100",
  57765=>"111111001",
  57766=>"101010010",
  57767=>"100111110",
  57768=>"010011110",
  57769=>"001101000",
  57770=>"000011110",
  57771=>"010001001",
  57772=>"100100111",
  57773=>"011110111",
  57774=>"000110100",
  57775=>"110001100",
  57776=>"111100011",
  57777=>"110110110",
  57778=>"010000101",
  57779=>"001101010",
  57780=>"000011001",
  57781=>"100101101",
  57782=>"000010000",
  57783=>"011011011",
  57784=>"000010000",
  57785=>"001000111",
  57786=>"100011100",
  57787=>"110110111",
  57788=>"100000000",
  57789=>"010000000",
  57790=>"100001111",
  57791=>"000000111",
  57792=>"000111010",
  57793=>"101101110",
  57794=>"111100010",
  57795=>"011000001",
  57796=>"101011111",
  57797=>"011000011",
  57798=>"000110111",
  57799=>"111011011",
  57800=>"110010000",
  57801=>"110100011",
  57802=>"000111000",
  57803=>"100001101",
  57804=>"000000010",
  57805=>"010001011",
  57806=>"111011011",
  57807=>"010110101",
  57808=>"100010010",
  57809=>"001110101",
  57810=>"101110000",
  57811=>"100001011",
  57812=>"101001111",
  57813=>"000101010",
  57814=>"101010000",
  57815=>"000000110",
  57816=>"101010010",
  57817=>"000110000",
  57818=>"110011000",
  57819=>"011110101",
  57820=>"101101011",
  57821=>"001000110",
  57822=>"010000000",
  57823=>"010011111",
  57824=>"100001010",
  57825=>"011101010",
  57826=>"110111010",
  57827=>"111000110",
  57828=>"111101101",
  57829=>"000011000",
  57830=>"000011000",
  57831=>"100111100",
  57832=>"010000100",
  57833=>"010111001",
  57834=>"001000001",
  57835=>"010100110",
  57836=>"011001011",
  57837=>"011110101",
  57838=>"111001110",
  57839=>"010111001",
  57840=>"111011011",
  57841=>"100001010",
  57842=>"100101111",
  57843=>"000011011",
  57844=>"110011101",
  57845=>"100111000",
  57846=>"001101011",
  57847=>"110110001",
  57848=>"010110010",
  57849=>"011011110",
  57850=>"111111011",
  57851=>"011010010",
  57852=>"001001100",
  57853=>"000000010",
  57854=>"000101101",
  57855=>"001000010",
  57856=>"100001010",
  57857=>"100000001",
  57858=>"011010011",
  57859=>"001010100",
  57860=>"101001000",
  57861=>"110001110",
  57862=>"100110010",
  57863=>"010011011",
  57864=>"100101000",
  57865=>"101100111",
  57866=>"010000110",
  57867=>"011110110",
  57868=>"111111001",
  57869=>"000000110",
  57870=>"000001011",
  57871=>"011100011",
  57872=>"100110101",
  57873=>"111011000",
  57874=>"000111101",
  57875=>"110101010",
  57876=>"111010100",
  57877=>"001111111",
  57878=>"001101000",
  57879=>"100011011",
  57880=>"111100011",
  57881=>"000010101",
  57882=>"101101110",
  57883=>"110101001",
  57884=>"101111111",
  57885=>"011100111",
  57886=>"011111100",
  57887=>"111101011",
  57888=>"000101001",
  57889=>"111000100",
  57890=>"000010100",
  57891=>"001010001",
  57892=>"110001000",
  57893=>"000110000",
  57894=>"101110101",
  57895=>"010101111",
  57896=>"110000000",
  57897=>"001010011",
  57898=>"110111110",
  57899=>"001101001",
  57900=>"011110100",
  57901=>"100100111",
  57902=>"100111100",
  57903=>"010000011",
  57904=>"000101001",
  57905=>"011011101",
  57906=>"000111011",
  57907=>"001011011",
  57908=>"011111010",
  57909=>"000001010",
  57910=>"010101100",
  57911=>"011011110",
  57912=>"010001000",
  57913=>"111011111",
  57914=>"000111110",
  57915=>"111001110",
  57916=>"110111101",
  57917=>"010001010",
  57918=>"001001011",
  57919=>"000000011",
  57920=>"000110010",
  57921=>"100101111",
  57922=>"111011100",
  57923=>"101110111",
  57924=>"111001001",
  57925=>"011101001",
  57926=>"001010011",
  57927=>"000101100",
  57928=>"010011010",
  57929=>"101111111",
  57930=>"110111111",
  57931=>"100110100",
  57932=>"100110101",
  57933=>"101000111",
  57934=>"111100100",
  57935=>"010111110",
  57936=>"001111001",
  57937=>"000010000",
  57938=>"111110001",
  57939=>"100101101",
  57940=>"010001101",
  57941=>"111000000",
  57942=>"000011110",
  57943=>"100010110",
  57944=>"100000011",
  57945=>"111100001",
  57946=>"001011110",
  57947=>"000100100",
  57948=>"111101001",
  57949=>"100100010",
  57950=>"110100110",
  57951=>"101000011",
  57952=>"101100111",
  57953=>"000010000",
  57954=>"101010000",
  57955=>"011100010",
  57956=>"000011111",
  57957=>"101011101",
  57958=>"100001100",
  57959=>"010001110",
  57960=>"110000010",
  57961=>"100101000",
  57962=>"100000111",
  57963=>"010101111",
  57964=>"010111110",
  57965=>"010011111",
  57966=>"101010001",
  57967=>"011010000",
  57968=>"001111110",
  57969=>"111110001",
  57970=>"011011111",
  57971=>"101010101",
  57972=>"001010001",
  57973=>"100101010",
  57974=>"100111010",
  57975=>"111001110",
  57976=>"000011000",
  57977=>"100001011",
  57978=>"011111101",
  57979=>"110100001",
  57980=>"001000100",
  57981=>"010101000",
  57982=>"001101101",
  57983=>"111110110",
  57984=>"101000001",
  57985=>"100000101",
  57986=>"011110000",
  57987=>"111101110",
  57988=>"000110001",
  57989=>"101111011",
  57990=>"101101000",
  57991=>"010100010",
  57992=>"000011000",
  57993=>"101000010",
  57994=>"000111101",
  57995=>"111011001",
  57996=>"000000011",
  57997=>"001110111",
  57998=>"111101111",
  57999=>"101000011",
  58000=>"111000000",
  58001=>"011010101",
  58002=>"010101111",
  58003=>"010111111",
  58004=>"101111000",
  58005=>"101011010",
  58006=>"011011111",
  58007=>"111100000",
  58008=>"011110101",
  58009=>"000010010",
  58010=>"010111100",
  58011=>"010101000",
  58012=>"011001110",
  58013=>"010001111",
  58014=>"101110001",
  58015=>"011000011",
  58016=>"110000110",
  58017=>"111110110",
  58018=>"001100111",
  58019=>"011110101",
  58020=>"111000000",
  58021=>"010100000",
  58022=>"110100011",
  58023=>"010011110",
  58024=>"000110100",
  58025=>"011111111",
  58026=>"101110100",
  58027=>"100100001",
  58028=>"110000110",
  58029=>"001000111",
  58030=>"000000101",
  58031=>"111101000",
  58032=>"011111111",
  58033=>"111100111",
  58034=>"001110110",
  58035=>"101110000",
  58036=>"010001000",
  58037=>"011111011",
  58038=>"010100100",
  58039=>"111111100",
  58040=>"100110101",
  58041=>"001010111",
  58042=>"001000100",
  58043=>"101111110",
  58044=>"111000010",
  58045=>"111010010",
  58046=>"100010100",
  58047=>"100010110",
  58048=>"011011000",
  58049=>"110101001",
  58050=>"100010011",
  58051=>"010100100",
  58052=>"010101101",
  58053=>"101001000",
  58054=>"110010111",
  58055=>"000011110",
  58056=>"110101111",
  58057=>"001111100",
  58058=>"101010000",
  58059=>"011000110",
  58060=>"011100111",
  58061=>"001001010",
  58062=>"010010010",
  58063=>"111111101",
  58064=>"111011000",
  58065=>"111011111",
  58066=>"101110111",
  58067=>"010101011",
  58068=>"010111010",
  58069=>"100111000",
  58070=>"000001001",
  58071=>"010010111",
  58072=>"011101000",
  58073=>"111001011",
  58074=>"110101101",
  58075=>"110101010",
  58076=>"111101100",
  58077=>"010010000",
  58078=>"111011001",
  58079=>"010010111",
  58080=>"010111000",
  58081=>"000110101",
  58082=>"011111000",
  58083=>"110011001",
  58084=>"101011011",
  58085=>"001001000",
  58086=>"111101001",
  58087=>"111100001",
  58088=>"010101100",
  58089=>"000101001",
  58090=>"100101011",
  58091=>"000011100",
  58092=>"000010110",
  58093=>"101011000",
  58094=>"110100101",
  58095=>"101000011",
  58096=>"111001101",
  58097=>"110011011",
  58098=>"000100101",
  58099=>"101110000",
  58100=>"011111111",
  58101=>"110101100",
  58102=>"110111010",
  58103=>"001101100",
  58104=>"100010100",
  58105=>"000110010",
  58106=>"011101000",
  58107=>"100010100",
  58108=>"111001011",
  58109=>"100100101",
  58110=>"000000110",
  58111=>"000101101",
  58112=>"001010111",
  58113=>"001001010",
  58114=>"001010101",
  58115=>"010000110",
  58116=>"001100011",
  58117=>"010001011",
  58118=>"010010100",
  58119=>"111000011",
  58120=>"010001000",
  58121=>"000001001",
  58122=>"010111101",
  58123=>"100010010",
  58124=>"001110110",
  58125=>"001111011",
  58126=>"001001011",
  58127=>"100011100",
  58128=>"001101100",
  58129=>"001111010",
  58130=>"001000000",
  58131=>"111101110",
  58132=>"100101110",
  58133=>"100111111",
  58134=>"101101001",
  58135=>"010000001",
  58136=>"010000011",
  58137=>"101001011",
  58138=>"101111111",
  58139=>"010111000",
  58140=>"000000101",
  58141=>"100001010",
  58142=>"101101101",
  58143=>"111100101",
  58144=>"001101001",
  58145=>"010001000",
  58146=>"110111000",
  58147=>"111110110",
  58148=>"010010000",
  58149=>"001000010",
  58150=>"010001000",
  58151=>"011001100",
  58152=>"011110010",
  58153=>"111110001",
  58154=>"001100010",
  58155=>"011110100",
  58156=>"110010011",
  58157=>"001100110",
  58158=>"000110101",
  58159=>"010011000",
  58160=>"100100101",
  58161=>"101001100",
  58162=>"111111100",
  58163=>"111001100",
  58164=>"011101110",
  58165=>"101000110",
  58166=>"111100111",
  58167=>"101011010",
  58168=>"001011110",
  58169=>"011101010",
  58170=>"111110111",
  58171=>"010010100",
  58172=>"111100000",
  58173=>"011110001",
  58174=>"110011000",
  58175=>"111110001",
  58176=>"110001010",
  58177=>"000111011",
  58178=>"111001110",
  58179=>"000001010",
  58180=>"010010011",
  58181=>"010011100",
  58182=>"000100111",
  58183=>"100000100",
  58184=>"111101101",
  58185=>"100010011",
  58186=>"111111111",
  58187=>"010000100",
  58188=>"100010010",
  58189=>"101110011",
  58190=>"011010011",
  58191=>"001101011",
  58192=>"000101011",
  58193=>"010001100",
  58194=>"011110001",
  58195=>"010111011",
  58196=>"011001101",
  58197=>"001000000",
  58198=>"000000100",
  58199=>"111010000",
  58200=>"111010101",
  58201=>"010010111",
  58202=>"111100010",
  58203=>"000101111",
  58204=>"110111110",
  58205=>"000001010",
  58206=>"111001000",
  58207=>"100000011",
  58208=>"000111101",
  58209=>"101100101",
  58210=>"010001110",
  58211=>"111100011",
  58212=>"101110011",
  58213=>"000001000",
  58214=>"101101110",
  58215=>"011110100",
  58216=>"001010001",
  58217=>"010101001",
  58218=>"011110011",
  58219=>"110101100",
  58220=>"000010100",
  58221=>"010000000",
  58222=>"100110110",
  58223=>"000111000",
  58224=>"011100000",
  58225=>"011110001",
  58226=>"001000101",
  58227=>"100011111",
  58228=>"000101111",
  58229=>"111101010",
  58230=>"110100000",
  58231=>"011011111",
  58232=>"001011000",
  58233=>"010001110",
  58234=>"011000000",
  58235=>"101110011",
  58236=>"110010101",
  58237=>"011010001",
  58238=>"001101100",
  58239=>"010010111",
  58240=>"101111111",
  58241=>"010101100",
  58242=>"111000011",
  58243=>"011000011",
  58244=>"101100110",
  58245=>"000101011",
  58246=>"111100111",
  58247=>"011011100",
  58248=>"101111100",
  58249=>"110100000",
  58250=>"000111001",
  58251=>"010100011",
  58252=>"111001010",
  58253=>"000101101",
  58254=>"101011000",
  58255=>"000001011",
  58256=>"110000100",
  58257=>"011000011",
  58258=>"000000011",
  58259=>"010100001",
  58260=>"111101110",
  58261=>"110000001",
  58262=>"010110010",
  58263=>"101011000",
  58264=>"101111011",
  58265=>"010011111",
  58266=>"000110111",
  58267=>"111111110",
  58268=>"000010010",
  58269=>"000110111",
  58270=>"001001010",
  58271=>"111000110",
  58272=>"000110010",
  58273=>"001010010",
  58274=>"101000101",
  58275=>"010101110",
  58276=>"011000001",
  58277=>"101101001",
  58278=>"001111010",
  58279=>"110010000",
  58280=>"111111101",
  58281=>"100010001",
  58282=>"011011010",
  58283=>"011100010",
  58284=>"010101010",
  58285=>"101000100",
  58286=>"011111000",
  58287=>"100101110",
  58288=>"011001011",
  58289=>"100111111",
  58290=>"010100100",
  58291=>"110000010",
  58292=>"000011111",
  58293=>"000011000",
  58294=>"100010001",
  58295=>"111001000",
  58296=>"110000001",
  58297=>"001010101",
  58298=>"010100100",
  58299=>"111001010",
  58300=>"010111100",
  58301=>"100101000",
  58302=>"001110110",
  58303=>"010001101",
  58304=>"010111010",
  58305=>"111001101",
  58306=>"110010000",
  58307=>"011001010",
  58308=>"110011101",
  58309=>"111001000",
  58310=>"011111011",
  58311=>"101001101",
  58312=>"011110011",
  58313=>"010011001",
  58314=>"101001111",
  58315=>"100000111",
  58316=>"011010011",
  58317=>"011000011",
  58318=>"010000001",
  58319=>"001011110",
  58320=>"010110111",
  58321=>"001110110",
  58322=>"011100001",
  58323=>"010111111",
  58324=>"010001110",
  58325=>"110000000",
  58326=>"000110100",
  58327=>"110101001",
  58328=>"101101001",
  58329=>"111110000",
  58330=>"000110100",
  58331=>"111101001",
  58332=>"010001010",
  58333=>"100111000",
  58334=>"111110001",
  58335=>"111100001",
  58336=>"001101010",
  58337=>"100010101",
  58338=>"000101101",
  58339=>"000101111",
  58340=>"010000010",
  58341=>"010001010",
  58342=>"010000111",
  58343=>"011111000",
  58344=>"100011000",
  58345=>"010001011",
  58346=>"101100000",
  58347=>"001000100",
  58348=>"110110110",
  58349=>"001011100",
  58350=>"010010001",
  58351=>"000101000",
  58352=>"010000000",
  58353=>"100110101",
  58354=>"110001001",
  58355=>"100000110",
  58356=>"011010110",
  58357=>"010010001",
  58358=>"101001010",
  58359=>"111010100",
  58360=>"000000100",
  58361=>"100000011",
  58362=>"100110110",
  58363=>"110110001",
  58364=>"111100011",
  58365=>"100010110",
  58366=>"101101000",
  58367=>"111010000",
  58368=>"110000011",
  58369=>"101000100",
  58370=>"010000111",
  58371=>"101000101",
  58372=>"101110011",
  58373=>"011101010",
  58374=>"010000111",
  58375=>"111010110",
  58376=>"011101110",
  58377=>"010110101",
  58378=>"000000110",
  58379=>"111111101",
  58380=>"100111001",
  58381=>"010110101",
  58382=>"011100110",
  58383=>"001111000",
  58384=>"011110101",
  58385=>"001111111",
  58386=>"101001101",
  58387=>"110111010",
  58388=>"000001001",
  58389=>"110000100",
  58390=>"011111011",
  58391=>"000111000",
  58392=>"001000000",
  58393=>"101010000",
  58394=>"110110110",
  58395=>"100101011",
  58396=>"100111110",
  58397=>"100111101",
  58398=>"001111010",
  58399=>"100110011",
  58400=>"111111111",
  58401=>"001011101",
  58402=>"000100100",
  58403=>"101000001",
  58404=>"111110010",
  58405=>"001010010",
  58406=>"111011101",
  58407=>"101000010",
  58408=>"111100000",
  58409=>"010100011",
  58410=>"001001111",
  58411=>"111101101",
  58412=>"000011110",
  58413=>"101100111",
  58414=>"011011111",
  58415=>"001000011",
  58416=>"110100101",
  58417=>"001011000",
  58418=>"101100111",
  58419=>"111111000",
  58420=>"100101011",
  58421=>"110110101",
  58422=>"110010100",
  58423=>"101001100",
  58424=>"001001110",
  58425=>"101101000",
  58426=>"011100001",
  58427=>"001111010",
  58428=>"011100001",
  58429=>"000111000",
  58430=>"111011110",
  58431=>"100110100",
  58432=>"010101010",
  58433=>"010000101",
  58434=>"000101101",
  58435=>"111101011",
  58436=>"000100000",
  58437=>"001010000",
  58438=>"001100010",
  58439=>"000000001",
  58440=>"100010010",
  58441=>"011111001",
  58442=>"111100001",
  58443=>"001001010",
  58444=>"110110011",
  58445=>"010010000",
  58446=>"011110001",
  58447=>"000011100",
  58448=>"110110101",
  58449=>"000000110",
  58450=>"001101101",
  58451=>"000111101",
  58452=>"001101110",
  58453=>"011110000",
  58454=>"011101000",
  58455=>"000100111",
  58456=>"001010011",
  58457=>"010100000",
  58458=>"000000001",
  58459=>"010100111",
  58460=>"110100110",
  58461=>"101001110",
  58462=>"000111011",
  58463=>"101000110",
  58464=>"011111100",
  58465=>"110111111",
  58466=>"100000110",
  58467=>"100000110",
  58468=>"110111101",
  58469=>"101001100",
  58470=>"011100011",
  58471=>"010100101",
  58472=>"010000110",
  58473=>"000010101",
  58474=>"011100011",
  58475=>"101011110",
  58476=>"001100111",
  58477=>"010110100",
  58478=>"101110001",
  58479=>"110011100",
  58480=>"011101000",
  58481=>"010011000",
  58482=>"000001111",
  58483=>"111001001",
  58484=>"101110000",
  58485=>"100011010",
  58486=>"111101010",
  58487=>"100011010",
  58488=>"111100001",
  58489=>"111101010",
  58490=>"100100000",
  58491=>"111111010",
  58492=>"011000101",
  58493=>"110000001",
  58494=>"000000011",
  58495=>"100110011",
  58496=>"111010110",
  58497=>"111011000",
  58498=>"000010000",
  58499=>"111000111",
  58500=>"100010101",
  58501=>"110001011",
  58502=>"100111100",
  58503=>"111111001",
  58504=>"010010010",
  58505=>"011110100",
  58506=>"100100110",
  58507=>"100001000",
  58508=>"111100100",
  58509=>"001001111",
  58510=>"011001010",
  58511=>"000010010",
  58512=>"010100001",
  58513=>"001100000",
  58514=>"000010100",
  58515=>"000110110",
  58516=>"011111011",
  58517=>"100001010",
  58518=>"100100000",
  58519=>"011000110",
  58520=>"101010110",
  58521=>"011010101",
  58522=>"011111001",
  58523=>"110100111",
  58524=>"101000011",
  58525=>"000010101",
  58526=>"110000001",
  58527=>"110110000",
  58528=>"110101011",
  58529=>"001010010",
  58530=>"000110111",
  58531=>"001111101",
  58532=>"010111111",
  58533=>"101001101",
  58534=>"110100110",
  58535=>"011010110",
  58536=>"010100011",
  58537=>"011001101",
  58538=>"010011011",
  58539=>"101110111",
  58540=>"101010111",
  58541=>"001101000",
  58542=>"001110111",
  58543=>"100010101",
  58544=>"000100100",
  58545=>"011010011",
  58546=>"011001011",
  58547=>"111011111",
  58548=>"101001111",
  58549=>"110001000",
  58550=>"111000011",
  58551=>"000100001",
  58552=>"001111011",
  58553=>"111101111",
  58554=>"001001000",
  58555=>"110000010",
  58556=>"101100111",
  58557=>"100110011",
  58558=>"000001111",
  58559=>"001111000",
  58560=>"101000100",
  58561=>"010010000",
  58562=>"010100110",
  58563=>"010111001",
  58564=>"100011011",
  58565=>"100000000",
  58566=>"110100111",
  58567=>"001001000",
  58568=>"110000101",
  58569=>"010100100",
  58570=>"100111011",
  58571=>"010111110",
  58572=>"001010110",
  58573=>"110000000",
  58574=>"001111010",
  58575=>"010011100",
  58576=>"010001110",
  58577=>"000011001",
  58578=>"010010110",
  58579=>"011011001",
  58580=>"010011000",
  58581=>"011110101",
  58582=>"011101110",
  58583=>"010100000",
  58584=>"010011000",
  58585=>"110110000",
  58586=>"101011011",
  58587=>"111110100",
  58588=>"110001001",
  58589=>"100001100",
  58590=>"111000010",
  58591=>"010011100",
  58592=>"000011110",
  58593=>"110110101",
  58594=>"110010011",
  58595=>"000000110",
  58596=>"010010111",
  58597=>"111000111",
  58598=>"011001000",
  58599=>"100111101",
  58600=>"011110101",
  58601=>"101101100",
  58602=>"011101100",
  58603=>"100000010",
  58604=>"100000001",
  58605=>"011001111",
  58606=>"011100000",
  58607=>"110100101",
  58608=>"111111101",
  58609=>"010001010",
  58610=>"000111110",
  58611=>"110111111",
  58612=>"001111001",
  58613=>"000001011",
  58614=>"110101100",
  58615=>"110011011",
  58616=>"011111000",
  58617=>"000111000",
  58618=>"100011101",
  58619=>"010110000",
  58620=>"010101001",
  58621=>"101101001",
  58622=>"100111100",
  58623=>"010001000",
  58624=>"000110011",
  58625=>"010010001",
  58626=>"100000111",
  58627=>"001001111",
  58628=>"101010110",
  58629=>"111110001",
  58630=>"010000110",
  58631=>"100000111",
  58632=>"000000011",
  58633=>"000111110",
  58634=>"111010101",
  58635=>"110100010",
  58636=>"010010000",
  58637=>"000010111",
  58638=>"011011001",
  58639=>"100010011",
  58640=>"110010010",
  58641=>"111001110",
  58642=>"101010111",
  58643=>"001000000",
  58644=>"110100000",
  58645=>"101011001",
  58646=>"001001101",
  58647=>"010100100",
  58648=>"011011110",
  58649=>"000000111",
  58650=>"110000110",
  58651=>"111011100",
  58652=>"010100001",
  58653=>"111001011",
  58654=>"011010110",
  58655=>"111111011",
  58656=>"100001000",
  58657=>"001111110",
  58658=>"011101000",
  58659=>"110101111",
  58660=>"001001000",
  58661=>"111100111",
  58662=>"100101111",
  58663=>"101101000",
  58664=>"100100010",
  58665=>"010101111",
  58666=>"111001010",
  58667=>"111111001",
  58668=>"011001111",
  58669=>"011100010",
  58670=>"111110111",
  58671=>"010000010",
  58672=>"100100011",
  58673=>"000010110",
  58674=>"101111011",
  58675=>"000111100",
  58676=>"111001101",
  58677=>"010011010",
  58678=>"111101111",
  58679=>"100101101",
  58680=>"101011100",
  58681=>"001001011",
  58682=>"000011010",
  58683=>"111000011",
  58684=>"111011000",
  58685=>"111111011",
  58686=>"000010100",
  58687=>"110101010",
  58688=>"011010100",
  58689=>"111101001",
  58690=>"000001010",
  58691=>"001111000",
  58692=>"101111101",
  58693=>"101100111",
  58694=>"101101101",
  58695=>"100101110",
  58696=>"010101110",
  58697=>"010100000",
  58698=>"010111011",
  58699=>"111010111",
  58700=>"110110111",
  58701=>"011110111",
  58702=>"011110010",
  58703=>"010101001",
  58704=>"010100110",
  58705=>"101100010",
  58706=>"101111111",
  58707=>"111001010",
  58708=>"101010100",
  58709=>"010010011",
  58710=>"100100100",
  58711=>"111110100",
  58712=>"001101000",
  58713=>"001000110",
  58714=>"111000010",
  58715=>"111101011",
  58716=>"010001010",
  58717=>"000001111",
  58718=>"011100010",
  58719=>"100000110",
  58720=>"110101110",
  58721=>"111011101",
  58722=>"101100111",
  58723=>"000001010",
  58724=>"011011100",
  58725=>"010011011",
  58726=>"000001011",
  58727=>"011111101",
  58728=>"100010010",
  58729=>"111100100",
  58730=>"110000011",
  58731=>"100100011",
  58732=>"111111111",
  58733=>"110001100",
  58734=>"111100101",
  58735=>"100111011",
  58736=>"100101101",
  58737=>"110110000",
  58738=>"110010000",
  58739=>"010110011",
  58740=>"000110010",
  58741=>"010000101",
  58742=>"010111111",
  58743=>"001000000",
  58744=>"111101110",
  58745=>"011101101",
  58746=>"010001010",
  58747=>"001111000",
  58748=>"010001001",
  58749=>"001111110",
  58750=>"001001111",
  58751=>"000101110",
  58752=>"000001000",
  58753=>"010110010",
  58754=>"011011000",
  58755=>"001011100",
  58756=>"000110001",
  58757=>"011010110",
  58758=>"000000110",
  58759=>"110101000",
  58760=>"111010010",
  58761=>"100110111",
  58762=>"111101100",
  58763=>"100001110",
  58764=>"110001010",
  58765=>"110010101",
  58766=>"101110011",
  58767=>"111111111",
  58768=>"111000010",
  58769=>"111100101",
  58770=>"101010101",
  58771=>"101011010",
  58772=>"000111100",
  58773=>"110101110",
  58774=>"101110101",
  58775=>"101110111",
  58776=>"101110011",
  58777=>"110100100",
  58778=>"110100111",
  58779=>"110000010",
  58780=>"110000001",
  58781=>"110110100",
  58782=>"000011111",
  58783=>"001111010",
  58784=>"101011110",
  58785=>"000010100",
  58786=>"010000000",
  58787=>"101010111",
  58788=>"010100001",
  58789=>"110000001",
  58790=>"101101100",
  58791=>"100111000",
  58792=>"001100000",
  58793=>"111101010",
  58794=>"101001010",
  58795=>"011010110",
  58796=>"010101100",
  58797=>"001100010",
  58798=>"011111001",
  58799=>"000110000",
  58800=>"010001100",
  58801=>"001001011",
  58802=>"011000111",
  58803=>"110010101",
  58804=>"001101100",
  58805=>"100001010",
  58806=>"001001101",
  58807=>"111001101",
  58808=>"101011011",
  58809=>"000011101",
  58810=>"111000001",
  58811=>"101101001",
  58812=>"001101001",
  58813=>"101010001",
  58814=>"000000000",
  58815=>"110010111",
  58816=>"110000010",
  58817=>"110101100",
  58818=>"000000111",
  58819=>"110010101",
  58820=>"000101000",
  58821=>"011000100",
  58822=>"100110001",
  58823=>"011100101",
  58824=>"101011101",
  58825=>"000111011",
  58826=>"101001001",
  58827=>"100011101",
  58828=>"001101011",
  58829=>"001111100",
  58830=>"000010000",
  58831=>"010111111",
  58832=>"111101001",
  58833=>"011000111",
  58834=>"000111101",
  58835=>"010000100",
  58836=>"100110011",
  58837=>"111111111",
  58838=>"111001100",
  58839=>"101100111",
  58840=>"011000111",
  58841=>"111001001",
  58842=>"100011101",
  58843=>"110010101",
  58844=>"111000010",
  58845=>"111001101",
  58846=>"001111001",
  58847=>"011010101",
  58848=>"111001010",
  58849=>"101110111",
  58850=>"000110011",
  58851=>"100001100",
  58852=>"111110100",
  58853=>"110110011",
  58854=>"000011001",
  58855=>"010000001",
  58856=>"101001001",
  58857=>"100011110",
  58858=>"010000111",
  58859=>"000111101",
  58860=>"000100001",
  58861=>"110110001",
  58862=>"000011001",
  58863=>"111110111",
  58864=>"010011100",
  58865=>"110001101",
  58866=>"000101110",
  58867=>"011101110",
  58868=>"111000000",
  58869=>"111111110",
  58870=>"010111100",
  58871=>"001111111",
  58872=>"001111000",
  58873=>"000011000",
  58874=>"011001001",
  58875=>"011111111",
  58876=>"010111000",
  58877=>"000100010",
  58878=>"001001101",
  58879=>"110111111",
  58880=>"011110011",
  58881=>"010111000",
  58882=>"010111011",
  58883=>"011100110",
  58884=>"111000100",
  58885=>"010010111",
  58886=>"110111111",
  58887=>"010000111",
  58888=>"000010100",
  58889=>"111011101",
  58890=>"101000111",
  58891=>"011110001",
  58892=>"000000011",
  58893=>"011100111",
  58894=>"110110000",
  58895=>"000010000",
  58896=>"100000000",
  58897=>"010111000",
  58898=>"010011100",
  58899=>"110001110",
  58900=>"100010010",
  58901=>"010000100",
  58902=>"111101000",
  58903=>"011010111",
  58904=>"101101011",
  58905=>"111111011",
  58906=>"100001001",
  58907=>"001010111",
  58908=>"000011111",
  58909=>"110010011",
  58910=>"010100000",
  58911=>"101010011",
  58912=>"110001110",
  58913=>"111111111",
  58914=>"000001001",
  58915=>"000000110",
  58916=>"001000000",
  58917=>"100101001",
  58918=>"001110010",
  58919=>"101000111",
  58920=>"000010011",
  58921=>"101000011",
  58922=>"001000101",
  58923=>"011011001",
  58924=>"111011101",
  58925=>"101100110",
  58926=>"000000100",
  58927=>"101110011",
  58928=>"010010000",
  58929=>"011100101",
  58930=>"000010101",
  58931=>"001011000",
  58932=>"001110000",
  58933=>"101001110",
  58934=>"100110000",
  58935=>"000011100",
  58936=>"010000101",
  58937=>"011010101",
  58938=>"111010001",
  58939=>"100101010",
  58940=>"100010110",
  58941=>"010100110",
  58942=>"011111100",
  58943=>"011111000",
  58944=>"010101011",
  58945=>"111110011",
  58946=>"010000010",
  58947=>"100110100",
  58948=>"110100110",
  58949=>"001100011",
  58950=>"000110010",
  58951=>"101000101",
  58952=>"110111111",
  58953=>"010100110",
  58954=>"101110000",
  58955=>"110010110",
  58956=>"001101001",
  58957=>"010101111",
  58958=>"001110100",
  58959=>"010111110",
  58960=>"010010101",
  58961=>"010101110",
  58962=>"000110100",
  58963=>"011000001",
  58964=>"110000101",
  58965=>"010100010",
  58966=>"101111100",
  58967=>"010000101",
  58968=>"101101001",
  58969=>"110101100",
  58970=>"100100110",
  58971=>"001001110",
  58972=>"100111000",
  58973=>"101011110",
  58974=>"101010110",
  58975=>"100100111",
  58976=>"100010100",
  58977=>"010011110",
  58978=>"110001010",
  58979=>"011011011",
  58980=>"000111000",
  58981=>"000011110",
  58982=>"000010011",
  58983=>"001011011",
  58984=>"010110100",
  58985=>"111001000",
  58986=>"011000101",
  58987=>"101101111",
  58988=>"011011111",
  58989=>"111000001",
  58990=>"001011110",
  58991=>"100001000",
  58992=>"100100000",
  58993=>"101011111",
  58994=>"001100100",
  58995=>"111001100",
  58996=>"110101000",
  58997=>"011100110",
  58998=>"111000101",
  58999=>"111000000",
  59000=>"110010000",
  59001=>"000011000",
  59002=>"101000001",
  59003=>"001001110",
  59004=>"011101111",
  59005=>"010100011",
  59006=>"011000011",
  59007=>"111011111",
  59008=>"110110101",
  59009=>"000110000",
  59010=>"101100011",
  59011=>"100001011",
  59012=>"110011101",
  59013=>"101110000",
  59014=>"111100110",
  59015=>"101111000",
  59016=>"101011011",
  59017=>"010100110",
  59018=>"111111111",
  59019=>"001000000",
  59020=>"011011101",
  59021=>"010100101",
  59022=>"100000010",
  59023=>"001000001",
  59024=>"110001100",
  59025=>"100111111",
  59026=>"001101110",
  59027=>"011001010",
  59028=>"111001110",
  59029=>"010010110",
  59030=>"111011010",
  59031=>"111010101",
  59032=>"111110100",
  59033=>"111010000",
  59034=>"101101111",
  59035=>"011001110",
  59036=>"010110010",
  59037=>"010101000",
  59038=>"001101111",
  59039=>"001010101",
  59040=>"000011100",
  59041=>"111111111",
  59042=>"000111000",
  59043=>"011011110",
  59044=>"110101011",
  59045=>"111110001",
  59046=>"011101010",
  59047=>"000011110",
  59048=>"100101010",
  59049=>"101101100",
  59050=>"001111001",
  59051=>"001011011",
  59052=>"000011000",
  59053=>"100111101",
  59054=>"001001101",
  59055=>"000100000",
  59056=>"000001011",
  59057=>"100010000",
  59058=>"011100101",
  59059=>"011010110",
  59060=>"010011001",
  59061=>"011111001",
  59062=>"100101111",
  59063=>"100011011",
  59064=>"011101000",
  59065=>"111101100",
  59066=>"110010001",
  59067=>"101111101",
  59068=>"000011110",
  59069=>"110000001",
  59070=>"111000111",
  59071=>"000010010",
  59072=>"111010011",
  59073=>"001010001",
  59074=>"111111110",
  59075=>"100100101",
  59076=>"101101101",
  59077=>"111111001",
  59078=>"111011101",
  59079=>"111111100",
  59080=>"101000110",
  59081=>"010010101",
  59082=>"110010101",
  59083=>"101011011",
  59084=>"000010110",
  59085=>"010000001",
  59086=>"000000100",
  59087=>"101010100",
  59088=>"010001001",
  59089=>"100110101",
  59090=>"000011000",
  59091=>"110100110",
  59092=>"100001111",
  59093=>"011011000",
  59094=>"101000011",
  59095=>"111110000",
  59096=>"110000000",
  59097=>"000101001",
  59098=>"011101111",
  59099=>"000100010",
  59100=>"001010111",
  59101=>"000001000",
  59102=>"010100111",
  59103=>"000100100",
  59104=>"001100110",
  59105=>"111000010",
  59106=>"100010011",
  59107=>"100100110",
  59108=>"110010110",
  59109=>"101111011",
  59110=>"011111100",
  59111=>"000101101",
  59112=>"010010100",
  59113=>"010011111",
  59114=>"110110100",
  59115=>"100010111",
  59116=>"111110111",
  59117=>"111010010",
  59118=>"100111000",
  59119=>"101110100",
  59120=>"011000100",
  59121=>"011100110",
  59122=>"111110001",
  59123=>"111111111",
  59124=>"100010100",
  59125=>"100110010",
  59126=>"101111110",
  59127=>"001001001",
  59128=>"010111111",
  59129=>"010110000",
  59130=>"011111010",
  59131=>"000110101",
  59132=>"101001100",
  59133=>"101100010",
  59134=>"000000110",
  59135=>"010011010",
  59136=>"100010001",
  59137=>"011111111",
  59138=>"011011100",
  59139=>"000100001",
  59140=>"111110001",
  59141=>"110101101",
  59142=>"000111100",
  59143=>"110110000",
  59144=>"111111101",
  59145=>"111000010",
  59146=>"000000101",
  59147=>"010101011",
  59148=>"101001011",
  59149=>"001110010",
  59150=>"010011101",
  59151=>"100001100",
  59152=>"100101001",
  59153=>"000001111",
  59154=>"101010010",
  59155=>"011011100",
  59156=>"111010100",
  59157=>"101011011",
  59158=>"101101000",
  59159=>"000111001",
  59160=>"010101001",
  59161=>"101111010",
  59162=>"101001000",
  59163=>"001000011",
  59164=>"111110000",
  59165=>"110100001",
  59166=>"011100110",
  59167=>"010101110",
  59168=>"011011011",
  59169=>"100000011",
  59170=>"000100101",
  59171=>"111011011",
  59172=>"110011111",
  59173=>"011100001",
  59174=>"101011101",
  59175=>"100010010",
  59176=>"100010000",
  59177=>"111001011",
  59178=>"101000001",
  59179=>"111000101",
  59180=>"110001100",
  59181=>"111000111",
  59182=>"001011100",
  59183=>"010111010",
  59184=>"010001010",
  59185=>"101111011",
  59186=>"011010010",
  59187=>"111100011",
  59188=>"011011101",
  59189=>"111001000",
  59190=>"010100000",
  59191=>"101101001",
  59192=>"001111001",
  59193=>"000010001",
  59194=>"111100111",
  59195=>"000101110",
  59196=>"100101010",
  59197=>"001000111",
  59198=>"001011111",
  59199=>"111000101",
  59200=>"001010010",
  59201=>"010111010",
  59202=>"000001110",
  59203=>"001000111",
  59204=>"111000000",
  59205=>"110010010",
  59206=>"011100001",
  59207=>"010110010",
  59208=>"100110101",
  59209=>"001010000",
  59210=>"101100000",
  59211=>"101111011",
  59212=>"001000110",
  59213=>"000110010",
  59214=>"111101111",
  59215=>"100111011",
  59216=>"011000101",
  59217=>"010001001",
  59218=>"111101110",
  59219=>"010001001",
  59220=>"010011011",
  59221=>"011001010",
  59222=>"111001110",
  59223=>"001010010",
  59224=>"100000011",
  59225=>"011011110",
  59226=>"100100011",
  59227=>"011111100",
  59228=>"011011111",
  59229=>"110101000",
  59230=>"011011001",
  59231=>"101000000",
  59232=>"101001111",
  59233=>"001001011",
  59234=>"111110110",
  59235=>"001000000",
  59236=>"100100001",
  59237=>"010100101",
  59238=>"111000100",
  59239=>"011011001",
  59240=>"110010111",
  59241=>"111110110",
  59242=>"111000110",
  59243=>"101110110",
  59244=>"011101000",
  59245=>"011010010",
  59246=>"110100000",
  59247=>"100111000",
  59248=>"100110001",
  59249=>"001001001",
  59250=>"100101010",
  59251=>"110111000",
  59252=>"010001111",
  59253=>"011110010",
  59254=>"110101000",
  59255=>"101000111",
  59256=>"000101100",
  59257=>"011111101",
  59258=>"010100100",
  59259=>"011101100",
  59260=>"010001010",
  59261=>"101010111",
  59262=>"111010110",
  59263=>"101010011",
  59264=>"010011001",
  59265=>"001000100",
  59266=>"101100011",
  59267=>"111001100",
  59268=>"111100000",
  59269=>"111111101",
  59270=>"100111100",
  59271=>"111010100",
  59272=>"010110011",
  59273=>"000100110",
  59274=>"110100000",
  59275=>"111111100",
  59276=>"111110111",
  59277=>"010010110",
  59278=>"100000101",
  59279=>"000000010",
  59280=>"011111000",
  59281=>"011110010",
  59282=>"010000010",
  59283=>"110001001",
  59284=>"111101111",
  59285=>"111000011",
  59286=>"110000110",
  59287=>"111000000",
  59288=>"110110011",
  59289=>"000011000",
  59290=>"111001101",
  59291=>"001101011",
  59292=>"011101000",
  59293=>"010101010",
  59294=>"010110110",
  59295=>"110000110",
  59296=>"001100011",
  59297=>"000001001",
  59298=>"111000010",
  59299=>"100110000",
  59300=>"100111010",
  59301=>"001101101",
  59302=>"110001100",
  59303=>"011100111",
  59304=>"000101011",
  59305=>"111100111",
  59306=>"001110001",
  59307=>"101001101",
  59308=>"101110001",
  59309=>"001010101",
  59310=>"010000011",
  59311=>"101100100",
  59312=>"101111011",
  59313=>"111001101",
  59314=>"101100000",
  59315=>"111100100",
  59316=>"111101111",
  59317=>"000001011",
  59318=>"001101010",
  59319=>"010111110",
  59320=>"110111101",
  59321=>"001011000",
  59322=>"110101011",
  59323=>"100010001",
  59324=>"111100001",
  59325=>"001001000",
  59326=>"101000110",
  59327=>"001000110",
  59328=>"001100110",
  59329=>"110111100",
  59330=>"110000100",
  59331=>"000000001",
  59332=>"010001110",
  59333=>"001111101",
  59334=>"000100011",
  59335=>"111011001",
  59336=>"001111011",
  59337=>"100100100",
  59338=>"001011110",
  59339=>"111110011",
  59340=>"011110101",
  59341=>"101000110",
  59342=>"011101111",
  59343=>"100000001",
  59344=>"100000100",
  59345=>"001010011",
  59346=>"101100011",
  59347=>"111110110",
  59348=>"100100110",
  59349=>"011010100",
  59350=>"010101101",
  59351=>"111111000",
  59352=>"101110111",
  59353=>"110000111",
  59354=>"001001011",
  59355=>"000011111",
  59356=>"011000111",
  59357=>"000001011",
  59358=>"000101001",
  59359=>"111110101",
  59360=>"011110100",
  59361=>"110000101",
  59362=>"110010010",
  59363=>"100100010",
  59364=>"010001101",
  59365=>"000011101",
  59366=>"011101010",
  59367=>"010111010",
  59368=>"101110110",
  59369=>"101001101",
  59370=>"000100110",
  59371=>"000111101",
  59372=>"101110010",
  59373=>"011001110",
  59374=>"100000100",
  59375=>"010011110",
  59376=>"100011110",
  59377=>"011110110",
  59378=>"101011000",
  59379=>"000101100",
  59380=>"100110111",
  59381=>"101001001",
  59382=>"111001111",
  59383=>"010011111",
  59384=>"100101011",
  59385=>"010100100",
  59386=>"110101111",
  59387=>"000010011",
  59388=>"010111010",
  59389=>"000010100",
  59390=>"001100010",
  59391=>"101000000",
  59392=>"001011101",
  59393=>"011101101",
  59394=>"100110111",
  59395=>"100011010",
  59396=>"010111110",
  59397=>"100000111",
  59398=>"001000000",
  59399=>"110100000",
  59400=>"011010010",
  59401=>"110011011",
  59402=>"111110011",
  59403=>"000011010",
  59404=>"000011000",
  59405=>"100100001",
  59406=>"001010000",
  59407=>"101000001",
  59408=>"010111100",
  59409=>"100111101",
  59410=>"100101111",
  59411=>"000100001",
  59412=>"100111100",
  59413=>"110111001",
  59414=>"101101000",
  59415=>"001011001",
  59416=>"100101110",
  59417=>"111011010",
  59418=>"110001100",
  59419=>"111001001",
  59420=>"101011100",
  59421=>"100101010",
  59422=>"110101000",
  59423=>"111111011",
  59424=>"111100101",
  59425=>"000111111",
  59426=>"110011110",
  59427=>"100001011",
  59428=>"101010101",
  59429=>"001001100",
  59430=>"000010001",
  59431=>"110100101",
  59432=>"101100010",
  59433=>"100000000",
  59434=>"000100110",
  59435=>"000101110",
  59436=>"100111000",
  59437=>"010001111",
  59438=>"011011011",
  59439=>"011111111",
  59440=>"111111111",
  59441=>"111010010",
  59442=>"001000111",
  59443=>"000100101",
  59444=>"110111100",
  59445=>"000101001",
  59446=>"011001101",
  59447=>"111001110",
  59448=>"000110001",
  59449=>"101111111",
  59450=>"010100011",
  59451=>"100111111",
  59452=>"001111010",
  59453=>"000011010",
  59454=>"011111101",
  59455=>"000100100",
  59456=>"010101101",
  59457=>"010011001",
  59458=>"011110100",
  59459=>"010000000",
  59460=>"101000011",
  59461=>"001101100",
  59462=>"011010100",
  59463=>"001100001",
  59464=>"111001001",
  59465=>"010001100",
  59466=>"001101101",
  59467=>"110001110",
  59468=>"100100110",
  59469=>"000011110",
  59470=>"100000010",
  59471=>"010100110",
  59472=>"100111101",
  59473=>"001001101",
  59474=>"100011000",
  59475=>"011100101",
  59476=>"010000000",
  59477=>"110000000",
  59478=>"010010010",
  59479=>"101111111",
  59480=>"100101001",
  59481=>"111100101",
  59482=>"111001000",
  59483=>"101001100",
  59484=>"000010101",
  59485=>"100001010",
  59486=>"111001100",
  59487=>"110001100",
  59488=>"001111000",
  59489=>"001001000",
  59490=>"101000100",
  59491=>"000001010",
  59492=>"011011000",
  59493=>"100111001",
  59494=>"010010101",
  59495=>"011010100",
  59496=>"100110010",
  59497=>"110110100",
  59498=>"010100000",
  59499=>"000001000",
  59500=>"100001101",
  59501=>"101100111",
  59502=>"111110000",
  59503=>"111000011",
  59504=>"001111111",
  59505=>"111111100",
  59506=>"110110101",
  59507=>"000000010",
  59508=>"101111101",
  59509=>"011111100",
  59510=>"100001110",
  59511=>"010100100",
  59512=>"001001011",
  59513=>"101001110",
  59514=>"001000011",
  59515=>"110000001",
  59516=>"100011000",
  59517=>"111011110",
  59518=>"101111001",
  59519=>"000010110",
  59520=>"110111111",
  59521=>"111110000",
  59522=>"010001000",
  59523=>"101111111",
  59524=>"101110111",
  59525=>"010111101",
  59526=>"101111010",
  59527=>"011101000",
  59528=>"001000000",
  59529=>"011111001",
  59530=>"111110111",
  59531=>"011001000",
  59532=>"110000101",
  59533=>"010001101",
  59534=>"110010000",
  59535=>"111101000",
  59536=>"001010001",
  59537=>"101100110",
  59538=>"010001101",
  59539=>"011011011",
  59540=>"110010010",
  59541=>"011010110",
  59542=>"101110101",
  59543=>"011101111",
  59544=>"011011100",
  59545=>"101000111",
  59546=>"110001010",
  59547=>"111011010",
  59548=>"001000000",
  59549=>"000001010",
  59550=>"010011010",
  59551=>"111000110",
  59552=>"101101011",
  59553=>"111001010",
  59554=>"011001001",
  59555=>"001101100",
  59556=>"001000011",
  59557=>"011010100",
  59558=>"001010110",
  59559=>"100101010",
  59560=>"101000000",
  59561=>"101111111",
  59562=>"010100000",
  59563=>"011000110",
  59564=>"010110011",
  59565=>"001111110",
  59566=>"000101100",
  59567=>"111111001",
  59568=>"000011001",
  59569=>"100000001",
  59570=>"010000000",
  59571=>"100011010",
  59572=>"101001001",
  59573=>"110011000",
  59574=>"100111010",
  59575=>"100100000",
  59576=>"111100111",
  59577=>"110110010",
  59578=>"110101001",
  59579=>"001100011",
  59580=>"011000000",
  59581=>"101010011",
  59582=>"111001110",
  59583=>"010101000",
  59584=>"000000000",
  59585=>"011101001",
  59586=>"011111111",
  59587=>"101111101",
  59588=>"101110100",
  59589=>"111010000",
  59590=>"111001000",
  59591=>"111011110",
  59592=>"000101111",
  59593=>"010010010",
  59594=>"101000110",
  59595=>"010011111",
  59596=>"111110111",
  59597=>"011011000",
  59598=>"100001111",
  59599=>"111001111",
  59600=>"010010101",
  59601=>"000100111",
  59602=>"100011000",
  59603=>"001110010",
  59604=>"110111111",
  59605=>"100011110",
  59606=>"001111010",
  59607=>"100000010",
  59608=>"001110101",
  59609=>"011100110",
  59610=>"101111010",
  59611=>"010100010",
  59612=>"111110101",
  59613=>"000010010",
  59614=>"110101001",
  59615=>"110110010",
  59616=>"110011101",
  59617=>"011010011",
  59618=>"111101001",
  59619=>"001101011",
  59620=>"001110000",
  59621=>"100001000",
  59622=>"001011010",
  59623=>"011111011",
  59624=>"111110100",
  59625=>"111100001",
  59626=>"011101111",
  59627=>"000000011",
  59628=>"010110111",
  59629=>"110011000",
  59630=>"111100100",
  59631=>"101110111",
  59632=>"000111101",
  59633=>"101110110",
  59634=>"110000001",
  59635=>"000000011",
  59636=>"010100010",
  59637=>"001000000",
  59638=>"111101000",
  59639=>"000001000",
  59640=>"001001011",
  59641=>"100001001",
  59642=>"100000011",
  59643=>"000011010",
  59644=>"111000001",
  59645=>"101001000",
  59646=>"110000100",
  59647=>"100100101",
  59648=>"011100101",
  59649=>"101011001",
  59650=>"111100000",
  59651=>"111010010",
  59652=>"001001001",
  59653=>"100111010",
  59654=>"100111111",
  59655=>"010000001",
  59656=>"000101011",
  59657=>"101011011",
  59658=>"110010010",
  59659=>"101100001",
  59660=>"001101000",
  59661=>"110001100",
  59662=>"111101011",
  59663=>"101000010",
  59664=>"000100000",
  59665=>"011110001",
  59666=>"001011110",
  59667=>"100011011",
  59668=>"100100111",
  59669=>"101001111",
  59670=>"011000000",
  59671=>"000010111",
  59672=>"101010101",
  59673=>"101100101",
  59674=>"000000010",
  59675=>"111100011",
  59676=>"000000001",
  59677=>"010110001",
  59678=>"101110011",
  59679=>"111001010",
  59680=>"110000101",
  59681=>"001010110",
  59682=>"011001001",
  59683=>"001001110",
  59684=>"100110110",
  59685=>"111001101",
  59686=>"011001011",
  59687=>"101101001",
  59688=>"111011110",
  59689=>"101110010",
  59690=>"100111011",
  59691=>"011111110",
  59692=>"001000111",
  59693=>"011111111",
  59694=>"110110001",
  59695=>"110001101",
  59696=>"101111000",
  59697=>"111000110",
  59698=>"001101100",
  59699=>"101010000",
  59700=>"010010001",
  59701=>"110110000",
  59702=>"111001011",
  59703=>"111111111",
  59704=>"110000100",
  59705=>"110011111",
  59706=>"001010000",
  59707=>"010010011",
  59708=>"010100001",
  59709=>"100000010",
  59710=>"011011000",
  59711=>"110100100",
  59712=>"001101001",
  59713=>"000100100",
  59714=>"111010000",
  59715=>"100001101",
  59716=>"011011010",
  59717=>"011000010",
  59718=>"111101111",
  59719=>"101010010",
  59720=>"100011010",
  59721=>"101111011",
  59722=>"000010001",
  59723=>"111111111",
  59724=>"101101110",
  59725=>"100110110",
  59726=>"101111101",
  59727=>"110110000",
  59728=>"111010000",
  59729=>"100100011",
  59730=>"111001110",
  59731=>"111011100",
  59732=>"000110100",
  59733=>"110101001",
  59734=>"001101001",
  59735=>"001101111",
  59736=>"000000010",
  59737=>"101100100",
  59738=>"100000101",
  59739=>"110111001",
  59740=>"011110000",
  59741=>"011011100",
  59742=>"010110000",
  59743=>"000111100",
  59744=>"001010100",
  59745=>"111110011",
  59746=>"000011111",
  59747=>"101110111",
  59748=>"111111111",
  59749=>"110100001",
  59750=>"001110010",
  59751=>"110010000",
  59752=>"010111111",
  59753=>"011011111",
  59754=>"001010001",
  59755=>"100010000",
  59756=>"001011111",
  59757=>"110011101",
  59758=>"001000001",
  59759=>"010010000",
  59760=>"010001001",
  59761=>"010010111",
  59762=>"101111100",
  59763=>"010000000",
  59764=>"000001101",
  59765=>"101011001",
  59766=>"100110100",
  59767=>"101011001",
  59768=>"010110000",
  59769=>"001111111",
  59770=>"001010010",
  59771=>"001010001",
  59772=>"111110011",
  59773=>"111010101",
  59774=>"101110010",
  59775=>"001010110",
  59776=>"001111000",
  59777=>"101001011",
  59778=>"001101101",
  59779=>"001011001",
  59780=>"100111001",
  59781=>"011101100",
  59782=>"011010111",
  59783=>"011010001",
  59784=>"100011110",
  59785=>"000111011",
  59786=>"011111000",
  59787=>"111100101",
  59788=>"001011000",
  59789=>"101010000",
  59790=>"110000100",
  59791=>"111101011",
  59792=>"010101110",
  59793=>"111111010",
  59794=>"010011100",
  59795=>"110011010",
  59796=>"111001101",
  59797=>"001000111",
  59798=>"000001001",
  59799=>"010011010",
  59800=>"001001010",
  59801=>"001000001",
  59802=>"010101100",
  59803=>"110000101",
  59804=>"111111111",
  59805=>"001101010",
  59806=>"110011010",
  59807=>"100111010",
  59808=>"000101001",
  59809=>"001101111",
  59810=>"011111011",
  59811=>"110110001",
  59812=>"100100111",
  59813=>"000101101",
  59814=>"100110000",
  59815=>"000110111",
  59816=>"000110100",
  59817=>"101011010",
  59818=>"111001000",
  59819=>"010010101",
  59820=>"100010101",
  59821=>"001011100",
  59822=>"100001001",
  59823=>"001010001",
  59824=>"011001111",
  59825=>"001000100",
  59826=>"111100000",
  59827=>"000011000",
  59828=>"101100100",
  59829=>"101011001",
  59830=>"010001011",
  59831=>"110110111",
  59832=>"101001111",
  59833=>"000000001",
  59834=>"011101101",
  59835=>"110000011",
  59836=>"000010001",
  59837=>"111000011",
  59838=>"101000001",
  59839=>"010101001",
  59840=>"001001111",
  59841=>"010101001",
  59842=>"111010110",
  59843=>"010101110",
  59844=>"001100001",
  59845=>"110001111",
  59846=>"110000111",
  59847=>"110111111",
  59848=>"110101001",
  59849=>"100100100",
  59850=>"000110000",
  59851=>"011011111",
  59852=>"000000011",
  59853=>"110000001",
  59854=>"100011111",
  59855=>"100001110",
  59856=>"000100000",
  59857=>"011101000",
  59858=>"111010001",
  59859=>"011000100",
  59860=>"000001100",
  59861=>"011100110",
  59862=>"100000001",
  59863=>"011010100",
  59864=>"110000110",
  59865=>"001000011",
  59866=>"111011001",
  59867=>"011111011",
  59868=>"101000000",
  59869=>"111100011",
  59870=>"111111110",
  59871=>"001010001",
  59872=>"110011010",
  59873=>"100101011",
  59874=>"011000001",
  59875=>"100010111",
  59876=>"001101101",
  59877=>"110100110",
  59878=>"100111001",
  59879=>"011111011",
  59880=>"011000101",
  59881=>"010110000",
  59882=>"000111101",
  59883=>"010001101",
  59884=>"010101001",
  59885=>"001011011",
  59886=>"000100010",
  59887=>"110101110",
  59888=>"100000010",
  59889=>"101111000",
  59890=>"000000100",
  59891=>"111111001",
  59892=>"100001000",
  59893=>"101000100",
  59894=>"100111100",
  59895=>"111111010",
  59896=>"010100010",
  59897=>"000110011",
  59898=>"101010101",
  59899=>"010110001",
  59900=>"001100110",
  59901=>"000101110",
  59902=>"010111010",
  59903=>"100110111",
  59904=>"111110011",
  59905=>"110010010",
  59906=>"001111011",
  59907=>"110001011",
  59908=>"011010011",
  59909=>"100100000",
  59910=>"001110101",
  59911=>"110001000",
  59912=>"010101011",
  59913=>"011110010",
  59914=>"101000111",
  59915=>"111110110",
  59916=>"110001001",
  59917=>"001110000",
  59918=>"111010110",
  59919=>"011011110",
  59920=>"000011101",
  59921=>"111000101",
  59922=>"101100111",
  59923=>"010101010",
  59924=>"111000110",
  59925=>"000110010",
  59926=>"101011111",
  59927=>"010101000",
  59928=>"001001101",
  59929=>"111011110",
  59930=>"111001111",
  59931=>"111101100",
  59932=>"111000001",
  59933=>"101110010",
  59934=>"110000100",
  59935=>"110000100",
  59936=>"111101011",
  59937=>"000100100",
  59938=>"101111000",
  59939=>"011111111",
  59940=>"000101011",
  59941=>"001100000",
  59942=>"110111111",
  59943=>"000011101",
  59944=>"111001010",
  59945=>"000010010",
  59946=>"101001100",
  59947=>"110000010",
  59948=>"010101110",
  59949=>"111101100",
  59950=>"010010111",
  59951=>"001111011",
  59952=>"010011010",
  59953=>"001111110",
  59954=>"011000111",
  59955=>"010000010",
  59956=>"011101100",
  59957=>"110010010",
  59958=>"110000000",
  59959=>"010010010",
  59960=>"011100111",
  59961=>"101001011",
  59962=>"010111000",
  59963=>"101101111",
  59964=>"110111110",
  59965=>"111011001",
  59966=>"100111100",
  59967=>"010101011",
  59968=>"001001000",
  59969=>"101100001",
  59970=>"111111111",
  59971=>"010001011",
  59972=>"110101001",
  59973=>"001100110",
  59974=>"011111011",
  59975=>"111111101",
  59976=>"100011101",
  59977=>"011011011",
  59978=>"111111000",
  59979=>"001011001",
  59980=>"111001101",
  59981=>"000000001",
  59982=>"111011101",
  59983=>"101011001",
  59984=>"101011110",
  59985=>"010100110",
  59986=>"100101110",
  59987=>"111001110",
  59988=>"011010010",
  59989=>"101100100",
  59990=>"011100111",
  59991=>"000010000",
  59992=>"011000110",
  59993=>"011011010",
  59994=>"101001111",
  59995=>"101100100",
  59996=>"000101111",
  59997=>"010000000",
  59998=>"010100111",
  59999=>"000100011",
  60000=>"101110101",
  60001=>"001101100",
  60002=>"001010011",
  60003=>"110011000",
  60004=>"100101101",
  60005=>"101101110",
  60006=>"111010000",
  60007=>"100100010",
  60008=>"100110110",
  60009=>"011001110",
  60010=>"010110111",
  60011=>"111001111",
  60012=>"100001000",
  60013=>"100010010",
  60014=>"011000111",
  60015=>"111001111",
  60016=>"111110111",
  60017=>"101110111",
  60018=>"011000111",
  60019=>"001000100",
  60020=>"011111011",
  60021=>"111100000",
  60022=>"000011010",
  60023=>"001010001",
  60024=>"010111011",
  60025=>"100001110",
  60026=>"011110010",
  60027=>"010100111",
  60028=>"111101101",
  60029=>"011010011",
  60030=>"000010010",
  60031=>"000011111",
  60032=>"010010000",
  60033=>"111010001",
  60034=>"011111011",
  60035=>"110001011",
  60036=>"000110010",
  60037=>"011000110",
  60038=>"111010011",
  60039=>"100010101",
  60040=>"100110010",
  60041=>"111101001",
  60042=>"011110010",
  60043=>"011010111",
  60044=>"000010000",
  60045=>"010011100",
  60046=>"011110001",
  60047=>"011111010",
  60048=>"101000000",
  60049=>"011111001",
  60050=>"001000001",
  60051=>"111001110",
  60052=>"001110111",
  60053=>"011111001",
  60054=>"001001111",
  60055=>"101011101",
  60056=>"100010100",
  60057=>"111111100",
  60058=>"011010111",
  60059=>"001000111",
  60060=>"111101010",
  60061=>"110010001",
  60062=>"000100110",
  60063=>"110111100",
  60064=>"011010011",
  60065=>"011000101",
  60066=>"011111111",
  60067=>"000011000",
  60068=>"011001011",
  60069=>"110011101",
  60070=>"010001001",
  60071=>"001101100",
  60072=>"010110100",
  60073=>"111001101",
  60074=>"111000001",
  60075=>"101010000",
  60076=>"100010101",
  60077=>"110001000",
  60078=>"000100010",
  60079=>"000101000",
  60080=>"000010000",
  60081=>"001000001",
  60082=>"110011101",
  60083=>"001001011",
  60084=>"101001001",
  60085=>"010110000",
  60086=>"110110001",
  60087=>"101001111",
  60088=>"110110110",
  60089=>"000001011",
  60090=>"110000110",
  60091=>"010011101",
  60092=>"111101000",
  60093=>"111101111",
  60094=>"111111110",
  60095=>"010110011",
  60096=>"111011101",
  60097=>"011010000",
  60098=>"111000111",
  60099=>"110010001",
  60100=>"101101001",
  60101=>"000001011",
  60102=>"111111110",
  60103=>"110111001",
  60104=>"010111010",
  60105=>"110100111",
  60106=>"010010100",
  60107=>"111111010",
  60108=>"010011111",
  60109=>"001100010",
  60110=>"110111101",
  60111=>"011111101",
  60112=>"101111110",
  60113=>"111010011",
  60114=>"110011011",
  60115=>"101101110",
  60116=>"101101000",
  60117=>"111010101",
  60118=>"100001010",
  60119=>"010000011",
  60120=>"100101111",
  60121=>"101101101",
  60122=>"001110101",
  60123=>"111001001",
  60124=>"110001101",
  60125=>"000110010",
  60126=>"110001101",
  60127=>"100010101",
  60128=>"011011001",
  60129=>"101110000",
  60130=>"010011000",
  60131=>"011101100",
  60132=>"100101001",
  60133=>"001110010",
  60134=>"111010111",
  60135=>"011000111",
  60136=>"001000100",
  60137=>"001000100",
  60138=>"100111110",
  60139=>"000011011",
  60140=>"110110001",
  60141=>"010100011",
  60142=>"101011101",
  60143=>"111100111",
  60144=>"101011010",
  60145=>"010010100",
  60146=>"110011100",
  60147=>"100110000",
  60148=>"000010001",
  60149=>"101110011",
  60150=>"110011000",
  60151=>"011111111",
  60152=>"100110101",
  60153=>"011011010",
  60154=>"110001111",
  60155=>"110000000",
  60156=>"101100001",
  60157=>"111000010",
  60158=>"000111010",
  60159=>"001111001",
  60160=>"111111011",
  60161=>"110111110",
  60162=>"010101000",
  60163=>"011110111",
  60164=>"101010000",
  60165=>"101001000",
  60166=>"000010010",
  60167=>"101111110",
  60168=>"001101000",
  60169=>"010011101",
  60170=>"110001110",
  60171=>"111110100",
  60172=>"011011010",
  60173=>"001010110",
  60174=>"100011011",
  60175=>"001111010",
  60176=>"100011111",
  60177=>"011010001",
  60178=>"001101000",
  60179=>"011011110",
  60180=>"011111001",
  60181=>"011001010",
  60182=>"001000011",
  60183=>"001000000",
  60184=>"101101101",
  60185=>"100101010",
  60186=>"110010101",
  60187=>"001010010",
  60188=>"100111011",
  60189=>"001001011",
  60190=>"001000000",
  60191=>"111010000",
  60192=>"100100000",
  60193=>"101010011",
  60194=>"100100101",
  60195=>"001000000",
  60196=>"101001001",
  60197=>"011101001",
  60198=>"000010111",
  60199=>"001010001",
  60200=>"010111010",
  60201=>"111101100",
  60202=>"101001011",
  60203=>"110011010",
  60204=>"100100110",
  60205=>"011011111",
  60206=>"100100101",
  60207=>"001100010",
  60208=>"011111010",
  60209=>"011001001",
  60210=>"100110110",
  60211=>"110111000",
  60212=>"101100011",
  60213=>"011000011",
  60214=>"001111001",
  60215=>"101010111",
  60216=>"001100100",
  60217=>"101010011",
  60218=>"001100100",
  60219=>"101100010",
  60220=>"110101111",
  60221=>"101001001",
  60222=>"101101110",
  60223=>"000101011",
  60224=>"101111000",
  60225=>"111111111",
  60226=>"100111110",
  60227=>"001001000",
  60228=>"101000000",
  60229=>"111110001",
  60230=>"111100001",
  60231=>"011110011",
  60232=>"111110111",
  60233=>"110111011",
  60234=>"000101111",
  60235=>"011101110",
  60236=>"001001011",
  60237=>"010010010",
  60238=>"011111011",
  60239=>"100101110",
  60240=>"000000000",
  60241=>"101010000",
  60242=>"111001110",
  60243=>"101011100",
  60244=>"011111011",
  60245=>"100011000",
  60246=>"101111111",
  60247=>"111001000",
  60248=>"110000000",
  60249=>"000100000",
  60250=>"110101010",
  60251=>"000101000",
  60252=>"111011100",
  60253=>"100100111",
  60254=>"110101011",
  60255=>"111101111",
  60256=>"101100010",
  60257=>"011101111",
  60258=>"000000001",
  60259=>"011101101",
  60260=>"101100010",
  60261=>"110101011",
  60262=>"100101111",
  60263=>"101111000",
  60264=>"110011000",
  60265=>"101011110",
  60266=>"001000100",
  60267=>"110000001",
  60268=>"010001011",
  60269=>"001010000",
  60270=>"010001100",
  60271=>"000001110",
  60272=>"111000101",
  60273=>"000001111",
  60274=>"110101001",
  60275=>"001000000",
  60276=>"001101110",
  60277=>"010010010",
  60278=>"110111001",
  60279=>"100010101",
  60280=>"101010111",
  60281=>"010110000",
  60282=>"111001001",
  60283=>"101011111",
  60284=>"010000011",
  60285=>"110011111",
  60286=>"000100100",
  60287=>"000010010",
  60288=>"000000011",
  60289=>"101111011",
  60290=>"010100100",
  60291=>"010111010",
  60292=>"001100001",
  60293=>"001010001",
  60294=>"111100111",
  60295=>"101110100",
  60296=>"110100000",
  60297=>"100111011",
  60298=>"000001000",
  60299=>"011101001",
  60300=>"101111111",
  60301=>"111111111",
  60302=>"101011011",
  60303=>"111010000",
  60304=>"001001000",
  60305=>"000011100",
  60306=>"101011000",
  60307=>"111110011",
  60308=>"010110100",
  60309=>"010000000",
  60310=>"011010010",
  60311=>"101000010",
  60312=>"110100111",
  60313=>"001000010",
  60314=>"100110101",
  60315=>"010000110",
  60316=>"010100111",
  60317=>"010011000",
  60318=>"101000010",
  60319=>"001100001",
  60320=>"110011101",
  60321=>"011000011",
  60322=>"010000101",
  60323=>"001110110",
  60324=>"111011010",
  60325=>"000001110",
  60326=>"001101111",
  60327=>"011001110",
  60328=>"110100011",
  60329=>"101111000",
  60330=>"000101000",
  60331=>"011101111",
  60332=>"101111011",
  60333=>"111011010",
  60334=>"010000010",
  60335=>"000100000",
  60336=>"000001001",
  60337=>"010010100",
  60338=>"110011011",
  60339=>"111010010",
  60340=>"011000100",
  60341=>"011111110",
  60342=>"011011011",
  60343=>"000110010",
  60344=>"110110110",
  60345=>"000010011",
  60346=>"101001111",
  60347=>"110100001",
  60348=>"111110101",
  60349=>"001111101",
  60350=>"010010100",
  60351=>"101011000",
  60352=>"101001101",
  60353=>"111101010",
  60354=>"001110101",
  60355=>"010110100",
  60356=>"110001010",
  60357=>"101001001",
  60358=>"010011001",
  60359=>"101101000",
  60360=>"010100011",
  60361=>"011101111",
  60362=>"101110110",
  60363=>"011011000",
  60364=>"000100100",
  60365=>"000111100",
  60366=>"001101001",
  60367=>"011100101",
  60368=>"011100001",
  60369=>"011101111",
  60370=>"000001011",
  60371=>"111011111",
  60372=>"101101111",
  60373=>"001011011",
  60374=>"111101101",
  60375=>"000001101",
  60376=>"010011011",
  60377=>"101101011",
  60378=>"100010111",
  60379=>"011001111",
  60380=>"111001101",
  60381=>"000001110",
  60382=>"101010010",
  60383=>"100011000",
  60384=>"010110000",
  60385=>"001110011",
  60386=>"011010011",
  60387=>"011001111",
  60388=>"001001011",
  60389=>"111011100",
  60390=>"110101110",
  60391=>"111010110",
  60392=>"010100001",
  60393=>"000000100",
  60394=>"111100111",
  60395=>"111100011",
  60396=>"010011110",
  60397=>"100111000",
  60398=>"111000100",
  60399=>"100111100",
  60400=>"111100111",
  60401=>"111000011",
  60402=>"111010001",
  60403=>"000000110",
  60404=>"110111011",
  60405=>"010110110",
  60406=>"000101100",
  60407=>"000001100",
  60408=>"100110111",
  60409=>"101101101",
  60410=>"100100111",
  60411=>"000100010",
  60412=>"001101000",
  60413=>"111001101",
  60414=>"011010000",
  60415=>"000011010",
  60416=>"011000001",
  60417=>"110111110",
  60418=>"010000011",
  60419=>"110110001",
  60420=>"111000100",
  60421=>"011101000",
  60422=>"001000111",
  60423=>"110101010",
  60424=>"000111110",
  60425=>"110001011",
  60426=>"101100111",
  60427=>"001010110",
  60428=>"001011111",
  60429=>"010111001",
  60430=>"111101101",
  60431=>"111001111",
  60432=>"001011110",
  60433=>"101110010",
  60434=>"101001101",
  60435=>"000111110",
  60436=>"110100010",
  60437=>"101010101",
  60438=>"000000101",
  60439=>"111001000",
  60440=>"010010010",
  60441=>"011001111",
  60442=>"000010101",
  60443=>"100110111",
  60444=>"101110000",
  60445=>"101111111",
  60446=>"011110111",
  60447=>"101110011",
  60448=>"101000001",
  60449=>"001000010",
  60450=>"111001101",
  60451=>"111101101",
  60452=>"100110010",
  60453=>"110101110",
  60454=>"001000100",
  60455=>"110111100",
  60456=>"111101001",
  60457=>"110000101",
  60458=>"001010100",
  60459=>"001110111",
  60460=>"011111010",
  60461=>"011111001",
  60462=>"100010100",
  60463=>"101011011",
  60464=>"010000100",
  60465=>"110111111",
  60466=>"101110100",
  60467=>"111011101",
  60468=>"100000100",
  60469=>"011011100",
  60470=>"000111101",
  60471=>"001001011",
  60472=>"001001000",
  60473=>"000100110",
  60474=>"100110010",
  60475=>"001101111",
  60476=>"011111110",
  60477=>"001100010",
  60478=>"010010000",
  60479=>"000100011",
  60480=>"100011001",
  60481=>"000000100",
  60482=>"101101011",
  60483=>"011110011",
  60484=>"011001110",
  60485=>"000001100",
  60486=>"101101000",
  60487=>"011010111",
  60488=>"110111010",
  60489=>"010001010",
  60490=>"101010111",
  60491=>"101100000",
  60492=>"101000111",
  60493=>"011001110",
  60494=>"101100111",
  60495=>"110111111",
  60496=>"000000010",
  60497=>"100000101",
  60498=>"000100101",
  60499=>"110001100",
  60500=>"001101000",
  60501=>"101101111",
  60502=>"111101011",
  60503=>"010000000",
  60504=>"111110000",
  60505=>"101000010",
  60506=>"110111101",
  60507=>"101001010",
  60508=>"111001011",
  60509=>"000000110",
  60510=>"000000110",
  60511=>"000111010",
  60512=>"101110101",
  60513=>"001010111",
  60514=>"101011101",
  60515=>"010110100",
  60516=>"001001000",
  60517=>"000001111",
  60518=>"010001000",
  60519=>"110101011",
  60520=>"100011001",
  60521=>"111011010",
  60522=>"001000101",
  60523=>"011101011",
  60524=>"111001110",
  60525=>"101000110",
  60526=>"010010111",
  60527=>"001111111",
  60528=>"101101100",
  60529=>"100001111",
  60530=>"000100100",
  60531=>"001110111",
  60532=>"011110111",
  60533=>"110010100",
  60534=>"001000011",
  60535=>"001010011",
  60536=>"001100100",
  60537=>"011111101",
  60538=>"101010011",
  60539=>"010001111",
  60540=>"000010010",
  60541=>"100111010",
  60542=>"100010110",
  60543=>"111001000",
  60544=>"110100101",
  60545=>"111111101",
  60546=>"111000000",
  60547=>"100001100",
  60548=>"011000000",
  60549=>"001101100",
  60550=>"110001010",
  60551=>"000010001",
  60552=>"111010111",
  60553=>"011010010",
  60554=>"001001011",
  60555=>"001100011",
  60556=>"111110101",
  60557=>"011111110",
  60558=>"000001101",
  60559=>"011011101",
  60560=>"111110101",
  60561=>"011101110",
  60562=>"110111000",
  60563=>"011111110",
  60564=>"000100011",
  60565=>"110110001",
  60566=>"010000000",
  60567=>"001000110",
  60568=>"000000001",
  60569=>"000000011",
  60570=>"111110000",
  60571=>"101111001",
  60572=>"010100011",
  60573=>"011101010",
  60574=>"100000100",
  60575=>"000000100",
  60576=>"110111010",
  60577=>"101100000",
  60578=>"010001011",
  60579=>"000111000",
  60580=>"010011110",
  60581=>"000100101",
  60582=>"100010100",
  60583=>"100000110",
  60584=>"111110010",
  60585=>"011101010",
  60586=>"111000001",
  60587=>"000001010",
  60588=>"000101000",
  60589=>"101010100",
  60590=>"101110100",
  60591=>"001011000",
  60592=>"001001101",
  60593=>"111011100",
  60594=>"110001000",
  60595=>"000001111",
  60596=>"110100011",
  60597=>"010110010",
  60598=>"110111000",
  60599=>"001011001",
  60600=>"111110111",
  60601=>"100001100",
  60602=>"010100110",
  60603=>"111111101",
  60604=>"010010010",
  60605=>"101001100",
  60606=>"010110110",
  60607=>"100010100",
  60608=>"000000111",
  60609=>"111110010",
  60610=>"110111000",
  60611=>"000010110",
  60612=>"111111010",
  60613=>"111010110",
  60614=>"001110111",
  60615=>"100000000",
  60616=>"011100111",
  60617=>"100001101",
  60618=>"010101001",
  60619=>"001001111",
  60620=>"010011011",
  60621=>"011011110",
  60622=>"011100110",
  60623=>"000011100",
  60624=>"001000100",
  60625=>"111111111",
  60626=>"010000000",
  60627=>"100110110",
  60628=>"001000010",
  60629=>"100111111",
  60630=>"011101100",
  60631=>"101000110",
  60632=>"000001010",
  60633=>"000000010",
  60634=>"011010001",
  60635=>"010001100",
  60636=>"110001001",
  60637=>"101100110",
  60638=>"000100000",
  60639=>"111101111",
  60640=>"000000111",
  60641=>"011010000",
  60642=>"101111100",
  60643=>"010000100",
  60644=>"011111001",
  60645=>"000100111",
  60646=>"000010111",
  60647=>"111111101",
  60648=>"011000010",
  60649=>"100100111",
  60650=>"101000100",
  60651=>"110000010",
  60652=>"011110101",
  60653=>"111110111",
  60654=>"011001111",
  60655=>"110010001",
  60656=>"001010110",
  60657=>"101001100",
  60658=>"000010100",
  60659=>"101011011",
  60660=>"100001100",
  60661=>"001101011",
  60662=>"101000011",
  60663=>"011100000",
  60664=>"001011101",
  60665=>"010010000",
  60666=>"100101001",
  60667=>"000001011",
  60668=>"001101100",
  60669=>"001110000",
  60670=>"111010001",
  60671=>"010000011",
  60672=>"100010011",
  60673=>"000111011",
  60674=>"000010110",
  60675=>"100001010",
  60676=>"111110110",
  60677=>"111111110",
  60678=>"010011101",
  60679=>"010101111",
  60680=>"111100000",
  60681=>"000101011",
  60682=>"101010010",
  60683=>"110000010",
  60684=>"101110111",
  60685=>"010001101",
  60686=>"100111001",
  60687=>"000010001",
  60688=>"100011011",
  60689=>"010111000",
  60690=>"000100011",
  60691=>"000001000",
  60692=>"010001011",
  60693=>"101001000",
  60694=>"110000111",
  60695=>"011001101",
  60696=>"101001101",
  60697=>"110101001",
  60698=>"011011111",
  60699=>"001000000",
  60700=>"010011011",
  60701=>"110100000",
  60702=>"101010110",
  60703=>"100011010",
  60704=>"000100100",
  60705=>"110101111",
  60706=>"111101100",
  60707=>"100101011",
  60708=>"010001101",
  60709=>"110101011",
  60710=>"110000000",
  60711=>"010011100",
  60712=>"010011111",
  60713=>"001000000",
  60714=>"010000011",
  60715=>"010011011",
  60716=>"010101111",
  60717=>"001000101",
  60718=>"000000111",
  60719=>"101000101",
  60720=>"000010111",
  60721=>"101000000",
  60722=>"001110111",
  60723=>"110010011",
  60724=>"110101010",
  60725=>"011011011",
  60726=>"001101100",
  60727=>"101110000",
  60728=>"010001101",
  60729=>"100000010",
  60730=>"111001000",
  60731=>"110010001",
  60732=>"100000001",
  60733=>"101001100",
  60734=>"101001100",
  60735=>"100101111",
  60736=>"101101111",
  60737=>"000001000",
  60738=>"101101111",
  60739=>"001100001",
  60740=>"010001110",
  60741=>"111101001",
  60742=>"000111101",
  60743=>"111100101",
  60744=>"100110111",
  60745=>"110001100",
  60746=>"111011001",
  60747=>"111000101",
  60748=>"101111101",
  60749=>"000110101",
  60750=>"001101100",
  60751=>"001101110",
  60752=>"101111000",
  60753=>"010111111",
  60754=>"010110010",
  60755=>"001100000",
  60756=>"000100010",
  60757=>"011111000",
  60758=>"010111111",
  60759=>"001110110",
  60760=>"010101110",
  60761=>"111100010",
  60762=>"111111010",
  60763=>"000110100",
  60764=>"101111010",
  60765=>"010111000",
  60766=>"011101111",
  60767=>"110100100",
  60768=>"101011010",
  60769=>"111110111",
  60770=>"111000001",
  60771=>"111000000",
  60772=>"101010110",
  60773=>"100011011",
  60774=>"000000000",
  60775=>"101101001",
  60776=>"001111110",
  60777=>"111000101",
  60778=>"011100000",
  60779=>"001001101",
  60780=>"000110001",
  60781=>"011001111",
  60782=>"101000111",
  60783=>"110001100",
  60784=>"101000011",
  60785=>"101011011",
  60786=>"010111001",
  60787=>"100001100",
  60788=>"000000110",
  60789=>"010001011",
  60790=>"101001100",
  60791=>"001110110",
  60792=>"000011000",
  60793=>"010010110",
  60794=>"111010111",
  60795=>"001100100",
  60796=>"110101010",
  60797=>"000100101",
  60798=>"101100010",
  60799=>"111100111",
  60800=>"100101011",
  60801=>"111001000",
  60802=>"010001000",
  60803=>"101110100",
  60804=>"010001000",
  60805=>"000011001",
  60806=>"001011011",
  60807=>"000110001",
  60808=>"001101110",
  60809=>"111011001",
  60810=>"100111011",
  60811=>"011000011",
  60812=>"101011111",
  60813=>"010011001",
  60814=>"010010111",
  60815=>"101110101",
  60816=>"011100000",
  60817=>"011000110",
  60818=>"110000100",
  60819=>"100100001",
  60820=>"100001001",
  60821=>"001110010",
  60822=>"111110111",
  60823=>"100010001",
  60824=>"000011111",
  60825=>"010111110",
  60826=>"100011000",
  60827=>"001001110",
  60828=>"011101100",
  60829=>"010010100",
  60830=>"010111111",
  60831=>"001110110",
  60832=>"010000000",
  60833=>"101101010",
  60834=>"101111001",
  60835=>"000000000",
  60836=>"101001111",
  60837=>"000000000",
  60838=>"001010011",
  60839=>"100110011",
  60840=>"111011001",
  60841=>"100111111",
  60842=>"111011000",
  60843=>"111001101",
  60844=>"100001110",
  60845=>"011011000",
  60846=>"011100010",
  60847=>"110100111",
  60848=>"011100111",
  60849=>"011111011",
  60850=>"001011010",
  60851=>"111010110",
  60852=>"000111101",
  60853=>"001001010",
  60854=>"110111100",
  60855=>"000100101",
  60856=>"101001010",
  60857=>"001101011",
  60858=>"001011010",
  60859=>"110010000",
  60860=>"000011010",
  60861=>"010111111",
  60862=>"000010001",
  60863=>"100001011",
  60864=>"100000000",
  60865=>"100110000",
  60866=>"011010101",
  60867=>"011101001",
  60868=>"110110100",
  60869=>"000110000",
  60870=>"110000001",
  60871=>"010001111",
  60872=>"011011110",
  60873=>"000111011",
  60874=>"101010011",
  60875=>"010111101",
  60876=>"101001000",
  60877=>"011110000",
  60878=>"101000001",
  60879=>"110110010",
  60880=>"100101111",
  60881=>"001100011",
  60882=>"000000101",
  60883=>"000001011",
  60884=>"011110110",
  60885=>"001011000",
  60886=>"011010010",
  60887=>"001000100",
  60888=>"001100110",
  60889=>"111000100",
  60890=>"111110101",
  60891=>"110100100",
  60892=>"011011100",
  60893=>"100110110",
  60894=>"010101000",
  60895=>"000100101",
  60896=>"111110011",
  60897=>"001011001",
  60898=>"011001101",
  60899=>"111001100",
  60900=>"001010010",
  60901=>"000100101",
  60902=>"000100001",
  60903=>"111000101",
  60904=>"010001101",
  60905=>"000011101",
  60906=>"100101100",
  60907=>"100000000",
  60908=>"101101010",
  60909=>"100001100",
  60910=>"110111101",
  60911=>"001001100",
  60912=>"101000111",
  60913=>"011001000",
  60914=>"110001000",
  60915=>"000001111",
  60916=>"001100111",
  60917=>"010011101",
  60918=>"110001011",
  60919=>"011101101",
  60920=>"011010001",
  60921=>"101110011",
  60922=>"100010010",
  60923=>"001100000",
  60924=>"111110110",
  60925=>"110000101",
  60926=>"000111001",
  60927=>"111000111",
  60928=>"011111000",
  60929=>"010001110",
  60930=>"001011100",
  60931=>"000000001",
  60932=>"001011101",
  60933=>"110101110",
  60934=>"011010110",
  60935=>"111101011",
  60936=>"111001001",
  60937=>"101111011",
  60938=>"000101011",
  60939=>"000000010",
  60940=>"111101001",
  60941=>"010101001",
  60942=>"110110010",
  60943=>"000100111",
  60944=>"001000001",
  60945=>"011000111",
  60946=>"011001001",
  60947=>"001111111",
  60948=>"000100110",
  60949=>"010110010",
  60950=>"010101000",
  60951=>"100100101",
  60952=>"000000101",
  60953=>"000110110",
  60954=>"100000101",
  60955=>"110110101",
  60956=>"101000101",
  60957=>"110001100",
  60958=>"100100111",
  60959=>"010101100",
  60960=>"000010011",
  60961=>"101101001",
  60962=>"011000001",
  60963=>"010100100",
  60964=>"101100011",
  60965=>"110101000",
  60966=>"010010000",
  60967=>"111101111",
  60968=>"011011001",
  60969=>"011000000",
  60970=>"011100001",
  60971=>"110100101",
  60972=>"000101101",
  60973=>"000010010",
  60974=>"111011000",
  60975=>"101000000",
  60976=>"111100010",
  60977=>"000011001",
  60978=>"000101101",
  60979=>"101011010",
  60980=>"101001011",
  60981=>"011100010",
  60982=>"110001001",
  60983=>"011001001",
  60984=>"111010010",
  60985=>"110101001",
  60986=>"111111000",
  60987=>"001000110",
  60988=>"001111101",
  60989=>"100100010",
  60990=>"000000100",
  60991=>"110010000",
  60992=>"101100111",
  60993=>"001001001",
  60994=>"100000000",
  60995=>"111000010",
  60996=>"110110000",
  60997=>"101100000",
  60998=>"010000100",
  60999=>"101010010",
  61000=>"100010011",
  61001=>"011010001",
  61002=>"111010101",
  61003=>"001101111",
  61004=>"110010100",
  61005=>"000000101",
  61006=>"011011101",
  61007=>"000101110",
  61008=>"001010010",
  61009=>"111110110",
  61010=>"101101100",
  61011=>"101001100",
  61012=>"110001110",
  61013=>"000001111",
  61014=>"110100011",
  61015=>"000101100",
  61016=>"010110011",
  61017=>"011001110",
  61018=>"001101111",
  61019=>"110100101",
  61020=>"111000010",
  61021=>"011000011",
  61022=>"001000000",
  61023=>"000001110",
  61024=>"001100000",
  61025=>"101011010",
  61026=>"000100000",
  61027=>"100000000",
  61028=>"011100010",
  61029=>"100100001",
  61030=>"001101000",
  61031=>"101000011",
  61032=>"000000100",
  61033=>"011111110",
  61034=>"011110010",
  61035=>"111000110",
  61036=>"111101111",
  61037=>"000111010",
  61038=>"010111011",
  61039=>"111001101",
  61040=>"101101101",
  61041=>"000001010",
  61042=>"100100101",
  61043=>"001010110",
  61044=>"100000001",
  61045=>"111010111",
  61046=>"101011111",
  61047=>"011010001",
  61048=>"110100101",
  61049=>"110000110",
  61050=>"111111110",
  61051=>"001011101",
  61052=>"000000010",
  61053=>"101010111",
  61054=>"001110011",
  61055=>"001011001",
  61056=>"000110011",
  61057=>"101111001",
  61058=>"011001101",
  61059=>"001000000",
  61060=>"011000111",
  61061=>"100110110",
  61062=>"110111110",
  61063=>"011011010",
  61064=>"100010000",
  61065=>"000000000",
  61066=>"000110100",
  61067=>"000001000",
  61068=>"001011001",
  61069=>"111100101",
  61070=>"111111011",
  61071=>"111000100",
  61072=>"110011001",
  61073=>"011010010",
  61074=>"111011111",
  61075=>"011101110",
  61076=>"100000011",
  61077=>"110101000",
  61078=>"000010001",
  61079=>"110000011",
  61080=>"010010001",
  61081=>"010101000",
  61082=>"000100001",
  61083=>"101101010",
  61084=>"111001011",
  61085=>"100011111",
  61086=>"110010011",
  61087=>"110110000",
  61088=>"100101110",
  61089=>"001111000",
  61090=>"100000101",
  61091=>"110110101",
  61092=>"010001001",
  61093=>"110001001",
  61094=>"100001110",
  61095=>"100001110",
  61096=>"100010001",
  61097=>"011000010",
  61098=>"000000011",
  61099=>"001001001",
  61100=>"101100000",
  61101=>"111010010",
  61102=>"100110111",
  61103=>"100000110",
  61104=>"001111000",
  61105=>"100110011",
  61106=>"000001011",
  61107=>"000101100",
  61108=>"010101101",
  61109=>"010100001",
  61110=>"110000111",
  61111=>"010100010",
  61112=>"111000001",
  61113=>"111000110",
  61114=>"011110011",
  61115=>"010100011",
  61116=>"111000011",
  61117=>"110011111",
  61118=>"000000011",
  61119=>"111100000",
  61120=>"010110011",
  61121=>"111001000",
  61122=>"101010100",
  61123=>"001010101",
  61124=>"110111111",
  61125=>"010010010",
  61126=>"110011100",
  61127=>"000100100",
  61128=>"110011100",
  61129=>"110100001",
  61130=>"011011111",
  61131=>"011001000",
  61132=>"110010010",
  61133=>"000000000",
  61134=>"011110110",
  61135=>"011011110",
  61136=>"100000011",
  61137=>"001000001",
  61138=>"110010001",
  61139=>"001011111",
  61140=>"101010100",
  61141=>"011100010",
  61142=>"000000010",
  61143=>"100001000",
  61144=>"001110111",
  61145=>"100110000",
  61146=>"100101100",
  61147=>"010011110",
  61148=>"101001110",
  61149=>"100000111",
  61150=>"001111111",
  61151=>"001001001",
  61152=>"110001110",
  61153=>"001111100",
  61154=>"010010010",
  61155=>"011000111",
  61156=>"000001100",
  61157=>"111010001",
  61158=>"100010111",
  61159=>"100011111",
  61160=>"111111010",
  61161=>"001010111",
  61162=>"111111110",
  61163=>"010001111",
  61164=>"001001011",
  61165=>"000001110",
  61166=>"110100000",
  61167=>"000010011",
  61168=>"010010010",
  61169=>"110100101",
  61170=>"100011000",
  61171=>"111001001",
  61172=>"111000010",
  61173=>"010111101",
  61174=>"110001100",
  61175=>"010100000",
  61176=>"011101100",
  61177=>"111011010",
  61178=>"011010111",
  61179=>"100101101",
  61180=>"100011000",
  61181=>"101111011",
  61182=>"010001001",
  61183=>"111101101",
  61184=>"100111100",
  61185=>"010011110",
  61186=>"000010111",
  61187=>"110000000",
  61188=>"010001001",
  61189=>"001011111",
  61190=>"101101110",
  61191=>"001111101",
  61192=>"110111000",
  61193=>"111000101",
  61194=>"011000011",
  61195=>"111110101",
  61196=>"111110101",
  61197=>"001101110",
  61198=>"000011100",
  61199=>"001010000",
  61200=>"110000111",
  61201=>"101111110",
  61202=>"111001000",
  61203=>"101111001",
  61204=>"011000101",
  61205=>"101101101",
  61206=>"011101001",
  61207=>"010110111",
  61208=>"000000001",
  61209=>"011101110",
  61210=>"000000000",
  61211=>"010011110",
  61212=>"100001100",
  61213=>"110000011",
  61214=>"110101110",
  61215=>"110100011",
  61216=>"001001001",
  61217=>"100010010",
  61218=>"000001110",
  61219=>"001000101",
  61220=>"100011101",
  61221=>"100001001",
  61222=>"110001101",
  61223=>"101010010",
  61224=>"111000000",
  61225=>"100000100",
  61226=>"101011110",
  61227=>"010111001",
  61228=>"100101001",
  61229=>"000110111",
  61230=>"111001011",
  61231=>"101111100",
  61232=>"000111111",
  61233=>"010111011",
  61234=>"111111000",
  61235=>"111000101",
  61236=>"100111111",
  61237=>"100000001",
  61238=>"011001010",
  61239=>"110000101",
  61240=>"011110101",
  61241=>"110110001",
  61242=>"111000001",
  61243=>"110000001",
  61244=>"000010100",
  61245=>"111011111",
  61246=>"100000000",
  61247=>"000000111",
  61248=>"000010101",
  61249=>"001001000",
  61250=>"010100010",
  61251=>"101101011",
  61252=>"010001101",
  61253=>"010100001",
  61254=>"110101111",
  61255=>"000000000",
  61256=>"101101001",
  61257=>"010111011",
  61258=>"101111010",
  61259=>"111110110",
  61260=>"010001011",
  61261=>"101101100",
  61262=>"100010111",
  61263=>"111010100",
  61264=>"111101000",
  61265=>"010001000",
  61266=>"001100010",
  61267=>"110011100",
  61268=>"111110101",
  61269=>"011000011",
  61270=>"000001111",
  61271=>"111011111",
  61272=>"110111100",
  61273=>"000111100",
  61274=>"000001000",
  61275=>"001010110",
  61276=>"011110111",
  61277=>"000010000",
  61278=>"001100011",
  61279=>"111001001",
  61280=>"000000010",
  61281=>"001111011",
  61282=>"000010100",
  61283=>"111100111",
  61284=>"011111000",
  61285=>"010010000",
  61286=>"100000000",
  61287=>"000000110",
  61288=>"111011110",
  61289=>"001000101",
  61290=>"101001110",
  61291=>"011101011",
  61292=>"011110100",
  61293=>"010000100",
  61294=>"101100100",
  61295=>"010000101",
  61296=>"100111100",
  61297=>"010011001",
  61298=>"101111110",
  61299=>"000010010",
  61300=>"011000101",
  61301=>"001000111",
  61302=>"111111111",
  61303=>"010001010",
  61304=>"011100100",
  61305=>"100111001",
  61306=>"101011101",
  61307=>"100111001",
  61308=>"010010001",
  61309=>"110000110",
  61310=>"000100011",
  61311=>"111101111",
  61312=>"100011111",
  61313=>"001010010",
  61314=>"001001000",
  61315=>"101110101",
  61316=>"000001111",
  61317=>"100010101",
  61318=>"100100100",
  61319=>"111011100",
  61320=>"111111110",
  61321=>"110000011",
  61322=>"000101011",
  61323=>"100001111",
  61324=>"100001110",
  61325=>"011000010",
  61326=>"011010000",
  61327=>"111110110",
  61328=>"100000100",
  61329=>"010010110",
  61330=>"110111100",
  61331=>"101010001",
  61332=>"000101100",
  61333=>"010001001",
  61334=>"001100001",
  61335=>"110000010",
  61336=>"110010101",
  61337=>"000110101",
  61338=>"001100111",
  61339=>"100000010",
  61340=>"010111011",
  61341=>"111001110",
  61342=>"010110000",
  61343=>"010100100",
  61344=>"011110110",
  61345=>"010001001",
  61346=>"110110000",
  61347=>"010001001",
  61348=>"011011001",
  61349=>"110001011",
  61350=>"101100110",
  61351=>"001000011",
  61352=>"101111111",
  61353=>"101010111",
  61354=>"000111001",
  61355=>"100110110",
  61356=>"101100101",
  61357=>"101110111",
  61358=>"010011000",
  61359=>"111111111",
  61360=>"000001100",
  61361=>"111111101",
  61362=>"001001000",
  61363=>"111000100",
  61364=>"010111001",
  61365=>"101010010",
  61366=>"100100010",
  61367=>"111010000",
  61368=>"101000010",
  61369=>"100101111",
  61370=>"000111101",
  61371=>"001000010",
  61372=>"011100110",
  61373=>"010000000",
  61374=>"000110000",
  61375=>"000100000",
  61376=>"110010010",
  61377=>"011111100",
  61378=>"000111000",
  61379=>"000000101",
  61380=>"110001011",
  61381=>"110101101",
  61382=>"000011000",
  61383=>"000110010",
  61384=>"000010010",
  61385=>"111011010",
  61386=>"101110010",
  61387=>"011110110",
  61388=>"100111110",
  61389=>"100000011",
  61390=>"000010010",
  61391=>"101000111",
  61392=>"001011101",
  61393=>"101100001",
  61394=>"010011010",
  61395=>"100001000",
  61396=>"101111111",
  61397=>"010000111",
  61398=>"001111110",
  61399=>"111000101",
  61400=>"110010111",
  61401=>"010100011",
  61402=>"111001100",
  61403=>"110100010",
  61404=>"110001100",
  61405=>"001101101",
  61406=>"000001101",
  61407=>"000001010",
  61408=>"000001011",
  61409=>"110110101",
  61410=>"011010001",
  61411=>"010001100",
  61412=>"101000111",
  61413=>"110000010",
  61414=>"111100010",
  61415=>"111000010",
  61416=>"000111000",
  61417=>"010100010",
  61418=>"010111110",
  61419=>"111011001",
  61420=>"100101000",
  61421=>"110000100",
  61422=>"011000010",
  61423=>"010010011",
  61424=>"000000111",
  61425=>"001010001",
  61426=>"110011011",
  61427=>"111101011",
  61428=>"101111010",
  61429=>"110001010",
  61430=>"101101001",
  61431=>"000001010",
  61432=>"011100111",
  61433=>"110111111",
  61434=>"111010010",
  61435=>"011010001",
  61436=>"100010011",
  61437=>"100010001",
  61438=>"000000110",
  61439=>"010110000",
  61440=>"011000000",
  61441=>"111110010",
  61442=>"110100010",
  61443=>"100101111",
  61444=>"000011100",
  61445=>"010100100",
  61446=>"100010001",
  61447=>"000000011",
  61448=>"010111100",
  61449=>"010010111",
  61450=>"000100101",
  61451=>"010011001",
  61452=>"101101110",
  61453=>"010011111",
  61454=>"101000100",
  61455=>"101101000",
  61456=>"110000001",
  61457=>"110111000",
  61458=>"000101000",
  61459=>"010110010",
  61460=>"010010001",
  61461=>"100100000",
  61462=>"011101110",
  61463=>"010100001",
  61464=>"110110101",
  61465=>"110101111",
  61466=>"111110000",
  61467=>"011001001",
  61468=>"000010010",
  61469=>"000111001",
  61470=>"011100100",
  61471=>"011011000",
  61472=>"010110110",
  61473=>"101100000",
  61474=>"011101101",
  61475=>"001110010",
  61476=>"001000100",
  61477=>"001010100",
  61478=>"110001001",
  61479=>"100011111",
  61480=>"110001111",
  61481=>"001101001",
  61482=>"000100101",
  61483=>"001001001",
  61484=>"000011000",
  61485=>"111100010",
  61486=>"010000001",
  61487=>"110101110",
  61488=>"011001000",
  61489=>"011011101",
  61490=>"010100100",
  61491=>"000111100",
  61492=>"101100110",
  61493=>"011011000",
  61494=>"100111100",
  61495=>"001011010",
  61496=>"000111001",
  61497=>"011000100",
  61498=>"100011101",
  61499=>"001111101",
  61500=>"111000000",
  61501=>"011000100",
  61502=>"110010011",
  61503=>"000101101",
  61504=>"100010001",
  61505=>"000010100",
  61506=>"011011001",
  61507=>"011011001",
  61508=>"101111001",
  61509=>"000111110",
  61510=>"011001001",
  61511=>"011100101",
  61512=>"100010101",
  61513=>"010100100",
  61514=>"000110110",
  61515=>"100110101",
  61516=>"011101000",
  61517=>"111101000",
  61518=>"111111101",
  61519=>"001101101",
  61520=>"100000110",
  61521=>"111111110",
  61522=>"011010111",
  61523=>"110010010",
  61524=>"110001101",
  61525=>"001110110",
  61526=>"110101111",
  61527=>"011111000",
  61528=>"001001101",
  61529=>"011010011",
  61530=>"101010101",
  61531=>"001010100",
  61532=>"101001111",
  61533=>"101100001",
  61534=>"100011011",
  61535=>"011101010",
  61536=>"101001000",
  61537=>"101001110",
  61538=>"010111110",
  61539=>"001100000",
  61540=>"010111110",
  61541=>"000101111",
  61542=>"111101011",
  61543=>"000110010",
  61544=>"000010101",
  61545=>"101010100",
  61546=>"110110110",
  61547=>"110000100",
  61548=>"111111001",
  61549=>"110101111",
  61550=>"010000000",
  61551=>"111110001",
  61552=>"010001010",
  61553=>"001100010",
  61554=>"111111000",
  61555=>"111100100",
  61556=>"110010111",
  61557=>"100000101",
  61558=>"100101111",
  61559=>"000111101",
  61560=>"110110111",
  61561=>"110101101",
  61562=>"010001000",
  61563=>"001001110",
  61564=>"010000010",
  61565=>"011110100",
  61566=>"111000110",
  61567=>"001110101",
  61568=>"110001101",
  61569=>"000010010",
  61570=>"000110000",
  61571=>"100001100",
  61572=>"000001011",
  61573=>"010101111",
  61574=>"000000101",
  61575=>"111101101",
  61576=>"010110010",
  61577=>"100111101",
  61578=>"100001100",
  61579=>"111010111",
  61580=>"110000001",
  61581=>"110100111",
  61582=>"110101011",
  61583=>"000001111",
  61584=>"110000101",
  61585=>"110010000",
  61586=>"000100011",
  61587=>"000101000",
  61588=>"101001100",
  61589=>"111000001",
  61590=>"111111101",
  61591=>"110001011",
  61592=>"011110010",
  61593=>"000011100",
  61594=>"001011101",
  61595=>"111010111",
  61596=>"101010100",
  61597=>"011101111",
  61598=>"101110010",
  61599=>"101110111",
  61600=>"101111000",
  61601=>"001101110",
  61602=>"111100100",
  61603=>"111010010",
  61604=>"001101001",
  61605=>"111011010",
  61606=>"010010010",
  61607=>"111111110",
  61608=>"011000000",
  61609=>"111110011",
  61610=>"101110010",
  61611=>"001100011",
  61612=>"100111111",
  61613=>"010111100",
  61614=>"101001100",
  61615=>"011101001",
  61616=>"100000101",
  61617=>"001000101",
  61618=>"101101111",
  61619=>"000111100",
  61620=>"000101000",
  61621=>"111001100",
  61622=>"000010100",
  61623=>"000001101",
  61624=>"010001100",
  61625=>"100011000",
  61626=>"011000101",
  61627=>"101010110",
  61628=>"011011111",
  61629=>"111111001",
  61630=>"000110011",
  61631=>"100011110",
  61632=>"101000110",
  61633=>"110011010",
  61634=>"001110111",
  61635=>"111101000",
  61636=>"001000110",
  61637=>"111111010",
  61638=>"111101101",
  61639=>"000010001",
  61640=>"000010001",
  61641=>"001010111",
  61642=>"101100101",
  61643=>"000111000",
  61644=>"010001101",
  61645=>"010101001",
  61646=>"011011011",
  61647=>"001011110",
  61648=>"000010100",
  61649=>"011110100",
  61650=>"110010001",
  61651=>"111100000",
  61652=>"001110010",
  61653=>"100110010",
  61654=>"100100001",
  61655=>"000100111",
  61656=>"100110011",
  61657=>"011010100",
  61658=>"100011001",
  61659=>"111011111",
  61660=>"110100111",
  61661=>"101101101",
  61662=>"001011100",
  61663=>"101000011",
  61664=>"111011101",
  61665=>"101010110",
  61666=>"010101111",
  61667=>"110000110",
  61668=>"100011100",
  61669=>"110111000",
  61670=>"101111000",
  61671=>"010101101",
  61672=>"101011010",
  61673=>"010011110",
  61674=>"010100011",
  61675=>"010111111",
  61676=>"110111000",
  61677=>"111100111",
  61678=>"110010111",
  61679=>"010111101",
  61680=>"001101100",
  61681=>"000101001",
  61682=>"101000010",
  61683=>"001010010",
  61684=>"011001101",
  61685=>"010000100",
  61686=>"110001001",
  61687=>"111001111",
  61688=>"000000110",
  61689=>"001000111",
  61690=>"001010111",
  61691=>"011101010",
  61692=>"001110101",
  61693=>"010100101",
  61694=>"101100000",
  61695=>"111000000",
  61696=>"010000011",
  61697=>"111110001",
  61698=>"001000001",
  61699=>"101111001",
  61700=>"000100111",
  61701=>"101001001",
  61702=>"100101011",
  61703=>"101000100",
  61704=>"101011000",
  61705=>"010001001",
  61706=>"001000010",
  61707=>"100100110",
  61708=>"101100001",
  61709=>"001110100",
  61710=>"011100101",
  61711=>"000001001",
  61712=>"101000000",
  61713=>"100101100",
  61714=>"010000111",
  61715=>"001010011",
  61716=>"111111010",
  61717=>"010010101",
  61718=>"110100000",
  61719=>"010100100",
  61720=>"001101000",
  61721=>"001100111",
  61722=>"001011111",
  61723=>"101011011",
  61724=>"110011111",
  61725=>"000000100",
  61726=>"111110111",
  61727=>"010000111",
  61728=>"111011101",
  61729=>"010010100",
  61730=>"001111001",
  61731=>"010001000",
  61732=>"111000111",
  61733=>"010011010",
  61734=>"000000110",
  61735=>"100000111",
  61736=>"011011011",
  61737=>"111111011",
  61738=>"000000000",
  61739=>"000001000",
  61740=>"010111111",
  61741=>"110011011",
  61742=>"001111111",
  61743=>"100101000",
  61744=>"011100010",
  61745=>"111100101",
  61746=>"011001000",
  61747=>"100000100",
  61748=>"001111010",
  61749=>"010010001",
  61750=>"010011011",
  61751=>"010110100",
  61752=>"110101101",
  61753=>"001111111",
  61754=>"001010110",
  61755=>"011101111",
  61756=>"001000001",
  61757=>"101111010",
  61758=>"101100010",
  61759=>"101001011",
  61760=>"101111000",
  61761=>"110110010",
  61762=>"111111110",
  61763=>"101111101",
  61764=>"101010010",
  61765=>"001111111",
  61766=>"000011010",
  61767=>"100000000",
  61768=>"001100100",
  61769=>"000000111",
  61770=>"010111001",
  61771=>"000110111",
  61772=>"001010011",
  61773=>"010111000",
  61774=>"011111001",
  61775=>"001001011",
  61776=>"100001000",
  61777=>"101101000",
  61778=>"001111010",
  61779=>"111001100",
  61780=>"010110101",
  61781=>"001100011",
  61782=>"100100100",
  61783=>"101110100",
  61784=>"000100110",
  61785=>"100001101",
  61786=>"111001000",
  61787=>"101111000",
  61788=>"100110001",
  61789=>"110010001",
  61790=>"010100001",
  61791=>"000110111",
  61792=>"001111000",
  61793=>"111110110",
  61794=>"101000010",
  61795=>"000000011",
  61796=>"000011001",
  61797=>"000110000",
  61798=>"110001010",
  61799=>"000100010",
  61800=>"001101011",
  61801=>"111001100",
  61802=>"000100101",
  61803=>"011111110",
  61804=>"101110101",
  61805=>"101110111",
  61806=>"010011110",
  61807=>"110100000",
  61808=>"111111001",
  61809=>"100011010",
  61810=>"000101111",
  61811=>"101001110",
  61812=>"001011001",
  61813=>"010011001",
  61814=>"011111111",
  61815=>"001010110",
  61816=>"100000111",
  61817=>"101101001",
  61818=>"011100011",
  61819=>"101000111",
  61820=>"110001001",
  61821=>"000100000",
  61822=>"111100011",
  61823=>"001110001",
  61824=>"101110101",
  61825=>"011111011",
  61826=>"000100001",
  61827=>"101000011",
  61828=>"110001110",
  61829=>"010110111",
  61830=>"000011111",
  61831=>"011101111",
  61832=>"111011001",
  61833=>"000010010",
  61834=>"101111110",
  61835=>"111000101",
  61836=>"000000100",
  61837=>"001000001",
  61838=>"010001000",
  61839=>"011000110",
  61840=>"001000111",
  61841=>"110110000",
  61842=>"000010000",
  61843=>"011110001",
  61844=>"010110001",
  61845=>"010011101",
  61846=>"001011011",
  61847=>"111001111",
  61848=>"000001011",
  61849=>"001000000",
  61850=>"111101011",
  61851=>"101110111",
  61852=>"100001111",
  61853=>"001100011",
  61854=>"110100100",
  61855=>"110100101",
  61856=>"101110100",
  61857=>"101101100",
  61858=>"000000100",
  61859=>"101100101",
  61860=>"110100111",
  61861=>"010000110",
  61862=>"111010010",
  61863=>"001010111",
  61864=>"000010000",
  61865=>"101111101",
  61866=>"110100010",
  61867=>"110111111",
  61868=>"111110000",
  61869=>"111011000",
  61870=>"111001010",
  61871=>"011011100",
  61872=>"001101101",
  61873=>"010001010",
  61874=>"101100100",
  61875=>"100001101",
  61876=>"011010001",
  61877=>"000010110",
  61878=>"011001100",
  61879=>"000001101",
  61880=>"011110101",
  61881=>"111000111",
  61882=>"001010110",
  61883=>"011111110",
  61884=>"110100001",
  61885=>"100011010",
  61886=>"000001001",
  61887=>"100011000",
  61888=>"111111111",
  61889=>"010011001",
  61890=>"010100010",
  61891=>"111011100",
  61892=>"001101011",
  61893=>"101001101",
  61894=>"100000101",
  61895=>"111100101",
  61896=>"001111111",
  61897=>"000001011",
  61898=>"101011010",
  61899=>"100101000",
  61900=>"000111010",
  61901=>"101110100",
  61902=>"011000110",
  61903=>"111010010",
  61904=>"010010000",
  61905=>"010000000",
  61906=>"000111011",
  61907=>"001000000",
  61908=>"111011111",
  61909=>"100000111",
  61910=>"111001101",
  61911=>"010101010",
  61912=>"001101101",
  61913=>"111100010",
  61914=>"001001100",
  61915=>"111011111",
  61916=>"000100010",
  61917=>"111110011",
  61918=>"010001111",
  61919=>"111100100",
  61920=>"111011000",
  61921=>"000001010",
  61922=>"110000000",
  61923=>"101110101",
  61924=>"101101000",
  61925=>"111011001",
  61926=>"110000000",
  61927=>"000000001",
  61928=>"100101000",
  61929=>"011010010",
  61930=>"001100110",
  61931=>"110100101",
  61932=>"111110011",
  61933=>"101101100",
  61934=>"111111100",
  61935=>"001101000",
  61936=>"000010011",
  61937=>"001101100",
  61938=>"001101100",
  61939=>"000001111",
  61940=>"101110101",
  61941=>"011101100",
  61942=>"010111100",
  61943=>"110110111",
  61944=>"111111011",
  61945=>"000011111",
  61946=>"111111100",
  61947=>"001100110",
  61948=>"001000001",
  61949=>"001001110",
  61950=>"011001011",
  61951=>"011101111",
  61952=>"100101111",
  61953=>"011000000",
  61954=>"001000101",
  61955=>"010110001",
  61956=>"100001110",
  61957=>"100111001",
  61958=>"110001011",
  61959=>"101110000",
  61960=>"000010010",
  61961=>"111110000",
  61962=>"110111101",
  61963=>"001100101",
  61964=>"000000010",
  61965=>"110011100",
  61966=>"111001000",
  61967=>"001001111",
  61968=>"001011100",
  61969=>"011111110",
  61970=>"110110010",
  61971=>"100100011",
  61972=>"111011000",
  61973=>"101100110",
  61974=>"010011010",
  61975=>"000001011",
  61976=>"001000000",
  61977=>"011011000",
  61978=>"101001001",
  61979=>"000111000",
  61980=>"100010110",
  61981=>"100000010",
  61982=>"100100011",
  61983=>"101001000",
  61984=>"100111001",
  61985=>"010000000",
  61986=>"001101001",
  61987=>"010110100",
  61988=>"000111000",
  61989=>"100101011",
  61990=>"000111010",
  61991=>"010010110",
  61992=>"110000101",
  61993=>"011111110",
  61994=>"111101110",
  61995=>"010011110",
  61996=>"001011110",
  61997=>"010001000",
  61998=>"101011000",
  61999=>"000101100",
  62000=>"110001010",
  62001=>"010110111",
  62002=>"000100101",
  62003=>"010111110",
  62004=>"101111111",
  62005=>"000011100",
  62006=>"110001011",
  62007=>"011101001",
  62008=>"100001111",
  62009=>"001011011",
  62010=>"101010101",
  62011=>"101100110",
  62012=>"000000010",
  62013=>"100100001",
  62014=>"101010001",
  62015=>"000000000",
  62016=>"110110001",
  62017=>"110100110",
  62018=>"100111111",
  62019=>"101010000",
  62020=>"101010010",
  62021=>"100001110",
  62022=>"111101010",
  62023=>"111110011",
  62024=>"001100001",
  62025=>"110011110",
  62026=>"111001010",
  62027=>"010000110",
  62028=>"111010100",
  62029=>"111111011",
  62030=>"101001001",
  62031=>"001101110",
  62032=>"000010101",
  62033=>"001001100",
  62034=>"101110111",
  62035=>"100001000",
  62036=>"000011010",
  62037=>"100001010",
  62038=>"000100001",
  62039=>"110101000",
  62040=>"000001110",
  62041=>"010000010",
  62042=>"101010010",
  62043=>"100011000",
  62044=>"011001111",
  62045=>"110000000",
  62046=>"000000000",
  62047=>"110110101",
  62048=>"010011111",
  62049=>"001010011",
  62050=>"110111011",
  62051=>"001010101",
  62052=>"111001001",
  62053=>"110110111",
  62054=>"010111001",
  62055=>"001011010",
  62056=>"000100010",
  62057=>"111010010",
  62058=>"010110100",
  62059=>"000010110",
  62060=>"010001101",
  62061=>"010000101",
  62062=>"000000010",
  62063=>"010001000",
  62064=>"001111011",
  62065=>"100000111",
  62066=>"011000110",
  62067=>"111110111",
  62068=>"000011100",
  62069=>"111101010",
  62070=>"101111110",
  62071=>"101001111",
  62072=>"111101110",
  62073=>"101110011",
  62074=>"101001000",
  62075=>"111101101",
  62076=>"011001010",
  62077=>"001000110",
  62078=>"111010101",
  62079=>"011001011",
  62080=>"101010011",
  62081=>"111100010",
  62082=>"101111100",
  62083=>"001001010",
  62084=>"110101001",
  62085=>"110101001",
  62086=>"101011001",
  62087=>"100000000",
  62088=>"110101000",
  62089=>"011111111",
  62090=>"001000000",
  62091=>"111001000",
  62092=>"011100011",
  62093=>"100011110",
  62094=>"011101000",
  62095=>"011110000",
  62096=>"110001110",
  62097=>"010011101",
  62098=>"111010110",
  62099=>"011001110",
  62100=>"111000000",
  62101=>"000100101",
  62102=>"010010101",
  62103=>"101111001",
  62104=>"100100001",
  62105=>"010000000",
  62106=>"100111101",
  62107=>"011101110",
  62108=>"001101001",
  62109=>"010000101",
  62110=>"010111001",
  62111=>"001101110",
  62112=>"010001010",
  62113=>"001010001",
  62114=>"111100101",
  62115=>"111100001",
  62116=>"110011000",
  62117=>"101101001",
  62118=>"100101010",
  62119=>"101011101",
  62120=>"010000001",
  62121=>"110110100",
  62122=>"110100010",
  62123=>"010010001",
  62124=>"001010010",
  62125=>"111000101",
  62126=>"111011110",
  62127=>"111101011",
  62128=>"101110101",
  62129=>"101000000",
  62130=>"001111010",
  62131=>"011001100",
  62132=>"011110111",
  62133=>"000000010",
  62134=>"101100011",
  62135=>"011111010",
  62136=>"001110010",
  62137=>"011010111",
  62138=>"010001110",
  62139=>"001010010",
  62140=>"011111000",
  62141=>"001111111",
  62142=>"001111100",
  62143=>"010001011",
  62144=>"000110001",
  62145=>"000011011",
  62146=>"010100110",
  62147=>"110000111",
  62148=>"100110100",
  62149=>"101100010",
  62150=>"010101111",
  62151=>"000101111",
  62152=>"011110000",
  62153=>"010101110",
  62154=>"110110011",
  62155=>"000111110",
  62156=>"111001001",
  62157=>"101011011",
  62158=>"110011011",
  62159=>"001000001",
  62160=>"111101001",
  62161=>"100010011",
  62162=>"001000110",
  62163=>"110111000",
  62164=>"101011111",
  62165=>"100001001",
  62166=>"000100011",
  62167=>"101000011",
  62168=>"101000111",
  62169=>"110100110",
  62170=>"010101111",
  62171=>"101111001",
  62172=>"101010101",
  62173=>"000110111",
  62174=>"101100010",
  62175=>"010001110",
  62176=>"111010111",
  62177=>"100100001",
  62178=>"111110000",
  62179=>"010111111",
  62180=>"100011010",
  62181=>"100001101",
  62182=>"100010010",
  62183=>"111111011",
  62184=>"001001000",
  62185=>"001101001",
  62186=>"111111111",
  62187=>"111110100",
  62188=>"000111011",
  62189=>"011110110",
  62190=>"001010100",
  62191=>"100111010",
  62192=>"101000000",
  62193=>"110100000",
  62194=>"100000010",
  62195=>"001110000",
  62196=>"011101101",
  62197=>"010001101",
  62198=>"011111101",
  62199=>"010001010",
  62200=>"110111100",
  62201=>"100000101",
  62202=>"000001011",
  62203=>"011000100",
  62204=>"010000111",
  62205=>"100110100",
  62206=>"100110001",
  62207=>"110100010",
  62208=>"011011001",
  62209=>"101000000",
  62210=>"111111010",
  62211=>"111100110",
  62212=>"000001000",
  62213=>"100010111",
  62214=>"011111110",
  62215=>"010010100",
  62216=>"001101111",
  62217=>"011000110",
  62218=>"000001101",
  62219=>"010101111",
  62220=>"010010110",
  62221=>"011110100",
  62222=>"011010001",
  62223=>"110100001",
  62224=>"000010000",
  62225=>"010100000",
  62226=>"111011101",
  62227=>"100101111",
  62228=>"110110000",
  62229=>"101011100",
  62230=>"110111110",
  62231=>"101101101",
  62232=>"111001011",
  62233=>"111100010",
  62234=>"101011101",
  62235=>"111001101",
  62236=>"110001101",
  62237=>"001001100",
  62238=>"101110100",
  62239=>"001000011",
  62240=>"011011100",
  62241=>"000010110",
  62242=>"011110111",
  62243=>"100010111",
  62244=>"110100010",
  62245=>"101000000",
  62246=>"110000111",
  62247=>"111100101",
  62248=>"100011010",
  62249=>"100101110",
  62250=>"010001010",
  62251=>"010011110",
  62252=>"110110000",
  62253=>"100011100",
  62254=>"101111000",
  62255=>"111001100",
  62256=>"101000101",
  62257=>"110100101",
  62258=>"001001010",
  62259=>"100001111",
  62260=>"100101110",
  62261=>"011111111",
  62262=>"010011111",
  62263=>"010111111",
  62264=>"100101000",
  62265=>"111101101",
  62266=>"111110001",
  62267=>"100011111",
  62268=>"010010010",
  62269=>"111000000",
  62270=>"001011100",
  62271=>"000110010",
  62272=>"111011111",
  62273=>"001010111",
  62274=>"001000000",
  62275=>"111111001",
  62276=>"110111100",
  62277=>"100110011",
  62278=>"111000000",
  62279=>"110111101",
  62280=>"111111110",
  62281=>"001101101",
  62282=>"101001001",
  62283=>"001111110",
  62284=>"110110101",
  62285=>"000100101",
  62286=>"110110111",
  62287=>"110001010",
  62288=>"111000001",
  62289=>"111000001",
  62290=>"010011110",
  62291=>"111110011",
  62292=>"110101001",
  62293=>"110001110",
  62294=>"100110001",
  62295=>"100010111",
  62296=>"111101010",
  62297=>"111000010",
  62298=>"011101100",
  62299=>"010100111",
  62300=>"101110110",
  62301=>"111101101",
  62302=>"000000100",
  62303=>"011010101",
  62304=>"011011011",
  62305=>"010110110",
  62306=>"010000010",
  62307=>"110010100",
  62308=>"100010100",
  62309=>"001001100",
  62310=>"111100001",
  62311=>"110101110",
  62312=>"000010111",
  62313=>"000101000",
  62314=>"111100000",
  62315=>"101011001",
  62316=>"101111101",
  62317=>"000011001",
  62318=>"010110111",
  62319=>"001000110",
  62320=>"000011000",
  62321=>"101111000",
  62322=>"010010011",
  62323=>"101100101",
  62324=>"111010111",
  62325=>"000110100",
  62326=>"001110100",
  62327=>"101111010",
  62328=>"110101001",
  62329=>"001100111",
  62330=>"100001111",
  62331=>"100010011",
  62332=>"011111000",
  62333=>"100111011",
  62334=>"110000010",
  62335=>"100001001",
  62336=>"010011000",
  62337=>"110001100",
  62338=>"010110101",
  62339=>"101100010",
  62340=>"101000010",
  62341=>"111011010",
  62342=>"101001110",
  62343=>"001011111",
  62344=>"111010000",
  62345=>"011110101",
  62346=>"111001100",
  62347=>"100101011",
  62348=>"001000100",
  62349=>"010110010",
  62350=>"110110101",
  62351=>"100110011",
  62352=>"111101111",
  62353=>"010000000",
  62354=>"011110000",
  62355=>"010000001",
  62356=>"101100101",
  62357=>"111111011",
  62358=>"011001000",
  62359=>"010000111",
  62360=>"111011101",
  62361=>"111001000",
  62362=>"011000101",
  62363=>"010110110",
  62364=>"110000010",
  62365=>"100100000",
  62366=>"101000100",
  62367=>"110011101",
  62368=>"100111011",
  62369=>"000110000",
  62370=>"110010110",
  62371=>"100001101",
  62372=>"000111100",
  62373=>"001010110",
  62374=>"000011001",
  62375=>"111100111",
  62376=>"011100000",
  62377=>"101110011",
  62378=>"100101111",
  62379=>"101001011",
  62380=>"000111110",
  62381=>"111110100",
  62382=>"010011000",
  62383=>"001111011",
  62384=>"100111100",
  62385=>"101011101",
  62386=>"101010010",
  62387=>"011000101",
  62388=>"000101110",
  62389=>"111011111",
  62390=>"111110100",
  62391=>"101101001",
  62392=>"100000001",
  62393=>"001111010",
  62394=>"101001110",
  62395=>"011000110",
  62396=>"101101011",
  62397=>"000000000",
  62398=>"101111010",
  62399=>"001101010",
  62400=>"000101011",
  62401=>"010110101",
  62402=>"001111000",
  62403=>"101000100",
  62404=>"010100001",
  62405=>"110000000",
  62406=>"111010100",
  62407=>"011110111",
  62408=>"101111100",
  62409=>"000101101",
  62410=>"100001111",
  62411=>"011111111",
  62412=>"011011001",
  62413=>"010110110",
  62414=>"110110011",
  62415=>"001100011",
  62416=>"010100110",
  62417=>"001000110",
  62418=>"101111000",
  62419=>"001001101",
  62420=>"000001010",
  62421=>"101100001",
  62422=>"001110000",
  62423=>"101101010",
  62424=>"101010011",
  62425=>"001111001",
  62426=>"100100111",
  62427=>"011111111",
  62428=>"010101011",
  62429=>"001010010",
  62430=>"100110011",
  62431=>"001111011",
  62432=>"110001111",
  62433=>"110011001",
  62434=>"100000001",
  62435=>"100100001",
  62436=>"000100001",
  62437=>"101111000",
  62438=>"010001101",
  62439=>"000100001",
  62440=>"000000010",
  62441=>"010101110",
  62442=>"000001010",
  62443=>"110100100",
  62444=>"010000011",
  62445=>"010100000",
  62446=>"110110111",
  62447=>"001101010",
  62448=>"101000010",
  62449=>"111111011",
  62450=>"000110111",
  62451=>"111101101",
  62452=>"111001000",
  62453=>"010100100",
  62454=>"000100010",
  62455=>"111111110",
  62456=>"101000011",
  62457=>"111111011",
  62458=>"001000011",
  62459=>"001000110",
  62460=>"010111001",
  62461=>"011010000",
  62462=>"000101010",
  62463=>"000100101",
  62464=>"110100100",
  62465=>"000110101",
  62466=>"100111010",
  62467=>"001000100",
  62468=>"111101111",
  62469=>"011000011",
  62470=>"010001100",
  62471=>"000111011",
  62472=>"011100000",
  62473=>"010011110",
  62474=>"111101010",
  62475=>"101100111",
  62476=>"111000001",
  62477=>"001111010",
  62478=>"101000010",
  62479=>"010100010",
  62480=>"111101111",
  62481=>"111011001",
  62482=>"111110110",
  62483=>"001001111",
  62484=>"101111001",
  62485=>"011100110",
  62486=>"111111101",
  62487=>"001010110",
  62488=>"010110110",
  62489=>"100010110",
  62490=>"110110010",
  62491=>"101111001",
  62492=>"101100001",
  62493=>"011010101",
  62494=>"011000000",
  62495=>"011000100",
  62496=>"100100111",
  62497=>"100101000",
  62498=>"111011000",
  62499=>"000011111",
  62500=>"111110010",
  62501=>"000101001",
  62502=>"101101001",
  62503=>"101101001",
  62504=>"101001011",
  62505=>"000101101",
  62506=>"101011010",
  62507=>"000001111",
  62508=>"011011011",
  62509=>"111100010",
  62510=>"011010010",
  62511=>"011110011",
  62512=>"000010100",
  62513=>"000000010",
  62514=>"000101001",
  62515=>"110111110",
  62516=>"110100100",
  62517=>"110010011",
  62518=>"001010100",
  62519=>"000010100",
  62520=>"010110000",
  62521=>"111101101",
  62522=>"011100000",
  62523=>"101100000",
  62524=>"001010000",
  62525=>"100000000",
  62526=>"101111000",
  62527=>"100110101",
  62528=>"100000001",
  62529=>"101000111",
  62530=>"110101100",
  62531=>"001100100",
  62532=>"111110110",
  62533=>"100111111",
  62534=>"111011101",
  62535=>"011011100",
  62536=>"001110110",
  62537=>"110010010",
  62538=>"110011001",
  62539=>"100000000",
  62540=>"010100100",
  62541=>"010000110",
  62542=>"010000001",
  62543=>"101110100",
  62544=>"100111010",
  62545=>"101100000",
  62546=>"111000100",
  62547=>"101101100",
  62548=>"111001100",
  62549=>"011100101",
  62550=>"011011100",
  62551=>"001011011",
  62552=>"010101010",
  62553=>"110011010",
  62554=>"000010100",
  62555=>"010010000",
  62556=>"010111000",
  62557=>"100000111",
  62558=>"011000000",
  62559=>"110111111",
  62560=>"111000010",
  62561=>"100001000",
  62562=>"000010010",
  62563=>"011101110",
  62564=>"011010010",
  62565=>"001110011",
  62566=>"011011010",
  62567=>"001011110",
  62568=>"100000011",
  62569=>"010000111",
  62570=>"101100001",
  62571=>"001001000",
  62572=>"010010010",
  62573=>"110100010",
  62574=>"011001111",
  62575=>"100110010",
  62576=>"001110000",
  62577=>"111110111",
  62578=>"011001111",
  62579=>"111001011",
  62580=>"110001111",
  62581=>"001100100",
  62582=>"110010110",
  62583=>"111001100",
  62584=>"101011100",
  62585=>"110000011",
  62586=>"000010000",
  62587=>"101010111",
  62588=>"101101000",
  62589=>"000010100",
  62590=>"101000000",
  62591=>"001111111",
  62592=>"000111100",
  62593=>"011011101",
  62594=>"100100010",
  62595=>"100100010",
  62596=>"011100110",
  62597=>"111001111",
  62598=>"101000100",
  62599=>"010111000",
  62600=>"011110001",
  62601=>"110011101",
  62602=>"111110100",
  62603=>"100110110",
  62604=>"110000100",
  62605=>"011100010",
  62606=>"110000110",
  62607=>"101100011",
  62608=>"100000101",
  62609=>"111010101",
  62610=>"100111110",
  62611=>"111011110",
  62612=>"001100001",
  62613=>"010100000",
  62614=>"011111010",
  62615=>"010110110",
  62616=>"011001000",
  62617=>"111100110",
  62618=>"101101011",
  62619=>"010110110",
  62620=>"100010110",
  62621=>"000110001",
  62622=>"101110100",
  62623=>"111011011",
  62624=>"110101010",
  62625=>"000110110",
  62626=>"000000101",
  62627=>"111000110",
  62628=>"110110111",
  62629=>"101100001",
  62630=>"001011000",
  62631=>"101110010",
  62632=>"111111101",
  62633=>"101011111",
  62634=>"010110011",
  62635=>"110100011",
  62636=>"000101101",
  62637=>"100010001",
  62638=>"110000100",
  62639=>"000000000",
  62640=>"111111011",
  62641=>"011011001",
  62642=>"101100111",
  62643=>"100001100",
  62644=>"100010010",
  62645=>"101101001",
  62646=>"110110011",
  62647=>"010010100",
  62648=>"000101011",
  62649=>"001101001",
  62650=>"101101100",
  62651=>"000101111",
  62652=>"000110101",
  62653=>"111001010",
  62654=>"111111001",
  62655=>"001100001",
  62656=>"100111000",
  62657=>"001010010",
  62658=>"001101110",
  62659=>"110000110",
  62660=>"111111010",
  62661=>"111111011",
  62662=>"000000111",
  62663=>"101110110",
  62664=>"000111011",
  62665=>"110010101",
  62666=>"000010100",
  62667=>"010100010",
  62668=>"001100100",
  62669=>"001111100",
  62670=>"001111001",
  62671=>"000111101",
  62672=>"100011000",
  62673=>"001101010",
  62674=>"101000101",
  62675=>"000000001",
  62676=>"101101100",
  62677=>"000011111",
  62678=>"001010010",
  62679=>"101011110",
  62680=>"110100100",
  62681=>"111010110",
  62682=>"000000010",
  62683=>"110010011",
  62684=>"110101100",
  62685=>"001111111",
  62686=>"100110100",
  62687=>"111000010",
  62688=>"100011101",
  62689=>"111011111",
  62690=>"000010100",
  62691=>"110011111",
  62692=>"010000011",
  62693=>"000011011",
  62694=>"011111001",
  62695=>"011000011",
  62696=>"011010011",
  62697=>"011100100",
  62698=>"000010110",
  62699=>"101001101",
  62700=>"010110100",
  62701=>"101010110",
  62702=>"110110011",
  62703=>"011111000",
  62704=>"011110101",
  62705=>"011011110",
  62706=>"010100111",
  62707=>"110100100",
  62708=>"110100011",
  62709=>"011001101",
  62710=>"000101000",
  62711=>"010010100",
  62712=>"011011110",
  62713=>"111001000",
  62714=>"000010110",
  62715=>"110011010",
  62716=>"011000011",
  62717=>"000101010",
  62718=>"010011101",
  62719=>"011110111",
  62720=>"111101011",
  62721=>"110101011",
  62722=>"000111001",
  62723=>"110111011",
  62724=>"111011011",
  62725=>"011100011",
  62726=>"110000011",
  62727=>"011101000",
  62728=>"001011111",
  62729=>"111110101",
  62730=>"100100111",
  62731=>"010011011",
  62732=>"000000011",
  62733=>"011100001",
  62734=>"010111111",
  62735=>"101000011",
  62736=>"110001100",
  62737=>"000010000",
  62738=>"001111100",
  62739=>"100111000",
  62740=>"100100011",
  62741=>"000011101",
  62742=>"010100101",
  62743=>"100100100",
  62744=>"001110001",
  62745=>"010110001",
  62746=>"100110111",
  62747=>"101110110",
  62748=>"010010101",
  62749=>"110101110",
  62750=>"011100101",
  62751=>"101100000",
  62752=>"010110001",
  62753=>"010110001",
  62754=>"110010011",
  62755=>"111000101",
  62756=>"100011101",
  62757=>"010010011",
  62758=>"101001101",
  62759=>"000011100",
  62760=>"001110110",
  62761=>"101110100",
  62762=>"011001011",
  62763=>"110100001",
  62764=>"100100110",
  62765=>"000000111",
  62766=>"110110110",
  62767=>"001101001",
  62768=>"101000101",
  62769=>"000100010",
  62770=>"010110011",
  62771=>"001100110",
  62772=>"101100000",
  62773=>"100000101",
  62774=>"101001001",
  62775=>"010010001",
  62776=>"001011110",
  62777=>"100111001",
  62778=>"000000111",
  62779=>"010110110",
  62780=>"110111000",
  62781=>"101111110",
  62782=>"101111011",
  62783=>"100111011",
  62784=>"011110000",
  62785=>"111010001",
  62786=>"110101100",
  62787=>"100110101",
  62788=>"011010010",
  62789=>"011010110",
  62790=>"111101010",
  62791=>"011111110",
  62792=>"010101011",
  62793=>"010110010",
  62794=>"100001100",
  62795=>"000001100",
  62796=>"101100000",
  62797=>"000000111",
  62798=>"100010011",
  62799=>"001011001",
  62800=>"101100011",
  62801=>"111010110",
  62802=>"100110111",
  62803=>"110100001",
  62804=>"000100101",
  62805=>"101111110",
  62806=>"001011001",
  62807=>"111011111",
  62808=>"000010110",
  62809=>"110110011",
  62810=>"100110011",
  62811=>"010101001",
  62812=>"100110100",
  62813=>"011110011",
  62814=>"011110111",
  62815=>"110100000",
  62816=>"000110110",
  62817=>"111110011",
  62818=>"110000001",
  62819=>"001110101",
  62820=>"010000101",
  62821=>"111110000",
  62822=>"000110100",
  62823=>"000001010",
  62824=>"011000100",
  62825=>"100011111",
  62826=>"110101000",
  62827=>"011010101",
  62828=>"101101000",
  62829=>"111100110",
  62830=>"101101101",
  62831=>"000100001",
  62832=>"001011111",
  62833=>"101011100",
  62834=>"001000010",
  62835=>"101001111",
  62836=>"000001001",
  62837=>"110100000",
  62838=>"010100001",
  62839=>"110000110",
  62840=>"101011111",
  62841=>"101000100",
  62842=>"101111100",
  62843=>"000110001",
  62844=>"111110100",
  62845=>"110011101",
  62846=>"001000011",
  62847=>"111100100",
  62848=>"110011111",
  62849=>"001111101",
  62850=>"111101111",
  62851=>"110010111",
  62852=>"111010111",
  62853=>"111110001",
  62854=>"111110000",
  62855=>"010001101",
  62856=>"110110001",
  62857=>"010010100",
  62858=>"000010101",
  62859=>"111111100",
  62860=>"010010010",
  62861=>"001010100",
  62862=>"000001100",
  62863=>"101100001",
  62864=>"011100100",
  62865=>"111110000",
  62866=>"111001111",
  62867=>"100101100",
  62868=>"110001100",
  62869=>"000000111",
  62870=>"000000001",
  62871=>"111110110",
  62872=>"111100110",
  62873=>"001010111",
  62874=>"011111000",
  62875=>"101010010",
  62876=>"011011010",
  62877=>"011010011",
  62878=>"100110110",
  62879=>"101000111",
  62880=>"011010010",
  62881=>"111001000",
  62882=>"111100011",
  62883=>"100111010",
  62884=>"011111110",
  62885=>"000100111",
  62886=>"011101000",
  62887=>"110000011",
  62888=>"110111011",
  62889=>"001100000",
  62890=>"001001111",
  62891=>"111000111",
  62892=>"101101000",
  62893=>"011101011",
  62894=>"100100000",
  62895=>"010000111",
  62896=>"110000111",
  62897=>"000000100",
  62898=>"101011110",
  62899=>"111011011",
  62900=>"011100011",
  62901=>"111111011",
  62902=>"001000110",
  62903=>"111110111",
  62904=>"110111011",
  62905=>"011101000",
  62906=>"101111111",
  62907=>"111111110",
  62908=>"111011111",
  62909=>"111111101",
  62910=>"100101010",
  62911=>"110100010",
  62912=>"010111011",
  62913=>"101100111",
  62914=>"010111000",
  62915=>"110010010",
  62916=>"001010000",
  62917=>"011111110",
  62918=>"111010110",
  62919=>"011000000",
  62920=>"110111101",
  62921=>"101001100",
  62922=>"000101110",
  62923=>"101001000",
  62924=>"010010011",
  62925=>"110000011",
  62926=>"010000010",
  62927=>"011000000",
  62928=>"110101001",
  62929=>"011110011",
  62930=>"011110011",
  62931=>"110001001",
  62932=>"100101111",
  62933=>"001011010",
  62934=>"011010010",
  62935=>"111111110",
  62936=>"101110111",
  62937=>"010100000",
  62938=>"101001011",
  62939=>"010111000",
  62940=>"000011100",
  62941=>"111100110",
  62942=>"100000111",
  62943=>"010110110",
  62944=>"110100101",
  62945=>"010100011",
  62946=>"010011001",
  62947=>"101110010",
  62948=>"000110011",
  62949=>"110000111",
  62950=>"000001100",
  62951=>"000011000",
  62952=>"011101000",
  62953=>"011101010",
  62954=>"110110100",
  62955=>"010110101",
  62956=>"111110011",
  62957=>"001000010",
  62958=>"101110011",
  62959=>"001101011",
  62960=>"101001001",
  62961=>"111101011",
  62962=>"111011011",
  62963=>"110100011",
  62964=>"110101001",
  62965=>"001101101",
  62966=>"100001010",
  62967=>"111100101",
  62968=>"011010110",
  62969=>"101011011",
  62970=>"001000011",
  62971=>"111101011",
  62972=>"100110110",
  62973=>"000000111",
  62974=>"111111101",
  62975=>"100110000",
  62976=>"110000011",
  62977=>"100000011",
  62978=>"101100111",
  62979=>"001001001",
  62980=>"110001010",
  62981=>"101101110",
  62982=>"101100000",
  62983=>"111100001",
  62984=>"010000111",
  62985=>"000110111",
  62986=>"010011000",
  62987=>"001100011",
  62988=>"000101011",
  62989=>"110010101",
  62990=>"001101010",
  62991=>"011011110",
  62992=>"001011100",
  62993=>"111111000",
  62994=>"001011111",
  62995=>"100110100",
  62996=>"011110001",
  62997=>"100100110",
  62998=>"101000110",
  62999=>"110111011",
  63000=>"101111100",
  63001=>"010000000",
  63002=>"100111111",
  63003=>"110010100",
  63004=>"110011101",
  63005=>"100011000",
  63006=>"000001010",
  63007=>"111100010",
  63008=>"000010010",
  63009=>"111110010",
  63010=>"000101010",
  63011=>"111011111",
  63012=>"101000111",
  63013=>"001101101",
  63014=>"011000011",
  63015=>"001110000",
  63016=>"011001110",
  63017=>"010011100",
  63018=>"000100111",
  63019=>"101001111",
  63020=>"101000101",
  63021=>"001100100",
  63022=>"110110011",
  63023=>"010010011",
  63024=>"000110111",
  63025=>"101011011",
  63026=>"101000101",
  63027=>"001101100",
  63028=>"010010100",
  63029=>"110110011",
  63030=>"011010110",
  63031=>"111111000",
  63032=>"001111010",
  63033=>"110000011",
  63034=>"101000100",
  63035=>"110110100",
  63036=>"111100011",
  63037=>"000000101",
  63038=>"010001010",
  63039=>"111100010",
  63040=>"101011011",
  63041=>"111110100",
  63042=>"111000111",
  63043=>"000111100",
  63044=>"100000101",
  63045=>"100010001",
  63046=>"010001000",
  63047=>"010111000",
  63048=>"010011011",
  63049=>"111001001",
  63050=>"111001010",
  63051=>"000100110",
  63052=>"111101110",
  63053=>"001000101",
  63054=>"000010101",
  63055=>"100101110",
  63056=>"001010010",
  63057=>"011100010",
  63058=>"100010010",
  63059=>"000101110",
  63060=>"110001100",
  63061=>"001001101",
  63062=>"001000100",
  63063=>"010011000",
  63064=>"100011011",
  63065=>"011101110",
  63066=>"011101101",
  63067=>"111001010",
  63068=>"001101000",
  63069=>"001110000",
  63070=>"100001100",
  63071=>"111110000",
  63072=>"011000001",
  63073=>"010110001",
  63074=>"011111100",
  63075=>"011011101",
  63076=>"001110111",
  63077=>"011101001",
  63078=>"111110100",
  63079=>"000101000",
  63080=>"011011001",
  63081=>"001100100",
  63082=>"111011111",
  63083=>"010001010",
  63084=>"111101000",
  63085=>"000000111",
  63086=>"000100011",
  63087=>"001111100",
  63088=>"110011000",
  63089=>"101111110",
  63090=>"010010001",
  63091=>"000000001",
  63092=>"100110101",
  63093=>"100000010",
  63094=>"011000101",
  63095=>"110100101",
  63096=>"000010110",
  63097=>"010000010",
  63098=>"000011000",
  63099=>"110011010",
  63100=>"110010011",
  63101=>"000000101",
  63102=>"011100000",
  63103=>"101000101",
  63104=>"111011000",
  63105=>"001110111",
  63106=>"010110000",
  63107=>"001100100",
  63108=>"011011011",
  63109=>"000000000",
  63110=>"000110010",
  63111=>"111111010",
  63112=>"100011110",
  63113=>"010001110",
  63114=>"101011110",
  63115=>"100010011",
  63116=>"111111001",
  63117=>"010110010",
  63118=>"110100101",
  63119=>"001000100",
  63120=>"010110011",
  63121=>"110101001",
  63122=>"100100101",
  63123=>"111100010",
  63124=>"001010001",
  63125=>"011001010",
  63126=>"110010010",
  63127=>"000110000",
  63128=>"111010010",
  63129=>"001011101",
  63130=>"101011001",
  63131=>"101110100",
  63132=>"100110110",
  63133=>"000010111",
  63134=>"000001110",
  63135=>"011000011",
  63136=>"111100011",
  63137=>"011000010",
  63138=>"000010101",
  63139=>"110110011",
  63140=>"111111001",
  63141=>"001111101",
  63142=>"010111001",
  63143=>"110110000",
  63144=>"110100000",
  63145=>"000000011",
  63146=>"010101010",
  63147=>"111110110",
  63148=>"110000001",
  63149=>"000010111",
  63150=>"001110101",
  63151=>"111001111",
  63152=>"000111000",
  63153=>"111001000",
  63154=>"000001000",
  63155=>"111011011",
  63156=>"010111000",
  63157=>"100111011",
  63158=>"011110000",
  63159=>"011111110",
  63160=>"110001000",
  63161=>"010110001",
  63162=>"001101101",
  63163=>"000101001",
  63164=>"011010001",
  63165=>"100010001",
  63166=>"100011101",
  63167=>"111101100",
  63168=>"111100111",
  63169=>"010010101",
  63170=>"111000000",
  63171=>"111011101",
  63172=>"101101000",
  63173=>"000001110",
  63174=>"000100000",
  63175=>"100100101",
  63176=>"000011100",
  63177=>"100100001",
  63178=>"000001101",
  63179=>"010010000",
  63180=>"110100101",
  63181=>"111111101",
  63182=>"001011010",
  63183=>"010000100",
  63184=>"000101001",
  63185=>"110000101",
  63186=>"101010101",
  63187=>"011010111",
  63188=>"001011001",
  63189=>"100010010",
  63190=>"000010010",
  63191=>"001100100",
  63192=>"000000011",
  63193=>"110101000",
  63194=>"010011001",
  63195=>"100101111",
  63196=>"100000101",
  63197=>"000101010",
  63198=>"000110011",
  63199=>"100001111",
  63200=>"000100001",
  63201=>"111011011",
  63202=>"111001000",
  63203=>"011101010",
  63204=>"011010100",
  63205=>"111100010",
  63206=>"101111001",
  63207=>"101011010",
  63208=>"010000001",
  63209=>"010100000",
  63210=>"110111010",
  63211=>"001101010",
  63212=>"011101111",
  63213=>"010000001",
  63214=>"100111111",
  63215=>"001111101",
  63216=>"111110111",
  63217=>"101011001",
  63218=>"011101000",
  63219=>"111100010",
  63220=>"110110001",
  63221=>"010101001",
  63222=>"110111010",
  63223=>"110100001",
  63224=>"011010011",
  63225=>"011001001",
  63226=>"110001101",
  63227=>"100111111",
  63228=>"101100101",
  63229=>"000000011",
  63230=>"111110100",
  63231=>"100100011",
  63232=>"100011110",
  63233=>"001111110",
  63234=>"011001000",
  63235=>"100001001",
  63236=>"001011001",
  63237=>"110001000",
  63238=>"110111101",
  63239=>"111011101",
  63240=>"101011010",
  63241=>"000111010",
  63242=>"010000111",
  63243=>"011100101",
  63244=>"000001010",
  63245=>"100101000",
  63246=>"011010110",
  63247=>"001110011",
  63248=>"110011000",
  63249=>"000000111",
  63250=>"011000000",
  63251=>"111110011",
  63252=>"100000000",
  63253=>"001100011",
  63254=>"001011101",
  63255=>"011000011",
  63256=>"111100101",
  63257=>"000000010",
  63258=>"010111100",
  63259=>"000100011",
  63260=>"101010111",
  63261=>"111010000",
  63262=>"010011111",
  63263=>"001011000",
  63264=>"110111111",
  63265=>"000101111",
  63266=>"010001110",
  63267=>"111110101",
  63268=>"101001111",
  63269=>"010000000",
  63270=>"101011110",
  63271=>"000000101",
  63272=>"010100000",
  63273=>"001001010",
  63274=>"110110001",
  63275=>"111011111",
  63276=>"101110101",
  63277=>"001000000",
  63278=>"000011101",
  63279=>"011011111",
  63280=>"001000110",
  63281=>"110101001",
  63282=>"100110011",
  63283=>"110000101",
  63284=>"010000101",
  63285=>"000100110",
  63286=>"100101000",
  63287=>"000001010",
  63288=>"000011001",
  63289=>"010111010",
  63290=>"101001010",
  63291=>"110000001",
  63292=>"011101000",
  63293=>"100111111",
  63294=>"011111100",
  63295=>"001000111",
  63296=>"010011101",
  63297=>"110101110",
  63298=>"111111000",
  63299=>"111011000",
  63300=>"011010010",
  63301=>"010111001",
  63302=>"001001010",
  63303=>"001111011",
  63304=>"010101011",
  63305=>"000101011",
  63306=>"011101110",
  63307=>"001111011",
  63308=>"010110111",
  63309=>"101111100",
  63310=>"001100000",
  63311=>"010111001",
  63312=>"111011100",
  63313=>"001100111",
  63314=>"111100101",
  63315=>"100010110",
  63316=>"111010100",
  63317=>"110001000",
  63318=>"101011011",
  63319=>"101010110",
  63320=>"010001010",
  63321=>"100010100",
  63322=>"110111010",
  63323=>"100101010",
  63324=>"001001101",
  63325=>"001110100",
  63326=>"010111011",
  63327=>"000111100",
  63328=>"101001001",
  63329=>"101110100",
  63330=>"101101011",
  63331=>"001111000",
  63332=>"000010111",
  63333=>"110011101",
  63334=>"001101011",
  63335=>"001000101",
  63336=>"001100001",
  63337=>"111101010",
  63338=>"000000101",
  63339=>"000101101",
  63340=>"001001111",
  63341=>"111101001",
  63342=>"100000101",
  63343=>"011100101",
  63344=>"100010100",
  63345=>"110000101",
  63346=>"001001001",
  63347=>"000110111",
  63348=>"010010110",
  63349=>"111001001",
  63350=>"000000000",
  63351=>"100001110",
  63352=>"111101100",
  63353=>"000001111",
  63354=>"011001011",
  63355=>"010100001",
  63356=>"011000000",
  63357=>"101011101",
  63358=>"110011101",
  63359=>"110011011",
  63360=>"010001010",
  63361=>"100001101",
  63362=>"101111101",
  63363=>"110111000",
  63364=>"101000010",
  63365=>"000100110",
  63366=>"011000001",
  63367=>"000011011",
  63368=>"010110010",
  63369=>"110011010",
  63370=>"000000010",
  63371=>"110100010",
  63372=>"011010100",
  63373=>"100110101",
  63374=>"000001001",
  63375=>"100010000",
  63376=>"010111100",
  63377=>"000101111",
  63378=>"000000111",
  63379=>"010001000",
  63380=>"100101001",
  63381=>"100110101",
  63382=>"010110001",
  63383=>"101001110",
  63384=>"001111000",
  63385=>"000100100",
  63386=>"011101001",
  63387=>"001101011",
  63388=>"111000110",
  63389=>"011011110",
  63390=>"011001011",
  63391=>"101101101",
  63392=>"000001111",
  63393=>"000100010",
  63394=>"000100001",
  63395=>"100000000",
  63396=>"110000101",
  63397=>"101001101",
  63398=>"001101110",
  63399=>"011101101",
  63400=>"001010101",
  63401=>"110011000",
  63402=>"100100111",
  63403=>"110010110",
  63404=>"010000001",
  63405=>"100100000",
  63406=>"100111110",
  63407=>"110100000",
  63408=>"101100100",
  63409=>"100110000",
  63410=>"101011111",
  63411=>"001010100",
  63412=>"110000110",
  63413=>"011000101",
  63414=>"101011111",
  63415=>"101011010",
  63416=>"101000100",
  63417=>"100110101",
  63418=>"111010011",
  63419=>"101001100",
  63420=>"000110111",
  63421=>"101101000",
  63422=>"010011111",
  63423=>"011011111",
  63424=>"001010000",
  63425=>"000111010",
  63426=>"100011010",
  63427=>"000001101",
  63428=>"100100010",
  63429=>"000101110",
  63430=>"111101101",
  63431=>"011000001",
  63432=>"110010000",
  63433=>"100111111",
  63434=>"011101110",
  63435=>"010110010",
  63436=>"111000001",
  63437=>"110110000",
  63438=>"001000100",
  63439=>"001010111",
  63440=>"101111011",
  63441=>"000000110",
  63442=>"001011111",
  63443=>"011000000",
  63444=>"100010101",
  63445=>"110011000",
  63446=>"001101110",
  63447=>"011110100",
  63448=>"010111001",
  63449=>"100000000",
  63450=>"000000001",
  63451=>"100100100",
  63452=>"110100111",
  63453=>"000010001",
  63454=>"000010001",
  63455=>"110111001",
  63456=>"011100001",
  63457=>"100110110",
  63458=>"101110100",
  63459=>"000001100",
  63460=>"001000010",
  63461=>"110100000",
  63462=>"110101100",
  63463=>"100000100",
  63464=>"000001011",
  63465=>"101001001",
  63466=>"000010110",
  63467=>"111010000",
  63468=>"100100101",
  63469=>"111001011",
  63470=>"111000011",
  63471=>"010111111",
  63472=>"100000000",
  63473=>"011010101",
  63474=>"100100010",
  63475=>"111100110",
  63476=>"001011010",
  63477=>"111001100",
  63478=>"011001011",
  63479=>"001111101",
  63480=>"010101000",
  63481=>"001000010",
  63482=>"111110011",
  63483=>"000111001",
  63484=>"010011111",
  63485=>"111010110",
  63486=>"101100001",
  63487=>"111110011",
  63488=>"111110011",
  63489=>"001001000",
  63490=>"000100011",
  63491=>"100010001",
  63492=>"011010100",
  63493=>"100110000",
  63494=>"010000110",
  63495=>"101100010",
  63496=>"111111111",
  63497=>"100100101",
  63498=>"111111010",
  63499=>"011101001",
  63500=>"011100000",
  63501=>"000000100",
  63502=>"010000001",
  63503=>"100100101",
  63504=>"110001100",
  63505=>"011000111",
  63506=>"010010001",
  63507=>"000101100",
  63508=>"100100001",
  63509=>"100101101",
  63510=>"110110011",
  63511=>"000000000",
  63512=>"111001010",
  63513=>"010111000",
  63514=>"000011011",
  63515=>"001100111",
  63516=>"101110011",
  63517=>"110001100",
  63518=>"011101100",
  63519=>"010110101",
  63520=>"110011111",
  63521=>"010011011",
  63522=>"001010110",
  63523=>"001100011",
  63524=>"101110111",
  63525=>"101001111",
  63526=>"000111011",
  63527=>"111010111",
  63528=>"000100000",
  63529=>"000100001",
  63530=>"000010111",
  63531=>"110111111",
  63532=>"000101100",
  63533=>"010011101",
  63534=>"011111000",
  63535=>"010000010",
  63536=>"011000100",
  63537=>"100000101",
  63538=>"011001001",
  63539=>"011100001",
  63540=>"110101000",
  63541=>"000100110",
  63542=>"011101101",
  63543=>"110100100",
  63544=>"001101001",
  63545=>"011110011",
  63546=>"100001111",
  63547=>"110000011",
  63548=>"110101111",
  63549=>"111111111",
  63550=>"101101111",
  63551=>"000001100",
  63552=>"111011010",
  63553=>"110101111",
  63554=>"010111100",
  63555=>"111101111",
  63556=>"111111011",
  63557=>"000100010",
  63558=>"011110111",
  63559=>"001011011",
  63560=>"100001101",
  63561=>"111111000",
  63562=>"111100010",
  63563=>"011111000",
  63564=>"110111110",
  63565=>"011110101",
  63566=>"111110100",
  63567=>"101000011",
  63568=>"100010101",
  63569=>"111010010",
  63570=>"101010100",
  63571=>"111100001",
  63572=>"110010011",
  63573=>"110100000",
  63574=>"001000001",
  63575=>"100011011",
  63576=>"000010011",
  63577=>"100011001",
  63578=>"001110000",
  63579=>"101110011",
  63580=>"001001110",
  63581=>"011011011",
  63582=>"110110110",
  63583=>"110100001",
  63584=>"000010101",
  63585=>"101111111",
  63586=>"000011110",
  63587=>"010111000",
  63588=>"000001011",
  63589=>"010101011",
  63590=>"000000111",
  63591=>"100100111",
  63592=>"011110010",
  63593=>"101000010",
  63594=>"010011001",
  63595=>"001101000",
  63596=>"110001000",
  63597=>"010010100",
  63598=>"011111100",
  63599=>"011000100",
  63600=>"111111100",
  63601=>"011110110",
  63602=>"100000101",
  63603=>"010111000",
  63604=>"110000100",
  63605=>"111010011",
  63606=>"111010100",
  63607=>"010110010",
  63608=>"000000001",
  63609=>"111011100",
  63610=>"111011000",
  63611=>"011100010",
  63612=>"101111010",
  63613=>"100011001",
  63614=>"111100101",
  63615=>"100011001",
  63616=>"100001101",
  63617=>"001000111",
  63618=>"011101010",
  63619=>"010001101",
  63620=>"000101001",
  63621=>"001100100",
  63622=>"000011100",
  63623=>"010000010",
  63624=>"111011011",
  63625=>"001110111",
  63626=>"100001100",
  63627=>"010011100",
  63628=>"001001011",
  63629=>"000010011",
  63630=>"100100011",
  63631=>"011011001",
  63632=>"101010100",
  63633=>"111100111",
  63634=>"000101001",
  63635=>"011110111",
  63636=>"110011001",
  63637=>"000100101",
  63638=>"000000001",
  63639=>"001000001",
  63640=>"000100001",
  63641=>"101110101",
  63642=>"001110110",
  63643=>"010011010",
  63644=>"100101010",
  63645=>"000001000",
  63646=>"011011110",
  63647=>"101101111",
  63648=>"111111001",
  63649=>"110101111",
  63650=>"001110000",
  63651=>"111111011",
  63652=>"110111110",
  63653=>"101100111",
  63654=>"110111001",
  63655=>"000010111",
  63656=>"110101001",
  63657=>"011111110",
  63658=>"110010110",
  63659=>"101100010",
  63660=>"100010000",
  63661=>"101110011",
  63662=>"111100110",
  63663=>"011010000",
  63664=>"100100010",
  63665=>"101010011",
  63666=>"000010001",
  63667=>"000110110",
  63668=>"010000010",
  63669=>"111010101",
  63670=>"000011001",
  63671=>"000100110",
  63672=>"010001111",
  63673=>"101110010",
  63674=>"111001110",
  63675=>"101011011",
  63676=>"011011100",
  63677=>"010101011",
  63678=>"010100001",
  63679=>"011010110",
  63680=>"111000111",
  63681=>"001010100",
  63682=>"111000010",
  63683=>"111100011",
  63684=>"101101011",
  63685=>"001100110",
  63686=>"010001100",
  63687=>"110100000",
  63688=>"011110010",
  63689=>"000011110",
  63690=>"000101101",
  63691=>"001101111",
  63692=>"100011001",
  63693=>"011000101",
  63694=>"101100111",
  63695=>"000000100",
  63696=>"100100010",
  63697=>"101111011",
  63698=>"101011111",
  63699=>"010001100",
  63700=>"111000101",
  63701=>"110101000",
  63702=>"000011111",
  63703=>"001001010",
  63704=>"010101000",
  63705=>"101011000",
  63706=>"010101100",
  63707=>"001000101",
  63708=>"011110110",
  63709=>"010110110",
  63710=>"101101111",
  63711=>"001100000",
  63712=>"001110100",
  63713=>"101010111",
  63714=>"100000101",
  63715=>"001010000",
  63716=>"100101100",
  63717=>"110011110",
  63718=>"010111101",
  63719=>"100010110",
  63720=>"001100010",
  63721=>"110111011",
  63722=>"101001101",
  63723=>"110000111",
  63724=>"010100100",
  63725=>"101000110",
  63726=>"110110110",
  63727=>"010111011",
  63728=>"111100100",
  63729=>"101101010",
  63730=>"100111011",
  63731=>"000111111",
  63732=>"100011011",
  63733=>"101010111",
  63734=>"111011101",
  63735=>"101110000",
  63736=>"101101111",
  63737=>"100110100",
  63738=>"001001011",
  63739=>"011011001",
  63740=>"000100010",
  63741=>"101111100",
  63742=>"101011111",
  63743=>"011011111",
  63744=>"011101000",
  63745=>"001111010",
  63746=>"011101010",
  63747=>"011101000",
  63748=>"011001110",
  63749=>"001100001",
  63750=>"011011111",
  63751=>"001011011",
  63752=>"110100101",
  63753=>"111001010",
  63754=>"100100110",
  63755=>"011100101",
  63756=>"001100100",
  63757=>"010101000",
  63758=>"110110101",
  63759=>"100100111",
  63760=>"000110000",
  63761=>"001000111",
  63762=>"010111011",
  63763=>"100111000",
  63764=>"011110101",
  63765=>"110110110",
  63766=>"001010101",
  63767=>"001110111",
  63768=>"011111100",
  63769=>"100100110",
  63770=>"111100111",
  63771=>"100110111",
  63772=>"110010111",
  63773=>"001000010",
  63774=>"000000110",
  63775=>"011000000",
  63776=>"101100110",
  63777=>"001010000",
  63778=>"010000101",
  63779=>"101000000",
  63780=>"000010001",
  63781=>"010110000",
  63782=>"000111111",
  63783=>"110101000",
  63784=>"010000000",
  63785=>"000000100",
  63786=>"010000100",
  63787=>"001110011",
  63788=>"001000111",
  63789=>"001001110",
  63790=>"110111101",
  63791=>"010101110",
  63792=>"001110110",
  63793=>"011100001",
  63794=>"000110000",
  63795=>"000001101",
  63796=>"010001111",
  63797=>"100101001",
  63798=>"000110011",
  63799=>"111011011",
  63800=>"001001000",
  63801=>"010101101",
  63802=>"000100111",
  63803=>"001101110",
  63804=>"101000001",
  63805=>"001000101",
  63806=>"110100000",
  63807=>"010010011",
  63808=>"100010011",
  63809=>"001111101",
  63810=>"111001100",
  63811=>"010010101",
  63812=>"101111100",
  63813=>"001001010",
  63814=>"001111100",
  63815=>"010011110",
  63816=>"000100110",
  63817=>"100101010",
  63818=>"011111011",
  63819=>"110001010",
  63820=>"011101000",
  63821=>"101010001",
  63822=>"001100000",
  63823=>"111000101",
  63824=>"101100101",
  63825=>"110110110",
  63826=>"011111001",
  63827=>"011110010",
  63828=>"100000001",
  63829=>"110000110",
  63830=>"010010010",
  63831=>"000111000",
  63832=>"010010111",
  63833=>"110001101",
  63834=>"100011010",
  63835=>"111001100",
  63836=>"010011011",
  63837=>"000101000",
  63838=>"100000110",
  63839=>"000110111",
  63840=>"101101100",
  63841=>"000111001",
  63842=>"110001101",
  63843=>"101111001",
  63844=>"101101101",
  63845=>"011011100",
  63846=>"100010110",
  63847=>"001100010",
  63848=>"010001011",
  63849=>"111110111",
  63850=>"001101100",
  63851=>"110000110",
  63852=>"010100111",
  63853=>"110101101",
  63854=>"011101101",
  63855=>"110011011",
  63856=>"101100011",
  63857=>"101110100",
  63858=>"001000100",
  63859=>"111011000",
  63860=>"101100011",
  63861=>"101011011",
  63862=>"110001111",
  63863=>"111111100",
  63864=>"000001000",
  63865=>"010101000",
  63866=>"001100011",
  63867=>"111000010",
  63868=>"110010111",
  63869=>"000100011",
  63870=>"100101010",
  63871=>"101001110",
  63872=>"100110100",
  63873=>"001100010",
  63874=>"000011101",
  63875=>"010011000",
  63876=>"111110110",
  63877=>"100010111",
  63878=>"000010101",
  63879=>"010001010",
  63880=>"010100111",
  63881=>"000111011",
  63882=>"001110000",
  63883=>"101000011",
  63884=>"110011100",
  63885=>"110000010",
  63886=>"010110001",
  63887=>"100000111",
  63888=>"101100011",
  63889=>"100110100",
  63890=>"010101111",
  63891=>"110101000",
  63892=>"001011110",
  63893=>"000010100",
  63894=>"000001111",
  63895=>"101110010",
  63896=>"111010110",
  63897=>"100100111",
  63898=>"101011000",
  63899=>"100101000",
  63900=>"111101100",
  63901=>"001011100",
  63902=>"110001011",
  63903=>"111001100",
  63904=>"111111111",
  63905=>"001000000",
  63906=>"010111110",
  63907=>"000110110",
  63908=>"011100100",
  63909=>"111001000",
  63910=>"000111010",
  63911=>"101101001",
  63912=>"110000010",
  63913=>"110010000",
  63914=>"001101100",
  63915=>"000000011",
  63916=>"010110011",
  63917=>"110101000",
  63918=>"000011100",
  63919=>"111101100",
  63920=>"101100011",
  63921=>"000000001",
  63922=>"001101111",
  63923=>"000111111",
  63924=>"111111101",
  63925=>"011001001",
  63926=>"111110101",
  63927=>"110010111",
  63928=>"110110110",
  63929=>"111110000",
  63930=>"101010111",
  63931=>"110100110",
  63932=>"101011101",
  63933=>"001010011",
  63934=>"101110000",
  63935=>"101100101",
  63936=>"100000100",
  63937=>"111110000",
  63938=>"111001001",
  63939=>"010101000",
  63940=>"101101110",
  63941=>"101010111",
  63942=>"111100000",
  63943=>"101111000",
  63944=>"011011111",
  63945=>"011100101",
  63946=>"101001011",
  63947=>"101011110",
  63948=>"110101000",
  63949=>"101101011",
  63950=>"111000011",
  63951=>"101101011",
  63952=>"001100011",
  63953=>"010011000",
  63954=>"100010011",
  63955=>"101101111",
  63956=>"100000111",
  63957=>"110001111",
  63958=>"100100010",
  63959=>"000001110",
  63960=>"110111110",
  63961=>"101000000",
  63962=>"100011110",
  63963=>"001110101",
  63964=>"101100000",
  63965=>"010001100",
  63966=>"000001001",
  63967=>"110100110",
  63968=>"001110010",
  63969=>"001111000",
  63970=>"111000001",
  63971=>"011101100",
  63972=>"010110000",
  63973=>"100101000",
  63974=>"100010101",
  63975=>"101101110",
  63976=>"011000100",
  63977=>"110001110",
  63978=>"101111010",
  63979=>"110011111",
  63980=>"101110001",
  63981=>"110000111",
  63982=>"110101101",
  63983=>"011000000",
  63984=>"110001010",
  63985=>"100101111",
  63986=>"111000011",
  63987=>"010001010",
  63988=>"001000010",
  63989=>"111011011",
  63990=>"000010101",
  63991=>"111110010",
  63992=>"100101110",
  63993=>"010000011",
  63994=>"111000011",
  63995=>"001110111",
  63996=>"000110111",
  63997=>"001100111",
  63998=>"010011010",
  63999=>"100001100",
  64000=>"000001101",
  64001=>"110111001",
  64002=>"100000010",
  64003=>"101101011",
  64004=>"111001001",
  64005=>"111101110",
  64006=>"111000101",
  64007=>"101011011",
  64008=>"111010000",
  64009=>"100010110",
  64010=>"110101000",
  64011=>"110100010",
  64012=>"010110010",
  64013=>"010111101",
  64014=>"010111100",
  64015=>"011001111",
  64016=>"000010011",
  64017=>"000100001",
  64018=>"100101101",
  64019=>"011001001",
  64020=>"110011010",
  64021=>"110110111",
  64022=>"011001101",
  64023=>"110101001",
  64024=>"110100010",
  64025=>"101011001",
  64026=>"111111111",
  64027=>"110101111",
  64028=>"110001111",
  64029=>"011011000",
  64030=>"111101110",
  64031=>"111010111",
  64032=>"000000101",
  64033=>"010111100",
  64034=>"010001000",
  64035=>"001000100",
  64036=>"101110101",
  64037=>"101010101",
  64038=>"010000001",
  64039=>"010110001",
  64040=>"000100000",
  64041=>"111110000",
  64042=>"100110101",
  64043=>"000000000",
  64044=>"001000000",
  64045=>"001111111",
  64046=>"001101110",
  64047=>"000100011",
  64048=>"111010101",
  64049=>"110011011",
  64050=>"100110111",
  64051=>"010011111",
  64052=>"011111000",
  64053=>"100011111",
  64054=>"010011010",
  64055=>"010010111",
  64056=>"100010000",
  64057=>"001110110",
  64058=>"111001001",
  64059=>"001011011",
  64060=>"110111110",
  64061=>"101101101",
  64062=>"110100110",
  64063=>"001111011",
  64064=>"101100000",
  64065=>"000110000",
  64066=>"111111111",
  64067=>"000010100",
  64068=>"111111010",
  64069=>"111101100",
  64070=>"111001110",
  64071=>"100011111",
  64072=>"000111010",
  64073=>"000110000",
  64074=>"001101001",
  64075=>"000111101",
  64076=>"110011101",
  64077=>"100011010",
  64078=>"111111001",
  64079=>"101010100",
  64080=>"000011111",
  64081=>"100000111",
  64082=>"110110000",
  64083=>"010011001",
  64084=>"100101011",
  64085=>"011010001",
  64086=>"000101101",
  64087=>"100001101",
  64088=>"011110011",
  64089=>"001010101",
  64090=>"001000000",
  64091=>"110100010",
  64092=>"100110111",
  64093=>"000011111",
  64094=>"011111110",
  64095=>"001110111",
  64096=>"010101000",
  64097=>"100011011",
  64098=>"111101101",
  64099=>"010100101",
  64100=>"100011000",
  64101=>"000100000",
  64102=>"000100010",
  64103=>"010011100",
  64104=>"000101001",
  64105=>"011011111",
  64106=>"101010101",
  64107=>"000000010",
  64108=>"111110000",
  64109=>"010010111",
  64110=>"111011011",
  64111=>"011110100",
  64112=>"011100100",
  64113=>"100101111",
  64114=>"011001101",
  64115=>"100011100",
  64116=>"011011000",
  64117=>"101000011",
  64118=>"001100100",
  64119=>"101101001",
  64120=>"010010010",
  64121=>"111100111",
  64122=>"010000001",
  64123=>"100011000",
  64124=>"010001000",
  64125=>"110011100",
  64126=>"000111101",
  64127=>"101110001",
  64128=>"010000110",
  64129=>"100101001",
  64130=>"011111000",
  64131=>"100101000",
  64132=>"011000100",
  64133=>"010110001",
  64134=>"010011100",
  64135=>"110010101",
  64136=>"111011110",
  64137=>"110110101",
  64138=>"100010111",
  64139=>"111001010",
  64140=>"110101111",
  64141=>"111101011",
  64142=>"000100111",
  64143=>"100011011",
  64144=>"001110111",
  64145=>"110111111",
  64146=>"111101111",
  64147=>"110011111",
  64148=>"110011000",
  64149=>"010110000",
  64150=>"101011101",
  64151=>"000101100",
  64152=>"101001110",
  64153=>"100011111",
  64154=>"110010000",
  64155=>"101010100",
  64156=>"000110010",
  64157=>"110001110",
  64158=>"110001010",
  64159=>"011111111",
  64160=>"011001011",
  64161=>"000010101",
  64162=>"000100110",
  64163=>"011010100",
  64164=>"010011110",
  64165=>"110101101",
  64166=>"111100110",
  64167=>"000011010",
  64168=>"111010100",
  64169=>"000000100",
  64170=>"010101110",
  64171=>"110010101",
  64172=>"100000010",
  64173=>"011010001",
  64174=>"000000100",
  64175=>"100000101",
  64176=>"000100110",
  64177=>"011111001",
  64178=>"010010101",
  64179=>"001111001",
  64180=>"010110011",
  64181=>"000110000",
  64182=>"101001000",
  64183=>"011001110",
  64184=>"110101110",
  64185=>"101001111",
  64186=>"001101101",
  64187=>"010111001",
  64188=>"111111011",
  64189=>"000110111",
  64190=>"010010111",
  64191=>"100000100",
  64192=>"000100000",
  64193=>"100111110",
  64194=>"101000111",
  64195=>"000111110",
  64196=>"111010011",
  64197=>"010001011",
  64198=>"001110010",
  64199=>"001101110",
  64200=>"100001110",
  64201=>"011100111",
  64202=>"101010001",
  64203=>"110110011",
  64204=>"100010000",
  64205=>"010011000",
  64206=>"001001000",
  64207=>"100101000",
  64208=>"001101010",
  64209=>"110101001",
  64210=>"111010010",
  64211=>"010111111",
  64212=>"111001101",
  64213=>"111110010",
  64214=>"101101111",
  64215=>"010011100",
  64216=>"101110100",
  64217=>"011101110",
  64218=>"011111101",
  64219=>"101000101",
  64220=>"010110111",
  64221=>"000011000",
  64222=>"101001000",
  64223=>"000000110",
  64224=>"100101011",
  64225=>"111010110",
  64226=>"010111100",
  64227=>"000000101",
  64228=>"100010011",
  64229=>"111100110",
  64230=>"000100010",
  64231=>"110111000",
  64232=>"100101001",
  64233=>"111000101",
  64234=>"001000110",
  64235=>"010100100",
  64236=>"100100100",
  64237=>"000100010",
  64238=>"100010001",
  64239=>"101101001",
  64240=>"011000000",
  64241=>"011100100",
  64242=>"001111100",
  64243=>"000111011",
  64244=>"001100001",
  64245=>"010000111",
  64246=>"110111001",
  64247=>"101110110",
  64248=>"100100011",
  64249=>"000001010",
  64250=>"111111001",
  64251=>"100101110",
  64252=>"111000101",
  64253=>"010110101",
  64254=>"010000100",
  64255=>"110110100",
  64256=>"111001100",
  64257=>"011101000",
  64258=>"111000010",
  64259=>"100101000",
  64260=>"000001001",
  64261=>"010000110",
  64262=>"011101111",
  64263=>"111111010",
  64264=>"100100101",
  64265=>"100000110",
  64266=>"111111011",
  64267=>"000000101",
  64268=>"111010110",
  64269=>"111010101",
  64270=>"110010011",
  64271=>"111101010",
  64272=>"010111010",
  64273=>"111100000",
  64274=>"011110001",
  64275=>"011000001",
  64276=>"000100001",
  64277=>"000011001",
  64278=>"110010101",
  64279=>"011101010",
  64280=>"100101100",
  64281=>"011000010",
  64282=>"111010110",
  64283=>"110110011",
  64284=>"010111000",
  64285=>"001100000",
  64286=>"111000000",
  64287=>"100011001",
  64288=>"001110001",
  64289=>"111010111",
  64290=>"100100001",
  64291=>"110001010",
  64292=>"001100011",
  64293=>"100000001",
  64294=>"101111100",
  64295=>"000111001",
  64296=>"100001011",
  64297=>"001111100",
  64298=>"111100101",
  64299=>"111000110",
  64300=>"000110000",
  64301=>"011111101",
  64302=>"101010001",
  64303=>"111111000",
  64304=>"000000101",
  64305=>"010011010",
  64306=>"110101000",
  64307=>"101111000",
  64308=>"101000101",
  64309=>"011000001",
  64310=>"011111000",
  64311=>"111001110",
  64312=>"001000111",
  64313=>"010100111",
  64314=>"111010010",
  64315=>"111010111",
  64316=>"011010110",
  64317=>"110100011",
  64318=>"010010000",
  64319=>"010111001",
  64320=>"101000011",
  64321=>"010001110",
  64322=>"011010000",
  64323=>"010101001",
  64324=>"111001001",
  64325=>"000001000",
  64326=>"111101001",
  64327=>"011100110",
  64328=>"001001010",
  64329=>"001111011",
  64330=>"101101101",
  64331=>"111100101",
  64332=>"111111100",
  64333=>"011010000",
  64334=>"110101000",
  64335=>"110000101",
  64336=>"111100101",
  64337=>"000111110",
  64338=>"100100010",
  64339=>"100000110",
  64340=>"000110100",
  64341=>"101011110",
  64342=>"000011111",
  64343=>"001100101",
  64344=>"000100100",
  64345=>"110011000",
  64346=>"100101010",
  64347=>"111010110",
  64348=>"000100001",
  64349=>"110110001",
  64350=>"010001011",
  64351=>"000111100",
  64352=>"000000011",
  64353=>"110001110",
  64354=>"000000100",
  64355=>"100101001",
  64356=>"001011011",
  64357=>"010110001",
  64358=>"111011101",
  64359=>"000010111",
  64360=>"101000010",
  64361=>"100000001",
  64362=>"011100100",
  64363=>"000010010",
  64364=>"000110101",
  64365=>"101111101",
  64366=>"100111011",
  64367=>"011101111",
  64368=>"011100101",
  64369=>"010011110",
  64370=>"011011100",
  64371=>"000001110",
  64372=>"011111100",
  64373=>"011101100",
  64374=>"000111111",
  64375=>"101110100",
  64376=>"100010000",
  64377=>"111101010",
  64378=>"011100111",
  64379=>"101101000",
  64380=>"001110010",
  64381=>"100001111",
  64382=>"101101001",
  64383=>"010011111",
  64384=>"010010011",
  64385=>"110111010",
  64386=>"001000010",
  64387=>"100010110",
  64388=>"001100000",
  64389=>"001100010",
  64390=>"011010100",
  64391=>"000000001",
  64392=>"100111101",
  64393=>"110011111",
  64394=>"111110100",
  64395=>"101000011",
  64396=>"110001100",
  64397=>"000011001",
  64398=>"011110000",
  64399=>"001000111",
  64400=>"001010101",
  64401=>"110011010",
  64402=>"010000010",
  64403=>"001100111",
  64404=>"111100100",
  64405=>"111001101",
  64406=>"110001000",
  64407=>"110111010",
  64408=>"101001101",
  64409=>"010010000",
  64410=>"110000011",
  64411=>"010111110",
  64412=>"010010001",
  64413=>"101100000",
  64414=>"011001111",
  64415=>"001110110",
  64416=>"100011001",
  64417=>"000111100",
  64418=>"101010001",
  64419=>"000110101",
  64420=>"000011011",
  64421=>"101100000",
  64422=>"001111100",
  64423=>"011101011",
  64424=>"010000111",
  64425=>"001101001",
  64426=>"001101000",
  64427=>"110111111",
  64428=>"111001010",
  64429=>"100000001",
  64430=>"101101110",
  64431=>"111011010",
  64432=>"100101010",
  64433=>"110011001",
  64434=>"001010001",
  64435=>"101111111",
  64436=>"111100011",
  64437=>"100111100",
  64438=>"111101101",
  64439=>"110110010",
  64440=>"001000111",
  64441=>"000011110",
  64442=>"100010101",
  64443=>"110111101",
  64444=>"111110100",
  64445=>"111101011",
  64446=>"000001111",
  64447=>"111110000",
  64448=>"010011100",
  64449=>"110100100",
  64450=>"100011100",
  64451=>"100010000",
  64452=>"101000010",
  64453=>"110100000",
  64454=>"000101001",
  64455=>"100100000",
  64456=>"000100100",
  64457=>"001011101",
  64458=>"111101111",
  64459=>"110001010",
  64460=>"010110000",
  64461=>"111010100",
  64462=>"110101000",
  64463=>"110101001",
  64464=>"111101110",
  64465=>"100001000",
  64466=>"101001000",
  64467=>"001110111",
  64468=>"100100000",
  64469=>"000101000",
  64470=>"000000000",
  64471=>"101110011",
  64472=>"011001010",
  64473=>"000001110",
  64474=>"111101101",
  64475=>"100100110",
  64476=>"100100110",
  64477=>"100111010",
  64478=>"111001100",
  64479=>"010000011",
  64480=>"110100000",
  64481=>"101001111",
  64482=>"110111000",
  64483=>"110000100",
  64484=>"100001010",
  64485=>"100111111",
  64486=>"101111000",
  64487=>"011111010",
  64488=>"011110100",
  64489=>"101001001",
  64490=>"101010101",
  64491=>"011101110",
  64492=>"111110110",
  64493=>"100001000",
  64494=>"011000001",
  64495=>"110011000",
  64496=>"000111001",
  64497=>"101000111",
  64498=>"111111010",
  64499=>"010000110",
  64500=>"010110011",
  64501=>"011101100",
  64502=>"100100010",
  64503=>"100010011",
  64504=>"001001101",
  64505=>"100111011",
  64506=>"010110111",
  64507=>"110111111",
  64508=>"011110111",
  64509=>"010100011",
  64510=>"101100101",
  64511=>"000011001",
  64512=>"011110011",
  64513=>"000011100",
  64514=>"100010111",
  64515=>"010000110",
  64516=>"001100101",
  64517=>"110010101",
  64518=>"111001000",
  64519=>"111100101",
  64520=>"100100101",
  64521=>"001001111",
  64522=>"001110010",
  64523=>"111100100",
  64524=>"111100000",
  64525=>"100010001",
  64526=>"111010011",
  64527=>"001101011",
  64528=>"111011001",
  64529=>"001001001",
  64530=>"110010001",
  64531=>"100001001",
  64532=>"000001010",
  64533=>"010110011",
  64534=>"111010011",
  64535=>"011111001",
  64536=>"011000101",
  64537=>"101100001",
  64538=>"111010010",
  64539=>"111101101",
  64540=>"000001111",
  64541=>"111111010",
  64542=>"100111100",
  64543=>"000011011",
  64544=>"100100011",
  64545=>"101011110",
  64546=>"101110001",
  64547=>"111101111",
  64548=>"101101011",
  64549=>"010001010",
  64550=>"111010101",
  64551=>"010010100",
  64552=>"101001010",
  64553=>"100010101",
  64554=>"011100001",
  64555=>"111011001",
  64556=>"101010001",
  64557=>"011101001",
  64558=>"111101110",
  64559=>"011011111",
  64560=>"001101101",
  64561=>"010011000",
  64562=>"101001100",
  64563=>"100000101",
  64564=>"011000111",
  64565=>"010000010",
  64566=>"110001001",
  64567=>"100011000",
  64568=>"101100111",
  64569=>"100011110",
  64570=>"100101100",
  64571=>"010100000",
  64572=>"100000100",
  64573=>"101110000",
  64574=>"011100110",
  64575=>"000110001",
  64576=>"011000101",
  64577=>"000010100",
  64578=>"000111001",
  64579=>"001010001",
  64580=>"011000011",
  64581=>"000110001",
  64582=>"101010001",
  64583=>"101101001",
  64584=>"010011010",
  64585=>"011010000",
  64586=>"000011011",
  64587=>"101100010",
  64588=>"010000011",
  64589=>"111001101",
  64590=>"011101110",
  64591=>"011101000",
  64592=>"001101110",
  64593=>"101010100",
  64594=>"100110100",
  64595=>"001111110",
  64596=>"101111110",
  64597=>"100001010",
  64598=>"101000111",
  64599=>"100101100",
  64600=>"010011111",
  64601=>"001100000",
  64602=>"100101010",
  64603=>"100110001",
  64604=>"001110101",
  64605=>"101000000",
  64606=>"000011010",
  64607=>"001001000",
  64608=>"011110110",
  64609=>"000000000",
  64610=>"011101000",
  64611=>"100011110",
  64612=>"010010110",
  64613=>"100100110",
  64614=>"110110101",
  64615=>"000100110",
  64616=>"010111111",
  64617=>"101010111",
  64618=>"100000011",
  64619=>"110100000",
  64620=>"101101011",
  64621=>"101010100",
  64622=>"010000100",
  64623=>"001110000",
  64624=>"001010100",
  64625=>"111000111",
  64626=>"100011100",
  64627=>"111010011",
  64628=>"010010111",
  64629=>"010011110",
  64630=>"101000110",
  64631=>"010101000",
  64632=>"101111010",
  64633=>"101100101",
  64634=>"000000000",
  64635=>"010111010",
  64636=>"100010111",
  64637=>"001000110",
  64638=>"101100000",
  64639=>"000000001",
  64640=>"110001111",
  64641=>"101001100",
  64642=>"010010010",
  64643=>"001000001",
  64644=>"101110000",
  64645=>"001000111",
  64646=>"111000100",
  64647=>"010010100",
  64648=>"100001111",
  64649=>"100100100",
  64650=>"101110000",
  64651=>"111011110",
  64652=>"111110100",
  64653=>"111010111",
  64654=>"011011010",
  64655=>"000000011",
  64656=>"110110111",
  64657=>"110101110",
  64658=>"011111001",
  64659=>"011000000",
  64660=>"010001101",
  64661=>"010010111",
  64662=>"110101001",
  64663=>"111101000",
  64664=>"110111001",
  64665=>"011100101",
  64666=>"111101001",
  64667=>"101001011",
  64668=>"111110011",
  64669=>"011100110",
  64670=>"000101101",
  64671=>"000000111",
  64672=>"010100110",
  64673=>"010000100",
  64674=>"010100001",
  64675=>"001100000",
  64676=>"000000000",
  64677=>"000100001",
  64678=>"100000101",
  64679=>"011101001",
  64680=>"000011110",
  64681=>"010011000",
  64682=>"100001111",
  64683=>"110100110",
  64684=>"110110001",
  64685=>"101100100",
  64686=>"100110110",
  64687=>"011100110",
  64688=>"110001001",
  64689=>"101110010",
  64690=>"001110100",
  64691=>"011101101",
  64692=>"110000000",
  64693=>"101110000",
  64694=>"000110111",
  64695=>"011010001",
  64696=>"001101010",
  64697=>"110100001",
  64698=>"011011010",
  64699=>"100011101",
  64700=>"111111111",
  64701=>"110001100",
  64702=>"011101000",
  64703=>"111101010",
  64704=>"101101101",
  64705=>"100011100",
  64706=>"001100110",
  64707=>"000011011",
  64708=>"100010100",
  64709=>"110101010",
  64710=>"001100010",
  64711=>"011100110",
  64712=>"000011100",
  64713=>"101100101",
  64714=>"111110000",
  64715=>"111110001",
  64716=>"011010001",
  64717=>"111011110",
  64718=>"101001010",
  64719=>"001100110",
  64720=>"110000010",
  64721=>"101010000",
  64722=>"100100011",
  64723=>"110000000",
  64724=>"111001101",
  64725=>"011101100",
  64726=>"000001001",
  64727=>"011100001",
  64728=>"000011101",
  64729=>"101100111",
  64730=>"111001001",
  64731=>"010010001",
  64732=>"011111110",
  64733=>"011101100",
  64734=>"100111001",
  64735=>"001011001",
  64736=>"100000010",
  64737=>"000001101",
  64738=>"111110111",
  64739=>"010010100",
  64740=>"111011111",
  64741=>"010000100",
  64742=>"110000000",
  64743=>"111010111",
  64744=>"001110111",
  64745=>"000001111",
  64746=>"100010110",
  64747=>"111100010",
  64748=>"100101111",
  64749=>"110111110",
  64750=>"000001011",
  64751=>"001100111",
  64752=>"010001111",
  64753=>"010111000",
  64754=>"000110100",
  64755=>"100001110",
  64756=>"100011111",
  64757=>"001000101",
  64758=>"010010101",
  64759=>"100110101",
  64760=>"110111101",
  64761=>"100100111",
  64762=>"000000010",
  64763=>"010111001",
  64764=>"100100010",
  64765=>"010001001",
  64766=>"111111010",
  64767=>"111111111",
  64768=>"111000000",
  64769=>"111101000",
  64770=>"101001111",
  64771=>"100100111",
  64772=>"111010001",
  64773=>"111100010",
  64774=>"001000001",
  64775=>"111111101",
  64776=>"101011001",
  64777=>"011110001",
  64778=>"110110111",
  64779=>"110000001",
  64780=>"101110110",
  64781=>"110001001",
  64782=>"000000001",
  64783=>"010010010",
  64784=>"011001110",
  64785=>"100001101",
  64786=>"100100100",
  64787=>"001111100",
  64788=>"001010101",
  64789=>"011010110",
  64790=>"000011100",
  64791=>"011111101",
  64792=>"111101000",
  64793=>"100101000",
  64794=>"000110010",
  64795=>"000100000",
  64796=>"011101111",
  64797=>"000000100",
  64798=>"111110001",
  64799=>"011110010",
  64800=>"100001100",
  64801=>"110101000",
  64802=>"100010101",
  64803=>"100011001",
  64804=>"110111001",
  64805=>"101110011",
  64806=>"010001011",
  64807=>"000000011",
  64808=>"100110100",
  64809=>"100001011",
  64810=>"100111011",
  64811=>"011011010",
  64812=>"100001010",
  64813=>"010111110",
  64814=>"001001101",
  64815=>"011111010",
  64816=>"000000100",
  64817=>"001110010",
  64818=>"001011100",
  64819=>"001100010",
  64820=>"010010101",
  64821=>"011100001",
  64822=>"001010010",
  64823=>"110101101",
  64824=>"000011101",
  64825=>"110110010",
  64826=>"101111001",
  64827=>"100010111",
  64828=>"000001100",
  64829=>"010001000",
  64830=>"101100111",
  64831=>"000001010",
  64832=>"001100011",
  64833=>"110000000",
  64834=>"000100111",
  64835=>"100001000",
  64836=>"001001000",
  64837=>"111011000",
  64838=>"001011000",
  64839=>"100111100",
  64840=>"000000101",
  64841=>"001110010",
  64842=>"100011010",
  64843=>"000001111",
  64844=>"110000010",
  64845=>"110111111",
  64846=>"000110111",
  64847=>"111110100",
  64848=>"011101111",
  64849=>"011100111",
  64850=>"011110001",
  64851=>"000101110",
  64852=>"110010110",
  64853=>"101011100",
  64854=>"011001000",
  64855=>"010001100",
  64856=>"000111100",
  64857=>"000100101",
  64858=>"001010111",
  64859=>"011111011",
  64860=>"100111011",
  64861=>"100001010",
  64862=>"000011111",
  64863=>"100101000",
  64864=>"110100100",
  64865=>"110100000",
  64866=>"100000110",
  64867=>"001000101",
  64868=>"100011011",
  64869=>"110100011",
  64870=>"000000110",
  64871=>"011001000",
  64872=>"011000011",
  64873=>"100000101",
  64874=>"011100000",
  64875=>"001110101",
  64876=>"011101010",
  64877=>"001010100",
  64878=>"111000110",
  64879=>"000101100",
  64880=>"001100010",
  64881=>"100000011",
  64882=>"000111011",
  64883=>"001010001",
  64884=>"100101010",
  64885=>"011100111",
  64886=>"011011001",
  64887=>"011100101",
  64888=>"100111010",
  64889=>"001011111",
  64890=>"100000010",
  64891=>"111001101",
  64892=>"101110110",
  64893=>"110100110",
  64894=>"100011100",
  64895=>"110000000",
  64896=>"011000001",
  64897=>"011111110",
  64898=>"111100111",
  64899=>"011001110",
  64900=>"001010110",
  64901=>"000101010",
  64902=>"111001011",
  64903=>"100011011",
  64904=>"010101101",
  64905=>"111001100",
  64906=>"000001110",
  64907=>"011100010",
  64908=>"110111101",
  64909=>"110111101",
  64910=>"111010111",
  64911=>"100000111",
  64912=>"110111100",
  64913=>"001000110",
  64914=>"101001101",
  64915=>"011111100",
  64916=>"100100010",
  64917=>"001000010",
  64918=>"010110101",
  64919=>"010100010",
  64920=>"000110010",
  64921=>"000111010",
  64922=>"011000111",
  64923=>"110001010",
  64924=>"101001001",
  64925=>"100010000",
  64926=>"111001111",
  64927=>"100110110",
  64928=>"010011010",
  64929=>"110101100",
  64930=>"100010100",
  64931=>"011001001",
  64932=>"110101110",
  64933=>"101111110",
  64934=>"011011001",
  64935=>"101000010",
  64936=>"010101001",
  64937=>"001110010",
  64938=>"110010101",
  64939=>"011000010",
  64940=>"001010111",
  64941=>"101111000",
  64942=>"000001111",
  64943=>"001011001",
  64944=>"010100000",
  64945=>"110001000",
  64946=>"101110000",
  64947=>"000001001",
  64948=>"111000100",
  64949=>"111111000",
  64950=>"110000001",
  64951=>"011100101",
  64952=>"001000000",
  64953=>"111010111",
  64954=>"001111000",
  64955=>"101001000",
  64956=>"111110011",
  64957=>"110010101",
  64958=>"110100010",
  64959=>"111101000",
  64960=>"010001010",
  64961=>"101000111",
  64962=>"101010011",
  64963=>"101010011",
  64964=>"000010100",
  64965=>"010010110",
  64966=>"000010011",
  64967=>"000000110",
  64968=>"100000000",
  64969=>"100100110",
  64970=>"000100011",
  64971=>"100011111",
  64972=>"000011110",
  64973=>"110010000",
  64974=>"110110110",
  64975=>"101100010",
  64976=>"101100101",
  64977=>"110000011",
  64978=>"000000000",
  64979=>"100111010",
  64980=>"101100111",
  64981=>"110000000",
  64982=>"110000110",
  64983=>"101100010",
  64984=>"111011100",
  64985=>"111010100",
  64986=>"010000000",
  64987=>"000101100",
  64988=>"101000111",
  64989=>"100100010",
  64990=>"101010010",
  64991=>"001101110",
  64992=>"101111010",
  64993=>"010111010",
  64994=>"001110000",
  64995=>"001000000",
  64996=>"001101110",
  64997=>"000010001",
  64998=>"001111111",
  64999=>"101001010",
  65000=>"110010101",
  65001=>"011000111",
  65002=>"011111110",
  65003=>"110111101",
  65004=>"000101101",
  65005=>"011001100",
  65006=>"111111111",
  65007=>"101001100",
  65008=>"010000111",
  65009=>"011010001",
  65010=>"000111101",
  65011=>"000010111",
  65012=>"011110001",
  65013=>"100010100",
  65014=>"001110001",
  65015=>"011000110",
  65016=>"011000011",
  65017=>"011101000",
  65018=>"000010010",
  65019=>"111111010",
  65020=>"101110101",
  65021=>"101110000",
  65022=>"101111110",
  65023=>"100110100",
  65024=>"000111010",
  65025=>"101101111",
  65026=>"011011001",
  65027=>"000000010",
  65028=>"010111011",
  65029=>"101100010",
  65030=>"001001010",
  65031=>"000110000",
  65032=>"100000101",
  65033=>"001110011",
  65034=>"000011000",
  65035=>"101001010",
  65036=>"100101011",
  65037=>"011001010",
  65038=>"011010100",
  65039=>"000101011",
  65040=>"000110111",
  65041=>"011111001",
  65042=>"111010010",
  65043=>"100110101",
  65044=>"011101010",
  65045=>"001001100",
  65046=>"111000011",
  65047=>"110111010",
  65048=>"100011011",
  65049=>"101100101",
  65050=>"100000011",
  65051=>"011011011",
  65052=>"110000011",
  65053=>"101000010",
  65054=>"011101000",
  65055=>"010110001",
  65056=>"111111011",
  65057=>"000100110",
  65058=>"011100101",
  65059=>"000011101",
  65060=>"100011101",
  65061=>"000000001",
  65062=>"101101111",
  65063=>"101000001",
  65064=>"100101011",
  65065=>"111010100",
  65066=>"110101111",
  65067=>"110111001",
  65068=>"101010001",
  65069=>"011111101",
  65070=>"010010100",
  65071=>"000111000",
  65072=>"100010010",
  65073=>"111101000",
  65074=>"011011111",
  65075=>"111000110",
  65076=>"011001001",
  65077=>"000111101",
  65078=>"101010111",
  65079=>"101001010",
  65080=>"111111101",
  65081=>"101110011",
  65082=>"110111010",
  65083=>"010000101",
  65084=>"111011001",
  65085=>"110001010",
  65086=>"001100101",
  65087=>"010001010",
  65088=>"001110010",
  65089=>"110000010",
  65090=>"111000101",
  65091=>"001001100",
  65092=>"001101101",
  65093=>"001010001",
  65094=>"011000101",
  65095=>"101111111",
  65096=>"000000110",
  65097=>"011101101",
  65098=>"100011010",
  65099=>"100101100",
  65100=>"001111111",
  65101=>"000000010",
  65102=>"011011100",
  65103=>"111101110",
  65104=>"000011001",
  65105=>"111010001",
  65106=>"010011100",
  65107=>"011100101",
  65108=>"110010110",
  65109=>"000000001",
  65110=>"010000000",
  65111=>"101010101",
  65112=>"111001010",
  65113=>"110100001",
  65114=>"110111000",
  65115=>"010010000",
  65116=>"110101001",
  65117=>"010000000",
  65118=>"100100000",
  65119=>"010101111",
  65120=>"100100011",
  65121=>"011000101",
  65122=>"010001010",
  65123=>"011101000",
  65124=>"000111101",
  65125=>"000001011",
  65126=>"001001001",
  65127=>"000100100",
  65128=>"010011001",
  65129=>"100100011",
  65130=>"011111100",
  65131=>"000011111",
  65132=>"001010111",
  65133=>"011100010",
  65134=>"011011000",
  65135=>"010100100",
  65136=>"011100011",
  65137=>"001000010",
  65138=>"110000000",
  65139=>"001001111",
  65140=>"000101011",
  65141=>"100111011",
  65142=>"001101010",
  65143=>"111000111",
  65144=>"000001100",
  65145=>"000000011",
  65146=>"101111101",
  65147=>"110001010",
  65148=>"100100001",
  65149=>"001101100",
  65150=>"100000111",
  65151=>"110101001",
  65152=>"000100001",
  65153=>"111011101",
  65154=>"001100100",
  65155=>"000000001",
  65156=>"111011000",
  65157=>"110111001",
  65158=>"101111000",
  65159=>"111100111",
  65160=>"001101010",
  65161=>"100110110",
  65162=>"011111010",
  65163=>"010010000",
  65164=>"000000110",
  65165=>"001001011",
  65166=>"110001001",
  65167=>"010110101",
  65168=>"000111101",
  65169=>"011111011",
  65170=>"010100101",
  65171=>"010101011",
  65172=>"100101111",
  65173=>"001001010",
  65174=>"110000101",
  65175=>"010000000",
  65176=>"110110011",
  65177=>"101010001",
  65178=>"111100001",
  65179=>"001001110",
  65180=>"000100000",
  65181=>"111111010",
  65182=>"001111110",
  65183=>"011010010",
  65184=>"000001111",
  65185=>"011101001",
  65186=>"010001001",
  65187=>"101101011",
  65188=>"001110001",
  65189=>"000111011",
  65190=>"000100001",
  65191=>"011011100",
  65192=>"111000001",
  65193=>"000000001",
  65194=>"010110000",
  65195=>"100010110",
  65196=>"000101010",
  65197=>"110000110",
  65198=>"000010111",
  65199=>"111011110",
  65200=>"011000110",
  65201=>"100111011",
  65202=>"111100010",
  65203=>"000011010",
  65204=>"011010111",
  65205=>"011000111",
  65206=>"000100110",
  65207=>"110001110",
  65208=>"111100010",
  65209=>"100010111",
  65210=>"000000011",
  65211=>"100101000",
  65212=>"101000010",
  65213=>"001000101",
  65214=>"000101100",
  65215=>"110111111",
  65216=>"010100110",
  65217=>"111110000",
  65218=>"000000111",
  65219=>"010000011",
  65220=>"000101101",
  65221=>"100100000",
  65222=>"110000001",
  65223=>"010101101",
  65224=>"110000000",
  65225=>"101111011",
  65226=>"110101010",
  65227=>"110101110",
  65228=>"110000100",
  65229=>"111101101",
  65230=>"101100111",
  65231=>"110100110",
  65232=>"011100011",
  65233=>"111101001",
  65234=>"101010101",
  65235=>"101010000",
  65236=>"000000101",
  65237=>"111100101",
  65238=>"110111011",
  65239=>"111000111",
  65240=>"101101110",
  65241=>"100001101",
  65242=>"010111000",
  65243=>"111011001",
  65244=>"101100010",
  65245=>"011111001",
  65246=>"101111110",
  65247=>"010010001",
  65248=>"001010100",
  65249=>"111001001",
  65250=>"011000111",
  65251=>"100100011",
  65252=>"110111110",
  65253=>"101000110",
  65254=>"101100011",
  65255=>"001001000",
  65256=>"110011111",
  65257=>"001101001",
  65258=>"001010010",
  65259=>"110010001",
  65260=>"100101010",
  65261=>"000011101",
  65262=>"111011010",
  65263=>"011111000",
  65264=>"111010011",
  65265=>"010101010",
  65266=>"111001100",
  65267=>"101100101",
  65268=>"110100011",
  65269=>"100000000",
  65270=>"000001110",
  65271=>"110110000",
  65272=>"011111011",
  65273=>"100101001",
  65274=>"001011100",
  65275=>"111011110",
  65276=>"000000100",
  65277=>"010001010",
  65278=>"101000100",
  65279=>"100010010",
  65280=>"010011101",
  65281=>"010010011",
  65282=>"101000001",
  65283=>"001110110",
  65284=>"100110001",
  65285=>"101001000",
  65286=>"010111010",
  65287=>"001000111",
  65288=>"111100110",
  65289=>"111010001",
  65290=>"011000010",
  65291=>"010000011",
  65292=>"011110100",
  65293=>"111111000",
  65294=>"001100101",
  65295=>"111001011",
  65296=>"111100101",
  65297=>"000010000",
  65298=>"100011011",
  65299=>"011110111",
  65300=>"101110101",
  65301=>"000100110",
  65302=>"111101010",
  65303=>"100000010",
  65304=>"000001000",
  65305=>"100101100",
  65306=>"001000110",
  65307=>"110110001",
  65308=>"110010011",
  65309=>"010001011",
  65310=>"010111111",
  65311=>"011111010",
  65312=>"011010001",
  65313=>"100010101",
  65314=>"111010011",
  65315=>"010001001",
  65316=>"010100011",
  65317=>"001100110",
  65318=>"101101111",
  65319=>"111101111",
  65320=>"001100001",
  65321=>"110010101",
  65322=>"000101101",
  65323=>"101001011",
  65324=>"101001100",
  65325=>"001101100",
  65326=>"100010100",
  65327=>"100011001",
  65328=>"111100010",
  65329=>"011000010",
  65330=>"110001011",
  65331=>"100111110",
  65332=>"100001001",
  65333=>"011110011",
  65334=>"101100110",
  65335=>"100100100",
  65336=>"101111010",
  65337=>"010010010",
  65338=>"000101101",
  65339=>"000001011",
  65340=>"010001100",
  65341=>"011100111",
  65342=>"111010000",
  65343=>"110010000",
  65344=>"001000010",
  65345=>"010000100",
  65346=>"010010100",
  65347=>"111011101",
  65348=>"100010010",
  65349=>"011011101",
  65350=>"011000100",
  65351=>"000000100",
  65352=>"000111101",
  65353=>"001100011",
  65354=>"110100001",
  65355=>"111010001",
  65356=>"010100111",
  65357=>"100111111",
  65358=>"010111010",
  65359=>"011011011",
  65360=>"101001011",
  65361=>"010100111",
  65362=>"101010000",
  65363=>"000010101",
  65364=>"000000001",
  65365=>"101100111",
  65366=>"011110110",
  65367=>"010101110",
  65368=>"000101001",
  65369=>"010011001",
  65370=>"001000101",
  65371=>"010010110",
  65372=>"010100101",
  65373=>"100010001",
  65374=>"010001111",
  65375=>"110110111",
  65376=>"011001010",
  65377=>"111111111",
  65378=>"100001111",
  65379=>"111010011",
  65380=>"100100111",
  65381=>"010101100",
  65382=>"101110111",
  65383=>"100011011",
  65384=>"101001100",
  65385=>"101001100",
  65386=>"110000011",
  65387=>"000111100",
  65388=>"101000100",
  65389=>"001110111",
  65390=>"000100001",
  65391=>"010010101",
  65392=>"001111011",
  65393=>"010010011",
  65394=>"101100110",
  65395=>"011110000",
  65396=>"001110010",
  65397=>"000000111",
  65398=>"010111010",
  65399=>"100111010",
  65400=>"111001001",
  65401=>"101010111",
  65402=>"010101010",
  65403=>"100001110",
  65404=>"010010001",
  65405=>"110110001",
  65406=>"101001000",
  65407=>"111001110",
  65408=>"111000111",
  65409=>"010011011",
  65410=>"110011010",
  65411=>"100000110",
  65412=>"110110101",
  65413=>"101001101",
  65414=>"101100000",
  65415=>"001010001",
  65416=>"100000010",
  65417=>"101010000",
  65418=>"001101101",
  65419=>"010001011",
  65420=>"000111110",
  65421=>"111010101",
  65422=>"000011010",
  65423=>"001111010",
  65424=>"100001000",
  65425=>"100111110",
  65426=>"100001101",
  65427=>"100001010",
  65428=>"111101010",
  65429=>"011000100",
  65430=>"010011111",
  65431=>"000110011",
  65432=>"100000110",
  65433=>"000000100",
  65434=>"000000110",
  65435=>"100010101",
  65436=>"101000100",
  65437=>"000101100",
  65438=>"011011111",
  65439=>"011001100",
  65440=>"000000111",
  65441=>"110100011",
  65442=>"001000011",
  65443=>"010000111",
  65444=>"010000000",
  65445=>"110101010",
  65446=>"011010001",
  65447=>"011100001",
  65448=>"110011000",
  65449=>"101110110",
  65450=>"110101100",
  65451=>"110000111",
  65452=>"011000001",
  65453=>"010110111",
  65454=>"101110101",
  65455=>"000111100",
  65456=>"100001111",
  65457=>"010100110",
  65458=>"111001110",
  65459=>"001001110",
  65460=>"101000001",
  65461=>"111111101",
  65462=>"111001111",
  65463=>"000011011",
  65464=>"101001001",
  65465=>"111101010",
  65466=>"001010101",
  65467=>"101110100",
  65468=>"110010011",
  65469=>"010001100",
  65470=>"110101001",
  65471=>"100101001",
  65472=>"010000100",
  65473=>"101001111",
  65474=>"000000000",
  65475=>"001111101",
  65476=>"010000100",
  65477=>"010101000",
  65478=>"110111100",
  65479=>"100110111",
  65480=>"000100001",
  65481=>"001010011",
  65482=>"110101000",
  65483=>"111000111",
  65484=>"111000001",
  65485=>"101000100",
  65486=>"000100110",
  65487=>"110100010",
  65488=>"110101011",
  65489=>"100111001",
  65490=>"010111100",
  65491=>"111001010",
  65492=>"000001111",
  65493=>"100111001",
  65494=>"100001000",
  65495=>"111001111",
  65496=>"001000011",
  65497=>"011101111",
  65498=>"110111110",
  65499=>"001001011",
  65500=>"011010111",
  65501=>"111100000",
  65502=>"110011110",
  65503=>"101010000",
  65504=>"100111010",
  65505=>"110010011",
  65506=>"011000011",
  65507=>"000110100",
  65508=>"001101000",
  65509=>"110111000",
  65510=>"001010010",
  65511=>"010001000",
  65512=>"101000010",
  65513=>"011000001",
  65514=>"011010100",
  65515=>"100100000",
  65516=>"110001100",
  65517=>"100110001",
  65518=>"000110011",
  65519=>"000111110",
  65520=>"110110000",
  65521=>"000011011",
  65522=>"110000000",
  65523=>"111111011",
  65524=>"011000111",
  65525=>"011110101",
  65526=>"011000010",
  65527=>"111111110",
  65528=>"101101001",
  65529=>"101010110",
  65530=>"001110000",
  65531=>"010011000",
  65532=>"010001111",
  65533=>"111011110",
  65534=>"001101110",
  65535=>"011100001");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;