LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_14_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(8)-1 DOWNTO 0));
END L8_14_WROM;

ARCHITECTURE RTL OF L8_14_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"101100111",
  1=>"110111110",
  2=>"101001101",
  3=>"101001000",
  4=>"010101100",
  5=>"011100011",
  6=>"001100011",
  7=>"001000010",
  8=>"111010101",
  9=>"110111100",
  10=>"100000011",
  11=>"000001101",
  12=>"110111000",
  13=>"110010011",
  14=>"111101001",
  15=>"100101111",
  16=>"010010011",
  17=>"101111110",
  18=>"000000001",
  19=>"000001111",
  20=>"100111011",
  21=>"111100010",
  22=>"111100101",
  23=>"110011100",
  24=>"101001000",
  25=>"111111001",
  26=>"010010101",
  27=>"001100101",
  28=>"111100011",
  29=>"001111011",
  30=>"111110010",
  31=>"001000001",
  32=>"011111110",
  33=>"100011011",
  34=>"000110100",
  35=>"010010111",
  36=>"111111010",
  37=>"100100100",
  38=>"000110110",
  39=>"111101001",
  40=>"101101110",
  41=>"000110001",
  42=>"001100110",
  43=>"010001001",
  44=>"010011101",
  45=>"010011101",
  46=>"110100011",
  47=>"111000100",
  48=>"101111111",
  49=>"111001100",
  50=>"011101001",
  51=>"110010000",
  52=>"101111110",
  53=>"011110010",
  54=>"000100001",
  55=>"001001011",
  56=>"001000110",
  57=>"000000100",
  58=>"001010111",
  59=>"000100101",
  60=>"011110111",
  61=>"101000111",
  62=>"010101101",
  63=>"111111100",
  64=>"111000111",
  65=>"100101101",
  66=>"100001001",
  67=>"111000010",
  68=>"110011010",
  69=>"101101110",
  70=>"010110110",
  71=>"010001110",
  72=>"111110000",
  73=>"000011111",
  74=>"100010011",
  75=>"111101010",
  76=>"101000011",
  77=>"011100110",
  78=>"111100110",
  79=>"001110000",
  80=>"000001111",
  81=>"111111111",
  82=>"110110100",
  83=>"110001001",
  84=>"001110001",
  85=>"111011000",
  86=>"101100111",
  87=>"000000000",
  88=>"010100111",
  89=>"010111101",
  90=>"000100110",
  91=>"001000101",
  92=>"011100000",
  93=>"101101000",
  94=>"000110111",
  95=>"111011010",
  96=>"101001110",
  97=>"110110011",
  98=>"001010100",
  99=>"000000100",
  100=>"000011110",
  101=>"011101101",
  102=>"010101100",
  103=>"111011010",
  104=>"101000001",
  105=>"110101101",
  106=>"001011110",
  107=>"100101010",
  108=>"111111111",
  109=>"000100110",
  110=>"010100110",
  111=>"100111000",
  112=>"011001010",
  113=>"101111111",
  114=>"011101010",
  115=>"011101001",
  116=>"000001001",
  117=>"010101111",
  118=>"001100001",
  119=>"101110001",
  120=>"001101001",
  121=>"010011000",
  122=>"111001001",
  123=>"100100100",
  124=>"001001100",
  125=>"011100001",
  126=>"011001000",
  127=>"110111101",
  128=>"010000010",
  129=>"101001000",
  130=>"010001001",
  131=>"101111000",
  132=>"000110100",
  133=>"001101111",
  134=>"101100111",
  135=>"001000000",
  136=>"000110101",
  137=>"100110000",
  138=>"110110000",
  139=>"111101100",
  140=>"010110000",
  141=>"001110010",
  142=>"000011111",
  143=>"111110100",
  144=>"011001001",
  145=>"001011101",
  146=>"000011000",
  147=>"000111100",
  148=>"100111101",
  149=>"010101101",
  150=>"000011010",
  151=>"111100000",
  152=>"100011100",
  153=>"000101100",
  154=>"000001000",
  155=>"100101100",
  156=>"111101001",
  157=>"100111100",
  158=>"010001110",
  159=>"010000000",
  160=>"111110111",
  161=>"011110001",
  162=>"110000001",
  163=>"010011111",
  164=>"100001001",
  165=>"101001101",
  166=>"010111001",
  167=>"110010100",
  168=>"011111100",
  169=>"011000111",
  170=>"110011011",
  171=>"011111010",
  172=>"010110110",
  173=>"010100001",
  174=>"101100110",
  175=>"001100011",
  176=>"001000111",
  177=>"111010000",
  178=>"011001011",
  179=>"110101010",
  180=>"000010000",
  181=>"001010001",
  182=>"101101111",
  183=>"000000110",
  184=>"001110110",
  185=>"110110100",
  186=>"011101011",
  187=>"010111110",
  188=>"100011110",
  189=>"110100100",
  190=>"001100001",
  191=>"110110010",
  192=>"011001111",
  193=>"001110110",
  194=>"011111010",
  195=>"111010001",
  196=>"011100101",
  197=>"101101000",
  198=>"000010010",
  199=>"100101110",
  200=>"011011111",
  201=>"001000110",
  202=>"111001011",
  203=>"011011110",
  204=>"100000011",
  205=>"111100110",
  206=>"010110101",
  207=>"000010001",
  208=>"111001010",
  209=>"001011101",
  210=>"011110011",
  211=>"111111110",
  212=>"111011100",
  213=>"110101011",
  214=>"011001011",
  215=>"111111011",
  216=>"110100010",
  217=>"000100010",
  218=>"110100100",
  219=>"011101001",
  220=>"010111010",
  221=>"001100011",
  222=>"110111111",
  223=>"010101000",
  224=>"000110010",
  225=>"111111011",
  226=>"111000100",
  227=>"001110110",
  228=>"101101000",
  229=>"001011101",
  230=>"101100010",
  231=>"101110110",
  232=>"010101000",
  233=>"011111100",
  234=>"011001010",
  235=>"000010010",
  236=>"101110111",
  237=>"100010110",
  238=>"010111101",
  239=>"101100001",
  240=>"111100101",
  241=>"000000001",
  242=>"110110011",
  243=>"000000101",
  244=>"110000101",
  245=>"101101111",
  246=>"010110101",
  247=>"000010010",
  248=>"111010000",
  249=>"001000111",
  250=>"111111011",
  251=>"000111000",
  252=>"101101111",
  253=>"111000001",
  254=>"101001101",
  255=>"100011100",
  256=>"010011111",
  257=>"101111010",
  258=>"010101000",
  259=>"010101000",
  260=>"100110011",
  261=>"100110000",
  262=>"101101001",
  263=>"000000100",
  264=>"010000101",
  265=>"000011010",
  266=>"100101100",
  267=>"010000010",
  268=>"101100001",
  269=>"101001111",
  270=>"010110000",
  271=>"110111110",
  272=>"100101001",
  273=>"111010010",
  274=>"001111111",
  275=>"110000110",
  276=>"100001111",
  277=>"010001010",
  278=>"110100111",
  279=>"011011001",
  280=>"001100001",
  281=>"001000000",
  282=>"010010111",
  283=>"001000001",
  284=>"111101111",
  285=>"100110110",
  286=>"011100101",
  287=>"100101101",
  288=>"000001001",
  289=>"100000000",
  290=>"011110100",
  291=>"101111011",
  292=>"000000000",
  293=>"110110011",
  294=>"010100001",
  295=>"011010001",
  296=>"010100110",
  297=>"001101000",
  298=>"010001001",
  299=>"001001011",
  300=>"010110111",
  301=>"000000101",
  302=>"001000011",
  303=>"111010110",
  304=>"101101101",
  305=>"010011001",
  306=>"000100011",
  307=>"000111000",
  308=>"000110111",
  309=>"011101001",
  310=>"101100010",
  311=>"101001010",
  312=>"110100100",
  313=>"000100010",
  314=>"011010110",
  315=>"100001010",
  316=>"110111011",
  317=>"100110110",
  318=>"110010011",
  319=>"011000111",
  320=>"010101000",
  321=>"010100111",
  322=>"010000100",
  323=>"000001110",
  324=>"011111010",
  325=>"101011111",
  326=>"111000000",
  327=>"010000011",
  328=>"010000000",
  329=>"000100000",
  330=>"111011001",
  331=>"101011111",
  332=>"111001001",
  333=>"000010100",
  334=>"000011101",
  335=>"010010110",
  336=>"100001111",
  337=>"111100001",
  338=>"000100111",
  339=>"101011100",
  340=>"010101000",
  341=>"110111111",
  342=>"101000011",
  343=>"001001100",
  344=>"011000110",
  345=>"010111110",
  346=>"111101110",
  347=>"000001010",
  348=>"100001101",
  349=>"010000000",
  350=>"011001010",
  351=>"011000110",
  352=>"101001100",
  353=>"101110111",
  354=>"000010001",
  355=>"010111001",
  356=>"010111000",
  357=>"110000111",
  358=>"001101101",
  359=>"011000110",
  360=>"001100111",
  361=>"011011110",
  362=>"101010011",
  363=>"000001000",
  364=>"001001101",
  365=>"111101111",
  366=>"111001000",
  367=>"011000001",
  368=>"100001010",
  369=>"001111000",
  370=>"011111001",
  371=>"100101011",
  372=>"111000010",
  373=>"100001111",
  374=>"001000110",
  375=>"000000010",
  376=>"100100010",
  377=>"011100000",
  378=>"101010000",
  379=>"110100011",
  380=>"011011001",
  381=>"000100000",
  382=>"010001000",
  383=>"101000011",
  384=>"100111011",
  385=>"000001001",
  386=>"110111000",
  387=>"101100100",
  388=>"001011100",
  389=>"011010000",
  390=>"110101111",
  391=>"001010000",
  392=>"010001111",
  393=>"010011010",
  394=>"111100110",
  395=>"010000100",
  396=>"000000010",
  397=>"101101101",
  398=>"000101011",
  399=>"110001000",
  400=>"111101100",
  401=>"001000111",
  402=>"010000000",
  403=>"011000110",
  404=>"011101000",
  405=>"001010101",
  406=>"000110011",
  407=>"000111110",
  408=>"010001111",
  409=>"111011110",
  410=>"111011111",
  411=>"110111110",
  412=>"111101111",
  413=>"001010000",
  414=>"011111100",
  415=>"100100100",
  416=>"111110100",
  417=>"000111111",
  418=>"000001100",
  419=>"110011011",
  420=>"001010001",
  421=>"010100000",
  422=>"110110110",
  423=>"111101101",
  424=>"110111010",
  425=>"001000000",
  426=>"000010000",
  427=>"100001110",
  428=>"001100111",
  429=>"111011011",
  430=>"010001111",
  431=>"111011100",
  432=>"011111010",
  433=>"100110100",
  434=>"000011000",
  435=>"011011010",
  436=>"100011111",
  437=>"100010100",
  438=>"110010010",
  439=>"111001111",
  440=>"010101111",
  441=>"001111100",
  442=>"001011000",
  443=>"100010010",
  444=>"111010000",
  445=>"110010010",
  446=>"100101111",
  447=>"111100100",
  448=>"001100101",
  449=>"001101111",
  450=>"101001010",
  451=>"011011100",
  452=>"000001100",
  453=>"101100110",
  454=>"010110001",
  455=>"100001010",
  456=>"000011100",
  457=>"000101001",
  458=>"001010000",
  459=>"010001110",
  460=>"100110111",
  461=>"001111111",
  462=>"011010101",
  463=>"010010101",
  464=>"010110111",
  465=>"111010010",
  466=>"000110000",
  467=>"000100100",
  468=>"000111111",
  469=>"010101001",
  470=>"100101000",
  471=>"001111111",
  472=>"000011100",
  473=>"111110111",
  474=>"110111000",
  475=>"111001000",
  476=>"011100001",
  477=>"010001000",
  478=>"101001111",
  479=>"110011000",
  480=>"111101101",
  481=>"000000011",
  482=>"100101111",
  483=>"010101000",
  484=>"000111100",
  485=>"001100010",
  486=>"101110011",
  487=>"100100000",
  488=>"000000000",
  489=>"000110101",
  490=>"100101101",
  491=>"000000111",
  492=>"011100011",
  493=>"000011111",
  494=>"010000011",
  495=>"000010110",
  496=>"010000110",
  497=>"001111001",
  498=>"111011111",
  499=>"011100011",
  500=>"001111111",
  501=>"011000000",
  502=>"000010101",
  503=>"111100011",
  504=>"000101100",
  505=>"011101011",
  506=>"110000110",
  507=>"101111100",
  508=>"101111001",
  509=>"000001010",
  510=>"101111100",
  511=>"010000101",
  512=>"001110000",
  513=>"100111110",
  514=>"100110101",
  515=>"000000100",
  516=>"001111011",
  517=>"000101110",
  518=>"001111110",
  519=>"010011011",
  520=>"010001001",
  521=>"111010010",
  522=>"010001111",
  523=>"011001101",
  524=>"111100111",
  525=>"000101110",
  526=>"001111000",
  527=>"110111100",
  528=>"011000010",
  529=>"001000111",
  530=>"111101010",
  531=>"111110110",
  532=>"100011001",
  533=>"010101000",
  534=>"001000111",
  535=>"011010011",
  536=>"100101010",
  537=>"001001011",
  538=>"111011000",
  539=>"111111101",
  540=>"111010111",
  541=>"111111001",
  542=>"011100011",
  543=>"011110111",
  544=>"100110000",
  545=>"000000000",
  546=>"000000100",
  547=>"101010010",
  548=>"000001010",
  549=>"011011101",
  550=>"101001011",
  551=>"111101010",
  552=>"011000010",
  553=>"101000010",
  554=>"001110111",
  555=>"010100000",
  556=>"111100111",
  557=>"101110111",
  558=>"111010000",
  559=>"111000111",
  560=>"011011010",
  561=>"010111011",
  562=>"111001000",
  563=>"101011011",
  564=>"110000011",
  565=>"101101110",
  566=>"111111000",
  567=>"000000000",
  568=>"010111111",
  569=>"010000001",
  570=>"110000100",
  571=>"000101010",
  572=>"111101010",
  573=>"011010100",
  574=>"100001010",
  575=>"011011001",
  576=>"101001111",
  577=>"001001100",
  578=>"010100001",
  579=>"010011110",
  580=>"101010000",
  581=>"011111000",
  582=>"111011110",
  583=>"111101111",
  584=>"111110000",
  585=>"110000010",
  586=>"111101000",
  587=>"011111111",
  588=>"010001010",
  589=>"100011100",
  590=>"111100000",
  591=>"010000000",
  592=>"010110111",
  593=>"010100000",
  594=>"100110100",
  595=>"100110100",
  596=>"111101100",
  597=>"011011001",
  598=>"110111100",
  599=>"001001011",
  600=>"011010001",
  601=>"110100101",
  602=>"110011001",
  603=>"001100110",
  604=>"011010001",
  605=>"100001101",
  606=>"111001100",
  607=>"011110100",
  608=>"110001111",
  609=>"001001001",
  610=>"001010001",
  611=>"110010000",
  612=>"100011000",
  613=>"111001010",
  614=>"111011100",
  615=>"011111000",
  616=>"100000110",
  617=>"000010011",
  618=>"100111011",
  619=>"011010111",
  620=>"101011100",
  621=>"110101101",
  622=>"100000011",
  623=>"101100010",
  624=>"001000110",
  625=>"010001000",
  626=>"110000101",
  627=>"100010110",
  628=>"101011110",
  629=>"100111110",
  630=>"110011111",
  631=>"100000010",
  632=>"110101010",
  633=>"100010001",
  634=>"000001000",
  635=>"111001000",
  636=>"010000100",
  637=>"110001000",
  638=>"111011111",
  639=>"110011000",
  640=>"101001110",
  641=>"011110101",
  642=>"011000110",
  643=>"010111111",
  644=>"101111011",
  645=>"101110001",
  646=>"010101111",
  647=>"110100010",
  648=>"111000011",
  649=>"000010010",
  650=>"010101101",
  651=>"111000000",
  652=>"010000001",
  653=>"001110101",
  654=>"011011001",
  655=>"001100000",
  656=>"101010101",
  657=>"000110000",
  658=>"010110110",
  659=>"011100011",
  660=>"110110110",
  661=>"001000001",
  662=>"010111110",
  663=>"111010101",
  664=>"101101000",
  665=>"110001110",
  666=>"100110101",
  667=>"100111011",
  668=>"000011000",
  669=>"001111001",
  670=>"001010111",
  671=>"001110110",
  672=>"100100100",
  673=>"111011001",
  674=>"001011100",
  675=>"100000001",
  676=>"110111110",
  677=>"001100010",
  678=>"010010000",
  679=>"100111111",
  680=>"000101011",
  681=>"001010011",
  682=>"001011100",
  683=>"011101000",
  684=>"110101101",
  685=>"101100011",
  686=>"100010011",
  687=>"001011001",
  688=>"000111010",
  689=>"111110111",
  690=>"010110000",
  691=>"111100011",
  692=>"101010101",
  693=>"111111001",
  694=>"001100101",
  695=>"100101000",
  696=>"101100100",
  697=>"101011000",
  698=>"101001111",
  699=>"000101011",
  700=>"111011000",
  701=>"101110010",
  702=>"010101001",
  703=>"001110100",
  704=>"100010111",
  705=>"010010000",
  706=>"100110111",
  707=>"101110011",
  708=>"111010000",
  709=>"000001000",
  710=>"010000010",
  711=>"011001000",
  712=>"100111011",
  713=>"001010101",
  714=>"010011110",
  715=>"110101101",
  716=>"111000101",
  717=>"001100001",
  718=>"001010001",
  719=>"100110100",
  720=>"010000111",
  721=>"001001111",
  722=>"111110110",
  723=>"101011101",
  724=>"001111010",
  725=>"011111000",
  726=>"100010100",
  727=>"110011100",
  728=>"010111110",
  729=>"010110010",
  730=>"110101101",
  731=>"011100100",
  732=>"110001100",
  733=>"001000110",
  734=>"001111110",
  735=>"100000010",
  736=>"110010001",
  737=>"111000000",
  738=>"101100010",
  739=>"010111101",
  740=>"110000010",
  741=>"000001100",
  742=>"011011010",
  743=>"001011101",
  744=>"100101110",
  745=>"111110100",
  746=>"001110000",
  747=>"001111010",
  748=>"010100001",
  749=>"101110100",
  750=>"110101001",
  751=>"010111111",
  752=>"100110011",
  753=>"100110110",
  754=>"100011001",
  755=>"100100010",
  756=>"001000010",
  757=>"110110110",
  758=>"010010110",
  759=>"010100100",
  760=>"110100101",
  761=>"010000110",
  762=>"001010101",
  763=>"001100011",
  764=>"010001110",
  765=>"101110100",
  766=>"001101001",
  767=>"111101100",
  768=>"101011011",
  769=>"000110001",
  770=>"111110110",
  771=>"111110111",
  772=>"001000010",
  773=>"000010100",
  774=>"010001110",
  775=>"011111111",
  776=>"011000101",
  777=>"100101100",
  778=>"110111110",
  779=>"001101111",
  780=>"010100001",
  781=>"110001000",
  782=>"111010001",
  783=>"010100010",
  784=>"010010011",
  785=>"001000000",
  786=>"001111011",
  787=>"111101001",
  788=>"111011001",
  789=>"000111011",
  790=>"011001101",
  791=>"000000110",
  792=>"101101110",
  793=>"101111111",
  794=>"111000010",
  795=>"111001111",
  796=>"111101000",
  797=>"111000110",
  798=>"111000010",
  799=>"110101011",
  800=>"111111010",
  801=>"101100111",
  802=>"011110111",
  803=>"110000001",
  804=>"011001000",
  805=>"111101001",
  806=>"100010001",
  807=>"001001111",
  808=>"100010101",
  809=>"001001010",
  810=>"111110011",
  811=>"101101101",
  812=>"001101001",
  813=>"001101111",
  814=>"111010101",
  815=>"101100110",
  816=>"011011111",
  817=>"100100001",
  818=>"001001000",
  819=>"000100000",
  820=>"010101000",
  821=>"000110000",
  822=>"011011010",
  823=>"111010110",
  824=>"000000001",
  825=>"011110010",
  826=>"001100000",
  827=>"110000001",
  828=>"101010110",
  829=>"010001111",
  830=>"100010101",
  831=>"101100111",
  832=>"000001001",
  833=>"101001101",
  834=>"111010100",
  835=>"101101100",
  836=>"110110010",
  837=>"011111010",
  838=>"111111000",
  839=>"001110001",
  840=>"111110001",
  841=>"111000001",
  842=>"001001111",
  843=>"101100000",
  844=>"111011110",
  845=>"100100101",
  846=>"001000110",
  847=>"111110001",
  848=>"111111110",
  849=>"100001001",
  850=>"000010101",
  851=>"001101001",
  852=>"110101110",
  853=>"101011111",
  854=>"101100111",
  855=>"100101000",
  856=>"101101010",
  857=>"000101100",
  858=>"001001011",
  859=>"001001000",
  860=>"010011110",
  861=>"110110100",
  862=>"010110000",
  863=>"011110101",
  864=>"001010000",
  865=>"000101001",
  866=>"110111000",
  867=>"001010101",
  868=>"010000011",
  869=>"011101101",
  870=>"110100111",
  871=>"110111110",
  872=>"101111001",
  873=>"110001000",
  874=>"000010001",
  875=>"001011000",
  876=>"100100011",
  877=>"101111101",
  878=>"100000010",
  879=>"010000101",
  880=>"101000001",
  881=>"010100101",
  882=>"101100110",
  883=>"100101101",
  884=>"100111000",
  885=>"000101001",
  886=>"010110100",
  887=>"111001100",
  888=>"001011100",
  889=>"110001001",
  890=>"100001010",
  891=>"100101111",
  892=>"111101100",
  893=>"111011110",
  894=>"001001000",
  895=>"010100100",
  896=>"111100011",
  897=>"100110101",
  898=>"010100001",
  899=>"011001010",
  900=>"001001101",
  901=>"111001100",
  902=>"000001110",
  903=>"111100010",
  904=>"000001100",
  905=>"100011110",
  906=>"000001010",
  907=>"001000111",
  908=>"010100001",
  909=>"010001001",
  910=>"001101010",
  911=>"101011000",
  912=>"111111111",
  913=>"101010001",
  914=>"000111000",
  915=>"100001111",
  916=>"010101110",
  917=>"101101011",
  918=>"001111001",
  919=>"100001100",
  920=>"110010001",
  921=>"000001010",
  922=>"100011101",
  923=>"101011000",
  924=>"100000000",
  925=>"000000010",
  926=>"111101101",
  927=>"001000110",
  928=>"100011100",
  929=>"011000100",
  930=>"000010100",
  931=>"110000001",
  932=>"000011100",
  933=>"111001100",
  934=>"101010010",
  935=>"100110110",
  936=>"010000111",
  937=>"110110010",
  938=>"110001011",
  939=>"101100110",
  940=>"011100110",
  941=>"001010110",
  942=>"000111100",
  943=>"000010110",
  944=>"110110000",
  945=>"111000110",
  946=>"001000001",
  947=>"100000011",
  948=>"110110010",
  949=>"110101011",
  950=>"101011111",
  951=>"100110101",
  952=>"111001001",
  953=>"100011100",
  954=>"110001110",
  955=>"100101100",
  956=>"000111001",
  957=>"101110011",
  958=>"000101101",
  959=>"010010110",
  960=>"001111111",
  961=>"000011100",
  962=>"011000110",
  963=>"001110000",
  964=>"111100010",
  965=>"011100110",
  966=>"100001110",
  967=>"000010011",
  968=>"001000000",
  969=>"101000000",
  970=>"111101000",
  971=>"101111101",
  972=>"101011011",
  973=>"101111011",
  974=>"101110111",
  975=>"111011110",
  976=>"011100010",
  977=>"010110101",
  978=>"110000101",
  979=>"100000100",
  980=>"011110111",
  981=>"101101100",
  982=>"101110011",
  983=>"001111001",
  984=>"010111000",
  985=>"111111111",
  986=>"110100001",
  987=>"000110110",
  988=>"010110110",
  989=>"101001110",
  990=>"101110000",
  991=>"001001100",
  992=>"000011001",
  993=>"010001000",
  994=>"010100101",
  995=>"100001010",
  996=>"001100001",
  997=>"000000101",
  998=>"010000111",
  999=>"001111111",
  1000=>"000001101",
  1001=>"000101010",
  1002=>"011011001",
  1003=>"100100111",
  1004=>"110110110",
  1005=>"011001001",
  1006=>"010010000",
  1007=>"000111101",
  1008=>"111100110",
  1009=>"010100001",
  1010=>"110110101",
  1011=>"101001111",
  1012=>"000000000",
  1013=>"010000011",
  1014=>"010000010",
  1015=>"000000111",
  1016=>"000101011",
  1017=>"011101011",
  1018=>"010010011",
  1019=>"110101101",
  1020=>"111110111",
  1021=>"010101100",
  1022=>"010011100",
  1023=>"001011111",
  1024=>"100000000",
  1025=>"011000001",
  1026=>"000000110",
  1027=>"111001010",
  1028=>"010111111",
  1029=>"110110011",
  1030=>"010100101",
  1031=>"001010110",
  1032=>"011111111",
  1033=>"110001100",
  1034=>"110001010",
  1035=>"111011011",
  1036=>"011111110",
  1037=>"100101000",
  1038=>"110011010",
  1039=>"001000110",
  1040=>"110111111",
  1041=>"110111100",
  1042=>"000010011",
  1043=>"010100110",
  1044=>"001001101",
  1045=>"101100110",
  1046=>"010101110",
  1047=>"010101110",
  1048=>"010101100",
  1049=>"000001010",
  1050=>"011000110",
  1051=>"101001101",
  1052=>"010001000",
  1053=>"110110000",
  1054=>"101110000",
  1055=>"110000110",
  1056=>"001000111",
  1057=>"100110100",
  1058=>"101000010",
  1059=>"010100011",
  1060=>"100101100",
  1061=>"110011100",
  1062=>"010010111",
  1063=>"101110110",
  1064=>"110110000",
  1065=>"010011001",
  1066=>"011011010",
  1067=>"010101011",
  1068=>"001001110",
  1069=>"100110011",
  1070=>"101011000",
  1071=>"111010000",
  1072=>"001110101",
  1073=>"001101110",
  1074=>"011010001",
  1075=>"010111000",
  1076=>"100101000",
  1077=>"111101011",
  1078=>"011001110",
  1079=>"001001010",
  1080=>"011000001",
  1081=>"111110010",
  1082=>"100010111",
  1083=>"111011101",
  1084=>"000110000",
  1085=>"110111010",
  1086=>"011010011",
  1087=>"001011011",
  1088=>"100101100",
  1089=>"010000101",
  1090=>"111000010",
  1091=>"011000011",
  1092=>"010100010",
  1093=>"000010000",
  1094=>"101101101",
  1095=>"111000111",
  1096=>"100000110",
  1097=>"010001110",
  1098=>"011101110",
  1099=>"101101000",
  1100=>"010111000",
  1101=>"110101100",
  1102=>"111111111",
  1103=>"101001010",
  1104=>"011011001",
  1105=>"111101100",
  1106=>"001101100",
  1107=>"111011010",
  1108=>"101110111",
  1109=>"101011011",
  1110=>"000001000",
  1111=>"110010110",
  1112=>"111010010",
  1113=>"101110000",
  1114=>"111011110",
  1115=>"111001110",
  1116=>"111110001",
  1117=>"110110100",
  1118=>"011001010",
  1119=>"100011101",
  1120=>"100110010",
  1121=>"110111101",
  1122=>"000001000",
  1123=>"000000100",
  1124=>"101000011",
  1125=>"000100110",
  1126=>"101010011",
  1127=>"111100100",
  1128=>"110110100",
  1129=>"001110100",
  1130=>"001101111",
  1131=>"111100011",
  1132=>"000011011",
  1133=>"101010000",
  1134=>"110000101",
  1135=>"000001010",
  1136=>"100011100",
  1137=>"001110001",
  1138=>"000001011",
  1139=>"101010011",
  1140=>"101010110",
  1141=>"001010111",
  1142=>"010000111",
  1143=>"110011011",
  1144=>"001110000",
  1145=>"111001000",
  1146=>"001010100",
  1147=>"100111011",
  1148=>"100110000",
  1149=>"010001010",
  1150=>"011010000",
  1151=>"111001001",
  1152=>"011110001",
  1153=>"011010011",
  1154=>"000001011",
  1155=>"011101001",
  1156=>"111000101",
  1157=>"001110001",
  1158=>"100110000",
  1159=>"011010000",
  1160=>"010011011",
  1161=>"010011101",
  1162=>"110011001",
  1163=>"101111001",
  1164=>"001101000",
  1165=>"110111101",
  1166=>"111001011",
  1167=>"111010010",
  1168=>"000110110",
  1169=>"101110010",
  1170=>"011111101",
  1171=>"101011101",
  1172=>"100000001",
  1173=>"111111110",
  1174=>"100010100",
  1175=>"110010110",
  1176=>"100011011",
  1177=>"100110110",
  1178=>"010010011",
  1179=>"001000010",
  1180=>"011110101",
  1181=>"001001110",
  1182=>"110111010",
  1183=>"011011111",
  1184=>"000000111",
  1185=>"100111011",
  1186=>"111100111",
  1187=>"000100001",
  1188=>"111111111",
  1189=>"000000001",
  1190=>"000011010",
  1191=>"110110000",
  1192=>"000111000",
  1193=>"101011111",
  1194=>"001100110",
  1195=>"001111110",
  1196=>"010110010",
  1197=>"001011110",
  1198=>"100010100",
  1199=>"111101100",
  1200=>"010000000",
  1201=>"011010001",
  1202=>"110100111",
  1203=>"111000011",
  1204=>"110100101",
  1205=>"000001010",
  1206=>"111101101",
  1207=>"100110110",
  1208=>"111111110",
  1209=>"000111101",
  1210=>"010001101",
  1211=>"110010101",
  1212=>"101101111",
  1213=>"001011110",
  1214=>"111000111",
  1215=>"101100010",
  1216=>"010100100",
  1217=>"000011110",
  1218=>"111010100",
  1219=>"110111111",
  1220=>"000011100",
  1221=>"010010011",
  1222=>"000001011",
  1223=>"100111011",
  1224=>"101010010",
  1225=>"101000100",
  1226=>"010011100",
  1227=>"101000000",
  1228=>"110100010",
  1229=>"101010001",
  1230=>"010011011",
  1231=>"100111100",
  1232=>"110111010",
  1233=>"100100000",
  1234=>"100100110",
  1235=>"001111110",
  1236=>"001110110",
  1237=>"001000100",
  1238=>"011101001",
  1239=>"001011000",
  1240=>"000101010",
  1241=>"110101010",
  1242=>"000110011",
  1243=>"100000110",
  1244=>"000000010",
  1245=>"010011010",
  1246=>"111111100",
  1247=>"110010000",
  1248=>"100000011",
  1249=>"101011101",
  1250=>"111101110",
  1251=>"100111100",
  1252=>"101101001",
  1253=>"101011010",
  1254=>"001101001",
  1255=>"001110001",
  1256=>"000000100",
  1257=>"111100000",
  1258=>"011011001",
  1259=>"011010011",
  1260=>"011110101",
  1261=>"101011010",
  1262=>"001100000",
  1263=>"101111111",
  1264=>"010110100",
  1265=>"000100110",
  1266=>"101100111",
  1267=>"001011001",
  1268=>"101100001",
  1269=>"010111011",
  1270=>"101110101",
  1271=>"010000001",
  1272=>"011111000",
  1273=>"000001100",
  1274=>"111100101",
  1275=>"100111100",
  1276=>"001110111",
  1277=>"000110000",
  1278=>"100100110",
  1279=>"001100011",
  1280=>"010110010",
  1281=>"001011000",
  1282=>"101010111",
  1283=>"111000010",
  1284=>"101101001",
  1285=>"111100101",
  1286=>"100010100",
  1287=>"010000011",
  1288=>"000111100",
  1289=>"110100110",
  1290=>"011110101",
  1291=>"011111111",
  1292=>"101101000",
  1293=>"101000010",
  1294=>"000011000",
  1295=>"110001000",
  1296=>"100000100",
  1297=>"011000101",
  1298=>"111111100",
  1299=>"110110011",
  1300=>"110111100",
  1301=>"110100001",
  1302=>"010111000",
  1303=>"000101111",
  1304=>"111000001",
  1305=>"001011000",
  1306=>"000011000",
  1307=>"100001000",
  1308=>"010101101",
  1309=>"011100000",
  1310=>"000001011",
  1311=>"001001101",
  1312=>"111001011",
  1313=>"101101111",
  1314=>"001001000",
  1315=>"010100110",
  1316=>"111001010",
  1317=>"101100100",
  1318=>"000010101",
  1319=>"001100000",
  1320=>"110001001",
  1321=>"011000111",
  1322=>"110111011",
  1323=>"010011010",
  1324=>"011100001",
  1325=>"000010000",
  1326=>"001011100",
  1327=>"010000110",
  1328=>"001000000",
  1329=>"111100100",
  1330=>"001111011",
  1331=>"010011111",
  1332=>"000000100",
  1333=>"011000001",
  1334=>"101000000",
  1335=>"011101100",
  1336=>"100001011",
  1337=>"011000000",
  1338=>"010010110",
  1339=>"111111110",
  1340=>"101001011",
  1341=>"110110010",
  1342=>"001110011",
  1343=>"111111110",
  1344=>"000010101",
  1345=>"110110110",
  1346=>"110110011",
  1347=>"001011000",
  1348=>"011010000",
  1349=>"111110010",
  1350=>"101100010",
  1351=>"111100001",
  1352=>"010000100",
  1353=>"000001011",
  1354=>"111010100",
  1355=>"101110000",
  1356=>"001000010",
  1357=>"100110101",
  1358=>"111011111",
  1359=>"111101010",
  1360=>"010010100",
  1361=>"100111011",
  1362=>"111001011",
  1363=>"010000010",
  1364=>"100000111",
  1365=>"110011000",
  1366=>"100100010",
  1367=>"000010100",
  1368=>"010100011",
  1369=>"011111100",
  1370=>"000011111",
  1371=>"011001110",
  1372=>"101101001",
  1373=>"001110001",
  1374=>"011111001",
  1375=>"001111011",
  1376=>"000111101",
  1377=>"111110010",
  1378=>"100100010",
  1379=>"000000001",
  1380=>"101101110",
  1381=>"101111000",
  1382=>"101000001",
  1383=>"010100111",
  1384=>"000000000",
  1385=>"001010010",
  1386=>"111101101",
  1387=>"000111000",
  1388=>"000000010",
  1389=>"100100110",
  1390=>"000110000",
  1391=>"110111101",
  1392=>"001010111",
  1393=>"100011010",
  1394=>"101111001",
  1395=>"001000111",
  1396=>"000101001",
  1397=>"110101000",
  1398=>"101011011",
  1399=>"000101001",
  1400=>"101001001",
  1401=>"010011110",
  1402=>"001000111",
  1403=>"011110100",
  1404=>"011011001",
  1405=>"011001011",
  1406=>"000011000",
  1407=>"001100000",
  1408=>"100111011",
  1409=>"101111000",
  1410=>"101011100",
  1411=>"111111100",
  1412=>"100100011",
  1413=>"000000001",
  1414=>"100110111",
  1415=>"011101100",
  1416=>"101101111",
  1417=>"010011010",
  1418=>"101011101",
  1419=>"110111000",
  1420=>"110011111",
  1421=>"010100001",
  1422=>"001010111",
  1423=>"101111101",
  1424=>"110000111",
  1425=>"111010010",
  1426=>"111100011",
  1427=>"110101110",
  1428=>"100011000",
  1429=>"000101001",
  1430=>"101000110",
  1431=>"001110010",
  1432=>"111011110",
  1433=>"101110001",
  1434=>"111100101",
  1435=>"111100010",
  1436=>"001010101",
  1437=>"110000001",
  1438=>"011101100",
  1439=>"101101010",
  1440=>"110100110",
  1441=>"011010010",
  1442=>"000001111",
  1443=>"110001111",
  1444=>"111010100",
  1445=>"010011101",
  1446=>"001110001",
  1447=>"110110010",
  1448=>"100010010",
  1449=>"100110110",
  1450=>"111000100",
  1451=>"111010110",
  1452=>"101110101",
  1453=>"011010101",
  1454=>"010011010",
  1455=>"000010010",
  1456=>"111011100",
  1457=>"000100010",
  1458=>"001010000",
  1459=>"011001010",
  1460=>"001111111",
  1461=>"010011011",
  1462=>"000111000",
  1463=>"001110010",
  1464=>"101111010",
  1465=>"010100010",
  1466=>"111011101",
  1467=>"100111110",
  1468=>"011011111",
  1469=>"010011110",
  1470=>"101000000",
  1471=>"010001011",
  1472=>"100001010",
  1473=>"010111011",
  1474=>"100000010",
  1475=>"000110111",
  1476=>"111001010",
  1477=>"011010011",
  1478=>"001101111",
  1479=>"000000100",
  1480=>"010000001",
  1481=>"101011101",
  1482=>"000100001",
  1483=>"001101011",
  1484=>"000011111",
  1485=>"011111111",
  1486=>"001000000",
  1487=>"100100100",
  1488=>"101100000",
  1489=>"000110111",
  1490=>"100000110",
  1491=>"011011000",
  1492=>"010010010",
  1493=>"010010000",
  1494=>"010100011",
  1495=>"010001100",
  1496=>"010000101",
  1497=>"111011001",
  1498=>"110110110",
  1499=>"011111111",
  1500=>"001000000",
  1501=>"111100011",
  1502=>"001110111",
  1503=>"001110100",
  1504=>"100101000",
  1505=>"000101010",
  1506=>"100100001",
  1507=>"001000101",
  1508=>"011101111",
  1509=>"011111100",
  1510=>"100110111",
  1511=>"101010000",
  1512=>"110100001",
  1513=>"000010001",
  1514=>"001100110",
  1515=>"011111011",
  1516=>"000001000",
  1517=>"011000110",
  1518=>"011101111",
  1519=>"110100001",
  1520=>"101010010",
  1521=>"010010010",
  1522=>"000101010",
  1523=>"110010110",
  1524=>"010001101",
  1525=>"111110100",
  1526=>"111101010",
  1527=>"100100100",
  1528=>"111100100",
  1529=>"000110011",
  1530=>"000111111",
  1531=>"011010001",
  1532=>"111001111",
  1533=>"000110000",
  1534=>"101000101",
  1535=>"100010100",
  1536=>"000100010",
  1537=>"011011001",
  1538=>"110111101",
  1539=>"101010000",
  1540=>"110010101",
  1541=>"001101011",
  1542=>"101101000",
  1543=>"011110110",
  1544=>"100101000",
  1545=>"001000101",
  1546=>"110000000",
  1547=>"011010101",
  1548=>"010000000",
  1549=>"100111111",
  1550=>"100011100",
  1551=>"010100010",
  1552=>"101111101",
  1553=>"111010011",
  1554=>"111001001",
  1555=>"001111011",
  1556=>"001101111",
  1557=>"101111111",
  1558=>"000001101",
  1559=>"100101101",
  1560=>"010010010",
  1561=>"100100011",
  1562=>"011100100",
  1563=>"110000100",
  1564=>"011110101",
  1565=>"110101010",
  1566=>"111010110",
  1567=>"011010001",
  1568=>"011110110",
  1569=>"100010111",
  1570=>"000010011",
  1571=>"000000011",
  1572=>"011001111",
  1573=>"111010101",
  1574=>"011001011",
  1575=>"001001110",
  1576=>"110001110",
  1577=>"011110111",
  1578=>"101111111",
  1579=>"100000001",
  1580=>"001100100",
  1581=>"000100110",
  1582=>"011000100",
  1583=>"010111010",
  1584=>"100001000",
  1585=>"011101110",
  1586=>"101000101",
  1587=>"110000101",
  1588=>"011001000",
  1589=>"111110111",
  1590=>"010110111",
  1591=>"010110100",
  1592=>"100100101",
  1593=>"111001110",
  1594=>"110011010",
  1595=>"111011000",
  1596=>"110010010",
  1597=>"100001111",
  1598=>"000000101",
  1599=>"111101011",
  1600=>"000100111",
  1601=>"000000011",
  1602=>"000001010",
  1603=>"000000111",
  1604=>"000010111",
  1605=>"001111111",
  1606=>"011011001",
  1607=>"001110100",
  1608=>"010100001",
  1609=>"101111110",
  1610=>"011100010",
  1611=>"010011010",
  1612=>"010001000",
  1613=>"110001011",
  1614=>"011011010",
  1615=>"100111100",
  1616=>"001101101",
  1617=>"101100010",
  1618=>"011110111",
  1619=>"111000011",
  1620=>"111100001",
  1621=>"100100100",
  1622=>"101111101",
  1623=>"011100100",
  1624=>"110100101",
  1625=>"010110010",
  1626=>"000000000",
  1627=>"111100111",
  1628=>"011101001",
  1629=>"000011010",
  1630=>"000101110",
  1631=>"110100100",
  1632=>"001010000",
  1633=>"001000000",
  1634=>"110101010",
  1635=>"111111111",
  1636=>"101100111",
  1637=>"001110111",
  1638=>"111111111",
  1639=>"111011110",
  1640=>"000100100",
  1641=>"111011110",
  1642=>"111011110",
  1643=>"111011010",
  1644=>"110100001",
  1645=>"010000110",
  1646=>"000000110",
  1647=>"111001111",
  1648=>"111110111",
  1649=>"010111011",
  1650=>"010111110",
  1651=>"011110101",
  1652=>"001111100",
  1653=>"010000001",
  1654=>"010001110",
  1655=>"101101000",
  1656=>"101000010",
  1657=>"001101011",
  1658=>"000110001",
  1659=>"011011110",
  1660=>"001011010",
  1661=>"111101011",
  1662=>"000100110",
  1663=>"010010001",
  1664=>"100001111",
  1665=>"101111101",
  1666=>"011001011",
  1667=>"100001101",
  1668=>"101101110",
  1669=>"010010110",
  1670=>"100011100",
  1671=>"100111011",
  1672=>"001010110",
  1673=>"011100000",
  1674=>"001111101",
  1675=>"011011110",
  1676=>"010011001",
  1677=>"010011010",
  1678=>"101100010",
  1679=>"000111110",
  1680=>"001010011",
  1681=>"100011010",
  1682=>"111100100",
  1683=>"000100001",
  1684=>"011101011",
  1685=>"001010001",
  1686=>"100110100",
  1687=>"000100101",
  1688=>"011001101",
  1689=>"011100001",
  1690=>"110100000",
  1691=>"111101001",
  1692=>"001001111",
  1693=>"111001001",
  1694=>"111101111",
  1695=>"110110000",
  1696=>"010101101",
  1697=>"110101101",
  1698=>"011110000",
  1699=>"010110110",
  1700=>"011000001",
  1701=>"011010111",
  1702=>"101001011",
  1703=>"101000111",
  1704=>"001000100",
  1705=>"111011011",
  1706=>"000111000",
  1707=>"111000000",
  1708=>"111001110",
  1709=>"010011011",
  1710=>"011001011",
  1711=>"011101010",
  1712=>"101011111",
  1713=>"001101000",
  1714=>"001000101",
  1715=>"000100010",
  1716=>"101001011",
  1717=>"111100101",
  1718=>"101110101",
  1719=>"010100011",
  1720=>"110111010",
  1721=>"101011010",
  1722=>"101010101",
  1723=>"001100110",
  1724=>"101011101",
  1725=>"000110100",
  1726=>"000010010",
  1727=>"111110011",
  1728=>"101010100",
  1729=>"011010000",
  1730=>"100111100",
  1731=>"101111101",
  1732=>"100110111",
  1733=>"111001101",
  1734=>"110110100",
  1735=>"010101001",
  1736=>"010010000",
  1737=>"010110111",
  1738=>"100111000",
  1739=>"000100000",
  1740=>"010011000",
  1741=>"001010001",
  1742=>"101100010",
  1743=>"101100011",
  1744=>"111001000",
  1745=>"011101100",
  1746=>"110100111",
  1747=>"110110101",
  1748=>"100011111",
  1749=>"100111010",
  1750=>"001101011",
  1751=>"110100110",
  1752=>"111111100",
  1753=>"111110110",
  1754=>"100101111",
  1755=>"010100011",
  1756=>"100001101",
  1757=>"001001110",
  1758=>"101000000",
  1759=>"001001011",
  1760=>"010100000",
  1761=>"010010010",
  1762=>"110101101",
  1763=>"010010101",
  1764=>"111001111",
  1765=>"011001100",
  1766=>"010001111",
  1767=>"000100100",
  1768=>"101000011",
  1769=>"011001001",
  1770=>"010100111",
  1771=>"110010001",
  1772=>"001010010",
  1773=>"101100000",
  1774=>"001100000",
  1775=>"101100000",
  1776=>"011100000",
  1777=>"111110000",
  1778=>"111001110",
  1779=>"010101010",
  1780=>"101010011",
  1781=>"001111011",
  1782=>"011100011",
  1783=>"001111000",
  1784=>"001000011",
  1785=>"101101100",
  1786=>"101101111",
  1787=>"011010000",
  1788=>"010011001",
  1789=>"111110000",
  1790=>"010011000",
  1791=>"001110000",
  1792=>"101101110",
  1793=>"110001001",
  1794=>"110001001",
  1795=>"001011000",
  1796=>"101010011",
  1797=>"000011001",
  1798=>"100010000",
  1799=>"001001111",
  1800=>"001100000",
  1801=>"010011111",
  1802=>"101001100",
  1803=>"111101000",
  1804=>"101000101",
  1805=>"001111011",
  1806=>"010011010",
  1807=>"000001010",
  1808=>"001001001",
  1809=>"001010010",
  1810=>"000101011",
  1811=>"010000011",
  1812=>"001000111",
  1813=>"001000111",
  1814=>"000000000",
  1815=>"110010010",
  1816=>"100110000",
  1817=>"110000000",
  1818=>"000111101",
  1819=>"010011101",
  1820=>"111001111",
  1821=>"000110110",
  1822=>"101011000",
  1823=>"010110100",
  1824=>"100100100",
  1825=>"001110111",
  1826=>"001001101",
  1827=>"101101111",
  1828=>"011001111",
  1829=>"000100011",
  1830=>"000110110",
  1831=>"100000110",
  1832=>"110110111",
  1833=>"000110010",
  1834=>"011011110",
  1835=>"101100100",
  1836=>"001100100",
  1837=>"001010010",
  1838=>"101010011",
  1839=>"101010101",
  1840=>"001001011",
  1841=>"011001110",
  1842=>"001010111",
  1843=>"110010000",
  1844=>"001110000",
  1845=>"110000011",
  1846=>"001000000",
  1847=>"101101101",
  1848=>"000100101",
  1849=>"101101111",
  1850=>"100010011",
  1851=>"101010110",
  1852=>"000111001",
  1853=>"111111111",
  1854=>"110111110",
  1855=>"111111111",
  1856=>"010010101",
  1857=>"000000000",
  1858=>"010100110",
  1859=>"001010110",
  1860=>"101010000",
  1861=>"000010011",
  1862=>"111100101",
  1863=>"010011101",
  1864=>"001001011",
  1865=>"101010110",
  1866=>"101001110",
  1867=>"000101010",
  1868=>"011010111",
  1869=>"101000111",
  1870=>"111111010",
  1871=>"100010011",
  1872=>"010001110",
  1873=>"101000110",
  1874=>"011110111",
  1875=>"110010110",
  1876=>"110101101",
  1877=>"011001110",
  1878=>"110110000",
  1879=>"101001111",
  1880=>"010010001",
  1881=>"101010000",
  1882=>"110101111",
  1883=>"001001111",
  1884=>"001111011",
  1885=>"000010111",
  1886=>"110001010",
  1887=>"100010010",
  1888=>"010010010",
  1889=>"111101011",
  1890=>"011010001",
  1891=>"111110110",
  1892=>"001000001",
  1893=>"111111000",
  1894=>"001010010",
  1895=>"100111100",
  1896=>"000001110",
  1897=>"001100010",
  1898=>"011100110",
  1899=>"000011111",
  1900=>"111011000",
  1901=>"111101111",
  1902=>"001010010",
  1903=>"010101011",
  1904=>"111110000",
  1905=>"101100101",
  1906=>"111010010",
  1907=>"000010101",
  1908=>"110000001",
  1909=>"111001101",
  1910=>"000111101",
  1911=>"011110100",
  1912=>"001110110",
  1913=>"111010100",
  1914=>"000100001",
  1915=>"100011100",
  1916=>"101000100",
  1917=>"000010001",
  1918=>"110000010",
  1919=>"100101110",
  1920=>"111011000",
  1921=>"111100110",
  1922=>"000000111",
  1923=>"011110110",
  1924=>"110111001",
  1925=>"111011001",
  1926=>"111101010",
  1927=>"100110010",
  1928=>"110101001",
  1929=>"010001010",
  1930=>"011110110",
  1931=>"001001000",
  1932=>"001110011",
  1933=>"110110111",
  1934=>"000100111",
  1935=>"001101110",
  1936=>"110000001",
  1937=>"100011100",
  1938=>"010100100",
  1939=>"000001100",
  1940=>"111110101",
  1941=>"110110110",
  1942=>"000110001",
  1943=>"001001010",
  1944=>"010001001",
  1945=>"010110010",
  1946=>"000101111",
  1947=>"011001001",
  1948=>"101001001",
  1949=>"111111111",
  1950=>"010000000",
  1951=>"000000101",
  1952=>"010001110",
  1953=>"111100011",
  1954=>"010101001",
  1955=>"010001100",
  1956=>"001111000",
  1957=>"101011100",
  1958=>"110101110",
  1959=>"010001010",
  1960=>"001010001",
  1961=>"101110111",
  1962=>"101110100",
  1963=>"110000110",
  1964=>"010100010",
  1965=>"111001101",
  1966=>"100011010",
  1967=>"011110011",
  1968=>"101110001",
  1969=>"111111100",
  1970=>"100100100",
  1971=>"100010100",
  1972=>"011110001",
  1973=>"111000100",
  1974=>"011011001",
  1975=>"011010110",
  1976=>"011010000",
  1977=>"101101110",
  1978=>"000101111",
  1979=>"100010100",
  1980=>"000010111",
  1981=>"000011000",
  1982=>"101011101",
  1983=>"100111011",
  1984=>"110111000",
  1985=>"101101110",
  1986=>"101010010",
  1987=>"110010100",
  1988=>"000000000",
  1989=>"111101011",
  1990=>"000000000",
  1991=>"100111001",
  1992=>"101001101",
  1993=>"100111011",
  1994=>"000100011",
  1995=>"010010011",
  1996=>"111100010",
  1997=>"100000001",
  1998=>"101111110",
  1999=>"011100111",
  2000=>"001011000",
  2001=>"011101100",
  2002=>"111110111",
  2003=>"011111000",
  2004=>"000010111",
  2005=>"111011111",
  2006=>"001000100",
  2007=>"000101010",
  2008=>"111000000",
  2009=>"001011110",
  2010=>"010001010",
  2011=>"000001110",
  2012=>"101111011",
  2013=>"000101110",
  2014=>"101001011",
  2015=>"111111110",
  2016=>"011000111",
  2017=>"011001000",
  2018=>"110100011",
  2019=>"100010011",
  2020=>"000011110",
  2021=>"101101111",
  2022=>"010011010",
  2023=>"001101010",
  2024=>"010111001",
  2025=>"101111100",
  2026=>"100111111",
  2027=>"111110001",
  2028=>"111001010",
  2029=>"110011111",
  2030=>"101111011",
  2031=>"110101011",
  2032=>"110110011",
  2033=>"100000111",
  2034=>"101001010",
  2035=>"000100001",
  2036=>"101001001",
  2037=>"101011100",
  2038=>"110110000",
  2039=>"011010111",
  2040=>"011011111",
  2041=>"001110111",
  2042=>"111100000",
  2043=>"010110101",
  2044=>"010101111",
  2045=>"001101011",
  2046=>"100001111",
  2047=>"101101101",
  2048=>"101001010",
  2049=>"100110101",
  2050=>"101100011",
  2051=>"110100010",
  2052=>"000010110",
  2053=>"111101011",
  2054=>"100101100",
  2055=>"001101101",
  2056=>"111010111",
  2057=>"101110111",
  2058=>"110111100",
  2059=>"110010011",
  2060=>"000100010",
  2061=>"001101000",
  2062=>"010100010",
  2063=>"011101000",
  2064=>"111100101",
  2065=>"011100011",
  2066=>"111101001",
  2067=>"001001110",
  2068=>"010100111",
  2069=>"111101011",
  2070=>"101000000",
  2071=>"000000000",
  2072=>"100000011",
  2073=>"011011011",
  2074=>"000101010",
  2075=>"011011001",
  2076=>"110010110",
  2077=>"011100010",
  2078=>"110100111",
  2079=>"001110010",
  2080=>"101101101",
  2081=>"100000101",
  2082=>"111001000",
  2083=>"101101010",
  2084=>"010001110",
  2085=>"111110101",
  2086=>"000011011",
  2087=>"001010111",
  2088=>"101110101",
  2089=>"011100110",
  2090=>"101100011",
  2091=>"000000010",
  2092=>"010011000",
  2093=>"101001010",
  2094=>"011110100",
  2095=>"001111001",
  2096=>"111100110",
  2097=>"111111110",
  2098=>"110011010",
  2099=>"111010110",
  2100=>"001011010",
  2101=>"001101100",
  2102=>"101101000",
  2103=>"001100110",
  2104=>"111000110",
  2105=>"011100100",
  2106=>"001111110",
  2107=>"101101101",
  2108=>"110001011",
  2109=>"101010010",
  2110=>"000001100",
  2111=>"101001101",
  2112=>"011000010",
  2113=>"101000001",
  2114=>"101011101",
  2115=>"111000011",
  2116=>"111111101",
  2117=>"100011001",
  2118=>"011001010",
  2119=>"011001000",
  2120=>"111111011",
  2121=>"101001001",
  2122=>"011101010",
  2123=>"010111010",
  2124=>"110110001",
  2125=>"101111000",
  2126=>"111111000",
  2127=>"110011001",
  2128=>"111000000",
  2129=>"101001001",
  2130=>"101000011",
  2131=>"010101010",
  2132=>"110111011",
  2133=>"100111101",
  2134=>"110110101",
  2135=>"110111100",
  2136=>"011001000",
  2137=>"011100001",
  2138=>"000111110",
  2139=>"010100001",
  2140=>"110001111",
  2141=>"111100100",
  2142=>"100101001",
  2143=>"110100100",
  2144=>"001001001",
  2145=>"011111101",
  2146=>"101000011",
  2147=>"010101110",
  2148=>"010000101",
  2149=>"010001011",
  2150=>"111010101",
  2151=>"011001111",
  2152=>"110101000",
  2153=>"111001110",
  2154=>"101010000",
  2155=>"110110100",
  2156=>"111000000",
  2157=>"010111000",
  2158=>"100000101",
  2159=>"100111111",
  2160=>"101001010",
  2161=>"001011110",
  2162=>"100000000",
  2163=>"100010010",
  2164=>"110010000",
  2165=>"011110110",
  2166=>"000001000",
  2167=>"110010101",
  2168=>"001001011",
  2169=>"011111111",
  2170=>"100001100",
  2171=>"111101100",
  2172=>"000001010",
  2173=>"011111001",
  2174=>"010010010",
  2175=>"010101010",
  2176=>"010111010",
  2177=>"001101001",
  2178=>"000000110",
  2179=>"001011001",
  2180=>"111011110",
  2181=>"110011100",
  2182=>"111100111",
  2183=>"100110111",
  2184=>"011100010",
  2185=>"100110110",
  2186=>"111010101",
  2187=>"011100101",
  2188=>"000011111",
  2189=>"000110101",
  2190=>"100000001",
  2191=>"101101001",
  2192=>"110011100",
  2193=>"111110101",
  2194=>"010100000",
  2195=>"001010001",
  2196=>"010110100",
  2197=>"100100100",
  2198=>"011111001",
  2199=>"010010101",
  2200=>"010010111",
  2201=>"101001111",
  2202=>"110000011",
  2203=>"100111111",
  2204=>"100110101",
  2205=>"000110001",
  2206=>"010011011",
  2207=>"000101011",
  2208=>"010010011",
  2209=>"100011110",
  2210=>"011001110",
  2211=>"011001101",
  2212=>"100110101",
  2213=>"111000000",
  2214=>"000010001",
  2215=>"111000100",
  2216=>"111110001",
  2217=>"101001000",
  2218=>"100011000",
  2219=>"000000100",
  2220=>"010110010",
  2221=>"110001110",
  2222=>"111100011",
  2223=>"000001110",
  2224=>"001101010",
  2225=>"000010110",
  2226=>"111101110",
  2227=>"010111001",
  2228=>"010011001",
  2229=>"000100011",
  2230=>"001111101",
  2231=>"001011101",
  2232=>"000001111",
  2233=>"101000111",
  2234=>"011000001",
  2235=>"101111011",
  2236=>"100111111",
  2237=>"111010000",
  2238=>"111110001",
  2239=>"011111111",
  2240=>"101011100",
  2241=>"111000111",
  2242=>"100101011",
  2243=>"110000000",
  2244=>"011000011",
  2245=>"000000011",
  2246=>"001100111",
  2247=>"011000100",
  2248=>"001111111",
  2249=>"001001100",
  2250=>"010110100",
  2251=>"000001111",
  2252=>"110101000",
  2253=>"000001111",
  2254=>"111110000",
  2255=>"110010100",
  2256=>"111111111",
  2257=>"101110101",
  2258=>"001101010",
  2259=>"011110000",
  2260=>"011101110",
  2261=>"101110011",
  2262=>"011010000",
  2263=>"110111111",
  2264=>"001111001",
  2265=>"110011110",
  2266=>"001010010",
  2267=>"001010101",
  2268=>"100001000",
  2269=>"000101110",
  2270=>"001111000",
  2271=>"000011001",
  2272=>"010010110",
  2273=>"001001010",
  2274=>"010101111",
  2275=>"111111101",
  2276=>"100001111",
  2277=>"000100010",
  2278=>"100000011",
  2279=>"110110101",
  2280=>"001011101",
  2281=>"101000100",
  2282=>"110111000",
  2283=>"100011000",
  2284=>"111111001",
  2285=>"010111011",
  2286=>"011100011",
  2287=>"110011111",
  2288=>"011000100",
  2289=>"001010000",
  2290=>"000011011",
  2291=>"010100000",
  2292=>"101010010",
  2293=>"111100110",
  2294=>"110011110",
  2295=>"100101111",
  2296=>"100000101",
  2297=>"000011001",
  2298=>"001001110",
  2299=>"100000100",
  2300=>"000100010",
  2301=>"001011110",
  2302=>"011101010",
  2303=>"000011110",
  2304=>"010101101",
  2305=>"011100001",
  2306=>"000001111",
  2307=>"010100110",
  2308=>"000010100",
  2309=>"011111100",
  2310=>"110001110",
  2311=>"110110000",
  2312=>"011110011",
  2313=>"001001001",
  2314=>"001010010",
  2315=>"100010000",
  2316=>"111011111",
  2317=>"100111010",
  2318=>"100001110",
  2319=>"010000010",
  2320=>"110100011",
  2321=>"101000100",
  2322=>"001101010",
  2323=>"100101010",
  2324=>"110010011",
  2325=>"011110110",
  2326=>"001111111",
  2327=>"011101110",
  2328=>"010101111",
  2329=>"000110000",
  2330=>"010000111",
  2331=>"110110100",
  2332=>"010100011",
  2333=>"100011000",
  2334=>"000011000",
  2335=>"101100110",
  2336=>"010101011",
  2337=>"111000001",
  2338=>"100000100",
  2339=>"011100001",
  2340=>"100100100",
  2341=>"000001110",
  2342=>"010010110",
  2343=>"000100000",
  2344=>"001010101",
  2345=>"110010010",
  2346=>"001111100",
  2347=>"001111101",
  2348=>"101000101",
  2349=>"001000010",
  2350=>"011110010",
  2351=>"000100000",
  2352=>"000001110",
  2353=>"101000010",
  2354=>"100000110",
  2355=>"001010101",
  2356=>"111110000",
  2357=>"011101110",
  2358=>"000101110",
  2359=>"110110000",
  2360=>"000100110",
  2361=>"111110001",
  2362=>"011111010",
  2363=>"101111010",
  2364=>"111101100",
  2365=>"001000110",
  2366=>"101010101",
  2367=>"111101101",
  2368=>"010000100",
  2369=>"000111010",
  2370=>"011011101",
  2371=>"111011001",
  2372=>"110010101",
  2373=>"001110001",
  2374=>"110101111",
  2375=>"111111111",
  2376=>"100101001",
  2377=>"100000101",
  2378=>"111000000",
  2379=>"010010000",
  2380=>"110001010",
  2381=>"110110111",
  2382=>"100111111",
  2383=>"010001000",
  2384=>"110011010",
  2385=>"101110100",
  2386=>"011000001",
  2387=>"011011011",
  2388=>"010000010",
  2389=>"111111000",
  2390=>"101010010",
  2391=>"001101010",
  2392=>"000111001",
  2393=>"111011101",
  2394=>"011011010",
  2395=>"111001010",
  2396=>"011111111",
  2397=>"011000110",
  2398=>"111011101",
  2399=>"110010011",
  2400=>"010101000",
  2401=>"101101100",
  2402=>"000010000",
  2403=>"001010000",
  2404=>"011000000",
  2405=>"101001111",
  2406=>"101110110",
  2407=>"001110101",
  2408=>"000110011",
  2409=>"000100111",
  2410=>"011011111",
  2411=>"011101111",
  2412=>"000101111",
  2413=>"011110100",
  2414=>"000001101",
  2415=>"101101111",
  2416=>"111010010",
  2417=>"000110111",
  2418=>"110111001",
  2419=>"111010110",
  2420=>"000010100",
  2421=>"000010001",
  2422=>"111001000",
  2423=>"000010100",
  2424=>"111101001",
  2425=>"010010001",
  2426=>"100011000",
  2427=>"111011111",
  2428=>"010010000",
  2429=>"100011000",
  2430=>"011001011",
  2431=>"100010011",
  2432=>"010110110",
  2433=>"010001111",
  2434=>"101100011",
  2435=>"000100011",
  2436=>"010010100",
  2437=>"000110100",
  2438=>"101101001",
  2439=>"001111011",
  2440=>"001011111",
  2441=>"011100000",
  2442=>"101110111",
  2443=>"010011001",
  2444=>"001101010",
  2445=>"100001001",
  2446=>"011110000",
  2447=>"010010011",
  2448=>"101100010",
  2449=>"010100001",
  2450=>"110001101",
  2451=>"000101110",
  2452=>"110110010",
  2453=>"010000010",
  2454=>"000110010",
  2455=>"000101111",
  2456=>"101000100",
  2457=>"110111000",
  2458=>"001100100",
  2459=>"111010011",
  2460=>"110101111",
  2461=>"000110111",
  2462=>"011101010",
  2463=>"000001001",
  2464=>"111110100",
  2465=>"011000110",
  2466=>"100110011",
  2467=>"100101111",
  2468=>"011011100",
  2469=>"011111111",
  2470=>"111111111",
  2471=>"000101111",
  2472=>"111111111",
  2473=>"100101111",
  2474=>"110001000",
  2475=>"000111111",
  2476=>"110000000",
  2477=>"100111111",
  2478=>"100000000",
  2479=>"011000000",
  2480=>"111001011",
  2481=>"011000011",
  2482=>"110101001",
  2483=>"111110011",
  2484=>"000010111",
  2485=>"000001011",
  2486=>"000111001",
  2487=>"111001100",
  2488=>"010100001",
  2489=>"111111000",
  2490=>"011011011",
  2491=>"011000111",
  2492=>"000011111",
  2493=>"110100011",
  2494=>"011101001",
  2495=>"001111011",
  2496=>"110110000",
  2497=>"000001100",
  2498=>"011101100",
  2499=>"000101010",
  2500=>"111001000",
  2501=>"101001101",
  2502=>"111001010",
  2503=>"011011100",
  2504=>"100001011",
  2505=>"100110100",
  2506=>"101101010",
  2507=>"011011101",
  2508=>"001000010",
  2509=>"110101110",
  2510=>"001111111",
  2511=>"100011010",
  2512=>"000111101",
  2513=>"011001010",
  2514=>"000111000",
  2515=>"000000010",
  2516=>"011001110",
  2517=>"101100100",
  2518=>"110111000",
  2519=>"111111111",
  2520=>"100110011",
  2521=>"110101010",
  2522=>"011011111",
  2523=>"000010010",
  2524=>"100111001",
  2525=>"111010101",
  2526=>"100001110",
  2527=>"010110111",
  2528=>"010100011",
  2529=>"100100101",
  2530=>"100000001",
  2531=>"010000000",
  2532=>"011000010",
  2533=>"111011010",
  2534=>"110000101",
  2535=>"001111000",
  2536=>"110001110",
  2537=>"000110000",
  2538=>"000001011",
  2539=>"101111111",
  2540=>"111111111",
  2541=>"111101010",
  2542=>"111010001",
  2543=>"111001110",
  2544=>"000100010",
  2545=>"001111110",
  2546=>"100111000",
  2547=>"010001101",
  2548=>"101011101",
  2549=>"101011000",
  2550=>"011111111",
  2551=>"100011010",
  2552=>"111000011",
  2553=>"101000110",
  2554=>"001000011",
  2555=>"111011000",
  2556=>"001101100",
  2557=>"111101000",
  2558=>"101111001",
  2559=>"101101100",
  2560=>"100110100",
  2561=>"010001011",
  2562=>"011001000",
  2563=>"001000011",
  2564=>"001110001",
  2565=>"101001100",
  2566=>"111010010",
  2567=>"000111110",
  2568=>"011100000",
  2569=>"001100101",
  2570=>"111011111",
  2571=>"000101110",
  2572=>"100111111",
  2573=>"110011001",
  2574=>"110000101",
  2575=>"111100000",
  2576=>"111110010",
  2577=>"110110100",
  2578=>"001010101",
  2579=>"111101000",
  2580=>"100101010",
  2581=>"111111011",
  2582=>"010011011",
  2583=>"111011010",
  2584=>"111000000",
  2585=>"010111110",
  2586=>"111010010",
  2587=>"011011000",
  2588=>"110111110",
  2589=>"010001101",
  2590=>"000000110",
  2591=>"111110111",
  2592=>"111111001",
  2593=>"011100000",
  2594=>"111010100",
  2595=>"010010110",
  2596=>"010110100",
  2597=>"111110100",
  2598=>"001100101",
  2599=>"011001010",
  2600=>"001010011",
  2601=>"010110011",
  2602=>"001001101",
  2603=>"110111110",
  2604=>"111100011",
  2605=>"011110000",
  2606=>"001110000",
  2607=>"101100101",
  2608=>"000100100",
  2609=>"110010111",
  2610=>"010011111",
  2611=>"001111010",
  2612=>"000000000",
  2613=>"101101110",
  2614=>"001000101",
  2615=>"101101010",
  2616=>"000011000",
  2617=>"001110101",
  2618=>"000011110",
  2619=>"111111101",
  2620=>"100110010",
  2621=>"000000010",
  2622=>"101110101",
  2623=>"100010010",
  2624=>"111100011",
  2625=>"111111011",
  2626=>"010011001",
  2627=>"000111110",
  2628=>"001011101",
  2629=>"100011111",
  2630=>"011100110",
  2631=>"000110111",
  2632=>"100111100",
  2633=>"111011101",
  2634=>"111000001",
  2635=>"100111101",
  2636=>"001110110",
  2637=>"001111101",
  2638=>"110000001",
  2639=>"110000100",
  2640=>"010011111",
  2641=>"001010001",
  2642=>"001001000",
  2643=>"000001110",
  2644=>"011101001",
  2645=>"111010010",
  2646=>"111101000",
  2647=>"100001110",
  2648=>"101011011",
  2649=>"101101111",
  2650=>"100010010",
  2651=>"010000111",
  2652=>"111000100",
  2653=>"000010011",
  2654=>"000000001",
  2655=>"110100101",
  2656=>"100110110",
  2657=>"101110010",
  2658=>"100100000",
  2659=>"111010011",
  2660=>"110111100",
  2661=>"110111010",
  2662=>"110010110",
  2663=>"001101011",
  2664=>"101001101",
  2665=>"001111100",
  2666=>"001000011",
  2667=>"000101001",
  2668=>"000000100",
  2669=>"010001011",
  2670=>"010101001",
  2671=>"110100111",
  2672=>"000100000",
  2673=>"101011011",
  2674=>"110110001",
  2675=>"100110101",
  2676=>"000111000",
  2677=>"000101000",
  2678=>"000110001",
  2679=>"110000010",
  2680=>"101001000",
  2681=>"010111110",
  2682=>"010010010",
  2683=>"101100000",
  2684=>"111100111",
  2685=>"010010101",
  2686=>"001011011",
  2687=>"000100000",
  2688=>"111101011",
  2689=>"111010101",
  2690=>"100011101",
  2691=>"101101110",
  2692=>"001011011",
  2693=>"011001010",
  2694=>"011001110",
  2695=>"100100101",
  2696=>"100000100",
  2697=>"110011111",
  2698=>"011010010",
  2699=>"110000001",
  2700=>"100010000",
  2701=>"000110001",
  2702=>"001100000",
  2703=>"111000100",
  2704=>"100010011",
  2705=>"011100101",
  2706=>"101010001",
  2707=>"001001000",
  2708=>"101000001",
  2709=>"001111111",
  2710=>"011101100",
  2711=>"110101000",
  2712=>"111011011",
  2713=>"011111111",
  2714=>"001010100",
  2715=>"111101110",
  2716=>"000111111",
  2717=>"011111001",
  2718=>"110001100",
  2719=>"001111110",
  2720=>"101100011",
  2721=>"001111010",
  2722=>"100010100",
  2723=>"001010110",
  2724=>"001001001",
  2725=>"100100001",
  2726=>"100100111",
  2727=>"110011110",
  2728=>"100111010",
  2729=>"000110011",
  2730=>"000101000",
  2731=>"100100010",
  2732=>"100101000",
  2733=>"101000100",
  2734=>"001100000",
  2735=>"101101101",
  2736=>"101101110",
  2737=>"100011010",
  2738=>"010100001",
  2739=>"101000100",
  2740=>"110010100",
  2741=>"101100100",
  2742=>"011100111",
  2743=>"111010010",
  2744=>"100000010",
  2745=>"111000000",
  2746=>"010111000",
  2747=>"101100110",
  2748=>"010000110",
  2749=>"111010011",
  2750=>"011000001",
  2751=>"000110001",
  2752=>"010111001",
  2753=>"010100101",
  2754=>"100111001",
  2755=>"001001011",
  2756=>"010110110",
  2757=>"000000110",
  2758=>"011000000",
  2759=>"101111101",
  2760=>"001000100",
  2761=>"011101011",
  2762=>"010110001",
  2763=>"000110110",
  2764=>"001111100",
  2765=>"110011101",
  2766=>"010010010",
  2767=>"001101111",
  2768=>"111100110",
  2769=>"111010010",
  2770=>"111100110",
  2771=>"000100111",
  2772=>"011110011",
  2773=>"101110110",
  2774=>"011110010",
  2775=>"111001011",
  2776=>"000110110",
  2777=>"110011111",
  2778=>"010010000",
  2779=>"100000000",
  2780=>"111010000",
  2781=>"101001101",
  2782=>"001001001",
  2783=>"010101000",
  2784=>"111001011",
  2785=>"011111001",
  2786=>"100111000",
  2787=>"111111110",
  2788=>"000101001",
  2789=>"011010110",
  2790=>"010000100",
  2791=>"110100000",
  2792=>"111101001",
  2793=>"111101010",
  2794=>"110101000",
  2795=>"000100010",
  2796=>"000000111",
  2797=>"100001001",
  2798=>"101010110",
  2799=>"001010010",
  2800=>"000000001",
  2801=>"001010011",
  2802=>"000001001",
  2803=>"001010100",
  2804=>"011100101",
  2805=>"111001110",
  2806=>"111101011",
  2807=>"000101110",
  2808=>"110100010",
  2809=>"001100111",
  2810=>"011110110",
  2811=>"110111010",
  2812=>"000111000",
  2813=>"111001011",
  2814=>"010110110",
  2815=>"000011000",
  2816=>"000000000",
  2817=>"000100010",
  2818=>"011010000",
  2819=>"101000110",
  2820=>"110011111",
  2821=>"111100101",
  2822=>"110010011",
  2823=>"000100010",
  2824=>"100111011",
  2825=>"010000010",
  2826=>"100011111",
  2827=>"010111100",
  2828=>"000011100",
  2829=>"100111101",
  2830=>"001001010",
  2831=>"100110011",
  2832=>"011010100",
  2833=>"011101000",
  2834=>"010000000",
  2835=>"010110101",
  2836=>"010101011",
  2837=>"001010101",
  2838=>"100001100",
  2839=>"100000010",
  2840=>"010111010",
  2841=>"100100101",
  2842=>"000100101",
  2843=>"111010010",
  2844=>"110011010",
  2845=>"000011011",
  2846=>"100001001",
  2847=>"100000100",
  2848=>"111100000",
  2849=>"011100010",
  2850=>"011100001",
  2851=>"111101011",
  2852=>"111000101",
  2853=>"101000100",
  2854=>"010111000",
  2855=>"011111111",
  2856=>"011000111",
  2857=>"001000100",
  2858=>"000111000",
  2859=>"000000010",
  2860=>"001110111",
  2861=>"100000111",
  2862=>"000000101",
  2863=>"000011111",
  2864=>"000101101",
  2865=>"111001110",
  2866=>"100101001",
  2867=>"001100100",
  2868=>"110111000",
  2869=>"111001011",
  2870=>"011110000",
  2871=>"101111110",
  2872=>"110111111",
  2873=>"001101101",
  2874=>"111000000",
  2875=>"101101111",
  2876=>"000001101",
  2877=>"111010001",
  2878=>"001110100",
  2879=>"011000011",
  2880=>"101101100",
  2881=>"101111110",
  2882=>"000000001",
  2883=>"110001001",
  2884=>"110010100",
  2885=>"011001100",
  2886=>"110010001",
  2887=>"010011010",
  2888=>"111111011",
  2889=>"001000100",
  2890=>"100101111",
  2891=>"111100011",
  2892=>"001001101",
  2893=>"110011011",
  2894=>"000001101",
  2895=>"101011111",
  2896=>"100000101",
  2897=>"011001101",
  2898=>"011000011",
  2899=>"011100010",
  2900=>"011001110",
  2901=>"000000111",
  2902=>"100100101",
  2903=>"100000000",
  2904=>"000011101",
  2905=>"110010110",
  2906=>"000101010",
  2907=>"100001101",
  2908=>"110111011",
  2909=>"111111000",
  2910=>"011001111",
  2911=>"110010001",
  2912=>"010010111",
  2913=>"100101100",
  2914=>"011000010",
  2915=>"000010011",
  2916=>"011001001",
  2917=>"001011011",
  2918=>"000011111",
  2919=>"111110101",
  2920=>"010011000",
  2921=>"000111001",
  2922=>"010111011",
  2923=>"110111001",
  2924=>"100100010",
  2925=>"100000111",
  2926=>"001011010",
  2927=>"011101000",
  2928=>"000010010",
  2929=>"100110010",
  2930=>"111111111",
  2931=>"111101010",
  2932=>"000110100",
  2933=>"111010100",
  2934=>"100010110",
  2935=>"110001011",
  2936=>"101001101",
  2937=>"001111011",
  2938=>"111101011",
  2939=>"110011011",
  2940=>"011000001",
  2941=>"001010110",
  2942=>"011011110",
  2943=>"010011000",
  2944=>"010011100",
  2945=>"111001000",
  2946=>"110000001",
  2947=>"010001001",
  2948=>"111101111",
  2949=>"110100110",
  2950=>"110101111",
  2951=>"101111110",
  2952=>"011000001",
  2953=>"110111111",
  2954=>"111110000",
  2955=>"000011110",
  2956=>"000110010",
  2957=>"111101111",
  2958=>"000111111",
  2959=>"111111111",
  2960=>"001011100",
  2961=>"000011100",
  2962=>"011000101",
  2963=>"101001110",
  2964=>"111110001",
  2965=>"111001100",
  2966=>"000000111",
  2967=>"000111111",
  2968=>"101111111",
  2969=>"111011101",
  2970=>"010101011",
  2971=>"111011001",
  2972=>"101000010",
  2973=>"000000100",
  2974=>"100001010",
  2975=>"111001110",
  2976=>"001001110",
  2977=>"100111111",
  2978=>"110011000",
  2979=>"000100001",
  2980=>"000010000",
  2981=>"100000011",
  2982=>"010000000",
  2983=>"011111010",
  2984=>"100100101",
  2985=>"010110000",
  2986=>"001100010",
  2987=>"011100100",
  2988=>"011110011",
  2989=>"011001111",
  2990=>"011001011",
  2991=>"010111111",
  2992=>"001101011",
  2993=>"010010110",
  2994=>"010001101",
  2995=>"010011000",
  2996=>"111101100",
  2997=>"000010000",
  2998=>"011100010",
  2999=>"001011111",
  3000=>"110011111",
  3001=>"100010100",
  3002=>"100011101",
  3003=>"000001110",
  3004=>"000010011",
  3005=>"101000101",
  3006=>"000111011",
  3007=>"000011000",
  3008=>"110001010",
  3009=>"101101110",
  3010=>"000100010",
  3011=>"111011000",
  3012=>"011000111",
  3013=>"000101100",
  3014=>"011111010",
  3015=>"101000110",
  3016=>"000110010",
  3017=>"001010011",
  3018=>"011111010",
  3019=>"111111001",
  3020=>"010111000",
  3021=>"111101001",
  3022=>"001000010",
  3023=>"001100110",
  3024=>"100011111",
  3025=>"110110001",
  3026=>"001101010",
  3027=>"110101010",
  3028=>"001101110",
  3029=>"001111111",
  3030=>"000100001",
  3031=>"110001000",
  3032=>"100100000",
  3033=>"110011011",
  3034=>"111010111",
  3035=>"000001001",
  3036=>"000100111",
  3037=>"010100101",
  3038=>"110011101",
  3039=>"001010001",
  3040=>"100110110",
  3041=>"101010000",
  3042=>"100001010",
  3043=>"101011100",
  3044=>"111001001",
  3045=>"000100011",
  3046=>"100011100",
  3047=>"000100000",
  3048=>"000010110",
  3049=>"101001101",
  3050=>"110000100",
  3051=>"111000110",
  3052=>"101110100",
  3053=>"100110111",
  3054=>"001100001",
  3055=>"010010010",
  3056=>"000000110",
  3057=>"111010100",
  3058=>"111010000",
  3059=>"111110111",
  3060=>"000001001",
  3061=>"010111001",
  3062=>"000000010",
  3063=>"110111101",
  3064=>"101111100",
  3065=>"101110101",
  3066=>"010001001",
  3067=>"101011011",
  3068=>"001000111",
  3069=>"110010100",
  3070=>"000000000",
  3071=>"000101001",
  3072=>"111000110",
  3073=>"110101010",
  3074=>"110011010",
  3075=>"100111000",
  3076=>"111100101",
  3077=>"010110111",
  3078=>"110110001",
  3079=>"111101000",
  3080=>"111100011",
  3081=>"100000001",
  3082=>"000001001",
  3083=>"000011110",
  3084=>"110011111",
  3085=>"000011001",
  3086=>"010010011",
  3087=>"111001010",
  3088=>"001011000",
  3089=>"111111000",
  3090=>"000000111",
  3091=>"000111011",
  3092=>"011100101",
  3093=>"000011100",
  3094=>"011100001",
  3095=>"000110111",
  3096=>"010111000",
  3097=>"110100111",
  3098=>"001000100",
  3099=>"111100100",
  3100=>"001111011",
  3101=>"010001101",
  3102=>"011011001",
  3103=>"011111001",
  3104=>"111111001",
  3105=>"110010001",
  3106=>"100111011",
  3107=>"000001011",
  3108=>"111111101",
  3109=>"011000000",
  3110=>"011101010",
  3111=>"001101110",
  3112=>"111011000",
  3113=>"001000001",
  3114=>"011011011",
  3115=>"111010110",
  3116=>"111101111",
  3117=>"000111001",
  3118=>"001001000",
  3119=>"111111011",
  3120=>"000101001",
  3121=>"111100110",
  3122=>"110000001",
  3123=>"110110010",
  3124=>"111110111",
  3125=>"110000011",
  3126=>"100001111",
  3127=>"010100100",
  3128=>"011110010",
  3129=>"000001011",
  3130=>"100000100",
  3131=>"000010101",
  3132=>"001111100",
  3133=>"000000010",
  3134=>"111111010",
  3135=>"000011100",
  3136=>"100101010",
  3137=>"011011100",
  3138=>"100010001",
  3139=>"011010101",
  3140=>"110010001",
  3141=>"110111111",
  3142=>"101001011",
  3143=>"000011001",
  3144=>"101101010",
  3145=>"111101101",
  3146=>"110000110",
  3147=>"000011111",
  3148=>"101010110",
  3149=>"111001001",
  3150=>"111111011",
  3151=>"110110110",
  3152=>"101000010",
  3153=>"111100100",
  3154=>"100001010",
  3155=>"100101110",
  3156=>"011110001",
  3157=>"001100000",
  3158=>"000101000",
  3159=>"100101101",
  3160=>"001110111",
  3161=>"101011101",
  3162=>"101001010",
  3163=>"111011101",
  3164=>"100101100",
  3165=>"001110110",
  3166=>"100001011",
  3167=>"011010110",
  3168=>"000001101",
  3169=>"011101100",
  3170=>"110000000",
  3171=>"010010110",
  3172=>"100000010",
  3173=>"011000011",
  3174=>"110011010",
  3175=>"110011101",
  3176=>"011001010",
  3177=>"011111110",
  3178=>"100000010",
  3179=>"011011001",
  3180=>"111011110",
  3181=>"011101011",
  3182=>"011000110",
  3183=>"101000000",
  3184=>"101111110",
  3185=>"100001010",
  3186=>"110000111",
  3187=>"110011000",
  3188=>"110000011",
  3189=>"011100110",
  3190=>"100001000",
  3191=>"011100111",
  3192=>"001001110",
  3193=>"011110100",
  3194=>"111010101",
  3195=>"110010010",
  3196=>"011011100",
  3197=>"111000101",
  3198=>"111101111",
  3199=>"000000001",
  3200=>"100001101",
  3201=>"111001010",
  3202=>"010110001",
  3203=>"000010010",
  3204=>"101101111",
  3205=>"001000111",
  3206=>"100100001",
  3207=>"010010100",
  3208=>"011000110",
  3209=>"100100001",
  3210=>"000101001",
  3211=>"100110110",
  3212=>"100000011",
  3213=>"011011010",
  3214=>"001110111",
  3215=>"111010010",
  3216=>"001010110",
  3217=>"000000000",
  3218=>"000011111",
  3219=>"101010111",
  3220=>"001110100",
  3221=>"101011011",
  3222=>"011011110",
  3223=>"101110101",
  3224=>"101000101",
  3225=>"110000101",
  3226=>"100101111",
  3227=>"101110110",
  3228=>"111110110",
  3229=>"010101010",
  3230=>"010111110",
  3231=>"100111000",
  3232=>"000111101",
  3233=>"001000100",
  3234=>"111001001",
  3235=>"000110101",
  3236=>"000001110",
  3237=>"011110101",
  3238=>"011110110",
  3239=>"001011110",
  3240=>"110000011",
  3241=>"101100100",
  3242=>"101000101",
  3243=>"111101001",
  3244=>"001110101",
  3245=>"011001000",
  3246=>"000011110",
  3247=>"101001000",
  3248=>"101101111",
  3249=>"000010110",
  3250=>"111100011",
  3251=>"100011101",
  3252=>"010011000",
  3253=>"010000100",
  3254=>"000000100",
  3255=>"000010101",
  3256=>"010010101",
  3257=>"101010100",
  3258=>"011010010",
  3259=>"111010111",
  3260=>"000000111",
  3261=>"100001011",
  3262=>"111111011",
  3263=>"111010011",
  3264=>"111010110",
  3265=>"100011110",
  3266=>"110001110",
  3267=>"010101110",
  3268=>"001111101",
  3269=>"000010100",
  3270=>"111111011",
  3271=>"111100100",
  3272=>"000011010",
  3273=>"001100100",
  3274=>"001011111",
  3275=>"100110010",
  3276=>"000100011",
  3277=>"011111110",
  3278=>"011011111",
  3279=>"110000011",
  3280=>"110000111",
  3281=>"101111010",
  3282=>"000101001",
  3283=>"111000110",
  3284=>"000010100",
  3285=>"001100000",
  3286=>"101110001",
  3287=>"010011010",
  3288=>"110100110",
  3289=>"101010100",
  3290=>"110011011",
  3291=>"111001000",
  3292=>"001001001",
  3293=>"010011011",
  3294=>"001000000",
  3295=>"001010000",
  3296=>"000100010",
  3297=>"001110101",
  3298=>"000100100",
  3299=>"110100010",
  3300=>"111100101",
  3301=>"001010010",
  3302=>"111101001",
  3303=>"100110000",
  3304=>"000010001",
  3305=>"011110100",
  3306=>"101110110",
  3307=>"111000100",
  3308=>"010101110",
  3309=>"101010010",
  3310=>"001001010",
  3311=>"101000001",
  3312=>"111010100",
  3313=>"100111010",
  3314=>"011010011",
  3315=>"101110010",
  3316=>"110101000",
  3317=>"110011111",
  3318=>"000110010",
  3319=>"110001100",
  3320=>"100100001",
  3321=>"101101111",
  3322=>"111110100",
  3323=>"000011011",
  3324=>"011010010",
  3325=>"001111001",
  3326=>"001111001",
  3327=>"000100110",
  3328=>"110011011",
  3329=>"101110101",
  3330=>"101000101",
  3331=>"000001101",
  3332=>"111001000",
  3333=>"011101110",
  3334=>"010011100",
  3335=>"011000101",
  3336=>"111110111",
  3337=>"000000100",
  3338=>"110111010",
  3339=>"100111111",
  3340=>"011110011",
  3341=>"010001101",
  3342=>"111100000",
  3343=>"000001010",
  3344=>"100010100",
  3345=>"010010001",
  3346=>"101000010",
  3347=>"100110111",
  3348=>"011010011",
  3349=>"010111111",
  3350=>"110111000",
  3351=>"000001111",
  3352=>"011010111",
  3353=>"000110010",
  3354=>"010100001",
  3355=>"101110000",
  3356=>"011011011",
  3357=>"100110101",
  3358=>"001000110",
  3359=>"100100110",
  3360=>"110111100",
  3361=>"000101010",
  3362=>"101111010",
  3363=>"011001010",
  3364=>"111101010",
  3365=>"001010011",
  3366=>"011000001",
  3367=>"001111011",
  3368=>"100011011",
  3369=>"010111111",
  3370=>"001001001",
  3371=>"101001101",
  3372=>"000000000",
  3373=>"000000011",
  3374=>"011101101",
  3375=>"111000110",
  3376=>"110011110",
  3377=>"101001000",
  3378=>"111111110",
  3379=>"100010100",
  3380=>"011100001",
  3381=>"000100001",
  3382=>"011011101",
  3383=>"100010111",
  3384=>"101110000",
  3385=>"100000101",
  3386=>"100000001",
  3387=>"111110101",
  3388=>"110100001",
  3389=>"000000101",
  3390=>"110101010",
  3391=>"001000010",
  3392=>"111000010",
  3393=>"010101101",
  3394=>"110010110",
  3395=>"001110100",
  3396=>"010111110",
  3397=>"101110111",
  3398=>"011010010",
  3399=>"111110101",
  3400=>"101001100",
  3401=>"110001001",
  3402=>"110111000",
  3403=>"000010110",
  3404=>"010100100",
  3405=>"001101000",
  3406=>"110000000",
  3407=>"000011101",
  3408=>"111111111",
  3409=>"110110100",
  3410=>"010000000",
  3411=>"000011011",
  3412=>"110100000",
  3413=>"000100111",
  3414=>"000010000",
  3415=>"000100001",
  3416=>"001111000",
  3417=>"000101001",
  3418=>"011110010",
  3419=>"000011100",
  3420=>"100111111",
  3421=>"110000101",
  3422=>"001111010",
  3423=>"111000101",
  3424=>"010100010",
  3425=>"011011111",
  3426=>"010001000",
  3427=>"110011010",
  3428=>"000101010",
  3429=>"011100101",
  3430=>"100111111",
  3431=>"111001000",
  3432=>"001110101",
  3433=>"101101111",
  3434=>"010010000",
  3435=>"010011000",
  3436=>"101001011",
  3437=>"001111101",
  3438=>"001101011",
  3439=>"000100010",
  3440=>"011100100",
  3441=>"010100111",
  3442=>"111010100",
  3443=>"111011100",
  3444=>"000011001",
  3445=>"101110101",
  3446=>"110000000",
  3447=>"100010111",
  3448=>"000100000",
  3449=>"111110011",
  3450=>"010111111",
  3451=>"000001100",
  3452=>"110000001",
  3453=>"000000111",
  3454=>"111001101",
  3455=>"001000000",
  3456=>"000001110",
  3457=>"001001011",
  3458=>"110101011",
  3459=>"100100011",
  3460=>"011000011",
  3461=>"100100100",
  3462=>"011000110",
  3463=>"011100000",
  3464=>"000111010",
  3465=>"100111110",
  3466=>"011101001",
  3467=>"100010010",
  3468=>"101110100",
  3469=>"111111100",
  3470=>"110111110",
  3471=>"010110000",
  3472=>"101111110",
  3473=>"110101001",
  3474=>"000000000",
  3475=>"111101101",
  3476=>"000111100",
  3477=>"101000011",
  3478=>"101010111",
  3479=>"100010011",
  3480=>"010111101",
  3481=>"111001011",
  3482=>"110100011",
  3483=>"111001100",
  3484=>"101110101",
  3485=>"111111011",
  3486=>"010111000",
  3487=>"110101000",
  3488=>"101001111",
  3489=>"011100111",
  3490=>"111001101",
  3491=>"100000000",
  3492=>"110010110",
  3493=>"001000001",
  3494=>"110111100",
  3495=>"101101100",
  3496=>"111010101",
  3497=>"011011000",
  3498=>"000001001",
  3499=>"000111101",
  3500=>"001111110",
  3501=>"000101010",
  3502=>"010001001",
  3503=>"011001110",
  3504=>"010110011",
  3505=>"110000001",
  3506=>"110010110",
  3507=>"111100110",
  3508=>"011111111",
  3509=>"010001101",
  3510=>"101110011",
  3511=>"000100000",
  3512=>"001001001",
  3513=>"010010101",
  3514=>"110011110",
  3515=>"101101101",
  3516=>"110101101",
  3517=>"110111001",
  3518=>"110010100",
  3519=>"001001101",
  3520=>"000010011",
  3521=>"110110110",
  3522=>"111000011",
  3523=>"100110001",
  3524=>"100000011",
  3525=>"000011000",
  3526=>"001100111",
  3527=>"001000001",
  3528=>"000000111",
  3529=>"011100100",
  3530=>"100001001",
  3531=>"011000100",
  3532=>"100110101",
  3533=>"110001011",
  3534=>"111001111",
  3535=>"000101010",
  3536=>"011001011",
  3537=>"010011000",
  3538=>"110111011",
  3539=>"111010101",
  3540=>"000010111",
  3541=>"001110001",
  3542=>"111111011",
  3543=>"111000101",
  3544=>"111101111",
  3545=>"100111000",
  3546=>"010001110",
  3547=>"100110011",
  3548=>"001101001",
  3549=>"110001001",
  3550=>"010010110",
  3551=>"110001001",
  3552=>"000001000",
  3553=>"110110011",
  3554=>"011000011",
  3555=>"011000000",
  3556=>"010011000",
  3557=>"100011001",
  3558=>"111010011",
  3559=>"000100011",
  3560=>"100010100",
  3561=>"000011101",
  3562=>"001010101",
  3563=>"100000111",
  3564=>"101100011",
  3565=>"011001111",
  3566=>"100001110",
  3567=>"000000000",
  3568=>"000110011",
  3569=>"110011111",
  3570=>"000010010",
  3571=>"010000110",
  3572=>"100010001",
  3573=>"110001110",
  3574=>"100000010",
  3575=>"010111111",
  3576=>"010110010",
  3577=>"111000010",
  3578=>"111100000",
  3579=>"101000101",
  3580=>"101000101",
  3581=>"111111111",
  3582=>"111101001",
  3583=>"010100000",
  3584=>"100000111",
  3585=>"110011100",
  3586=>"001010011",
  3587=>"001000001",
  3588=>"110000001",
  3589=>"011011110",
  3590=>"110000011",
  3591=>"110001111",
  3592=>"110011001",
  3593=>"111010001",
  3594=>"000000001",
  3595=>"110010100",
  3596=>"010100110",
  3597=>"100100000",
  3598=>"101101110",
  3599=>"000010101",
  3600=>"000101010",
  3601=>"000111111",
  3602=>"001010001",
  3603=>"000011001",
  3604=>"000010001",
  3605=>"010011110",
  3606=>"011101100",
  3607=>"001001001",
  3608=>"100001101",
  3609=>"000101001",
  3610=>"000100011",
  3611=>"000110101",
  3612=>"110101110",
  3613=>"101111101",
  3614=>"001011010",
  3615=>"100100110",
  3616=>"110010100",
  3617=>"000010110",
  3618=>"000001100",
  3619=>"001001100",
  3620=>"011000110",
  3621=>"000010100",
  3622=>"111100100",
  3623=>"000111011",
  3624=>"000010000",
  3625=>"100010110",
  3626=>"011101101",
  3627=>"110111001",
  3628=>"111100010",
  3629=>"001111001",
  3630=>"101011111",
  3631=>"111010110",
  3632=>"111100111",
  3633=>"010011011",
  3634=>"110010101",
  3635=>"111100010",
  3636=>"001011110",
  3637=>"010111000",
  3638=>"000001110",
  3639=>"001010010",
  3640=>"001001101",
  3641=>"001110011",
  3642=>"001011011",
  3643=>"100101111",
  3644=>"000010000",
  3645=>"011110001",
  3646=>"111000110",
  3647=>"110101100",
  3648=>"101010100",
  3649=>"000000110",
  3650=>"110101111",
  3651=>"010011010",
  3652=>"110101000",
  3653=>"011111001",
  3654=>"110110001",
  3655=>"011001110",
  3656=>"100110001",
  3657=>"011101001",
  3658=>"001010001",
  3659=>"101110011",
  3660=>"000101100",
  3661=>"000101001",
  3662=>"000100100",
  3663=>"001001001",
  3664=>"000000110",
  3665=>"001101000",
  3666=>"110100110",
  3667=>"100100000",
  3668=>"111100001",
  3669=>"011001111",
  3670=>"010001010",
  3671=>"100110101",
  3672=>"100001001",
  3673=>"101100010",
  3674=>"100010111",
  3675=>"110010100",
  3676=>"101000010",
  3677=>"000100110",
  3678=>"010101111",
  3679=>"011010000",
  3680=>"010110111",
  3681=>"001001000",
  3682=>"001001111",
  3683=>"111110000",
  3684=>"001000001",
  3685=>"011000100",
  3686=>"000111111",
  3687=>"110000111",
  3688=>"110000101",
  3689=>"110110100",
  3690=>"010110110",
  3691=>"110010110",
  3692=>"100010101",
  3693=>"111111001",
  3694=>"000010101",
  3695=>"111110000",
  3696=>"111011110",
  3697=>"000001100",
  3698=>"110100000",
  3699=>"000100000",
  3700=>"110111010",
  3701=>"100001110",
  3702=>"011000010",
  3703=>"000110111",
  3704=>"100100111",
  3705=>"000110111",
  3706=>"101001101",
  3707=>"101110000",
  3708=>"100011000",
  3709=>"101001100",
  3710=>"111110010",
  3711=>"011101100",
  3712=>"010010000",
  3713=>"001110001",
  3714=>"100110000",
  3715=>"011101101",
  3716=>"110001110",
  3717=>"101110001",
  3718=>"011111001",
  3719=>"010111011",
  3720=>"011101100",
  3721=>"101000110",
  3722=>"111110101",
  3723=>"100100000",
  3724=>"111100110",
  3725=>"101010011",
  3726=>"111001111",
  3727=>"100011010",
  3728=>"001100000",
  3729=>"110101011",
  3730=>"111111111",
  3731=>"100001110",
  3732=>"001010011",
  3733=>"011010011",
  3734=>"001001000",
  3735=>"011011101",
  3736=>"011011100",
  3737=>"001000110",
  3738=>"100001110",
  3739=>"110110000",
  3740=>"100001011",
  3741=>"011111010",
  3742=>"101100000",
  3743=>"000111100",
  3744=>"001000110",
  3745=>"100010111",
  3746=>"000110100",
  3747=>"101111010",
  3748=>"110010111",
  3749=>"111001111",
  3750=>"100011110",
  3751=>"011010010",
  3752=>"111101111",
  3753=>"000100000",
  3754=>"101111100",
  3755=>"000011111",
  3756=>"100000000",
  3757=>"010000000",
  3758=>"011111011",
  3759=>"111111110",
  3760=>"000100111",
  3761=>"001011101",
  3762=>"101000110",
  3763=>"111101000",
  3764=>"001101110",
  3765=>"111110000",
  3766=>"111110000",
  3767=>"001111011",
  3768=>"011101011",
  3769=>"010001001",
  3770=>"011101010",
  3771=>"101110001",
  3772=>"011110001",
  3773=>"110011010",
  3774=>"101100101",
  3775=>"000101001",
  3776=>"111001011",
  3777=>"010011000",
  3778=>"000011010",
  3779=>"010100000",
  3780=>"010011010",
  3781=>"001010101",
  3782=>"000110011",
  3783=>"111000101",
  3784=>"101110111",
  3785=>"010001110",
  3786=>"111011101",
  3787=>"011100101",
  3788=>"100110110",
  3789=>"110100111",
  3790=>"011111110",
  3791=>"111110001",
  3792=>"001000110",
  3793=>"100011101",
  3794=>"010111110",
  3795=>"001110000",
  3796=>"010101010",
  3797=>"110010000",
  3798=>"100100111",
  3799=>"101100100",
  3800=>"000100011",
  3801=>"100111111",
  3802=>"011011100",
  3803=>"000101111",
  3804=>"001111000",
  3805=>"100011110",
  3806=>"101100000",
  3807=>"000100010",
  3808=>"011100111",
  3809=>"110010111",
  3810=>"110010010",
  3811=>"110110111",
  3812=>"100010101",
  3813=>"110110110",
  3814=>"110000001",
  3815=>"010110010",
  3816=>"011000101",
  3817=>"100010001",
  3818=>"001100001",
  3819=>"001110011",
  3820=>"100000100",
  3821=>"000100011",
  3822=>"101110101",
  3823=>"010000010",
  3824=>"001001101",
  3825=>"011111110",
  3826=>"111010011",
  3827=>"110000111",
  3828=>"100100001",
  3829=>"011010011",
  3830=>"111001010",
  3831=>"110100111",
  3832=>"011011101",
  3833=>"110110000",
  3834=>"000011000",
  3835=>"101001011",
  3836=>"000100001",
  3837=>"000011101",
  3838=>"011100111",
  3839=>"010011101",
  3840=>"111110100",
  3841=>"110000000",
  3842=>"011111001",
  3843=>"000111010",
  3844=>"100110000",
  3845=>"001110000",
  3846=>"000110100",
  3847=>"001000110",
  3848=>"110000101",
  3849=>"010010000",
  3850=>"100001111",
  3851=>"000001001",
  3852=>"000101001",
  3853=>"110100100",
  3854=>"101000010",
  3855=>"001000000",
  3856=>"101011111",
  3857=>"110000011",
  3858=>"000110001",
  3859=>"111001010",
  3860=>"000010100",
  3861=>"100010100",
  3862=>"010110110",
  3863=>"111000010",
  3864=>"100001010",
  3865=>"111111110",
  3866=>"101001001",
  3867=>"001110100",
  3868=>"010001011",
  3869=>"110101110",
  3870=>"011001011",
  3871=>"010111101",
  3872=>"000100011",
  3873=>"110000101",
  3874=>"101110101",
  3875=>"000111011",
  3876=>"011111110",
  3877=>"011100111",
  3878=>"100100100",
  3879=>"000001110",
  3880=>"010001100",
  3881=>"000100000",
  3882=>"100111011",
  3883=>"001111011",
  3884=>"111111110",
  3885=>"000010001",
  3886=>"011110111",
  3887=>"010010011",
  3888=>"101011001",
  3889=>"111110010",
  3890=>"001110001",
  3891=>"011111111",
  3892=>"001010000",
  3893=>"111110111",
  3894=>"011001100",
  3895=>"010011101",
  3896=>"011011111",
  3897=>"000000000",
  3898=>"111000101",
  3899=>"000100011",
  3900=>"110000101",
  3901=>"001101001",
  3902=>"000000010",
  3903=>"101001011",
  3904=>"111110100",
  3905=>"011001010",
  3906=>"001110100",
  3907=>"111011001",
  3908=>"011101101",
  3909=>"001111011",
  3910=>"101110110",
  3911=>"010100111",
  3912=>"111110100",
  3913=>"010001100",
  3914=>"010100100",
  3915=>"010100010",
  3916=>"101110011",
  3917=>"011111100",
  3918=>"100000001",
  3919=>"111100001",
  3920=>"101010011",
  3921=>"101101011",
  3922=>"000001011",
  3923=>"001010001",
  3924=>"100111111",
  3925=>"110110100",
  3926=>"000000000",
  3927=>"110100110",
  3928=>"000001101",
  3929=>"101011101",
  3930=>"001001111",
  3931=>"000101110",
  3932=>"010111000",
  3933=>"011111101",
  3934=>"011110100",
  3935=>"110110101",
  3936=>"111101010",
  3937=>"011010111",
  3938=>"001000100",
  3939=>"101011001",
  3940=>"111011111",
  3941=>"000000010",
  3942=>"110101111",
  3943=>"000101110",
  3944=>"111010101",
  3945=>"010010100",
  3946=>"100101011",
  3947=>"110001000",
  3948=>"011100110",
  3949=>"101001101",
  3950=>"000001000",
  3951=>"000110001",
  3952=>"100100001",
  3953=>"101100110",
  3954=>"101000111",
  3955=>"001110110",
  3956=>"011011100",
  3957=>"000110010",
  3958=>"010110101",
  3959=>"101011111",
  3960=>"111011001",
  3961=>"011110111",
  3962=>"110111010",
  3963=>"100001011",
  3964=>"101110000",
  3965=>"011010011",
  3966=>"000000010",
  3967=>"010110000",
  3968=>"110110100",
  3969=>"101110010",
  3970=>"001100001",
  3971=>"010111010",
  3972=>"000100010",
  3973=>"100101000",
  3974=>"000010001",
  3975=>"011000010",
  3976=>"000101011",
  3977=>"110000110",
  3978=>"101101001",
  3979=>"111110111",
  3980=>"111111110",
  3981=>"001110101",
  3982=>"111001101",
  3983=>"010011000",
  3984=>"110010111",
  3985=>"100000011",
  3986=>"111011100",
  3987=>"101100101",
  3988=>"000100011",
  3989=>"010100111",
  3990=>"001110011",
  3991=>"001000000",
  3992=>"111100001",
  3993=>"011101100",
  3994=>"011110111",
  3995=>"100101110",
  3996=>"010011110",
  3997=>"000111100",
  3998=>"110111011",
  3999=>"000001010",
  4000=>"010101110",
  4001=>"111011000",
  4002=>"011111010",
  4003=>"110011110",
  4004=>"100101000",
  4005=>"110011111",
  4006=>"110011001",
  4007=>"000000001",
  4008=>"011011110",
  4009=>"000100001",
  4010=>"011100011",
  4011=>"101100011",
  4012=>"100111111",
  4013=>"110001011",
  4014=>"000011010",
  4015=>"011011101",
  4016=>"001001111",
  4017=>"011011111",
  4018=>"000011100",
  4019=>"110101000",
  4020=>"010101001",
  4021=>"110101111",
  4022=>"111110100",
  4023=>"111110000",
  4024=>"111111001",
  4025=>"110001010",
  4026=>"100100001",
  4027=>"100001110",
  4028=>"000001100",
  4029=>"101110010",
  4030=>"010000000",
  4031=>"101110001",
  4032=>"000000000",
  4033=>"011101000",
  4034=>"010111111",
  4035=>"001010111",
  4036=>"011001011",
  4037=>"001011110",
  4038=>"101100010",
  4039=>"100110110",
  4040=>"000100101",
  4041=>"010011001",
  4042=>"110001001",
  4043=>"010010110",
  4044=>"101111101",
  4045=>"111100101",
  4046=>"110010100",
  4047=>"101000111",
  4048=>"001100001",
  4049=>"000111001",
  4050=>"011110000",
  4051=>"100011001",
  4052=>"010001101",
  4053=>"101101011",
  4054=>"111000111",
  4055=>"011000110",
  4056=>"010111101",
  4057=>"011000101",
  4058=>"111100000",
  4059=>"001100000",
  4060=>"110101100",
  4061=>"001101001",
  4062=>"100001100",
  4063=>"011001100",
  4064=>"110101000",
  4065=>"001011100",
  4066=>"000101000",
  4067=>"100110000",
  4068=>"001001101",
  4069=>"011001010",
  4070=>"101101011",
  4071=>"000010010",
  4072=>"010100111",
  4073=>"110010110",
  4074=>"110011000",
  4075=>"010111111",
  4076=>"111011010",
  4077=>"111100000",
  4078=>"101010000",
  4079=>"110111111",
  4080=>"000011111",
  4081=>"000111001",
  4082=>"101101110",
  4083=>"100000110",
  4084=>"011100011",
  4085=>"110000100",
  4086=>"010010011",
  4087=>"101100101",
  4088=>"000100101",
  4089=>"101001010",
  4090=>"111110000",
  4091=>"100011111",
  4092=>"111001000",
  4093=>"101101110",
  4094=>"101111001",
  4095=>"111001010",
  4096=>"011000000",
  4097=>"000010010",
  4098=>"000101010",
  4099=>"010000111",
  4100=>"000000110",
  4101=>"110110110",
  4102=>"101001010",
  4103=>"011010000",
  4104=>"001101100",
  4105=>"000101110",
  4106=>"010101111",
  4107=>"110010001",
  4108=>"100011111",
  4109=>"000011010",
  4110=>"001101110",
  4111=>"011110001",
  4112=>"111101111",
  4113=>"001110001",
  4114=>"000100110",
  4115=>"110000010",
  4116=>"011110010",
  4117=>"101010101",
  4118=>"100111010",
  4119=>"010000110",
  4120=>"101110101",
  4121=>"101010011",
  4122=>"100011001",
  4123=>"111111101",
  4124=>"100111101",
  4125=>"100101000",
  4126=>"101110011",
  4127=>"010000010",
  4128=>"000100111",
  4129=>"010010000",
  4130=>"111011011",
  4131=>"101000010",
  4132=>"101011001",
  4133=>"100101101",
  4134=>"001001001",
  4135=>"101000011",
  4136=>"101010010",
  4137=>"011100010",
  4138=>"100101001",
  4139=>"100011010",
  4140=>"010001011",
  4141=>"110101111",
  4142=>"011101001",
  4143=>"110000000",
  4144=>"100001111",
  4145=>"001100100",
  4146=>"010001110",
  4147=>"000101111",
  4148=>"001101010",
  4149=>"000110100",
  4150=>"101110001",
  4151=>"110101001",
  4152=>"000000110",
  4153=>"100001000",
  4154=>"000110001",
  4155=>"110010000",
  4156=>"011000111",
  4157=>"011101001",
  4158=>"110000101",
  4159=>"010111111",
  4160=>"111101011",
  4161=>"000110001",
  4162=>"000101010",
  4163=>"000101011",
  4164=>"111010010",
  4165=>"110010111",
  4166=>"010011101",
  4167=>"110110100",
  4168=>"011011110",
  4169=>"101110110",
  4170=>"101000110",
  4171=>"000111110",
  4172=>"010011000",
  4173=>"111111110",
  4174=>"100101000",
  4175=>"011100111",
  4176=>"011101001",
  4177=>"011000000",
  4178=>"001101011",
  4179=>"000111000",
  4180=>"110011000",
  4181=>"010111001",
  4182=>"101010101",
  4183=>"001001111",
  4184=>"110001110",
  4185=>"011000111",
  4186=>"101110111",
  4187=>"100101100",
  4188=>"111000101",
  4189=>"111101101",
  4190=>"101101011",
  4191=>"110110010",
  4192=>"010111000",
  4193=>"010010110",
  4194=>"000010001",
  4195=>"101100101",
  4196=>"111010011",
  4197=>"100011110",
  4198=>"100101010",
  4199=>"011101001",
  4200=>"110011110",
  4201=>"000100010",
  4202=>"010011010",
  4203=>"011000010",
  4204=>"011000011",
  4205=>"101000100",
  4206=>"000111011",
  4207=>"100101111",
  4208=>"011000101",
  4209=>"010101100",
  4210=>"111000000",
  4211=>"001011010",
  4212=>"111110101",
  4213=>"011000010",
  4214=>"011000011",
  4215=>"000100001",
  4216=>"101001110",
  4217=>"110000111",
  4218=>"100101001",
  4219=>"001100101",
  4220=>"111111011",
  4221=>"101000110",
  4222=>"010011010",
  4223=>"101110100",
  4224=>"001100111",
  4225=>"001111101",
  4226=>"101001011",
  4227=>"111110110",
  4228=>"010010111",
  4229=>"100101001",
  4230=>"011101101",
  4231=>"101010000",
  4232=>"100101110",
  4233=>"101100011",
  4234=>"000010101",
  4235=>"110000101",
  4236=>"100110001",
  4237=>"011011011",
  4238=>"111111111",
  4239=>"101010101",
  4240=>"010000111",
  4241=>"011010010",
  4242=>"110100110",
  4243=>"111110110",
  4244=>"101110001",
  4245=>"001111100",
  4246=>"011000011",
  4247=>"111110001",
  4248=>"111000111",
  4249=>"110011110",
  4250=>"111101100",
  4251=>"111101111",
  4252=>"111110010",
  4253=>"110010011",
  4254=>"100000011",
  4255=>"111110010",
  4256=>"000001111",
  4257=>"010010010",
  4258=>"110010001",
  4259=>"000011000",
  4260=>"011101100",
  4261=>"011101110",
  4262=>"000101100",
  4263=>"011110000",
  4264=>"001011001",
  4265=>"101001111",
  4266=>"010100000",
  4267=>"111111101",
  4268=>"101101001",
  4269=>"011001101",
  4270=>"101100000",
  4271=>"001000000",
  4272=>"111111111",
  4273=>"000110100",
  4274=>"010010001",
  4275=>"000101101",
  4276=>"001000000",
  4277=>"111100111",
  4278=>"000000001",
  4279=>"010000100",
  4280=>"011011111",
  4281=>"001011011",
  4282=>"100000100",
  4283=>"100000101",
  4284=>"000001100",
  4285=>"110100011",
  4286=>"010001010",
  4287=>"000001010",
  4288=>"000100101",
  4289=>"001010000",
  4290=>"001000111",
  4291=>"101101000",
  4292=>"010001100",
  4293=>"110000001",
  4294=>"100111111",
  4295=>"010100110",
  4296=>"101111101",
  4297=>"001110011",
  4298=>"111000111",
  4299=>"110110101",
  4300=>"001101101",
  4301=>"111100010",
  4302=>"001010001",
  4303=>"100000011",
  4304=>"010111001",
  4305=>"000110110",
  4306=>"011111100",
  4307=>"000001000",
  4308=>"110010001",
  4309=>"100100101",
  4310=>"000000001",
  4311=>"010100100",
  4312=>"010111011",
  4313=>"000010111",
  4314=>"100111111",
  4315=>"010010101",
  4316=>"010000000",
  4317=>"111111110",
  4318=>"110111101",
  4319=>"000100110",
  4320=>"000101101",
  4321=>"100011001",
  4322=>"000000001",
  4323=>"101000111",
  4324=>"111111010",
  4325=>"110001110",
  4326=>"000110010",
  4327=>"110001110",
  4328=>"101101110",
  4329=>"011011111",
  4330=>"000110110",
  4331=>"000111111",
  4332=>"100111101",
  4333=>"010000111",
  4334=>"111010010",
  4335=>"110000001",
  4336=>"010001110",
  4337=>"101100100",
  4338=>"101000001",
  4339=>"011011011",
  4340=>"011001001",
  4341=>"010001000",
  4342=>"110001011",
  4343=>"111100110",
  4344=>"110110101",
  4345=>"101110000",
  4346=>"001111100",
  4347=>"101011101",
  4348=>"011100011",
  4349=>"001101011",
  4350=>"010000000",
  4351=>"101100100",
  4352=>"100010000",
  4353=>"011101000",
  4354=>"010111101",
  4355=>"011010110",
  4356=>"001001001",
  4357=>"100011111",
  4358=>"011101100",
  4359=>"000100001",
  4360=>"010101010",
  4361=>"100000000",
  4362=>"001111101",
  4363=>"001110011",
  4364=>"110011101",
  4365=>"001011000",
  4366=>"011010110",
  4367=>"001110000",
  4368=>"111110101",
  4369=>"111011111",
  4370=>"110010100",
  4371=>"110110100",
  4372=>"111110110",
  4373=>"000101100",
  4374=>"101011111",
  4375=>"100001111",
  4376=>"001001000",
  4377=>"110010011",
  4378=>"001101101",
  4379=>"101011010",
  4380=>"110110001",
  4381=>"011000010",
  4382=>"110110011",
  4383=>"111111111",
  4384=>"110101011",
  4385=>"111001000",
  4386=>"110110011",
  4387=>"101000111",
  4388=>"000000000",
  4389=>"111011001",
  4390=>"100100010",
  4391=>"100111111",
  4392=>"010100011",
  4393=>"000111110",
  4394=>"111001110",
  4395=>"011010001",
  4396=>"000001100",
  4397=>"010110000",
  4398=>"110000100",
  4399=>"010000101",
  4400=>"011000100",
  4401=>"000100000",
  4402=>"000100101",
  4403=>"000000011",
  4404=>"101111000",
  4405=>"001011111",
  4406=>"000100110",
  4407=>"100111010",
  4408=>"111111111",
  4409=>"111110010",
  4410=>"010000000",
  4411=>"101110010",
  4412=>"010101001",
  4413=>"100010011",
  4414=>"101011111",
  4415=>"001001010",
  4416=>"000111010",
  4417=>"000100000",
  4418=>"011100000",
  4419=>"010011111",
  4420=>"010001111",
  4421=>"001011001",
  4422=>"011111100",
  4423=>"111111001",
  4424=>"111100001",
  4425=>"011110101",
  4426=>"010111010",
  4427=>"001000110",
  4428=>"000101110",
  4429=>"001000001",
  4430=>"101011111",
  4431=>"011111111",
  4432=>"011111010",
  4433=>"100011011",
  4434=>"010110111",
  4435=>"011100000",
  4436=>"010100011",
  4437=>"111001110",
  4438=>"100110100",
  4439=>"110010000",
  4440=>"000000010",
  4441=>"110010001",
  4442=>"010111011",
  4443=>"001100110",
  4444=>"100111110",
  4445=>"001010000",
  4446=>"001111100",
  4447=>"110010111",
  4448=>"111010101",
  4449=>"010011000",
  4450=>"011011000",
  4451=>"011000010",
  4452=>"010011001",
  4453=>"101011101",
  4454=>"001101100",
  4455=>"111110110",
  4456=>"010110101",
  4457=>"101010000",
  4458=>"111100110",
  4459=>"001001101",
  4460=>"111101100",
  4461=>"010001000",
  4462=>"100100001",
  4463=>"001111111",
  4464=>"000101111",
  4465=>"101111101",
  4466=>"010100110",
  4467=>"001000110",
  4468=>"111101000",
  4469=>"110111010",
  4470=>"101110110",
  4471=>"100011010",
  4472=>"110111111",
  4473=>"010101001",
  4474=>"000111100",
  4475=>"100101111",
  4476=>"101011101",
  4477=>"111010011",
  4478=>"000100110",
  4479=>"111111000",
  4480=>"110101111",
  4481=>"010001111",
  4482=>"110001101",
  4483=>"001101011",
  4484=>"110100010",
  4485=>"101101001",
  4486=>"100011011",
  4487=>"001000000",
  4488=>"100100011",
  4489=>"010010001",
  4490=>"100011000",
  4491=>"111101110",
  4492=>"001101011",
  4493=>"011110001",
  4494=>"001100011",
  4495=>"010010011",
  4496=>"111000001",
  4497=>"010101111",
  4498=>"000000010",
  4499=>"111111011",
  4500=>"111110111",
  4501=>"010011000",
  4502=>"000101100",
  4503=>"110110000",
  4504=>"001100001",
  4505=>"011000101",
  4506=>"111100010",
  4507=>"010001001",
  4508=>"110010000",
  4509=>"101110100",
  4510=>"110010000",
  4511=>"011100011",
  4512=>"000000011",
  4513=>"000001001",
  4514=>"110011111",
  4515=>"010010000",
  4516=>"010001000",
  4517=>"001100000",
  4518=>"100010100",
  4519=>"001100100",
  4520=>"011100101",
  4521=>"001110000",
  4522=>"010110111",
  4523=>"101011011",
  4524=>"001001111",
  4525=>"101111101",
  4526=>"010000100",
  4527=>"001101110",
  4528=>"101011000",
  4529=>"101110110",
  4530=>"101111111",
  4531=>"000111100",
  4532=>"111011111",
  4533=>"110001100",
  4534=>"100110110",
  4535=>"000111000",
  4536=>"010000101",
  4537=>"100010001",
  4538=>"011101111",
  4539=>"111101010",
  4540=>"110010001",
  4541=>"110111000",
  4542=>"111001100",
  4543=>"001011000",
  4544=>"111100110",
  4545=>"111010010",
  4546=>"011011100",
  4547=>"100101111",
  4548=>"111010110",
  4549=>"110111001",
  4550=>"100110010",
  4551=>"100100001",
  4552=>"111000000",
  4553=>"111101100",
  4554=>"010000111",
  4555=>"111101000",
  4556=>"010101000",
  4557=>"010010001",
  4558=>"111000000",
  4559=>"101010001",
  4560=>"011011101",
  4561=>"011111000",
  4562=>"110011110",
  4563=>"101001010",
  4564=>"001100100",
  4565=>"001000000",
  4566=>"101110101",
  4567=>"000101000",
  4568=>"110111100",
  4569=>"010101101",
  4570=>"001100010",
  4571=>"100111011",
  4572=>"001011100",
  4573=>"101111010",
  4574=>"000110111",
  4575=>"110111100",
  4576=>"110111100",
  4577=>"110110100",
  4578=>"000101011",
  4579=>"101011111",
  4580=>"101011110",
  4581=>"000011001",
  4582=>"011010010",
  4583=>"001100100",
  4584=>"001000111",
  4585=>"000000111",
  4586=>"111011100",
  4587=>"001011110",
  4588=>"001111011",
  4589=>"010010110",
  4590=>"111111000",
  4591=>"111110011",
  4592=>"011101000",
  4593=>"001000110",
  4594=>"110010000",
  4595=>"110011010",
  4596=>"111111100",
  4597=>"000110001",
  4598=>"100111011",
  4599=>"001010110",
  4600=>"000000000",
  4601=>"000010010",
  4602=>"001000101",
  4603=>"010111101",
  4604=>"000110110",
  4605=>"100110000",
  4606=>"000000110",
  4607=>"011001010",
  4608=>"111001011",
  4609=>"001111000",
  4610=>"110110000",
  4611=>"000100001",
  4612=>"000010010",
  4613=>"100011001",
  4614=>"111100000",
  4615=>"001000110",
  4616=>"100000000",
  4617=>"001011111",
  4618=>"101110111",
  4619=>"000100100",
  4620=>"011010111",
  4621=>"111001010",
  4622=>"000110011",
  4623=>"100001111",
  4624=>"101111101",
  4625=>"110010000",
  4626=>"110101100",
  4627=>"101000100",
  4628=>"111011001",
  4629=>"011110100",
  4630=>"000111001",
  4631=>"111001111",
  4632=>"011001010",
  4633=>"010011111",
  4634=>"001001000",
  4635=>"110000010",
  4636=>"011000110",
  4637=>"001010000",
  4638=>"101100010",
  4639=>"111111100",
  4640=>"001000000",
  4641=>"110100101",
  4642=>"001010010",
  4643=>"010000110",
  4644=>"111101000",
  4645=>"000110000",
  4646=>"000010110",
  4647=>"110001101",
  4648=>"101110111",
  4649=>"101100011",
  4650=>"001100000",
  4651=>"111010000",
  4652=>"101011001",
  4653=>"010001011",
  4654=>"010110001",
  4655=>"110100000",
  4656=>"111101111",
  4657=>"110010111",
  4658=>"110101001",
  4659=>"101110101",
  4660=>"000111001",
  4661=>"001001011",
  4662=>"101011011",
  4663=>"000111001",
  4664=>"001110010",
  4665=>"110010110",
  4666=>"111000101",
  4667=>"111011011",
  4668=>"010000011",
  4669=>"111100010",
  4670=>"111100001",
  4671=>"100111110",
  4672=>"000101110",
  4673=>"000100010",
  4674=>"001000000",
  4675=>"000001101",
  4676=>"101010110",
  4677=>"010100110",
  4678=>"111000111",
  4679=>"010011111",
  4680=>"100010000",
  4681=>"001111111",
  4682=>"010010101",
  4683=>"000100100",
  4684=>"110000010",
  4685=>"111111001",
  4686=>"011011000",
  4687=>"011001100",
  4688=>"000001001",
  4689=>"111001100",
  4690=>"111110010",
  4691=>"101111110",
  4692=>"111100110",
  4693=>"000010000",
  4694=>"011010101",
  4695=>"000000111",
  4696=>"010111111",
  4697=>"010011000",
  4698=>"111000010",
  4699=>"110011100",
  4700=>"010101101",
  4701=>"100100111",
  4702=>"010100001",
  4703=>"001001000",
  4704=>"010001010",
  4705=>"001100001",
  4706=>"101101111",
  4707=>"011101100",
  4708=>"101100100",
  4709=>"011011111",
  4710=>"000000100",
  4711=>"010001100",
  4712=>"010000001",
  4713=>"111101001",
  4714=>"101010111",
  4715=>"000011010",
  4716=>"000000000",
  4717=>"011100000",
  4718=>"010011001",
  4719=>"001010101",
  4720=>"101010100",
  4721=>"101110110",
  4722=>"000101111",
  4723=>"101000100",
  4724=>"000100011",
  4725=>"111101010",
  4726=>"111100000",
  4727=>"101101100",
  4728=>"000001001",
  4729=>"101100100",
  4730=>"111010101",
  4731=>"110111100",
  4732=>"100000110",
  4733=>"111011000",
  4734=>"001011000",
  4735=>"011001001",
  4736=>"101111100",
  4737=>"001111100",
  4738=>"010110010",
  4739=>"000011011",
  4740=>"111100010",
  4741=>"000000100",
  4742=>"100010111",
  4743=>"010111100",
  4744=>"011010011",
  4745=>"111100101",
  4746=>"001100001",
  4747=>"001001100",
  4748=>"110000101",
  4749=>"011111011",
  4750=>"011111110",
  4751=>"011000110",
  4752=>"010010111",
  4753=>"111110010",
  4754=>"011101010",
  4755=>"100101101",
  4756=>"010011001",
  4757=>"011101111",
  4758=>"000010010",
  4759=>"000110101",
  4760=>"100110100",
  4761=>"010110010",
  4762=>"101000011",
  4763=>"010011001",
  4764=>"001100000",
  4765=>"000111011",
  4766=>"000100110",
  4767=>"101011010",
  4768=>"110000010",
  4769=>"100100011",
  4770=>"111100011",
  4771=>"011001111",
  4772=>"101010000",
  4773=>"111010001",
  4774=>"011010101",
  4775=>"111101111",
  4776=>"010001010",
  4777=>"110101011",
  4778=>"011000100",
  4779=>"100011010",
  4780=>"111011001",
  4781=>"000111001",
  4782=>"010101000",
  4783=>"011001110",
  4784=>"111011100",
  4785=>"110100111",
  4786=>"100101110",
  4787=>"001101000",
  4788=>"100001110",
  4789=>"110000111",
  4790=>"010100100",
  4791=>"111010010",
  4792=>"011010100",
  4793=>"110101001",
  4794=>"000011110",
  4795=>"001000110",
  4796=>"000001010",
  4797=>"010010000",
  4798=>"101000101",
  4799=>"000001111",
  4800=>"101100100",
  4801=>"000000010",
  4802=>"001101010",
  4803=>"101001111",
  4804=>"010000000",
  4805=>"011101010",
  4806=>"011110000",
  4807=>"000000010",
  4808=>"110000000",
  4809=>"010000001",
  4810=>"111011100",
  4811=>"111101000",
  4812=>"101000010",
  4813=>"111111001",
  4814=>"011010101",
  4815=>"010110010",
  4816=>"001011000",
  4817=>"101010111",
  4818=>"010101101",
  4819=>"101000011",
  4820=>"100111010",
  4821=>"110000010",
  4822=>"111000100",
  4823=>"100100110",
  4824=>"001101011",
  4825=>"001110101",
  4826=>"110011011",
  4827=>"111101100",
  4828=>"100101101",
  4829=>"111011010",
  4830=>"011100111",
  4831=>"111111100",
  4832=>"111011100",
  4833=>"011110111",
  4834=>"110110011",
  4835=>"101001100",
  4836=>"111010010",
  4837=>"010110000",
  4838=>"000100100",
  4839=>"111110010",
  4840=>"001101101",
  4841=>"001110111",
  4842=>"111101111",
  4843=>"100001110",
  4844=>"111001001",
  4845=>"110001001",
  4846=>"111100010",
  4847=>"110010010",
  4848=>"010100111",
  4849=>"101100000",
  4850=>"101000001",
  4851=>"000110011",
  4852=>"000001010",
  4853=>"100100101",
  4854=>"111100011",
  4855=>"100011011",
  4856=>"001110000",
  4857=>"110011111",
  4858=>"111010111",
  4859=>"111101010",
  4860=>"010000101",
  4861=>"110110000",
  4862=>"111010000",
  4863=>"001011001",
  4864=>"010010001",
  4865=>"010000011",
  4866=>"111101111",
  4867=>"000000100",
  4868=>"111110111",
  4869=>"010100110",
  4870=>"001110110",
  4871=>"011111001",
  4872=>"001101111",
  4873=>"001010111",
  4874=>"000100001",
  4875=>"100100000",
  4876=>"000000011",
  4877=>"110011101",
  4878=>"010000001",
  4879=>"111110100",
  4880=>"001010011",
  4881=>"101110111",
  4882=>"001110110",
  4883=>"100011011",
  4884=>"001011010",
  4885=>"111011000",
  4886=>"100101010",
  4887=>"010110110",
  4888=>"001100010",
  4889=>"001111110",
  4890=>"101100000",
  4891=>"010000111",
  4892=>"001000110",
  4893=>"110100101",
  4894=>"000010110",
  4895=>"110111101",
  4896=>"100000001",
  4897=>"001100011",
  4898=>"111000000",
  4899=>"110011010",
  4900=>"011100110",
  4901=>"010100000",
  4902=>"111110000",
  4903=>"000101001",
  4904=>"101100001",
  4905=>"110010111",
  4906=>"011111101",
  4907=>"011001010",
  4908=>"111000010",
  4909=>"011011000",
  4910=>"111000010",
  4911=>"111010100",
  4912=>"000101110",
  4913=>"010110011",
  4914=>"111010001",
  4915=>"001001100",
  4916=>"011001110",
  4917=>"001011101",
  4918=>"000101110",
  4919=>"110010000",
  4920=>"111100001",
  4921=>"010111010",
  4922=>"010011010",
  4923=>"000110001",
  4924=>"101101111",
  4925=>"000100010",
  4926=>"100110100",
  4927=>"110011001",
  4928=>"111110011",
  4929=>"110111110",
  4930=>"111101110",
  4931=>"010100101",
  4932=>"100111000",
  4933=>"110010011",
  4934=>"100001101",
  4935=>"011111001",
  4936=>"101001100",
  4937=>"100100111",
  4938=>"100010100",
  4939=>"101000100",
  4940=>"111011000",
  4941=>"111110111",
  4942=>"111100000",
  4943=>"001100000",
  4944=>"010010010",
  4945=>"000011100",
  4946=>"011001110",
  4947=>"010001101",
  4948=>"011001001",
  4949=>"110100110",
  4950=>"110110100",
  4951=>"101100001",
  4952=>"100100101",
  4953=>"110001011",
  4954=>"010110001",
  4955=>"101000010",
  4956=>"111000111",
  4957=>"001000011",
  4958=>"100010010",
  4959=>"111000101",
  4960=>"011101010",
  4961=>"100100110",
  4962=>"001011010",
  4963=>"100100000",
  4964=>"010001001",
  4965=>"110110100",
  4966=>"001001110",
  4967=>"101001010",
  4968=>"100000101",
  4969=>"010010001",
  4970=>"010001110",
  4971=>"100010010",
  4972=>"100011001",
  4973=>"101001111",
  4974=>"001001001",
  4975=>"110000000",
  4976=>"010000110",
  4977=>"100011001",
  4978=>"110010010",
  4979=>"101111010",
  4980=>"000110100",
  4981=>"111000000",
  4982=>"111000001",
  4983=>"001011111",
  4984=>"100110111",
  4985=>"001001010",
  4986=>"001001011",
  4987=>"011010001",
  4988=>"101000001",
  4989=>"101011110",
  4990=>"101011011",
  4991=>"101011111",
  4992=>"111110111",
  4993=>"001010111",
  4994=>"001001001",
  4995=>"010111000",
  4996=>"111110000",
  4997=>"000100000",
  4998=>"111101111",
  4999=>"000101101",
  5000=>"010110111",
  5001=>"110000111",
  5002=>"111110010",
  5003=>"011010010",
  5004=>"110111101",
  5005=>"010011111",
  5006=>"110001110",
  5007=>"001000000",
  5008=>"100011100",
  5009=>"110011111",
  5010=>"001110100",
  5011=>"101100101",
  5012=>"100011010",
  5013=>"001010011",
  5014=>"001011001",
  5015=>"000110011",
  5016=>"011011000",
  5017=>"001010111",
  5018=>"010000010",
  5019=>"101000010",
  5020=>"110001000",
  5021=>"001001111",
  5022=>"001010101",
  5023=>"000110100",
  5024=>"000110101",
  5025=>"110111000",
  5026=>"110001010",
  5027=>"111110011",
  5028=>"000010101",
  5029=>"011101010",
  5030=>"000011100",
  5031=>"101110000",
  5032=>"011101110",
  5033=>"101111111",
  5034=>"101100100",
  5035=>"000100000",
  5036=>"000010010",
  5037=>"111010010",
  5038=>"110110001",
  5039=>"011111001",
  5040=>"101000111",
  5041=>"111011101",
  5042=>"101011011",
  5043=>"101100001",
  5044=>"010011110",
  5045=>"100011000",
  5046=>"110001011",
  5047=>"111001000",
  5048=>"000110100",
  5049=>"101011000",
  5050=>"101011001",
  5051=>"100001011",
  5052=>"011001100",
  5053=>"110011001",
  5054=>"001000000",
  5055=>"101010110",
  5056=>"011111110",
  5057=>"010001101",
  5058=>"101010111",
  5059=>"011101100",
  5060=>"011111011",
  5061=>"110010001",
  5062=>"111011111",
  5063=>"001011011",
  5064=>"000100001",
  5065=>"101011010",
  5066=>"110000010",
  5067=>"110101000",
  5068=>"001001010",
  5069=>"100110100",
  5070=>"001001110",
  5071=>"100111010",
  5072=>"101011111",
  5073=>"110000000",
  5074=>"111001111",
  5075=>"010010000",
  5076=>"001011001",
  5077=>"101000001",
  5078=>"010001110",
  5079=>"001001111",
  5080=>"111101100",
  5081=>"011110101",
  5082=>"111101010",
  5083=>"001110110",
  5084=>"000001100",
  5085=>"111111001",
  5086=>"000011101",
  5087=>"110101010",
  5088=>"001111010",
  5089=>"011110001",
  5090=>"111110100",
  5091=>"111010111",
  5092=>"010010110",
  5093=>"010011000",
  5094=>"100110011",
  5095=>"011000000",
  5096=>"100111111",
  5097=>"111101001",
  5098=>"000000001",
  5099=>"010101100",
  5100=>"100011011",
  5101=>"101110001",
  5102=>"001111010",
  5103=>"100100010",
  5104=>"100101111",
  5105=>"010111110",
  5106=>"010001100",
  5107=>"010000100",
  5108=>"101110000",
  5109=>"100111100",
  5110=>"000100110",
  5111=>"111111100",
  5112=>"111010001",
  5113=>"010100111",
  5114=>"101110111",
  5115=>"101101000",
  5116=>"100001110",
  5117=>"111011101",
  5118=>"100001001",
  5119=>"100110001",
  5120=>"011000111",
  5121=>"100100010",
  5122=>"011011001",
  5123=>"001000111",
  5124=>"110101100",
  5125=>"101101100",
  5126=>"011100101",
  5127=>"111100100",
  5128=>"100011100",
  5129=>"110000000",
  5130=>"110100001",
  5131=>"100110011",
  5132=>"110010110",
  5133=>"100010111",
  5134=>"111101111",
  5135=>"100100001",
  5136=>"011010110",
  5137=>"101000100",
  5138=>"100010111",
  5139=>"111110100",
  5140=>"111111011",
  5141=>"110110110",
  5142=>"101001101",
  5143=>"011011100",
  5144=>"011000011",
  5145=>"011101010",
  5146=>"100100101",
  5147=>"000010111",
  5148=>"000010100",
  5149=>"111111011",
  5150=>"000010010",
  5151=>"110000101",
  5152=>"101010100",
  5153=>"101110111",
  5154=>"101001001",
  5155=>"100000100",
  5156=>"001010001",
  5157=>"111110010",
  5158=>"001101011",
  5159=>"110110111",
  5160=>"100110100",
  5161=>"100110111",
  5162=>"000011010",
  5163=>"101001101",
  5164=>"110011001",
  5165=>"101111010",
  5166=>"001100011",
  5167=>"000110101",
  5168=>"010010000",
  5169=>"010110110",
  5170=>"011010010",
  5171=>"000100011",
  5172=>"110100100",
  5173=>"001101101",
  5174=>"100100000",
  5175=>"010010111",
  5176=>"111001110",
  5177=>"100001000",
  5178=>"000010001",
  5179=>"011010010",
  5180=>"010001110",
  5181=>"101100010",
  5182=>"000001101",
  5183=>"010011011",
  5184=>"101001100",
  5185=>"000000100",
  5186=>"101000001",
  5187=>"111111111",
  5188=>"111110101",
  5189=>"101010010",
  5190=>"101101100",
  5191=>"010001100",
  5192=>"101111101",
  5193=>"111111110",
  5194=>"110011010",
  5195=>"111101010",
  5196=>"101111110",
  5197=>"101101100",
  5198=>"111100010",
  5199=>"110011001",
  5200=>"000011011",
  5201=>"010001000",
  5202=>"010111101",
  5203=>"000000000",
  5204=>"001111011",
  5205=>"101001010",
  5206=>"010101000",
  5207=>"001111110",
  5208=>"011111000",
  5209=>"000000111",
  5210=>"001010100",
  5211=>"100101101",
  5212=>"101010011",
  5213=>"100100111",
  5214=>"011010000",
  5215=>"010010011",
  5216=>"001011011",
  5217=>"101101110",
  5218=>"100010101",
  5219=>"101011001",
  5220=>"100110011",
  5221=>"011001011",
  5222=>"101100110",
  5223=>"000110110",
  5224=>"001100010",
  5225=>"101010011",
  5226=>"100000000",
  5227=>"101001000",
  5228=>"111101011",
  5229=>"100010101",
  5230=>"101011100",
  5231=>"100111111",
  5232=>"010000000",
  5233=>"101101111",
  5234=>"111101111",
  5235=>"111110100",
  5236=>"010011100",
  5237=>"010001111",
  5238=>"111100010",
  5239=>"100100001",
  5240=>"011001001",
  5241=>"000001111",
  5242=>"011011101",
  5243=>"101011001",
  5244=>"100111111",
  5245=>"100100011",
  5246=>"001000000",
  5247=>"100100001",
  5248=>"000000000",
  5249=>"110111101",
  5250=>"001000100",
  5251=>"101000000",
  5252=>"010010000",
  5253=>"001101000",
  5254=>"000101011",
  5255=>"110010101",
  5256=>"010010111",
  5257=>"111100010",
  5258=>"100111110",
  5259=>"110111101",
  5260=>"010111101",
  5261=>"111000001",
  5262=>"101100010",
  5263=>"110011000",
  5264=>"011000101",
  5265=>"110100100",
  5266=>"000001000",
  5267=>"011110010",
  5268=>"111110010",
  5269=>"001101110",
  5270=>"010101011",
  5271=>"000100111",
  5272=>"000011100",
  5273=>"101111111",
  5274=>"100101001",
  5275=>"001101100",
  5276=>"011100100",
  5277=>"000100100",
  5278=>"011110110",
  5279=>"000110111",
  5280=>"101001001",
  5281=>"110011100",
  5282=>"010000110",
  5283=>"100000000",
  5284=>"111100001",
  5285=>"000100110",
  5286=>"011100110",
  5287=>"101010110",
  5288=>"011111110",
  5289=>"101010001",
  5290=>"000101011",
  5291=>"110110101",
  5292=>"001100100",
  5293=>"111011101",
  5294=>"011000001",
  5295=>"011000110",
  5296=>"001010101",
  5297=>"000011011",
  5298=>"001100111",
  5299=>"100010010",
  5300=>"011000111",
  5301=>"111011010",
  5302=>"101010000",
  5303=>"110001011",
  5304=>"000110101",
  5305=>"000100100",
  5306=>"111010001",
  5307=>"000100100",
  5308=>"010010000",
  5309=>"111011110",
  5310=>"010011011",
  5311=>"100010101",
  5312=>"111010010",
  5313=>"111110000",
  5314=>"110011000",
  5315=>"101010110",
  5316=>"001001100",
  5317=>"101111011",
  5318=>"111100000",
  5319=>"101100110",
  5320=>"110001100",
  5321=>"100000101",
  5322=>"010110001",
  5323=>"010100100",
  5324=>"000100101",
  5325=>"110101111",
  5326=>"000111010",
  5327=>"001010110",
  5328=>"100000110",
  5329=>"110010110",
  5330=>"101101111",
  5331=>"100010110",
  5332=>"000011001",
  5333=>"110001100",
  5334=>"111010100",
  5335=>"111011100",
  5336=>"111110111",
  5337=>"011001001",
  5338=>"011011101",
  5339=>"111011010",
  5340=>"110011011",
  5341=>"011101111",
  5342=>"110100101",
  5343=>"011010101",
  5344=>"000110101",
  5345=>"100111101",
  5346=>"110101010",
  5347=>"001111000",
  5348=>"001011001",
  5349=>"101100111",
  5350=>"110010111",
  5351=>"110000100",
  5352=>"001001100",
  5353=>"101000000",
  5354=>"101101001",
  5355=>"011101111",
  5356=>"010100010",
  5357=>"101010010",
  5358=>"111001010",
  5359=>"110111000",
  5360=>"111110100",
  5361=>"111001101",
  5362=>"000101111",
  5363=>"000111100",
  5364=>"101100110",
  5365=>"000110010",
  5366=>"000100010",
  5367=>"100110111",
  5368=>"100101110",
  5369=>"000000001",
  5370=>"000101001",
  5371=>"000001101",
  5372=>"011100000",
  5373=>"001110011",
  5374=>"011010110",
  5375=>"100010000",
  5376=>"001110111",
  5377=>"010101100",
  5378=>"101011010",
  5379=>"100011111",
  5380=>"100011110",
  5381=>"001011000",
  5382=>"100000100",
  5383=>"001010011",
  5384=>"000011100",
  5385=>"000001000",
  5386=>"110001111",
  5387=>"110010101",
  5388=>"000111111",
  5389=>"000000101",
  5390=>"110011101",
  5391=>"111001100",
  5392=>"000111011",
  5393=>"011011000",
  5394=>"111101011",
  5395=>"100000000",
  5396=>"101110100",
  5397=>"000111100",
  5398=>"010111110",
  5399=>"100001001",
  5400=>"110111010",
  5401=>"110011111",
  5402=>"111100010",
  5403=>"001010000",
  5404=>"111111010",
  5405=>"011100010",
  5406=>"000110010",
  5407=>"001010111",
  5408=>"111001111",
  5409=>"001000101",
  5410=>"001011101",
  5411=>"011111011",
  5412=>"111011000",
  5413=>"000000110",
  5414=>"100101000",
  5415=>"110101011",
  5416=>"111101100",
  5417=>"011110101",
  5418=>"100001110",
  5419=>"101010010",
  5420=>"111100110",
  5421=>"110000011",
  5422=>"000000011",
  5423=>"111010101",
  5424=>"010001010",
  5425=>"110010100",
  5426=>"111111111",
  5427=>"011111001",
  5428=>"000000101",
  5429=>"101001011",
  5430=>"110011001",
  5431=>"111110100",
  5432=>"011011001",
  5433=>"011100000",
  5434=>"111111111",
  5435=>"101011100",
  5436=>"101010000",
  5437=>"001101011",
  5438=>"000111110",
  5439=>"111001110",
  5440=>"011101011",
  5441=>"000100000",
  5442=>"111000000",
  5443=>"101001110",
  5444=>"011000111",
  5445=>"111110001",
  5446=>"100000001",
  5447=>"101011011",
  5448=>"000101101",
  5449=>"011111111",
  5450=>"010100010",
  5451=>"110010011",
  5452=>"011110101",
  5453=>"000110111",
  5454=>"000111001",
  5455=>"101110000",
  5456=>"101110000",
  5457=>"000110000",
  5458=>"010011100",
  5459=>"001100011",
  5460=>"100101000",
  5461=>"100110111",
  5462=>"010011000",
  5463=>"010011111",
  5464=>"011000100",
  5465=>"101110000",
  5466=>"001011111",
  5467=>"100001000",
  5468=>"100101100",
  5469=>"000001010",
  5470=>"101111000",
  5471=>"000001101",
  5472=>"011100111",
  5473=>"010010000",
  5474=>"011010111",
  5475=>"001001111",
  5476=>"110010101",
  5477=>"110011100",
  5478=>"010110101",
  5479=>"010000110",
  5480=>"100001111",
  5481=>"001111110",
  5482=>"100000110",
  5483=>"010000111",
  5484=>"100011100",
  5485=>"111110001",
  5486=>"101100100",
  5487=>"011100111",
  5488=>"001111110",
  5489=>"100100000",
  5490=>"101000001",
  5491=>"000111101",
  5492=>"111101101",
  5493=>"011100111",
  5494=>"011010111",
  5495=>"000010111",
  5496=>"011110111",
  5497=>"101010000",
  5498=>"110001001",
  5499=>"110001101",
  5500=>"000011101",
  5501=>"010001000",
  5502=>"010000011",
  5503=>"010110110",
  5504=>"010000000",
  5505=>"011010110",
  5506=>"101010000",
  5507=>"110111100",
  5508=>"000010111",
  5509=>"001110001",
  5510=>"011001011",
  5511=>"111011100",
  5512=>"000110111",
  5513=>"111011011",
  5514=>"111010110",
  5515=>"111001011",
  5516=>"101011101",
  5517=>"000001110",
  5518=>"000011101",
  5519=>"000000010",
  5520=>"111100000",
  5521=>"100011011",
  5522=>"110001110",
  5523=>"001110011",
  5524=>"001100101",
  5525=>"001001011",
  5526=>"011011011",
  5527=>"010101111",
  5528=>"111100001",
  5529=>"011110100",
  5530=>"000110111",
  5531=>"010101001",
  5532=>"010111000",
  5533=>"001000110",
  5534=>"110001010",
  5535=>"100010001",
  5536=>"000001001",
  5537=>"101100111",
  5538=>"011111001",
  5539=>"001000101",
  5540=>"010100000",
  5541=>"001111001",
  5542=>"111000000",
  5543=>"101100110",
  5544=>"100000000",
  5545=>"101110011",
  5546=>"000001111",
  5547=>"001000101",
  5548=>"011001101",
  5549=>"000100011",
  5550=>"000111100",
  5551=>"110010001",
  5552=>"111010111",
  5553=>"000001100",
  5554=>"011100011",
  5555=>"010101011",
  5556=>"111001000",
  5557=>"101011001",
  5558=>"110111110",
  5559=>"110001000",
  5560=>"111000011",
  5561=>"111100111",
  5562=>"000100101",
  5563=>"110111010",
  5564=>"100111000",
  5565=>"011110000",
  5566=>"001010011",
  5567=>"001111011",
  5568=>"110011001",
  5569=>"000100111",
  5570=>"010110101",
  5571=>"000101001",
  5572=>"000110111",
  5573=>"100100100",
  5574=>"010001000",
  5575=>"001000010",
  5576=>"111010001",
  5577=>"000000100",
  5578=>"110000101",
  5579=>"011000010",
  5580=>"011001110",
  5581=>"110110110",
  5582=>"011010111",
  5583=>"011000101",
  5584=>"101110001",
  5585=>"000111010",
  5586=>"000001110",
  5587=>"001111010",
  5588=>"010001111",
  5589=>"100010111",
  5590=>"010110000",
  5591=>"110001100",
  5592=>"000010100",
  5593=>"110001010",
  5594=>"111010011",
  5595=>"010010000",
  5596=>"110111101",
  5597=>"010100110",
  5598=>"010111011",
  5599=>"100111011",
  5600=>"011100111",
  5601=>"110010001",
  5602=>"101011111",
  5603=>"111100010",
  5604=>"100101110",
  5605=>"101101011",
  5606=>"001011111",
  5607=>"101100011",
  5608=>"110010100",
  5609=>"110101000",
  5610=>"111111001",
  5611=>"001100001",
  5612=>"100000000",
  5613=>"110100011",
  5614=>"010001000",
  5615=>"111010111",
  5616=>"110001001",
  5617=>"111111111",
  5618=>"100111000",
  5619=>"101011111",
  5620=>"001010011",
  5621=>"000110111",
  5622=>"100110110",
  5623=>"000110100",
  5624=>"001001011",
  5625=>"011001010",
  5626=>"110111111",
  5627=>"011010000",
  5628=>"000101011",
  5629=>"110000000",
  5630=>"000111110",
  5631=>"110010111",
  5632=>"100100001",
  5633=>"110110110",
  5634=>"001101111",
  5635=>"001101011",
  5636=>"001011100",
  5637=>"000011011",
  5638=>"101000000",
  5639=>"111001011",
  5640=>"111010111",
  5641=>"100101110",
  5642=>"110100110",
  5643=>"111011000",
  5644=>"011011101",
  5645=>"010010110",
  5646=>"000100111",
  5647=>"010010101",
  5648=>"011111011",
  5649=>"001110111",
  5650=>"100110110",
  5651=>"100000001",
  5652=>"011101010",
  5653=>"110010111",
  5654=>"011011110",
  5655=>"101001111",
  5656=>"101101011",
  5657=>"000011010",
  5658=>"111000010",
  5659=>"111010010",
  5660=>"101010011",
  5661=>"001011001",
  5662=>"000011001",
  5663=>"100010100",
  5664=>"010010000",
  5665=>"110010000",
  5666=>"011101011",
  5667=>"110111110",
  5668=>"010001111",
  5669=>"001111000",
  5670=>"011010011",
  5671=>"100010111",
  5672=>"001101110",
  5673=>"101100111",
  5674=>"010011010",
  5675=>"100010111",
  5676=>"100100001",
  5677=>"100000011",
  5678=>"011100111",
  5679=>"100001111",
  5680=>"001111000",
  5681=>"001001111",
  5682=>"000100000",
  5683=>"011010011",
  5684=>"110011010",
  5685=>"110101101",
  5686=>"000000011",
  5687=>"111110111",
  5688=>"001111111",
  5689=>"001110101",
  5690=>"011000011",
  5691=>"101011011",
  5692=>"110100110",
  5693=>"110011010",
  5694=>"011000100",
  5695=>"010110000",
  5696=>"100111011",
  5697=>"111100101",
  5698=>"110100001",
  5699=>"010010000",
  5700=>"011011101",
  5701=>"001101011",
  5702=>"001100011",
  5703=>"101100100",
  5704=>"101111011",
  5705=>"111111011",
  5706=>"000011011",
  5707=>"110111010",
  5708=>"011111101",
  5709=>"100001101",
  5710=>"100010101",
  5711=>"010110110",
  5712=>"010101011",
  5713=>"111000101",
  5714=>"000111000",
  5715=>"011010101",
  5716=>"000000010",
  5717=>"001010111",
  5718=>"011000001",
  5719=>"101010110",
  5720=>"001110110",
  5721=>"101000010",
  5722=>"001111100",
  5723=>"110011100",
  5724=>"000011100",
  5725=>"000000100",
  5726=>"101111100",
  5727=>"000000110",
  5728=>"111110011",
  5729=>"110001101",
  5730=>"000010111",
  5731=>"010101110",
  5732=>"000101010",
  5733=>"100110111",
  5734=>"111000101",
  5735=>"101001010",
  5736=>"010011001",
  5737=>"010100100",
  5738=>"011111011",
  5739=>"001011100",
  5740=>"001000111",
  5741=>"111011010",
  5742=>"111000001",
  5743=>"101110000",
  5744=>"111011001",
  5745=>"110110100",
  5746=>"101101101",
  5747=>"001001111",
  5748=>"111101100",
  5749=>"101000010",
  5750=>"011110100",
  5751=>"000100110",
  5752=>"001000000",
  5753=>"110001101",
  5754=>"111010100",
  5755=>"111010000",
  5756=>"011000111",
  5757=>"000110010",
  5758=>"111101100",
  5759=>"101000110",
  5760=>"110001011",
  5761=>"101110110",
  5762=>"000010001",
  5763=>"110000100",
  5764=>"000110110",
  5765=>"011110010",
  5766=>"000111010",
  5767=>"111111111",
  5768=>"000111001",
  5769=>"000010110",
  5770=>"101110010",
  5771=>"111011000",
  5772=>"011010101",
  5773=>"001111110",
  5774=>"111110001",
  5775=>"000010000",
  5776=>"011100011",
  5777=>"000110110",
  5778=>"100101001",
  5779=>"101001101",
  5780=>"111101011",
  5781=>"000000110",
  5782=>"110000001",
  5783=>"101100001",
  5784=>"111000111",
  5785=>"100011001",
  5786=>"110110000",
  5787=>"101110010",
  5788=>"001000010",
  5789=>"011010001",
  5790=>"001001011",
  5791=>"010111101",
  5792=>"100011110",
  5793=>"110001011",
  5794=>"110001101",
  5795=>"011000001",
  5796=>"101000011",
  5797=>"111111001",
  5798=>"011000001",
  5799=>"100111000",
  5800=>"111011101",
  5801=>"101001110",
  5802=>"000110000",
  5803=>"011000110",
  5804=>"100101100",
  5805=>"101101001",
  5806=>"010101011",
  5807=>"100000000",
  5808=>"001110111",
  5809=>"010000110",
  5810=>"001100001",
  5811=>"111110001",
  5812=>"100000111",
  5813=>"000101000",
  5814=>"110100110",
  5815=>"101111010",
  5816=>"111011100",
  5817=>"111110101",
  5818=>"001111111",
  5819=>"010010101",
  5820=>"000111010",
  5821=>"001011011",
  5822=>"000100000",
  5823=>"000010010",
  5824=>"011101001",
  5825=>"010101000",
  5826=>"110100000",
  5827=>"011010011",
  5828=>"010101100",
  5829=>"001000000",
  5830=>"001000110",
  5831=>"011001011",
  5832=>"000010110",
  5833=>"011001000",
  5834=>"110110010",
  5835=>"011010000",
  5836=>"011011000",
  5837=>"111001000",
  5838=>"010111001",
  5839=>"011111111",
  5840=>"011101100",
  5841=>"100011001",
  5842=>"010101011",
  5843=>"000010111",
  5844=>"001000101",
  5845=>"110011111",
  5846=>"101000010",
  5847=>"101001010",
  5848=>"000011001",
  5849=>"110110110",
  5850=>"101111100",
  5851=>"001001111",
  5852=>"111000010",
  5853=>"010100000",
  5854=>"000110011",
  5855=>"101111010",
  5856=>"111101110",
  5857=>"000011011",
  5858=>"010111101",
  5859=>"000110101",
  5860=>"001001100",
  5861=>"000101000",
  5862=>"011100101",
  5863=>"010100110",
  5864=>"100110101",
  5865=>"111011000",
  5866=>"000100100",
  5867=>"001000001",
  5868=>"100000111",
  5869=>"010000101",
  5870=>"100000001",
  5871=>"010011101",
  5872=>"111110101",
  5873=>"010110010",
  5874=>"101011110",
  5875=>"100000010",
  5876=>"110110000",
  5877=>"110000011",
  5878=>"101000100",
  5879=>"110111010",
  5880=>"111101011",
  5881=>"111011111",
  5882=>"000000100",
  5883=>"011101101",
  5884=>"000011100",
  5885=>"010000000",
  5886=>"101000101",
  5887=>"011111110",
  5888=>"000110110",
  5889=>"001111010",
  5890=>"000000110",
  5891=>"001110111",
  5892=>"011010100",
  5893=>"110100001",
  5894=>"101111101",
  5895=>"010101101",
  5896=>"000010011",
  5897=>"110110010",
  5898=>"000100000",
  5899=>"100111011",
  5900=>"101011001",
  5901=>"111110111",
  5902=>"001001100",
  5903=>"000010101",
  5904=>"100111100",
  5905=>"101101010",
  5906=>"000111101",
  5907=>"111001010",
  5908=>"101000100",
  5909=>"111110011",
  5910=>"101111000",
  5911=>"110011110",
  5912=>"000011011",
  5913=>"001001001",
  5914=>"001000010",
  5915=>"111000111",
  5916=>"110110011",
  5917=>"011111110",
  5918=>"100101101",
  5919=>"111110000",
  5920=>"000100001",
  5921=>"001010100",
  5922=>"101010010",
  5923=>"110010001",
  5924=>"010010000",
  5925=>"001001011",
  5926=>"011100000",
  5927=>"010111101",
  5928=>"001011000",
  5929=>"100010000",
  5930=>"100001001",
  5931=>"001110001",
  5932=>"001100110",
  5933=>"111100110",
  5934=>"101001000",
  5935=>"110010000",
  5936=>"000100101",
  5937=>"101010101",
  5938=>"000000101",
  5939=>"001010011",
  5940=>"000100100",
  5941=>"111000111",
  5942=>"000011110",
  5943=>"001000110",
  5944=>"100110110",
  5945=>"110110001",
  5946=>"111001011",
  5947=>"001111010",
  5948=>"100100010",
  5949=>"000000100",
  5950=>"100011011",
  5951=>"110000011",
  5952=>"110110100",
  5953=>"101010000",
  5954=>"001101101",
  5955=>"010100010",
  5956=>"000100100",
  5957=>"110011101",
  5958=>"100011110",
  5959=>"110111011",
  5960=>"001101000",
  5961=>"101110001",
  5962=>"011110110",
  5963=>"011001110",
  5964=>"111001110",
  5965=>"101110000",
  5966=>"110101001",
  5967=>"101010010",
  5968=>"000000111",
  5969=>"001111111",
  5970=>"010000100",
  5971=>"000101111",
  5972=>"001101010",
  5973=>"101010000",
  5974=>"101000011",
  5975=>"101111010",
  5976=>"010111101",
  5977=>"101001101",
  5978=>"101011011",
  5979=>"000110110",
  5980=>"101001001",
  5981=>"001000101",
  5982=>"110010101",
  5983=>"110111111",
  5984=>"001001011",
  5985=>"000001000",
  5986=>"111111111",
  5987=>"001111110",
  5988=>"110100100",
  5989=>"111011100",
  5990=>"000000000",
  5991=>"011001011",
  5992=>"110001100",
  5993=>"100010011",
  5994=>"010010000",
  5995=>"010100111",
  5996=>"100101010",
  5997=>"011001001",
  5998=>"000100001",
  5999=>"000111110",
  6000=>"011001001",
  6001=>"111001010",
  6002=>"101100000",
  6003=>"001001111",
  6004=>"010011010",
  6005=>"111110101",
  6006=>"111111100",
  6007=>"011001001",
  6008=>"010000011",
  6009=>"110001101",
  6010=>"111100101",
  6011=>"111001010",
  6012=>"001011111",
  6013=>"011101010",
  6014=>"111110001",
  6015=>"010000110",
  6016=>"011010100",
  6017=>"101101010",
  6018=>"011010010",
  6019=>"110110111",
  6020=>"100101111",
  6021=>"010110010",
  6022=>"000111000",
  6023=>"101010110",
  6024=>"011101010",
  6025=>"100111100",
  6026=>"110101110",
  6027=>"101101101",
  6028=>"100011100",
  6029=>"111110100",
  6030=>"011101100",
  6031=>"000101110",
  6032=>"011110001",
  6033=>"001110101",
  6034=>"100101001",
  6035=>"110101001",
  6036=>"010101000",
  6037=>"111011110",
  6038=>"011101000",
  6039=>"000101001",
  6040=>"111001010",
  6041=>"011011011",
  6042=>"001001000",
  6043=>"100100101",
  6044=>"100110111",
  6045=>"011111110",
  6046=>"110111000",
  6047=>"000111110",
  6048=>"100100000",
  6049=>"000001100",
  6050=>"111110001",
  6051=>"011001001",
  6052=>"111001111",
  6053=>"010100100",
  6054=>"101110010",
  6055=>"011100110",
  6056=>"010001111",
  6057=>"010101100",
  6058=>"100001000",
  6059=>"101011001",
  6060=>"111100010",
  6061=>"100000111",
  6062=>"011110010",
  6063=>"100101001",
  6064=>"001001100",
  6065=>"111001011",
  6066=>"010111101",
  6067=>"110001001",
  6068=>"010010111",
  6069=>"000110001",
  6070=>"110101011",
  6071=>"110110011",
  6072=>"111000101",
  6073=>"000000100",
  6074=>"000000011",
  6075=>"111011011",
  6076=>"010111100",
  6077=>"111111100",
  6078=>"100101111",
  6079=>"010000000",
  6080=>"010011101",
  6081=>"001110100",
  6082=>"111011100",
  6083=>"000011110",
  6084=>"101011010",
  6085=>"111101110",
  6086=>"111111010",
  6087=>"110001110",
  6088=>"100011100",
  6089=>"001100011",
  6090=>"001100101",
  6091=>"001011100",
  6092=>"011100010",
  6093=>"110010100",
  6094=>"010100010",
  6095=>"000110000",
  6096=>"111011011",
  6097=>"100100000",
  6098=>"111111001",
  6099=>"010000001",
  6100=>"011101110",
  6101=>"111110111",
  6102=>"000011000",
  6103=>"111111110",
  6104=>"011110011",
  6105=>"001000011",
  6106=>"111100000",
  6107=>"011000001",
  6108=>"010010011",
  6109=>"001110000",
  6110=>"101101001",
  6111=>"110111010",
  6112=>"010011010",
  6113=>"011011001",
  6114=>"110010101",
  6115=>"001111001",
  6116=>"110110010",
  6117=>"001110001",
  6118=>"011000000",
  6119=>"100101110",
  6120=>"000110011",
  6121=>"010101100",
  6122=>"000000110",
  6123=>"000001100",
  6124=>"101111101",
  6125=>"100100000",
  6126=>"110101011",
  6127=>"000101110",
  6128=>"010110111",
  6129=>"000100010",
  6130=>"101010100",
  6131=>"110110111",
  6132=>"100111111",
  6133=>"100001010",
  6134=>"011110001",
  6135=>"010111001",
  6136=>"100010111",
  6137=>"101010100",
  6138=>"110100101",
  6139=>"100110000",
  6140=>"110110111",
  6141=>"000000010",
  6142=>"110010100",
  6143=>"010110101",
  6144=>"011110011",
  6145=>"000000111",
  6146=>"111110001",
  6147=>"001001100",
  6148=>"010101001",
  6149=>"100110110",
  6150=>"011111100",
  6151=>"001101001",
  6152=>"110100001",
  6153=>"001000000",
  6154=>"110101001",
  6155=>"100000011",
  6156=>"001001110",
  6157=>"010111100",
  6158=>"000011101",
  6159=>"101111110",
  6160=>"001101111",
  6161=>"111101011",
  6162=>"101100011",
  6163=>"100011000",
  6164=>"111111011",
  6165=>"010011100",
  6166=>"101101100",
  6167=>"100000111",
  6168=>"001101000",
  6169=>"000001111",
  6170=>"100000011",
  6171=>"000101001",
  6172=>"100110010",
  6173=>"010101001",
  6174=>"111011101",
  6175=>"111000101",
  6176=>"111010001",
  6177=>"010001111",
  6178=>"011000111",
  6179=>"101110011",
  6180=>"000000011",
  6181=>"011110001",
  6182=>"010110001",
  6183=>"101110011",
  6184=>"101000110",
  6185=>"000110101",
  6186=>"000011011",
  6187=>"111111001",
  6188=>"000001110",
  6189=>"111110010",
  6190=>"111100001",
  6191=>"000110100",
  6192=>"100011011",
  6193=>"011010011",
  6194=>"011000000",
  6195=>"000100101",
  6196=>"100000110",
  6197=>"011001001",
  6198=>"101011111",
  6199=>"000010101",
  6200=>"001000110",
  6201=>"001100001",
  6202=>"110100110",
  6203=>"001010000",
  6204=>"000011010",
  6205=>"001001011",
  6206=>"100011001",
  6207=>"000111010",
  6208=>"101101001",
  6209=>"111010100",
  6210=>"100011100",
  6211=>"100000011",
  6212=>"101101110",
  6213=>"110011000",
  6214=>"100011011",
  6215=>"111110111",
  6216=>"110100000",
  6217=>"010011110",
  6218=>"110000100",
  6219=>"110001100",
  6220=>"001000001",
  6221=>"110000100",
  6222=>"101011000",
  6223=>"100110110",
  6224=>"101100000",
  6225=>"000001101",
  6226=>"010000101",
  6227=>"011011001",
  6228=>"111001101",
  6229=>"001100001",
  6230=>"110010000",
  6231=>"101111010",
  6232=>"111111111",
  6233=>"111111010",
  6234=>"011011111",
  6235=>"010010000",
  6236=>"011111110",
  6237=>"010100100",
  6238=>"101001101",
  6239=>"111111110",
  6240=>"110011100",
  6241=>"111000111",
  6242=>"001000100",
  6243=>"100011101",
  6244=>"010010011",
  6245=>"010101001",
  6246=>"100110100",
  6247=>"010110001",
  6248=>"011111001",
  6249=>"110111100",
  6250=>"110001001",
  6251=>"000011000",
  6252=>"001000011",
  6253=>"101001001",
  6254=>"010000101",
  6255=>"000011101",
  6256=>"101000000",
  6257=>"111001001",
  6258=>"110111101",
  6259=>"011010001",
  6260=>"001111100",
  6261=>"010000100",
  6262=>"111100110",
  6263=>"001111101",
  6264=>"000110011",
  6265=>"001101010",
  6266=>"001100011",
  6267=>"010001010",
  6268=>"111001010",
  6269=>"111101110",
  6270=>"100101001",
  6271=>"111000010",
  6272=>"010001001",
  6273=>"001001111",
  6274=>"000001010",
  6275=>"001101110",
  6276=>"101010001",
  6277=>"000001010",
  6278=>"000100101",
  6279=>"001111111",
  6280=>"111101001",
  6281=>"011101111",
  6282=>"100000100",
  6283=>"110010001",
  6284=>"001010000",
  6285=>"100111101",
  6286=>"100111001",
  6287=>"101001000",
  6288=>"101010000",
  6289=>"100110110",
  6290=>"110011001",
  6291=>"100000010",
  6292=>"101001010",
  6293=>"010001111",
  6294=>"011111000",
  6295=>"001110000",
  6296=>"100100111",
  6297=>"011101000",
  6298=>"100101001",
  6299=>"000100110",
  6300=>"101101001",
  6301=>"111111000",
  6302=>"100010101",
  6303=>"100100111",
  6304=>"011100100",
  6305=>"001110101",
  6306=>"000110011",
  6307=>"100001000",
  6308=>"110010010",
  6309=>"001101001",
  6310=>"010111101",
  6311=>"101100111",
  6312=>"111110111",
  6313=>"010000010",
  6314=>"111101000",
  6315=>"100110101",
  6316=>"001111111",
  6317=>"001100011",
  6318=>"001010111",
  6319=>"101101101",
  6320=>"000001110",
  6321=>"001001010",
  6322=>"110010011",
  6323=>"101000010",
  6324=>"110010101",
  6325=>"100011000",
  6326=>"101001010",
  6327=>"010110110",
  6328=>"010101000",
  6329=>"111001011",
  6330=>"011000100",
  6331=>"001001101",
  6332=>"000100000",
  6333=>"101101010",
  6334=>"100011011",
  6335=>"000010000",
  6336=>"001000011",
  6337=>"100101000",
  6338=>"001111100",
  6339=>"010111011",
  6340=>"011110000",
  6341=>"010111101",
  6342=>"110011000",
  6343=>"110101000",
  6344=>"101111000",
  6345=>"101101101",
  6346=>"010011101",
  6347=>"011100101",
  6348=>"110110001",
  6349=>"010110101",
  6350=>"110100111",
  6351=>"001110111",
  6352=>"010001001",
  6353=>"000011011",
  6354=>"001100100",
  6355=>"011001001",
  6356=>"000110011",
  6357=>"100100000",
  6358=>"000001001",
  6359=>"101100101",
  6360=>"101101010",
  6361=>"101101110",
  6362=>"101001010",
  6363=>"110010000",
  6364=>"010000111",
  6365=>"011101001",
  6366=>"011001110",
  6367=>"000100011",
  6368=>"000000000",
  6369=>"010000100",
  6370=>"000110111",
  6371=>"110000110",
  6372=>"100000100",
  6373=>"101110101",
  6374=>"010110001",
  6375=>"001001100",
  6376=>"001111101",
  6377=>"101111010",
  6378=>"011011101",
  6379=>"100000111",
  6380=>"100001110",
  6381=>"001100110",
  6382=>"111110110",
  6383=>"100111001",
  6384=>"111001100",
  6385=>"010111110",
  6386=>"110000000",
  6387=>"000010111",
  6388=>"111001000",
  6389=>"100100011",
  6390=>"101010010",
  6391=>"100001000",
  6392=>"010010001",
  6393=>"111110111",
  6394=>"100110100",
  6395=>"101000110",
  6396=>"110110001",
  6397=>"010111010",
  6398=>"001100111",
  6399=>"000000111",
  6400=>"010100001",
  6401=>"110001111",
  6402=>"000111001",
  6403=>"001000111",
  6404=>"101001101",
  6405=>"000000101",
  6406=>"000010100",
  6407=>"000110101",
  6408=>"011100001",
  6409=>"001010010",
  6410=>"011111000",
  6411=>"101000001",
  6412=>"101011011",
  6413=>"010111101",
  6414=>"110110101",
  6415=>"010111110",
  6416=>"001111001",
  6417=>"101001000",
  6418=>"110110111",
  6419=>"100111100",
  6420=>"000100101",
  6421=>"010110000",
  6422=>"011011111",
  6423=>"001000100",
  6424=>"111111000",
  6425=>"010001001",
  6426=>"010000001",
  6427=>"101001111",
  6428=>"010101101",
  6429=>"100011001",
  6430=>"111101001",
  6431=>"001111001",
  6432=>"100101111",
  6433=>"101110011",
  6434=>"101100001",
  6435=>"000111011",
  6436=>"011101111",
  6437=>"100010010",
  6438=>"011111011",
  6439=>"100111010",
  6440=>"100100100",
  6441=>"111011111",
  6442=>"011010101",
  6443=>"110111101",
  6444=>"010111111",
  6445=>"000010111",
  6446=>"000100001",
  6447=>"100100101",
  6448=>"111101110",
  6449=>"110110001",
  6450=>"011000001",
  6451=>"001001110",
  6452=>"101000011",
  6453=>"001100101",
  6454=>"010000110",
  6455=>"111101000",
  6456=>"111011100",
  6457=>"011001001",
  6458=>"101100101",
  6459=>"110101101",
  6460=>"000101000",
  6461=>"000011011",
  6462=>"101011001",
  6463=>"101101100",
  6464=>"101111001",
  6465=>"110101111",
  6466=>"010110101",
  6467=>"001111111",
  6468=>"101000011",
  6469=>"001110101",
  6470=>"010100000",
  6471=>"011110110",
  6472=>"001001000",
  6473=>"001010001",
  6474=>"111111000",
  6475=>"111000101",
  6476=>"010110001",
  6477=>"001001110",
  6478=>"101111101",
  6479=>"010111101",
  6480=>"001110110",
  6481=>"010110000",
  6482=>"100001011",
  6483=>"010111110",
  6484=>"110000011",
  6485=>"011110110",
  6486=>"100111101",
  6487=>"010010010",
  6488=>"110100011",
  6489=>"011100101",
  6490=>"011011101",
  6491=>"110010100",
  6492=>"000111100",
  6493=>"101111110",
  6494=>"100100010",
  6495=>"000000100",
  6496=>"011111001",
  6497=>"011100000",
  6498=>"110110101",
  6499=>"001111111",
  6500=>"010000000",
  6501=>"111100010",
  6502=>"000011001",
  6503=>"000111010",
  6504=>"000101000",
  6505=>"000000000",
  6506=>"111010010",
  6507=>"011001110",
  6508=>"100110110",
  6509=>"001001101",
  6510=>"010100010",
  6511=>"000000110",
  6512=>"110000100",
  6513=>"001011111",
  6514=>"010011101",
  6515=>"111110111",
  6516=>"110001100",
  6517=>"111110100",
  6518=>"111010111",
  6519=>"001010011",
  6520=>"111111001",
  6521=>"100010110",
  6522=>"111111111",
  6523=>"111001000",
  6524=>"010000001",
  6525=>"101111110",
  6526=>"101110011",
  6527=>"011000101",
  6528=>"110100100",
  6529=>"111111111",
  6530=>"100001110",
  6531=>"001100000",
  6532=>"111111110",
  6533=>"010110101",
  6534=>"101111001",
  6535=>"111101101",
  6536=>"010010001",
  6537=>"010111000",
  6538=>"011100111",
  6539=>"110000011",
  6540=>"100011100",
  6541=>"011010010",
  6542=>"000101011",
  6543=>"001011010",
  6544=>"101010100",
  6545=>"101000001",
  6546=>"011011100",
  6547=>"101100101",
  6548=>"111011100",
  6549=>"010001001",
  6550=>"011000100",
  6551=>"011101011",
  6552=>"001011101",
  6553=>"101111110",
  6554=>"110011111",
  6555=>"000001011",
  6556=>"101111010",
  6557=>"000000100",
  6558=>"001010010",
  6559=>"101110110",
  6560=>"111000110",
  6561=>"000010010",
  6562=>"000110000",
  6563=>"011111010",
  6564=>"111110100",
  6565=>"000110100",
  6566=>"011010001",
  6567=>"001000010",
  6568=>"010100111",
  6569=>"011010101",
  6570=>"111111101",
  6571=>"100011001",
  6572=>"000000100",
  6573=>"000100111",
  6574=>"001100000",
  6575=>"101101010",
  6576=>"111111110",
  6577=>"101110110",
  6578=>"110111000",
  6579=>"011110001",
  6580=>"000011111",
  6581=>"000000001",
  6582=>"010001111",
  6583=>"111100000",
  6584=>"001100000",
  6585=>"010011010",
  6586=>"011111101",
  6587=>"110011101",
  6588=>"100011010",
  6589=>"000011101",
  6590=>"100001000",
  6591=>"101110111",
  6592=>"001100111",
  6593=>"011000010",
  6594=>"111011101",
  6595=>"111111010",
  6596=>"000100101",
  6597=>"111010100",
  6598=>"010110000",
  6599=>"101010011",
  6600=>"000000100",
  6601=>"010001110",
  6602=>"011010101",
  6603=>"011111110",
  6604=>"001000010",
  6605=>"010111011",
  6606=>"010011110",
  6607=>"101100011",
  6608=>"111110100",
  6609=>"101011011",
  6610=>"000011010",
  6611=>"000110001",
  6612=>"111100100",
  6613=>"001000000",
  6614=>"001000101",
  6615=>"000101001",
  6616=>"000000101",
  6617=>"001000111",
  6618=>"111110011",
  6619=>"110111011",
  6620=>"110000001",
  6621=>"111001101",
  6622=>"101101011",
  6623=>"000000000",
  6624=>"111101100",
  6625=>"000100000",
  6626=>"010110011",
  6627=>"110111001",
  6628=>"110110111",
  6629=>"111010010",
  6630=>"101001010",
  6631=>"010001010",
  6632=>"110011011",
  6633=>"101111001",
  6634=>"100000010",
  6635=>"100010000",
  6636=>"111101100",
  6637=>"100001111",
  6638=>"100010011",
  6639=>"011011101",
  6640=>"110010111",
  6641=>"110011110",
  6642=>"101101110",
  6643=>"000000001",
  6644=>"001010101",
  6645=>"011011010",
  6646=>"000101101",
  6647=>"001100111",
  6648=>"101101111",
  6649=>"011001101",
  6650=>"000000001",
  6651=>"011011100",
  6652=>"111100101",
  6653=>"001011001",
  6654=>"101000111",
  6655=>"110100100",
  6656=>"011110100",
  6657=>"010000111",
  6658=>"001000100",
  6659=>"010101111",
  6660=>"110111010",
  6661=>"011000100",
  6662=>"001001111",
  6663=>"111100001",
  6664=>"001010001",
  6665=>"100000101",
  6666=>"111000101",
  6667=>"100000000",
  6668=>"110100001",
  6669=>"100110011",
  6670=>"101001100",
  6671=>"001000101",
  6672=>"001100011",
  6673=>"111010101",
  6674=>"101101011",
  6675=>"110101101",
  6676=>"100110011",
  6677=>"110010010",
  6678=>"000110000",
  6679=>"101011000",
  6680=>"010000000",
  6681=>"111011111",
  6682=>"010110110",
  6683=>"001111010",
  6684=>"000101101",
  6685=>"010000001",
  6686=>"010011000",
  6687=>"101010000",
  6688=>"000110011",
  6689=>"011000110",
  6690=>"000011001",
  6691=>"110110001",
  6692=>"111010110",
  6693=>"001010110",
  6694=>"110101101",
  6695=>"010011001",
  6696=>"111101100",
  6697=>"100101110",
  6698=>"010011111",
  6699=>"001011111",
  6700=>"100001001",
  6701=>"101010001",
  6702=>"010101000",
  6703=>"010111000",
  6704=>"111100011",
  6705=>"100001111",
  6706=>"001111100",
  6707=>"000100011",
  6708=>"010000011",
  6709=>"100101110",
  6710=>"000001111",
  6711=>"111111101",
  6712=>"001000101",
  6713=>"111111000",
  6714=>"001001111",
  6715=>"001000110",
  6716=>"011000101",
  6717=>"010110010",
  6718=>"010101111",
  6719=>"101001101",
  6720=>"000011000",
  6721=>"000000001",
  6722=>"110111101",
  6723=>"000001000",
  6724=>"111001100",
  6725=>"100000110",
  6726=>"001000100",
  6727=>"111101111",
  6728=>"100111001",
  6729=>"000111001",
  6730=>"010111100",
  6731=>"001011011",
  6732=>"010100001",
  6733=>"111111010",
  6734=>"001010011",
  6735=>"111111000",
  6736=>"100111010",
  6737=>"111110101",
  6738=>"101101010",
  6739=>"100011010",
  6740=>"100011001",
  6741=>"011000110",
  6742=>"100000101",
  6743=>"010001110",
  6744=>"100010010",
  6745=>"010001000",
  6746=>"101000011",
  6747=>"000000011",
  6748=>"110010101",
  6749=>"000000100",
  6750=>"111110110",
  6751=>"001111011",
  6752=>"101011001",
  6753=>"010011001",
  6754=>"100001001",
  6755=>"110001011",
  6756=>"111111110",
  6757=>"111011111",
  6758=>"110001011",
  6759=>"010111001",
  6760=>"100010101",
  6761=>"000010011",
  6762=>"110110001",
  6763=>"101001101",
  6764=>"100111010",
  6765=>"100001101",
  6766=>"101000011",
  6767=>"100111000",
  6768=>"110000111",
  6769=>"001111101",
  6770=>"000000000",
  6771=>"101010010",
  6772=>"001010110",
  6773=>"000001101",
  6774=>"110010010",
  6775=>"111100101",
  6776=>"000011111",
  6777=>"010010001",
  6778=>"111101011",
  6779=>"110010111",
  6780=>"001010100",
  6781=>"111100111",
  6782=>"100110100",
  6783=>"000011100",
  6784=>"111110110",
  6785=>"101001111",
  6786=>"010000000",
  6787=>"110000101",
  6788=>"011011101",
  6789=>"101000000",
  6790=>"101100011",
  6791=>"001001101",
  6792=>"001111001",
  6793=>"110001100",
  6794=>"001101100",
  6795=>"100010100",
  6796=>"010000000",
  6797=>"110101000",
  6798=>"000010111",
  6799=>"011101110",
  6800=>"010100110",
  6801=>"110110101",
  6802=>"001000111",
  6803=>"011010110",
  6804=>"100111011",
  6805=>"111101000",
  6806=>"101001100",
  6807=>"111010010",
  6808=>"010101110",
  6809=>"110110011",
  6810=>"001001000",
  6811=>"100011000",
  6812=>"101011101",
  6813=>"010111000",
  6814=>"110010011",
  6815=>"000010000",
  6816=>"001100110",
  6817=>"011000100",
  6818=>"100111110",
  6819=>"101101111",
  6820=>"001000100",
  6821=>"010011001",
  6822=>"100111001",
  6823=>"101110110",
  6824=>"000000111",
  6825=>"110001100",
  6826=>"001100011",
  6827=>"010101110",
  6828=>"111110110",
  6829=>"011011000",
  6830=>"111001011",
  6831=>"011100111",
  6832=>"011110001",
  6833=>"010000100",
  6834=>"101000111",
  6835=>"011010000",
  6836=>"001000101",
  6837=>"100111111",
  6838=>"111110001",
  6839=>"001000010",
  6840=>"001011110",
  6841=>"000111001",
  6842=>"001011100",
  6843=>"101010111",
  6844=>"101011011",
  6845=>"011100100",
  6846=>"000111100",
  6847=>"101110000",
  6848=>"111011011",
  6849=>"000010100",
  6850=>"010000010",
  6851=>"110111011",
  6852=>"110101110",
  6853=>"011001000",
  6854=>"110000101",
  6855=>"111010101",
  6856=>"001100001",
  6857=>"011010101",
  6858=>"111100001",
  6859=>"010000110",
  6860=>"001111101",
  6861=>"001110011",
  6862=>"110111100",
  6863=>"011100001",
  6864=>"000100100",
  6865=>"011100110",
  6866=>"110110001",
  6867=>"010010010",
  6868=>"100100100",
  6869=>"011100001",
  6870=>"110001111",
  6871=>"101010111",
  6872=>"101011100",
  6873=>"100111100",
  6874=>"111101111",
  6875=>"110001011",
  6876=>"001100101",
  6877=>"000011010",
  6878=>"111110101",
  6879=>"101110001",
  6880=>"111101111",
  6881=>"110110101",
  6882=>"101100010",
  6883=>"100010010",
  6884=>"000111011",
  6885=>"010111001",
  6886=>"110111100",
  6887=>"101000001",
  6888=>"101000101",
  6889=>"100001111",
  6890=>"011110100",
  6891=>"001010010",
  6892=>"100011101",
  6893=>"101001101",
  6894=>"101001101",
  6895=>"110001100",
  6896=>"011111110",
  6897=>"001101001",
  6898=>"001101010",
  6899=>"100000011",
  6900=>"110010100",
  6901=>"011110101",
  6902=>"000001001",
  6903=>"111010010",
  6904=>"101010001",
  6905=>"100010001",
  6906=>"010010011",
  6907=>"101000111",
  6908=>"011000000",
  6909=>"110000100",
  6910=>"110100111",
  6911=>"010011000",
  6912=>"001011011",
  6913=>"001110101",
  6914=>"001110110",
  6915=>"010101010",
  6916=>"110101100",
  6917=>"011011111",
  6918=>"000011000",
  6919=>"011011001",
  6920=>"101001011",
  6921=>"010101101",
  6922=>"100100001",
  6923=>"001101111",
  6924=>"101001111",
  6925=>"010100000",
  6926=>"011110010",
  6927=>"110100100",
  6928=>"010001100",
  6929=>"000101000",
  6930=>"010111001",
  6931=>"010101110",
  6932=>"110100010",
  6933=>"100001100",
  6934=>"001111101",
  6935=>"101110110",
  6936=>"110010101",
  6937=>"110011110",
  6938=>"010111010",
  6939=>"100011011",
  6940=>"111011110",
  6941=>"010010111",
  6942=>"001110101",
  6943=>"100001101",
  6944=>"011110100",
  6945=>"101111001",
  6946=>"101110000",
  6947=>"110100010",
  6948=>"111111010",
  6949=>"110000000",
  6950=>"000100000",
  6951=>"101100111",
  6952=>"000000110",
  6953=>"010101000",
  6954=>"000101001",
  6955=>"011011111",
  6956=>"010100110",
  6957=>"111000100",
  6958=>"000011101",
  6959=>"000101111",
  6960=>"101001111",
  6961=>"001010011",
  6962=>"000100010",
  6963=>"011100111",
  6964=>"010110011",
  6965=>"010000111",
  6966=>"101000001",
  6967=>"000111000",
  6968=>"010100000",
  6969=>"110010100",
  6970=>"001111100",
  6971=>"111010010",
  6972=>"101011010",
  6973=>"011111100",
  6974=>"101001110",
  6975=>"000111010",
  6976=>"111001100",
  6977=>"111010100",
  6978=>"001101010",
  6979=>"010110111",
  6980=>"111001101",
  6981=>"101001101",
  6982=>"001010001",
  6983=>"100001010",
  6984=>"110111010",
  6985=>"110001001",
  6986=>"011001110",
  6987=>"000101011",
  6988=>"010110000",
  6989=>"111100101",
  6990=>"001001000",
  6991=>"001110010",
  6992=>"000000000",
  6993=>"111111011",
  6994=>"001010000",
  6995=>"111100011",
  6996=>"001000011",
  6997=>"101000011",
  6998=>"010000001",
  6999=>"001000010",
  7000=>"011010000",
  7001=>"000010001",
  7002=>"000111110",
  7003=>"111001000",
  7004=>"001110011",
  7005=>"000000001",
  7006=>"111111011",
  7007=>"010011011",
  7008=>"011001000",
  7009=>"010000001",
  7010=>"111011111",
  7011=>"010101101",
  7012=>"010101100",
  7013=>"001001100",
  7014=>"000110010",
  7015=>"101111100",
  7016=>"100111011",
  7017=>"100011110",
  7018=>"111010110",
  7019=>"111101110",
  7020=>"001100000",
  7021=>"010100110",
  7022=>"101010011",
  7023=>"010001001",
  7024=>"100010011",
  7025=>"110100000",
  7026=>"110011101",
  7027=>"011100000",
  7028=>"011110100",
  7029=>"111100100",
  7030=>"110010010",
  7031=>"101000000",
  7032=>"001110011",
  7033=>"100101011",
  7034=>"001011000",
  7035=>"011100011",
  7036=>"100011001",
  7037=>"010010000",
  7038=>"101100111",
  7039=>"001111111",
  7040=>"100011110",
  7041=>"000000001",
  7042=>"001001101",
  7043=>"101010011",
  7044=>"001011001",
  7045=>"100111011",
  7046=>"010000111",
  7047=>"101100001",
  7048=>"011011011",
  7049=>"101110111",
  7050=>"011111101",
  7051=>"001011010",
  7052=>"000110111",
  7053=>"111110011",
  7054=>"100011000",
  7055=>"100000100",
  7056=>"111101001",
  7057=>"100000100",
  7058=>"000100011",
  7059=>"001011001",
  7060=>"110000110",
  7061=>"001110010",
  7062=>"110000001",
  7063=>"110101101",
  7064=>"010101001",
  7065=>"101111011",
  7066=>"011010001",
  7067=>"111101000",
  7068=>"011100000",
  7069=>"100001000",
  7070=>"110110101",
  7071=>"011110000",
  7072=>"101101110",
  7073=>"111010100",
  7074=>"011100100",
  7075=>"111111011",
  7076=>"110110110",
  7077=>"100000101",
  7078=>"000100010",
  7079=>"010100001",
  7080=>"111010111",
  7081=>"111001011",
  7082=>"101100011",
  7083=>"000001001",
  7084=>"101101111",
  7085=>"101111101",
  7086=>"011111100",
  7087=>"100001011",
  7088=>"011011110",
  7089=>"000011101",
  7090=>"110001110",
  7091=>"011000100",
  7092=>"000011110",
  7093=>"111100111",
  7094=>"110101100",
  7095=>"011100111",
  7096=>"010100000",
  7097=>"111011011",
  7098=>"000010001",
  7099=>"000111000",
  7100=>"010010111",
  7101=>"101110001",
  7102=>"000110010",
  7103=>"111011010",
  7104=>"111100001",
  7105=>"001010011",
  7106=>"110111001",
  7107=>"110101110",
  7108=>"111100100",
  7109=>"111101111",
  7110=>"111000100",
  7111=>"011110101",
  7112=>"101010100",
  7113=>"101011110",
  7114=>"100110111",
  7115=>"101101001",
  7116=>"000110110",
  7117=>"010000110",
  7118=>"001101001",
  7119=>"010000111",
  7120=>"111011000",
  7121=>"101101101",
  7122=>"110110100",
  7123=>"010010010",
  7124=>"001110010",
  7125=>"000010001",
  7126=>"011111111",
  7127=>"000110100",
  7128=>"111100000",
  7129=>"010010101",
  7130=>"101111011",
  7131=>"101001100",
  7132=>"000011011",
  7133=>"110100001",
  7134=>"000101101",
  7135=>"101100110",
  7136=>"101011001",
  7137=>"011000111",
  7138=>"001110101",
  7139=>"100100111",
  7140=>"010010000",
  7141=>"000110101",
  7142=>"000100001",
  7143=>"110010011",
  7144=>"011000000",
  7145=>"011001011",
  7146=>"111001100",
  7147=>"110110100",
  7148=>"000011101",
  7149=>"110000110",
  7150=>"110111011",
  7151=>"000011111",
  7152=>"011100100",
  7153=>"100011010",
  7154=>"011110111",
  7155=>"111011001",
  7156=>"100110000",
  7157=>"001100100",
  7158=>"000111111",
  7159=>"110010010",
  7160=>"010011010",
  7161=>"000100100",
  7162=>"001010011",
  7163=>"011001111",
  7164=>"110101010",
  7165=>"011001000",
  7166=>"000010100",
  7167=>"100010010",
  7168=>"000000100",
  7169=>"110011010",
  7170=>"110011000",
  7171=>"011111000",
  7172=>"001001100",
  7173=>"111111110",
  7174=>"010101001",
  7175=>"001000110",
  7176=>"111110111",
  7177=>"001000101",
  7178=>"001010001",
  7179=>"000001101",
  7180=>"011000111",
  7181=>"001100100",
  7182=>"100011110",
  7183=>"111001001",
  7184=>"110101111",
  7185=>"101000110",
  7186=>"100111011",
  7187=>"100001011",
  7188=>"101101000",
  7189=>"001010001",
  7190=>"111101101",
  7191=>"000000010",
  7192=>"011011011",
  7193=>"011010110",
  7194=>"011000101",
  7195=>"110000011",
  7196=>"111001001",
  7197=>"110000001",
  7198=>"001101010",
  7199=>"011011100",
  7200=>"100000110",
  7201=>"111001010",
  7202=>"001110011",
  7203=>"001000100",
  7204=>"000111001",
  7205=>"011011000",
  7206=>"100101100",
  7207=>"101001001",
  7208=>"010011111",
  7209=>"100001100",
  7210=>"101111110",
  7211=>"011000001",
  7212=>"001000001",
  7213=>"101111101",
  7214=>"100100110",
  7215=>"110010110",
  7216=>"011110111",
  7217=>"100110111",
  7218=>"000011100",
  7219=>"000100001",
  7220=>"010001001",
  7221=>"101001011",
  7222=>"000100111",
  7223=>"000010111",
  7224=>"101000110",
  7225=>"101100000",
  7226=>"001000101",
  7227=>"111001010",
  7228=>"011110111",
  7229=>"101010010",
  7230=>"001101000",
  7231=>"110101100",
  7232=>"110110110",
  7233=>"111011010",
  7234=>"011011001",
  7235=>"000001000",
  7236=>"000000001",
  7237=>"000010100",
  7238=>"001011101",
  7239=>"001101010",
  7240=>"001000000",
  7241=>"100011000",
  7242=>"110101100",
  7243=>"010010010",
  7244=>"010001111",
  7245=>"011010100",
  7246=>"101110101",
  7247=>"101000111",
  7248=>"111010101",
  7249=>"100010101",
  7250=>"101100101",
  7251=>"001010111",
  7252=>"111101100",
  7253=>"001000000",
  7254=>"011011101",
  7255=>"001010001",
  7256=>"100010010",
  7257=>"010000100",
  7258=>"110011101",
  7259=>"101000011",
  7260=>"110011101",
  7261=>"100110001",
  7262=>"111010000",
  7263=>"011001111",
  7264=>"001000000",
  7265=>"000101000",
  7266=>"110110110",
  7267=>"110010101",
  7268=>"010011111",
  7269=>"100101010",
  7270=>"010101100",
  7271=>"000111111",
  7272=>"000101111",
  7273=>"111011111",
  7274=>"011100101",
  7275=>"100101001",
  7276=>"001010110",
  7277=>"101110000",
  7278=>"111011000",
  7279=>"110010001",
  7280=>"001000010",
  7281=>"111100101",
  7282=>"010000111",
  7283=>"111101001",
  7284=>"110100000",
  7285=>"111111001",
  7286=>"010111000",
  7287=>"111101000",
  7288=>"010111011",
  7289=>"110100111",
  7290=>"111111111",
  7291=>"011000100",
  7292=>"100011110",
  7293=>"110100100",
  7294=>"001010001",
  7295=>"111001011",
  7296=>"000001111",
  7297=>"100110010",
  7298=>"010111011",
  7299=>"011010100",
  7300=>"110111100",
  7301=>"111111010",
  7302=>"001001101",
  7303=>"111001110",
  7304=>"001000010",
  7305=>"000001011",
  7306=>"001101110",
  7307=>"101100010",
  7308=>"110111000",
  7309=>"101110000",
  7310=>"000010011",
  7311=>"011100001",
  7312=>"111100011",
  7313=>"100000000",
  7314=>"101010101",
  7315=>"110111111",
  7316=>"001111101",
  7317=>"100111010",
  7318=>"010011001",
  7319=>"101101001",
  7320=>"011000001",
  7321=>"101001100",
  7322=>"110001101",
  7323=>"101110011",
  7324=>"101100100",
  7325=>"000010011",
  7326=>"111000010",
  7327=>"101000010",
  7328=>"111001100",
  7329=>"100011011",
  7330=>"001100000",
  7331=>"100101101",
  7332=>"011010101",
  7333=>"011001110",
  7334=>"010001101",
  7335=>"011011000",
  7336=>"011010010",
  7337=>"010000101",
  7338=>"101110111",
  7339=>"011101000",
  7340=>"000100100",
  7341=>"001101010",
  7342=>"111000010",
  7343=>"101010110",
  7344=>"001101110",
  7345=>"001111001",
  7346=>"100001000",
  7347=>"100110001",
  7348=>"000010000",
  7349=>"000101000",
  7350=>"011100111",
  7351=>"110000101",
  7352=>"000110011",
  7353=>"101101111",
  7354=>"110010110",
  7355=>"111111111",
  7356=>"110011100",
  7357=>"110000001",
  7358=>"100001101",
  7359=>"000001010",
  7360=>"111101110",
  7361=>"100101100",
  7362=>"000000110",
  7363=>"011110111",
  7364=>"001000110",
  7365=>"100101001",
  7366=>"110110110",
  7367=>"010001101",
  7368=>"100011011",
  7369=>"100111011",
  7370=>"000010110",
  7371=>"111011111",
  7372=>"111011101",
  7373=>"100011100",
  7374=>"000100000",
  7375=>"001011101",
  7376=>"110001010",
  7377=>"010100010",
  7378=>"101110111",
  7379=>"110011100",
  7380=>"110011111",
  7381=>"101010010",
  7382=>"010001011",
  7383=>"101000000",
  7384=>"010000010",
  7385=>"110111010",
  7386=>"100100101",
  7387=>"011101110",
  7388=>"011001111",
  7389=>"111111011",
  7390=>"101001101",
  7391=>"110111001",
  7392=>"000110010",
  7393=>"111100000",
  7394=>"000110100",
  7395=>"011011100",
  7396=>"101001000",
  7397=>"110111110",
  7398=>"011000101",
  7399=>"111110100",
  7400=>"001010100",
  7401=>"010111110",
  7402=>"011101111",
  7403=>"000011010",
  7404=>"001000001",
  7405=>"011010101",
  7406=>"101101010",
  7407=>"011101110",
  7408=>"111000010",
  7409=>"110001101",
  7410=>"010000000",
  7411=>"111100110",
  7412=>"000011011",
  7413=>"001010110",
  7414=>"101110011",
  7415=>"001101000",
  7416=>"100101110",
  7417=>"100110000",
  7418=>"011000001",
  7419=>"100001010",
  7420=>"001001100",
  7421=>"111000011",
  7422=>"111111100",
  7423=>"111110100",
  7424=>"010110001",
  7425=>"110010100",
  7426=>"100011101",
  7427=>"011011111",
  7428=>"110000001",
  7429=>"000100100",
  7430=>"100010010",
  7431=>"111000110",
  7432=>"101111100",
  7433=>"000011101",
  7434=>"101010101",
  7435=>"000000110",
  7436=>"010001100",
  7437=>"101001100",
  7438=>"000101110",
  7439=>"001000110",
  7440=>"001101001",
  7441=>"111011101",
  7442=>"010111111",
  7443=>"110101100",
  7444=>"010011010",
  7445=>"001100011",
  7446=>"101100011",
  7447=>"011010101",
  7448=>"110001000",
  7449=>"101100110",
  7450=>"000000100",
  7451=>"101111011",
  7452=>"101100110",
  7453=>"110111101",
  7454=>"010110101",
  7455=>"000001000",
  7456=>"000101000",
  7457=>"110000110",
  7458=>"101100001",
  7459=>"111111111",
  7460=>"010111001",
  7461=>"101001110",
  7462=>"001110100",
  7463=>"011001001",
  7464=>"010011111",
  7465=>"101111111",
  7466=>"101001110",
  7467=>"100000100",
  7468=>"000110000",
  7469=>"011111111",
  7470=>"111011111",
  7471=>"110010011",
  7472=>"101100011",
  7473=>"001000101",
  7474=>"100010100",
  7475=>"101101011",
  7476=>"001100111",
  7477=>"001000101",
  7478=>"100110101",
  7479=>"111110110",
  7480=>"000100100",
  7481=>"101111110",
  7482=>"001110010",
  7483=>"011110101",
  7484=>"101011111",
  7485=>"100001100",
  7486=>"100111111",
  7487=>"101100001",
  7488=>"000011000",
  7489=>"111001100",
  7490=>"010101001",
  7491=>"101111111",
  7492=>"101101000",
  7493=>"100001110",
  7494=>"000100110",
  7495=>"111000000",
  7496=>"111011011",
  7497=>"001000101",
  7498=>"111011110",
  7499=>"110010110",
  7500=>"000001011",
  7501=>"100001100",
  7502=>"011011001",
  7503=>"110101111",
  7504=>"010100010",
  7505=>"100010000",
  7506=>"110010110",
  7507=>"101100110",
  7508=>"000010001",
  7509=>"100010000",
  7510=>"001111001",
  7511=>"011011001",
  7512=>"001001001",
  7513=>"111011000",
  7514=>"110100111",
  7515=>"111000001",
  7516=>"101101110",
  7517=>"001000000",
  7518=>"000110010",
  7519=>"100101011",
  7520=>"110011010",
  7521=>"100110100",
  7522=>"110010100",
  7523=>"110011000",
  7524=>"000000110",
  7525=>"011111111",
  7526=>"001111100",
  7527=>"110111001",
  7528=>"101010000",
  7529=>"100000011",
  7530=>"111101101",
  7531=>"101010101",
  7532=>"000110100",
  7533=>"101100111",
  7534=>"011101101",
  7535=>"011100111",
  7536=>"100101101",
  7537=>"011100001",
  7538=>"000001101",
  7539=>"111110001",
  7540=>"100001110",
  7541=>"101011011",
  7542=>"001101001",
  7543=>"001001000",
  7544=>"000011100",
  7545=>"111110000",
  7546=>"011101000",
  7547=>"000100110",
  7548=>"111000000",
  7549=>"011110010",
  7550=>"000010101",
  7551=>"101010001",
  7552=>"100001111",
  7553=>"111111010",
  7554=>"101101010",
  7555=>"010001011",
  7556=>"001000100",
  7557=>"001000111",
  7558=>"101110011",
  7559=>"110111100",
  7560=>"001010000",
  7561=>"001000101",
  7562=>"000110010",
  7563=>"100101111",
  7564=>"010100010",
  7565=>"101011101",
  7566=>"000101100",
  7567=>"110101111",
  7568=>"100111001",
  7569=>"101101110",
  7570=>"011110110",
  7571=>"111000110",
  7572=>"011011000",
  7573=>"111110001",
  7574=>"001111110",
  7575=>"101011110",
  7576=>"000110100",
  7577=>"000111110",
  7578=>"000111110",
  7579=>"110000011",
  7580=>"010000110",
  7581=>"111110011",
  7582=>"101110011",
  7583=>"010000000",
  7584=>"101000011",
  7585=>"001011010",
  7586=>"011001101",
  7587=>"010000010",
  7588=>"100111010",
  7589=>"100000100",
  7590=>"101010011",
  7591=>"101011000",
  7592=>"110011111",
  7593=>"110000101",
  7594=>"001001111",
  7595=>"101110111",
  7596=>"000100000",
  7597=>"111110111",
  7598=>"110110010",
  7599=>"001001100",
  7600=>"100001110",
  7601=>"111001101",
  7602=>"101011111",
  7603=>"101110010",
  7604=>"010001001",
  7605=>"111111010",
  7606=>"011010011",
  7607=>"101100110",
  7608=>"111011010",
  7609=>"100010011",
  7610=>"000100000",
  7611=>"000100010",
  7612=>"100001010",
  7613=>"011111010",
  7614=>"100000110",
  7615=>"101000101",
  7616=>"100001101",
  7617=>"011001011",
  7618=>"111001001",
  7619=>"001111000",
  7620=>"100101100",
  7621=>"011100000",
  7622=>"000100000",
  7623=>"000100001",
  7624=>"001001000",
  7625=>"111011001",
  7626=>"110101010",
  7627=>"001000111",
  7628=>"110101001",
  7629=>"010000011",
  7630=>"111111111",
  7631=>"010101000",
  7632=>"011110001",
  7633=>"111111111",
  7634=>"110111110",
  7635=>"110011111",
  7636=>"011011000",
  7637=>"010111100",
  7638=>"101111101",
  7639=>"110101110",
  7640=>"000001010",
  7641=>"111001011",
  7642=>"101101100",
  7643=>"110110101",
  7644=>"101000010",
  7645=>"100101111",
  7646=>"100111101",
  7647=>"001100100",
  7648=>"101000001",
  7649=>"101110101",
  7650=>"110011001",
  7651=>"110101111",
  7652=>"010000001",
  7653=>"101011100",
  7654=>"011001100",
  7655=>"001001000",
  7656=>"110100010",
  7657=>"100111011",
  7658=>"100000101",
  7659=>"010000011",
  7660=>"111110101",
  7661=>"010001100",
  7662=>"000110010",
  7663=>"000111111",
  7664=>"010101010",
  7665=>"110110011",
  7666=>"001111001",
  7667=>"001100001",
  7668=>"111000010",
  7669=>"001110111",
  7670=>"011010000",
  7671=>"010001101",
  7672=>"111100100",
  7673=>"111100001",
  7674=>"100111000",
  7675=>"011111111",
  7676=>"000000100",
  7677=>"110101101",
  7678=>"100000000",
  7679=>"111110011",
  7680=>"111000011",
  7681=>"111000101",
  7682=>"101100100",
  7683=>"110101000",
  7684=>"101010011",
  7685=>"001100001",
  7686=>"110011111",
  7687=>"010011001",
  7688=>"100001000",
  7689=>"100000011",
  7690=>"010000000",
  7691=>"110001010",
  7692=>"100111000",
  7693=>"001001101",
  7694=>"010000111",
  7695=>"111100001",
  7696=>"000111000",
  7697=>"100100111",
  7698=>"111100101",
  7699=>"111111111",
  7700=>"101000001",
  7701=>"111110100",
  7702=>"111010101",
  7703=>"011111011",
  7704=>"110111000",
  7705=>"111001101",
  7706=>"010110011",
  7707=>"001010010",
  7708=>"100011011",
  7709=>"011010000",
  7710=>"100000010",
  7711=>"011011111",
  7712=>"001011011",
  7713=>"010110101",
  7714=>"100000101",
  7715=>"111110101",
  7716=>"001100100",
  7717=>"011010011",
  7718=>"111001100",
  7719=>"110011110",
  7720=>"010111111",
  7721=>"100011110",
  7722=>"100111011",
  7723=>"110001011",
  7724=>"001011010",
  7725=>"011011011",
  7726=>"010010010",
  7727=>"010001000",
  7728=>"110010011",
  7729=>"100011110",
  7730=>"111011000",
  7731=>"100101000",
  7732=>"011110111",
  7733=>"111001101",
  7734=>"111100100",
  7735=>"001000001",
  7736=>"111000100",
  7737=>"111000011",
  7738=>"001110001",
  7739=>"111101000",
  7740=>"000110111",
  7741=>"100001111",
  7742=>"100100011",
  7743=>"000011010",
  7744=>"000000001",
  7745=>"000001111",
  7746=>"011111111",
  7747=>"100011010",
  7748=>"101010110",
  7749=>"001000100",
  7750=>"110001111",
  7751=>"101111011",
  7752=>"100011100",
  7753=>"101000111",
  7754=>"100010100",
  7755=>"101100110",
  7756=>"000001101",
  7757=>"101001111",
  7758=>"010010001",
  7759=>"000011011",
  7760=>"111100111",
  7761=>"111010100",
  7762=>"000100100",
  7763=>"100011010",
  7764=>"000101011",
  7765=>"101100011",
  7766=>"011111011",
  7767=>"001001100",
  7768=>"011000000",
  7769=>"110010111",
  7770=>"100101111",
  7771=>"001111011",
  7772=>"011101100",
  7773=>"101101110",
  7774=>"001111101",
  7775=>"100011001",
  7776=>"110110001",
  7777=>"000000001",
  7778=>"001010011",
  7779=>"010000001",
  7780=>"111010000",
  7781=>"111101110",
  7782=>"000011011",
  7783=>"000011101",
  7784=>"010011010",
  7785=>"101010011",
  7786=>"010101101",
  7787=>"101101110",
  7788=>"001000011",
  7789=>"101000110",
  7790=>"010000100",
  7791=>"001110101",
  7792=>"111101111",
  7793=>"001010111",
  7794=>"010111010",
  7795=>"101110010",
  7796=>"101110001",
  7797=>"010000100",
  7798=>"111111001",
  7799=>"111111101",
  7800=>"111110111",
  7801=>"110101010",
  7802=>"001100001",
  7803=>"000101001",
  7804=>"011001111",
  7805=>"011010111",
  7806=>"100101111",
  7807=>"001000010",
  7808=>"111101101",
  7809=>"110111101",
  7810=>"101101011",
  7811=>"011110010",
  7812=>"011110000",
  7813=>"110111001",
  7814=>"111001111",
  7815=>"000000010",
  7816=>"000010101",
  7817=>"001010110",
  7818=>"100110111",
  7819=>"111110010",
  7820=>"011011101",
  7821=>"111101101",
  7822=>"011110001",
  7823=>"100000000",
  7824=>"000110000",
  7825=>"101001100",
  7826=>"011110111",
  7827=>"000000111",
  7828=>"000111100",
  7829=>"101101000",
  7830=>"111011001",
  7831=>"101001100",
  7832=>"111101111",
  7833=>"100111011",
  7834=>"100010101",
  7835=>"001110011",
  7836=>"111001110",
  7837=>"110100101",
  7838=>"000000110",
  7839=>"000111011",
  7840=>"111001110",
  7841=>"000010111",
  7842=>"011011010",
  7843=>"010111101",
  7844=>"000001110",
  7845=>"000000011",
  7846=>"101101101",
  7847=>"011100110",
  7848=>"111011000",
  7849=>"001000001",
  7850=>"111011010",
  7851=>"011001001",
  7852=>"100010000",
  7853=>"001100100",
  7854=>"111110000",
  7855=>"000001001",
  7856=>"010011111",
  7857=>"010011011",
  7858=>"001100100",
  7859=>"110000100",
  7860=>"101001010",
  7861=>"001111100",
  7862=>"011111101",
  7863=>"010100001",
  7864=>"110111110",
  7865=>"110010110",
  7866=>"000010100",
  7867=>"010000001",
  7868=>"101000000",
  7869=>"101101110",
  7870=>"011000101",
  7871=>"100101101",
  7872=>"100000111",
  7873=>"010110001",
  7874=>"110111111",
  7875=>"001000000",
  7876=>"010000110",
  7877=>"000011100",
  7878=>"011110100",
  7879=>"111011100",
  7880=>"101001101",
  7881=>"000001001",
  7882=>"101110100",
  7883=>"111110111",
  7884=>"100101011",
  7885=>"010100100",
  7886=>"001010111",
  7887=>"011101000",
  7888=>"001001100",
  7889=>"010100000",
  7890=>"100001001",
  7891=>"001010100",
  7892=>"110101111",
  7893=>"001011011",
  7894=>"110110111",
  7895=>"110001100",
  7896=>"110000000",
  7897=>"100101111",
  7898=>"011000000",
  7899=>"001011001",
  7900=>"001100011",
  7901=>"010101000",
  7902=>"001101011",
  7903=>"100011001",
  7904=>"011110011",
  7905=>"011111000",
  7906=>"011011001",
  7907=>"110001101",
  7908=>"000111000",
  7909=>"011011000",
  7910=>"001110100",
  7911=>"101011000",
  7912=>"110000010",
  7913=>"110000110",
  7914=>"011111010",
  7915=>"101001111",
  7916=>"010110000",
  7917=>"000110101",
  7918=>"001101000",
  7919=>"001111011",
  7920=>"010010110",
  7921=>"000011111",
  7922=>"110100110",
  7923=>"111001000",
  7924=>"011000001",
  7925=>"100101110",
  7926=>"011001010",
  7927=>"000000100",
  7928=>"111010110",
  7929=>"010011100",
  7930=>"101110001",
  7931=>"010100110",
  7932=>"001111111",
  7933=>"111100101",
  7934=>"001101110",
  7935=>"000000100",
  7936=>"001111010",
  7937=>"010110101",
  7938=>"101101000",
  7939=>"000000110",
  7940=>"100100000",
  7941=>"000100011",
  7942=>"001111110",
  7943=>"010111100",
  7944=>"011010110",
  7945=>"000000111",
  7946=>"111001110",
  7947=>"101001101",
  7948=>"110101001",
  7949=>"001011001",
  7950=>"111111111",
  7951=>"011001101",
  7952=>"001001011",
  7953=>"111010010",
  7954=>"101101010",
  7955=>"100010101",
  7956=>"101000011",
  7957=>"110111000",
  7958=>"011011101",
  7959=>"111100010",
  7960=>"001001000",
  7961=>"010101001",
  7962=>"011001101",
  7963=>"000010010",
  7964=>"111101000",
  7965=>"010110100",
  7966=>"100001111",
  7967=>"110000000",
  7968=>"111010010",
  7969=>"110010011",
  7970=>"000001000",
  7971=>"000100101",
  7972=>"111100010",
  7973=>"010101101",
  7974=>"111111000",
  7975=>"010001100",
  7976=>"101111001",
  7977=>"100001000",
  7978=>"111010000",
  7979=>"011110101",
  7980=>"010000010",
  7981=>"010010100",
  7982=>"110001010",
  7983=>"101101001",
  7984=>"000010101",
  7985=>"010010101",
  7986=>"001111010",
  7987=>"110111101",
  7988=>"101000110",
  7989=>"000110001",
  7990=>"010111101",
  7991=>"111001110",
  7992=>"011011001",
  7993=>"111000100",
  7994=>"001101100",
  7995=>"000110011",
  7996=>"111100110",
  7997=>"101011010",
  7998=>"000000100",
  7999=>"110110100",
  8000=>"110111101",
  8001=>"000001110",
  8002=>"101101111",
  8003=>"001101001",
  8004=>"111101110",
  8005=>"011100000",
  8006=>"001100101",
  8007=>"001001110",
  8008=>"010101110",
  8009=>"101001111",
  8010=>"000110101",
  8011=>"110101111",
  8012=>"111101000",
  8013=>"000110100",
  8014=>"001110100",
  8015=>"100110010",
  8016=>"101100100",
  8017=>"000100000",
  8018=>"001101011",
  8019=>"000101110",
  8020=>"110101110",
  8021=>"110001101",
  8022=>"100011100",
  8023=>"100001111",
  8024=>"111001101",
  8025=>"011100011",
  8026=>"010011011",
  8027=>"001011110",
  8028=>"010110011",
  8029=>"100000100",
  8030=>"110011101",
  8031=>"010010100",
  8032=>"010100010",
  8033=>"001110011",
  8034=>"001110010",
  8035=>"000100110",
  8036=>"100000000",
  8037=>"110101011",
  8038=>"110110011",
  8039=>"001101110",
  8040=>"110011001",
  8041=>"110000110",
  8042=>"111010000",
  8043=>"100100000",
  8044=>"100100010",
  8045=>"011011011",
  8046=>"000100101",
  8047=>"001000110",
  8048=>"100101110",
  8049=>"011010111",
  8050=>"101110010",
  8051=>"000111001",
  8052=>"100000000",
  8053=>"101000110",
  8054=>"110000011",
  8055=>"100110111",
  8056=>"000010011",
  8057=>"010010000",
  8058=>"101001111",
  8059=>"111000110",
  8060=>"101111111",
  8061=>"011100010",
  8062=>"111111111",
  8063=>"110000000",
  8064=>"000110110",
  8065=>"110010101",
  8066=>"111101011",
  8067=>"101101000",
  8068=>"101111011",
  8069=>"110101011",
  8070=>"100011101",
  8071=>"010100100",
  8072=>"000001010",
  8073=>"110100010",
  8074=>"111110010",
  8075=>"111111111",
  8076=>"101011111",
  8077=>"001011111",
  8078=>"010100000",
  8079=>"100100000",
  8080=>"101101001",
  8081=>"111010111",
  8082=>"100001001",
  8083=>"111101011",
  8084=>"000100000",
  8085=>"000011110",
  8086=>"000011010",
  8087=>"101100000",
  8088=>"011000100",
  8089=>"110000100",
  8090=>"111110100",
  8091=>"100010010",
  8092=>"110110010",
  8093=>"001100110",
  8094=>"111001111",
  8095=>"011000001",
  8096=>"111100000",
  8097=>"000101010",
  8098=>"110011110",
  8099=>"011001111",
  8100=>"101110110",
  8101=>"110110011",
  8102=>"111010110",
  8103=>"000000110",
  8104=>"010000000",
  8105=>"000001110",
  8106=>"011010100",
  8107=>"110010011",
  8108=>"110101100",
  8109=>"101100110",
  8110=>"100000001",
  8111=>"100000101",
  8112=>"001110000",
  8113=>"111110110",
  8114=>"001100110",
  8115=>"100001000",
  8116=>"000110100",
  8117=>"100110001",
  8118=>"010110011",
  8119=>"100011100",
  8120=>"011011011",
  8121=>"101011001",
  8122=>"110110111",
  8123=>"100110101",
  8124=>"100100101",
  8125=>"110000111",
  8126=>"101110110",
  8127=>"100001110",
  8128=>"011000111",
  8129=>"010010100",
  8130=>"110111010",
  8131=>"110011111",
  8132=>"000010001",
  8133=>"110001010",
  8134=>"111111111",
  8135=>"010001101",
  8136=>"000000000",
  8137=>"111100110",
  8138=>"111101011",
  8139=>"101001000",
  8140=>"111001001",
  8141=>"111010000",
  8142=>"111101111",
  8143=>"010000111",
  8144=>"110001101",
  8145=>"110011110",
  8146=>"101101111",
  8147=>"010000000",
  8148=>"011110010",
  8149=>"110001110",
  8150=>"101010110",
  8151=>"000000000",
  8152=>"110100010",
  8153=>"001011101",
  8154=>"010011100",
  8155=>"101110011",
  8156=>"010011110",
  8157=>"010010100",
  8158=>"010010000",
  8159=>"111111111",
  8160=>"011000100",
  8161=>"110110111",
  8162=>"010111100",
  8163=>"110011111",
  8164=>"101101011",
  8165=>"000000010",
  8166=>"000001001",
  8167=>"111110110",
  8168=>"001011111",
  8169=>"100100110",
  8170=>"100001011",
  8171=>"000011111",
  8172=>"000001111",
  8173=>"001101011",
  8174=>"101100110",
  8175=>"000110011",
  8176=>"101101010",
  8177=>"000100111",
  8178=>"101100100",
  8179=>"011110110",
  8180=>"110000010",
  8181=>"111101010",
  8182=>"111111111",
  8183=>"100101110",
  8184=>"011001111",
  8185=>"101110000",
  8186=>"001110111",
  8187=>"000000010",
  8188=>"100100001",
  8189=>"110110010",
  8190=>"001100011",
  8191=>"000101110",
  8192=>"010101011",
  8193=>"100111011",
  8194=>"010001111",
  8195=>"011011010",
  8196=>"010011110",
  8197=>"011001111",
  8198=>"101010000",
  8199=>"111001000",
  8200=>"111101100",
  8201=>"111001100",
  8202=>"001100001",
  8203=>"011111100",
  8204=>"000110001",
  8205=>"010101011",
  8206=>"101000001",
  8207=>"010100011",
  8208=>"111001110",
  8209=>"000001110",
  8210=>"101010100",
  8211=>"101111101",
  8212=>"111010100",
  8213=>"011000111",
  8214=>"101101111",
  8215=>"011000110",
  8216=>"100001010",
  8217=>"000101101",
  8218=>"011010100",
  8219=>"011111010",
  8220=>"011110110",
  8221=>"100011001",
  8222=>"011101000",
  8223=>"000011001",
  8224=>"011001011",
  8225=>"111101010",
  8226=>"010111110",
  8227=>"011100000",
  8228=>"000011001",
  8229=>"101010001",
  8230=>"011111011",
  8231=>"000110101",
  8232=>"001000000",
  8233=>"110110111",
  8234=>"101100101",
  8235=>"101110100",
  8236=>"011010011",
  8237=>"001011000",
  8238=>"101111110",
  8239=>"101100000",
  8240=>"011000011",
  8241=>"000010000",
  8242=>"111000100",
  8243=>"011011100",
  8244=>"101101011",
  8245=>"011100101",
  8246=>"001000000",
  8247=>"000100001",
  8248=>"111000011",
  8249=>"100100001",
  8250=>"111011100",
  8251=>"001000100",
  8252=>"110011111",
  8253=>"100000110",
  8254=>"000111011",
  8255=>"010101110",
  8256=>"000011001",
  8257=>"110101011",
  8258=>"101010100",
  8259=>"000110010",
  8260=>"010101000",
  8261=>"000110001",
  8262=>"100010011",
  8263=>"111110011",
  8264=>"001011001",
  8265=>"110010111",
  8266=>"101110010",
  8267=>"100001010",
  8268=>"110100011",
  8269=>"000010110",
  8270=>"000110000",
  8271=>"100101010",
  8272=>"111000110",
  8273=>"000001000",
  8274=>"101001011",
  8275=>"000110001",
  8276=>"111100001",
  8277=>"001110000",
  8278=>"000110110",
  8279=>"110110000",
  8280=>"101011101",
  8281=>"110110100",
  8282=>"010010100",
  8283=>"110001110",
  8284=>"010101000",
  8285=>"101101111",
  8286=>"100011000",
  8287=>"110101001",
  8288=>"110011001",
  8289=>"111011011",
  8290=>"001111111",
  8291=>"011010110",
  8292=>"011010100",
  8293=>"100111000",
  8294=>"001110101",
  8295=>"111011101",
  8296=>"100111001",
  8297=>"001100101",
  8298=>"001011111",
  8299=>"011101000",
  8300=>"001010011",
  8301=>"001000001",
  8302=>"101111110",
  8303=>"010110100",
  8304=>"011001000",
  8305=>"000100100",
  8306=>"010000001",
  8307=>"100101100",
  8308=>"101110010",
  8309=>"101110010",
  8310=>"000011011",
  8311=>"000000110",
  8312=>"011101010",
  8313=>"011011011",
  8314=>"001000010",
  8315=>"100111001",
  8316=>"001001011",
  8317=>"000111011",
  8318=>"110111101",
  8319=>"101100011",
  8320=>"010011010",
  8321=>"100110111",
  8322=>"110000001",
  8323=>"000000100",
  8324=>"001011101",
  8325=>"100100100",
  8326=>"011111010",
  8327=>"000010010",
  8328=>"101100111",
  8329=>"110011101",
  8330=>"001110000",
  8331=>"100001111",
  8332=>"000100101",
  8333=>"111000000",
  8334=>"000001001",
  8335=>"000111101",
  8336=>"101010001",
  8337=>"001100000",
  8338=>"110111111",
  8339=>"001110111",
  8340=>"001010001",
  8341=>"011100010",
  8342=>"100110110",
  8343=>"110110111",
  8344=>"110001000",
  8345=>"100111101",
  8346=>"000011101",
  8347=>"101011001",
  8348=>"000010000",
  8349=>"000100000",
  8350=>"110011100",
  8351=>"010011000",
  8352=>"001010001",
  8353=>"111100000",
  8354=>"111010000",
  8355=>"100011101",
  8356=>"101111111",
  8357=>"011001011",
  8358=>"111111001",
  8359=>"011111011",
  8360=>"110010001",
  8361=>"100000010",
  8362=>"000000000",
  8363=>"011100000",
  8364=>"010101111",
  8365=>"011011000",
  8366=>"010111110",
  8367=>"101010001",
  8368=>"100100010",
  8369=>"011111100",
  8370=>"011110011",
  8371=>"010111010",
  8372=>"111111100",
  8373=>"000111001",
  8374=>"100110000",
  8375=>"111001101",
  8376=>"011000110",
  8377=>"101011101",
  8378=>"101000001",
  8379=>"101100001",
  8380=>"110110000",
  8381=>"010011011",
  8382=>"000000111",
  8383=>"001100000",
  8384=>"110101001",
  8385=>"101111011",
  8386=>"000011111",
  8387=>"011100111",
  8388=>"001001111",
  8389=>"101001101",
  8390=>"101110000",
  8391=>"110000011",
  8392=>"010100011",
  8393=>"010100011",
  8394=>"001110000",
  8395=>"101011000",
  8396=>"011111111",
  8397=>"001111111",
  8398=>"011010011",
  8399=>"100100000",
  8400=>"001101000",
  8401=>"000101110",
  8402=>"010010001",
  8403=>"111111110",
  8404=>"100000001",
  8405=>"011100101",
  8406=>"101000010",
  8407=>"011000100",
  8408=>"011110000",
  8409=>"000110001",
  8410=>"110010000",
  8411=>"001011011",
  8412=>"010000000",
  8413=>"000000110",
  8414=>"110010001",
  8415=>"111110101",
  8416=>"011100011",
  8417=>"000110010",
  8418=>"000001110",
  8419=>"000110000",
  8420=>"110000111",
  8421=>"011000100",
  8422=>"110111111",
  8423=>"011101011",
  8424=>"011001001",
  8425=>"000001101",
  8426=>"010111100",
  8427=>"000011101",
  8428=>"000000001",
  8429=>"001101101",
  8430=>"110101101",
  8431=>"010001000",
  8432=>"011010011",
  8433=>"100101011",
  8434=>"110101110",
  8435=>"000010110",
  8436=>"001000010",
  8437=>"010010000",
  8438=>"111000100",
  8439=>"000110100",
  8440=>"101101001",
  8441=>"011111011",
  8442=>"000010000",
  8443=>"010011010",
  8444=>"011110001",
  8445=>"011010000",
  8446=>"111100000",
  8447=>"111010100",
  8448=>"010001101",
  8449=>"000001101",
  8450=>"000000010",
  8451=>"111111011",
  8452=>"011010001",
  8453=>"011010001",
  8454=>"001000110",
  8455=>"001000010",
  8456=>"111100100",
  8457=>"111000010",
  8458=>"111101100",
  8459=>"001111111",
  8460=>"000100101",
  8461=>"010101011",
  8462=>"000100011",
  8463=>"010100001",
  8464=>"100011101",
  8465=>"101110101",
  8466=>"111010111",
  8467=>"110101110",
  8468=>"100010000",
  8469=>"111010000",
  8470=>"111001000",
  8471=>"001010001",
  8472=>"110001110",
  8473=>"000010001",
  8474=>"101111110",
  8475=>"101101110",
  8476=>"000100000",
  8477=>"110001100",
  8478=>"000111110",
  8479=>"001000100",
  8480=>"010001000",
  8481=>"000110000",
  8482=>"111000111",
  8483=>"100000001",
  8484=>"000000111",
  8485=>"110010011",
  8486=>"011101011",
  8487=>"100010110",
  8488=>"010001011",
  8489=>"110011111",
  8490=>"100001010",
  8491=>"101100011",
  8492=>"000110000",
  8493=>"011110111",
  8494=>"111110111",
  8495=>"110010100",
  8496=>"100001010",
  8497=>"011111101",
  8498=>"101110111",
  8499=>"000000001",
  8500=>"101100101",
  8501=>"010000000",
  8502=>"111101101",
  8503=>"110000110",
  8504=>"001001000",
  8505=>"100110000",
  8506=>"011100011",
  8507=>"010101100",
  8508=>"110101110",
  8509=>"101001100",
  8510=>"101100100",
  8511=>"101110001",
  8512=>"111111011",
  8513=>"110100011",
  8514=>"010010001",
  8515=>"111001101",
  8516=>"100001110",
  8517=>"000100101",
  8518=>"000110100",
  8519=>"101000110",
  8520=>"100101100",
  8521=>"100101001",
  8522=>"011110110",
  8523=>"011100101",
  8524=>"100010010",
  8525=>"010110101",
  8526=>"111010011",
  8527=>"111101101",
  8528=>"000111011",
  8529=>"000101101",
  8530=>"110001011",
  8531=>"111011110",
  8532=>"011011010",
  8533=>"100100110",
  8534=>"010001011",
  8535=>"100010110",
  8536=>"001110001",
  8537=>"000110010",
  8538=>"000110011",
  8539=>"001001011",
  8540=>"100000100",
  8541=>"101011001",
  8542=>"111001011",
  8543=>"001011000",
  8544=>"110101100",
  8545=>"011000010",
  8546=>"111001001",
  8547=>"101001000",
  8548=>"011100010",
  8549=>"101111101",
  8550=>"101000001",
  8551=>"011010101",
  8552=>"000010000",
  8553=>"000111100",
  8554=>"110110010",
  8555=>"111111111",
  8556=>"100010101",
  8557=>"100111011",
  8558=>"111110011",
  8559=>"000111110",
  8560=>"111101011",
  8561=>"100001101",
  8562=>"100111100",
  8563=>"100111111",
  8564=>"011110000",
  8565=>"110111001",
  8566=>"100010110",
  8567=>"001111111",
  8568=>"111111000",
  8569=>"001000000",
  8570=>"010111110",
  8571=>"011100101",
  8572=>"011110100",
  8573=>"100100010",
  8574=>"100101011",
  8575=>"000101111",
  8576=>"101001100",
  8577=>"000010000",
  8578=>"100111010",
  8579=>"000101101",
  8580=>"101011010",
  8581=>"010011110",
  8582=>"110111010",
  8583=>"101000001",
  8584=>"101001010",
  8585=>"010100101",
  8586=>"001000000",
  8587=>"011101000",
  8588=>"010110110",
  8589=>"111110000",
  8590=>"010111100",
  8591=>"011110010",
  8592=>"011100000",
  8593=>"011001011",
  8594=>"001101100",
  8595=>"000011000",
  8596=>"111101110",
  8597=>"000101010",
  8598=>"110011011",
  8599=>"000011100",
  8600=>"010000011",
  8601=>"100111101",
  8602=>"111111111",
  8603=>"011001010",
  8604=>"110000100",
  8605=>"101110111",
  8606=>"101010101",
  8607=>"111010101",
  8608=>"011010111",
  8609=>"111110011",
  8610=>"110100110",
  8611=>"000001100",
  8612=>"000101000",
  8613=>"001000111",
  8614=>"110100100",
  8615=>"101000111",
  8616=>"101100011",
  8617=>"111011011",
  8618=>"110010011",
  8619=>"000010101",
  8620=>"000000000",
  8621=>"111110110",
  8622=>"011100000",
  8623=>"100111111",
  8624=>"100100101",
  8625=>"011011010",
  8626=>"111101110",
  8627=>"000001001",
  8628=>"111101001",
  8629=>"010010010",
  8630=>"001010010",
  8631=>"100100110",
  8632=>"101010110",
  8633=>"011110101",
  8634=>"111010100",
  8635=>"101010010",
  8636=>"001111111",
  8637=>"101000001",
  8638=>"010000011",
  8639=>"110001101",
  8640=>"011100010",
  8641=>"000000011",
  8642=>"111101011",
  8643=>"100111101",
  8644=>"100110001",
  8645=>"010101110",
  8646=>"011010001",
  8647=>"011100001",
  8648=>"111010111",
  8649=>"101101110",
  8650=>"111100010",
  8651=>"000010001",
  8652=>"011010100",
  8653=>"100111001",
  8654=>"110101001",
  8655=>"001010100",
  8656=>"111001101",
  8657=>"111101101",
  8658=>"001010110",
  8659=>"010111010",
  8660=>"101010000",
  8661=>"001111011",
  8662=>"100100100",
  8663=>"110011101",
  8664=>"010010000",
  8665=>"110010100",
  8666=>"101011010",
  8667=>"100110000",
  8668=>"001001110",
  8669=>"000001011",
  8670=>"111010111",
  8671=>"111100000",
  8672=>"111100111",
  8673=>"000110000",
  8674=>"101011001",
  8675=>"001000111",
  8676=>"000110010",
  8677=>"100110011",
  8678=>"010010111",
  8679=>"110001010",
  8680=>"110100101",
  8681=>"111100110",
  8682=>"100001001",
  8683=>"011101010",
  8684=>"010011101",
  8685=>"111001000",
  8686=>"011100110",
  8687=>"011001100",
  8688=>"011110010",
  8689=>"101100000",
  8690=>"110100100",
  8691=>"001100010",
  8692=>"000000011",
  8693=>"001110010",
  8694=>"111110000",
  8695=>"010000100",
  8696=>"010101001",
  8697=>"110001101",
  8698=>"000001001",
  8699=>"110110001",
  8700=>"000000000",
  8701=>"000101101",
  8702=>"111110001",
  8703=>"110101001",
  8704=>"101101000",
  8705=>"101000111",
  8706=>"000010011",
  8707=>"000100011",
  8708=>"010010101",
  8709=>"011011010",
  8710=>"100001001",
  8711=>"111101110",
  8712=>"110010000",
  8713=>"010110011",
  8714=>"001111111",
  8715=>"011000001",
  8716=>"111101100",
  8717=>"001111111",
  8718=>"000000000",
  8719=>"011001001",
  8720=>"111010111",
  8721=>"100110010",
  8722=>"101000100",
  8723=>"110001001",
  8724=>"000001010",
  8725=>"101011110",
  8726=>"110111100",
  8727=>"101110110",
  8728=>"000110001",
  8729=>"000101001",
  8730=>"010110001",
  8731=>"100111101",
  8732=>"100000100",
  8733=>"100110111",
  8734=>"101100001",
  8735=>"101101010",
  8736=>"100101001",
  8737=>"011111100",
  8738=>"111001011",
  8739=>"110001000",
  8740=>"000000101",
  8741=>"000111000",
  8742=>"010101010",
  8743=>"011100101",
  8744=>"110000110",
  8745=>"110110010",
  8746=>"100000110",
  8747=>"010111101",
  8748=>"011011111",
  8749=>"110000011",
  8750=>"011111110",
  8751=>"000000111",
  8752=>"100000111",
  8753=>"010000011",
  8754=>"100111110",
  8755=>"111110010",
  8756=>"001011111",
  8757=>"110111110",
  8758=>"110110101",
  8759=>"010111101",
  8760=>"111001111",
  8761=>"111101100",
  8762=>"011100010",
  8763=>"000111011",
  8764=>"111100101",
  8765=>"011001011",
  8766=>"000001001",
  8767=>"001100101",
  8768=>"111111101",
  8769=>"101111010",
  8770=>"010101100",
  8771=>"100100111",
  8772=>"010001110",
  8773=>"110101010",
  8774=>"101100000",
  8775=>"010011111",
  8776=>"000100001",
  8777=>"001110010",
  8778=>"101110110",
  8779=>"001011111",
  8780=>"000000110",
  8781=>"010010011",
  8782=>"100111100",
  8783=>"100001001",
  8784=>"101110110",
  8785=>"001100000",
  8786=>"100000101",
  8787=>"010110110",
  8788=>"101110110",
  8789=>"110011000",
  8790=>"011110010",
  8791=>"101100101",
  8792=>"111010011",
  8793=>"100011111",
  8794=>"111101000",
  8795=>"010011001",
  8796=>"101110111",
  8797=>"110101010",
  8798=>"010010001",
  8799=>"010101101",
  8800=>"110001001",
  8801=>"001000000",
  8802=>"010001100",
  8803=>"100101111",
  8804=>"111111000",
  8805=>"001010101",
  8806=>"011110101",
  8807=>"011001101",
  8808=>"111000110",
  8809=>"001110101",
  8810=>"111001001",
  8811=>"000111101",
  8812=>"010101001",
  8813=>"011011011",
  8814=>"000001001",
  8815=>"110100011",
  8816=>"011101110",
  8817=>"100110110",
  8818=>"010010110",
  8819=>"001101100",
  8820=>"000011000",
  8821=>"000010010",
  8822=>"111011100",
  8823=>"101001111",
  8824=>"111000010",
  8825=>"100100000",
  8826=>"000100011",
  8827=>"010100100",
  8828=>"110101100",
  8829=>"110001000",
  8830=>"101111101",
  8831=>"110010111",
  8832=>"010010111",
  8833=>"001101111",
  8834=>"001100000",
  8835=>"011111101",
  8836=>"010101001",
  8837=>"010110011",
  8838=>"110000110",
  8839=>"010010100",
  8840=>"110000111",
  8841=>"001000001",
  8842=>"011101011",
  8843=>"010100010",
  8844=>"000010101",
  8845=>"000001100",
  8846=>"101000101",
  8847=>"100000101",
  8848=>"001011111",
  8849=>"001001010",
  8850=>"010011101",
  8851=>"100111110",
  8852=>"001110110",
  8853=>"111101011",
  8854=>"111101001",
  8855=>"110110011",
  8856=>"101111110",
  8857=>"110111110",
  8858=>"110001001",
  8859=>"110001000",
  8860=>"110001010",
  8861=>"100101110",
  8862=>"110111110",
  8863=>"010110000",
  8864=>"100101110",
  8865=>"011010011",
  8866=>"000010110",
  8867=>"110111001",
  8868=>"010010111",
  8869=>"000010100",
  8870=>"111001111",
  8871=>"100101001",
  8872=>"101011110",
  8873=>"110110110",
  8874=>"100000010",
  8875=>"000101110",
  8876=>"001101000",
  8877=>"111111010",
  8878=>"100010111",
  8879=>"000111110",
  8880=>"100010011",
  8881=>"011011110",
  8882=>"101100110",
  8883=>"111111010",
  8884=>"001101000",
  8885=>"110011001",
  8886=>"000110011",
  8887=>"111001011",
  8888=>"110010101",
  8889=>"110100000",
  8890=>"010010010",
  8891=>"001001000",
  8892=>"011010100",
  8893=>"101011001",
  8894=>"000011011",
  8895=>"001111001",
  8896=>"110011111",
  8897=>"101011100",
  8898=>"011101100",
  8899=>"000000001",
  8900=>"101111000",
  8901=>"000110111",
  8902=>"001110010",
  8903=>"001001111",
  8904=>"001010110",
  8905=>"101001000",
  8906=>"010000010",
  8907=>"110100000",
  8908=>"001111101",
  8909=>"110110011",
  8910=>"100001011",
  8911=>"011001101",
  8912=>"100111110",
  8913=>"111001000",
  8914=>"101111111",
  8915=>"110010101",
  8916=>"110111011",
  8917=>"100100010",
  8918=>"001001011",
  8919=>"011101010",
  8920=>"100110100",
  8921=>"001010011",
  8922=>"110011011",
  8923=>"111011101",
  8924=>"100100111",
  8925=>"001111000",
  8926=>"100011010",
  8927=>"011100001",
  8928=>"000000000",
  8929=>"001110001",
  8930=>"001100100",
  8931=>"101011010",
  8932=>"100000010",
  8933=>"010001110",
  8934=>"101011101",
  8935=>"111111111",
  8936=>"010100110",
  8937=>"101010101",
  8938=>"101011011",
  8939=>"101111111",
  8940=>"111101010",
  8941=>"111101011",
  8942=>"110110101",
  8943=>"001010110",
  8944=>"100010001",
  8945=>"111111100",
  8946=>"011101001",
  8947=>"001111101",
  8948=>"101000111",
  8949=>"000100001",
  8950=>"111000010",
  8951=>"010010001",
  8952=>"101111100",
  8953=>"010110100",
  8954=>"110110001",
  8955=>"100110111",
  8956=>"111110000",
  8957=>"110111011",
  8958=>"111110100",
  8959=>"101010011",
  8960=>"110101000",
  8961=>"110100111",
  8962=>"000010010",
  8963=>"110100111",
  8964=>"011110011",
  8965=>"001101111",
  8966=>"001010100",
  8967=>"110010110",
  8968=>"011010111",
  8969=>"001011100",
  8970=>"011000101",
  8971=>"001000000",
  8972=>"110001100",
  8973=>"000101010",
  8974=>"010010001",
  8975=>"110111000",
  8976=>"010101100",
  8977=>"110111001",
  8978=>"101000000",
  8979=>"000010000",
  8980=>"100001011",
  8981=>"000111111",
  8982=>"000011100",
  8983=>"001100100",
  8984=>"110000001",
  8985=>"011010001",
  8986=>"110100001",
  8987=>"110100100",
  8988=>"111010010",
  8989=>"011010110",
  8990=>"111010100",
  8991=>"110111001",
  8992=>"100110111",
  8993=>"100110001",
  8994=>"111111001",
  8995=>"001110010",
  8996=>"001110001",
  8997=>"010111111",
  8998=>"010001101",
  8999=>"011010011",
  9000=>"010010000",
  9001=>"011011101",
  9002=>"111100001",
  9003=>"001010111",
  9004=>"000011011",
  9005=>"111011011",
  9006=>"110100001",
  9007=>"000111011",
  9008=>"000110100",
  9009=>"111101110",
  9010=>"011110011",
  9011=>"011101010",
  9012=>"010100110",
  9013=>"000101001",
  9014=>"000100100",
  9015=>"000111000",
  9016=>"011111100",
  9017=>"000000000",
  9018=>"101000001",
  9019=>"000011100",
  9020=>"100011010",
  9021=>"000000001",
  9022=>"000100110",
  9023=>"010111011",
  9024=>"000101101",
  9025=>"111110011",
  9026=>"101111100",
  9027=>"010111011",
  9028=>"000001010",
  9029=>"111111110",
  9030=>"011001100",
  9031=>"011000000",
  9032=>"001101110",
  9033=>"011001011",
  9034=>"110000000",
  9035=>"011010000",
  9036=>"101101111",
  9037=>"000000100",
  9038=>"100001001",
  9039=>"100110111",
  9040=>"000011101",
  9041=>"110111011",
  9042=>"000110010",
  9043=>"010001000",
  9044=>"010010000",
  9045=>"000110010",
  9046=>"110001001",
  9047=>"001101101",
  9048=>"111111100",
  9049=>"100011000",
  9050=>"111010010",
  9051=>"000011000",
  9052=>"010101110",
  9053=>"111000011",
  9054=>"000010101",
  9055=>"011111010",
  9056=>"100101000",
  9057=>"000101010",
  9058=>"000001101",
  9059=>"100001011",
  9060=>"110001100",
  9061=>"011000000",
  9062=>"001111011",
  9063=>"011011011",
  9064=>"010011011",
  9065=>"001100001",
  9066=>"011010110",
  9067=>"000000010",
  9068=>"011111110",
  9069=>"111110001",
  9070=>"011000100",
  9071=>"010011000",
  9072=>"001011101",
  9073=>"011001111",
  9074=>"000011110",
  9075=>"011111101",
  9076=>"001001101",
  9077=>"110001010",
  9078=>"100010110",
  9079=>"100011000",
  9080=>"100011010",
  9081=>"000101100",
  9082=>"001010100",
  9083=>"100100101",
  9084=>"111111001",
  9085=>"111011100",
  9086=>"011000010",
  9087=>"111011111",
  9088=>"011111111",
  9089=>"010111100",
  9090=>"100101001",
  9091=>"011100111",
  9092=>"000101001",
  9093=>"011010000",
  9094=>"101110111",
  9095=>"001111000",
  9096=>"010110111",
  9097=>"010111001",
  9098=>"011101001",
  9099=>"111111111",
  9100=>"011101011",
  9101=>"100101000",
  9102=>"111000011",
  9103=>"001001100",
  9104=>"001101010",
  9105=>"110011001",
  9106=>"010111110",
  9107=>"110001111",
  9108=>"100111001",
  9109=>"001010110",
  9110=>"000101101",
  9111=>"001101101",
  9112=>"100000001",
  9113=>"111101111",
  9114=>"111010000",
  9115=>"100101111",
  9116=>"000010100",
  9117=>"001110100",
  9118=>"001100011",
  9119=>"111101100",
  9120=>"111001000",
  9121=>"010101111",
  9122=>"011111101",
  9123=>"011111001",
  9124=>"101011001",
  9125=>"001100001",
  9126=>"111001101",
  9127=>"111001100",
  9128=>"111111010",
  9129=>"100010100",
  9130=>"101111011",
  9131=>"110000101",
  9132=>"101111001",
  9133=>"001110000",
  9134=>"000001001",
  9135=>"010000000",
  9136=>"100010000",
  9137=>"011101101",
  9138=>"010000010",
  9139=>"111010101",
  9140=>"001000101",
  9141=>"100110100",
  9142=>"110110111",
  9143=>"011100001",
  9144=>"000000110",
  9145=>"111110011",
  9146=>"000011100",
  9147=>"010101001",
  9148=>"111000101",
  9149=>"101011011",
  9150=>"010000110",
  9151=>"000011110",
  9152=>"100100010",
  9153=>"010000110",
  9154=>"100110011",
  9155=>"001000001",
  9156=>"100010000",
  9157=>"110110101",
  9158=>"111110111",
  9159=>"101000100",
  9160=>"010001100",
  9161=>"101110110",
  9162=>"101110001",
  9163=>"111111101",
  9164=>"111011111",
  9165=>"000000010",
  9166=>"001110111",
  9167=>"111110011",
  9168=>"010111000",
  9169=>"001110111",
  9170=>"111100011",
  9171=>"010011000",
  9172=>"110001100",
  9173=>"100101010",
  9174=>"111011101",
  9175=>"100000000",
  9176=>"101011111",
  9177=>"100110101",
  9178=>"010010010",
  9179=>"011011001",
  9180=>"000100000",
  9181=>"110110101",
  9182=>"011111011",
  9183=>"010110011",
  9184=>"101101010",
  9185=>"111110100",
  9186=>"001000000",
  9187=>"100001011",
  9188=>"000010110",
  9189=>"110111110",
  9190=>"101101000",
  9191=>"111010000",
  9192=>"001000110",
  9193=>"010100000",
  9194=>"101111000",
  9195=>"101111100",
  9196=>"010011010",
  9197=>"100110100",
  9198=>"010001001",
  9199=>"001001100",
  9200=>"101111111",
  9201=>"001000111",
  9202=>"100000110",
  9203=>"001100011",
  9204=>"111011110",
  9205=>"001111110",
  9206=>"110001111",
  9207=>"110111000",
  9208=>"011000010",
  9209=>"010000010",
  9210=>"110110100",
  9211=>"010110111",
  9212=>"111010001",
  9213=>"111110101",
  9214=>"010100111",
  9215=>"001111111",
  9216=>"100101010",
  9217=>"011011001",
  9218=>"100000000",
  9219=>"000011000",
  9220=>"011000100",
  9221=>"011000101",
  9222=>"001011111",
  9223=>"111100111",
  9224=>"001110110",
  9225=>"111101110",
  9226=>"011001101",
  9227=>"010000110",
  9228=>"010011000",
  9229=>"011000001",
  9230=>"101001101",
  9231=>"000010101",
  9232=>"000101011",
  9233=>"110010010",
  9234=>"100010011",
  9235=>"001000000",
  9236=>"000100110",
  9237=>"100001110",
  9238=>"010100111",
  9239=>"101000101",
  9240=>"010111001",
  9241=>"101001001",
  9242=>"001111101",
  9243=>"100110000",
  9244=>"100100011",
  9245=>"111111101",
  9246=>"000001010",
  9247=>"010001000",
  9248=>"111011111",
  9249=>"010000000",
  9250=>"000101010",
  9251=>"001010011",
  9252=>"000000111",
  9253=>"101110111",
  9254=>"000100000",
  9255=>"100101010",
  9256=>"111011110",
  9257=>"100010000",
  9258=>"000010010",
  9259=>"010001111",
  9260=>"101101011",
  9261=>"001101011",
  9262=>"010100100",
  9263=>"100110011",
  9264=>"010101010",
  9265=>"111001010",
  9266=>"000100100",
  9267=>"100100100",
  9268=>"100110110",
  9269=>"110101010",
  9270=>"110101011",
  9271=>"101100001",
  9272=>"011100101",
  9273=>"001110111",
  9274=>"010101001",
  9275=>"101001011",
  9276=>"111011101",
  9277=>"101001001",
  9278=>"011000101",
  9279=>"100110010",
  9280=>"011111010",
  9281=>"000110111",
  9282=>"101000001",
  9283=>"101100101",
  9284=>"101100000",
  9285=>"011011110",
  9286=>"110111011",
  9287=>"101110001",
  9288=>"101011011",
  9289=>"010011101",
  9290=>"011010001",
  9291=>"000001101",
  9292=>"011010010",
  9293=>"011001010",
  9294=>"101010011",
  9295=>"101110011",
  9296=>"001101011",
  9297=>"001001010",
  9298=>"001100110",
  9299=>"111100100",
  9300=>"110010000",
  9301=>"110110010",
  9302=>"100111110",
  9303=>"001011000",
  9304=>"101110010",
  9305=>"101100011",
  9306=>"111111011",
  9307=>"001011010",
  9308=>"010000000",
  9309=>"000010100",
  9310=>"011100001",
  9311=>"111011110",
  9312=>"110100010",
  9313=>"101110100",
  9314=>"010101110",
  9315=>"000110101",
  9316=>"010011011",
  9317=>"110011010",
  9318=>"111011001",
  9319=>"001101010",
  9320=>"010100011",
  9321=>"011110111",
  9322=>"010000011",
  9323=>"100010001",
  9324=>"110011100",
  9325=>"111100101",
  9326=>"000101000",
  9327=>"000011011",
  9328=>"111110110",
  9329=>"011110010",
  9330=>"100111000",
  9331=>"000100000",
  9332=>"111000111",
  9333=>"111011000",
  9334=>"100111100",
  9335=>"100100100",
  9336=>"000001001",
  9337=>"111110011",
  9338=>"010011110",
  9339=>"001011001",
  9340=>"011100100",
  9341=>"110111100",
  9342=>"111011101",
  9343=>"000010011",
  9344=>"100010000",
  9345=>"000100001",
  9346=>"000001111",
  9347=>"010001010",
  9348=>"101010111",
  9349=>"011000100",
  9350=>"010011111",
  9351=>"001101001",
  9352=>"001111000",
  9353=>"110010000",
  9354=>"110110000",
  9355=>"011100101",
  9356=>"110001000",
  9357=>"011100110",
  9358=>"001111000",
  9359=>"100011000",
  9360=>"011111101",
  9361=>"011000111",
  9362=>"100110000",
  9363=>"011101000",
  9364=>"111101001",
  9365=>"001101110",
  9366=>"001101111",
  9367=>"001001011",
  9368=>"000010111",
  9369=>"100010001",
  9370=>"111001010",
  9371=>"001110001",
  9372=>"010010111",
  9373=>"000001000",
  9374=>"100100100",
  9375=>"010100011",
  9376=>"001000000",
  9377=>"000001000",
  9378=>"100100000",
  9379=>"001010111",
  9380=>"001000111",
  9381=>"101111010",
  9382=>"011011010",
  9383=>"110110100",
  9384=>"101011001",
  9385=>"000101111",
  9386=>"011110110",
  9387=>"111000011",
  9388=>"001010000",
  9389=>"000010111",
  9390=>"001101110",
  9391=>"110101111",
  9392=>"110011000",
  9393=>"000011100",
  9394=>"000010111",
  9395=>"000011111",
  9396=>"001001110",
  9397=>"111111001",
  9398=>"110110110",
  9399=>"000010101",
  9400=>"101111000",
  9401=>"011110000",
  9402=>"100101100",
  9403=>"001000110",
  9404=>"111001110",
  9405=>"001000101",
  9406=>"000110010",
  9407=>"011101011",
  9408=>"011011100",
  9409=>"011000101",
  9410=>"011101010",
  9411=>"101101111",
  9412=>"111111001",
  9413=>"000000111",
  9414=>"010011010",
  9415=>"110001011",
  9416=>"101101110",
  9417=>"010111111",
  9418=>"010110100",
  9419=>"000111110",
  9420=>"101110010",
  9421=>"001111001",
  9422=>"011100011",
  9423=>"101101101",
  9424=>"100100011",
  9425=>"011101000",
  9426=>"001001001",
  9427=>"001001001",
  9428=>"111010101",
  9429=>"011111001",
  9430=>"000101100",
  9431=>"100110001",
  9432=>"100010001",
  9433=>"111110110",
  9434=>"011101111",
  9435=>"101111011",
  9436=>"111001000",
  9437=>"010100010",
  9438=>"000100000",
  9439=>"011101000",
  9440=>"100011010",
  9441=>"011101010",
  9442=>"101100110",
  9443=>"011001100",
  9444=>"111101111",
  9445=>"011011100",
  9446=>"011001010",
  9447=>"011010000",
  9448=>"101001110",
  9449=>"111111111",
  9450=>"111001101",
  9451=>"000011000",
  9452=>"001000000",
  9453=>"111101011",
  9454=>"110111000",
  9455=>"101111111",
  9456=>"000010011",
  9457=>"001010010",
  9458=>"100100101",
  9459=>"111001111",
  9460=>"111011101",
  9461=>"010110000",
  9462=>"111011011",
  9463=>"011010010",
  9464=>"110011011",
  9465=>"110001110",
  9466=>"101001011",
  9467=>"000101011",
  9468=>"110000000",
  9469=>"111101001",
  9470=>"010110010",
  9471=>"101110011",
  9472=>"110111010",
  9473=>"100100011",
  9474=>"010111110",
  9475=>"010110110",
  9476=>"110100010",
  9477=>"010101111",
  9478=>"000100000",
  9479=>"101010010",
  9480=>"110000001",
  9481=>"000111110",
  9482=>"011111111",
  9483=>"000110101",
  9484=>"011101011",
  9485=>"010001110",
  9486=>"110011111",
  9487=>"110001000",
  9488=>"110111110",
  9489=>"011100011",
  9490=>"111011001",
  9491=>"001000011",
  9492=>"001010011",
  9493=>"110101101",
  9494=>"000000011",
  9495=>"000011000",
  9496=>"111101101",
  9497=>"100010111",
  9498=>"110000100",
  9499=>"111100001",
  9500=>"100011011",
  9501=>"000100111",
  9502=>"110011000",
  9503=>"111100011",
  9504=>"001100001",
  9505=>"111101111",
  9506=>"100000111",
  9507=>"100110011",
  9508=>"000001110",
  9509=>"111011011",
  9510=>"111000001",
  9511=>"111111111",
  9512=>"001000011",
  9513=>"110100111",
  9514=>"101100000",
  9515=>"111100010",
  9516=>"111111000",
  9517=>"100110111",
  9518=>"011001010",
  9519=>"001101101",
  9520=>"000000000",
  9521=>"011010100",
  9522=>"100110000",
  9523=>"000001010",
  9524=>"110100001",
  9525=>"000111100",
  9526=>"001101100",
  9527=>"110110111",
  9528=>"011000101",
  9529=>"010101010",
  9530=>"010000010",
  9531=>"111110011",
  9532=>"001010001",
  9533=>"101111101",
  9534=>"111011001",
  9535=>"000110100",
  9536=>"011010111",
  9537=>"100010101",
  9538=>"111101100",
  9539=>"011001101",
  9540=>"101111100",
  9541=>"001011001",
  9542=>"111110100",
  9543=>"111001011",
  9544=>"011111011",
  9545=>"010100111",
  9546=>"111011110",
  9547=>"010101011",
  9548=>"011111010",
  9549=>"001111100",
  9550=>"111111111",
  9551=>"010010011",
  9552=>"111111110",
  9553=>"111110100",
  9554=>"111100010",
  9555=>"011011110",
  9556=>"111000011",
  9557=>"001111100",
  9558=>"011011001",
  9559=>"100011101",
  9560=>"000100110",
  9561=>"100110111",
  9562=>"010100011",
  9563=>"000010110",
  9564=>"010101000",
  9565=>"011001010",
  9566=>"000101110",
  9567=>"000001010",
  9568=>"010000001",
  9569=>"000011111",
  9570=>"011111110",
  9571=>"100110110",
  9572=>"000101111",
  9573=>"010010111",
  9574=>"001001110",
  9575=>"010110011",
  9576=>"101110111",
  9577=>"011110000",
  9578=>"010010110",
  9579=>"011111100",
  9580=>"101100101",
  9581=>"101011101",
  9582=>"001101011",
  9583=>"111000101",
  9584=>"001101101",
  9585=>"101011000",
  9586=>"111011010",
  9587=>"011011011",
  9588=>"100001101",
  9589=>"101101110",
  9590=>"010100000",
  9591=>"001011100",
  9592=>"000011010",
  9593=>"111001011",
  9594=>"100101111",
  9595=>"000000110",
  9596=>"110001010",
  9597=>"111100101",
  9598=>"010111010",
  9599=>"101100010",
  9600=>"111101101",
  9601=>"001011100",
  9602=>"001101000",
  9603=>"000011111",
  9604=>"011011011",
  9605=>"001111100",
  9606=>"011111011",
  9607=>"111001001",
  9608=>"011101101",
  9609=>"010111001",
  9610=>"011001111",
  9611=>"010111101",
  9612=>"001101010",
  9613=>"001100100",
  9614=>"000000101",
  9615=>"000000101",
  9616=>"000101100",
  9617=>"111010011",
  9618=>"101110010",
  9619=>"110001111",
  9620=>"100010100",
  9621=>"011101110",
  9622=>"110111001",
  9623=>"110101010",
  9624=>"000011010",
  9625=>"100100100",
  9626=>"101001000",
  9627=>"101000011",
  9628=>"111101011",
  9629=>"111101000",
  9630=>"110010011",
  9631=>"001010110",
  9632=>"000100000",
  9633=>"010110101",
  9634=>"101111011",
  9635=>"001010010",
  9636=>"101101011",
  9637=>"001001110",
  9638=>"110001110",
  9639=>"001110000",
  9640=>"110010101",
  9641=>"100110101",
  9642=>"001111001",
  9643=>"000011011",
  9644=>"001000010",
  9645=>"111111100",
  9646=>"001111010",
  9647=>"100101011",
  9648=>"101110011",
  9649=>"010010010",
  9650=>"100010010",
  9651=>"001010110",
  9652=>"001101001",
  9653=>"100101111",
  9654=>"000110110",
  9655=>"110110111",
  9656=>"101010111",
  9657=>"110111100",
  9658=>"000010010",
  9659=>"111101111",
  9660=>"110011100",
  9661=>"110010111",
  9662=>"000011000",
  9663=>"010100000",
  9664=>"111010000",
  9665=>"110110001",
  9666=>"100000100",
  9667=>"001001000",
  9668=>"101110000",
  9669=>"110111010",
  9670=>"011110001",
  9671=>"100010011",
  9672=>"100110011",
  9673=>"010111000",
  9674=>"110011010",
  9675=>"010111011",
  9676=>"010001010",
  9677=>"001010011",
  9678=>"010000101",
  9679=>"111010010",
  9680=>"101001111",
  9681=>"001001001",
  9682=>"111010100",
  9683=>"001100001",
  9684=>"000110010",
  9685=>"001100011",
  9686=>"110110110",
  9687=>"111010111",
  9688=>"111001110",
  9689=>"100101101",
  9690=>"011010001",
  9691=>"111111011",
  9692=>"011100001",
  9693=>"011011001",
  9694=>"011101111",
  9695=>"100101110",
  9696=>"000101101",
  9697=>"110011010",
  9698=>"110001011",
  9699=>"001010000",
  9700=>"111001000",
  9701=>"011010000",
  9702=>"100011000",
  9703=>"000101111",
  9704=>"111101100",
  9705=>"010101010",
  9706=>"110000000",
  9707=>"110100000",
  9708=>"111001100",
  9709=>"001111110",
  9710=>"100011000",
  9711=>"111110110",
  9712=>"111111000",
  9713=>"001101111",
  9714=>"001111100",
  9715=>"000001111",
  9716=>"110011110",
  9717=>"011010000",
  9718=>"101000110",
  9719=>"010101000",
  9720=>"111100011",
  9721=>"100110101",
  9722=>"110110010",
  9723=>"011000011",
  9724=>"000100100",
  9725=>"011010101",
  9726=>"110111001",
  9727=>"000001100",
  9728=>"010001100",
  9729=>"111100101",
  9730=>"000010101",
  9731=>"111001000",
  9732=>"100000111",
  9733=>"111101000",
  9734=>"001101101",
  9735=>"100101000",
  9736=>"001111001",
  9737=>"011000000",
  9738=>"111101010",
  9739=>"000001001",
  9740=>"110000100",
  9741=>"000001000",
  9742=>"111100000",
  9743=>"001101011",
  9744=>"011001100",
  9745=>"000111111",
  9746=>"011111111",
  9747=>"101001100",
  9748=>"101111100",
  9749=>"001100111",
  9750=>"100001010",
  9751=>"000000111",
  9752=>"010010110",
  9753=>"000111001",
  9754=>"111010010",
  9755=>"100001000",
  9756=>"111011011",
  9757=>"100101110",
  9758=>"110011000",
  9759=>"110010010",
  9760=>"011101001",
  9761=>"111110111",
  9762=>"011101010",
  9763=>"100101110",
  9764=>"101011100",
  9765=>"100111101",
  9766=>"111101111",
  9767=>"111000110",
  9768=>"001101110",
  9769=>"111010110",
  9770=>"110010111",
  9771=>"000111001",
  9772=>"101110010",
  9773=>"001000101",
  9774=>"101100111",
  9775=>"001011110",
  9776=>"111001111",
  9777=>"001000111",
  9778=>"111111000",
  9779=>"101011011",
  9780=>"010111101",
  9781=>"111011111",
  9782=>"010110000",
  9783=>"000101001",
  9784=>"111111110",
  9785=>"110100111",
  9786=>"000000001",
  9787=>"100100101",
  9788=>"001100101",
  9789=>"011011000",
  9790=>"101001101",
  9791=>"110001001",
  9792=>"101001001",
  9793=>"101010101",
  9794=>"111101111",
  9795=>"011010010",
  9796=>"011011111",
  9797=>"010000110",
  9798=>"011011001",
  9799=>"010010001",
  9800=>"111011101",
  9801=>"101110110",
  9802=>"111010000",
  9803=>"010000010",
  9804=>"100011000",
  9805=>"000011111",
  9806=>"000010011",
  9807=>"000110000",
  9808=>"100011000",
  9809=>"000000010",
  9810=>"001111001",
  9811=>"001000101",
  9812=>"110110100",
  9813=>"000110001",
  9814=>"100111100",
  9815=>"100110100",
  9816=>"000110110",
  9817=>"000011000",
  9818=>"101011110",
  9819=>"100100000",
  9820=>"111010111",
  9821=>"000101001",
  9822=>"110011111",
  9823=>"011111011",
  9824=>"100111000",
  9825=>"111010010",
  9826=>"111011011",
  9827=>"010111101",
  9828=>"011001101",
  9829=>"011001011",
  9830=>"010110011",
  9831=>"010011000",
  9832=>"000110010",
  9833=>"000000001",
  9834=>"101110101",
  9835=>"000011001",
  9836=>"111000011",
  9837=>"000011110",
  9838=>"000001010",
  9839=>"100110110",
  9840=>"101001111",
  9841=>"010110111",
  9842=>"110010111",
  9843=>"101001000",
  9844=>"011001110",
  9845=>"111101000",
  9846=>"100100111",
  9847=>"111101100",
  9848=>"101100110",
  9849=>"101000100",
  9850=>"010100100",
  9851=>"001010010",
  9852=>"111111000",
  9853=>"010110111",
  9854=>"100000101",
  9855=>"100110110",
  9856=>"111101011",
  9857=>"110000001",
  9858=>"001011011",
  9859=>"010100100",
  9860=>"001011111",
  9861=>"111001001",
  9862=>"101000001",
  9863=>"001100111",
  9864=>"101100001",
  9865=>"001001000",
  9866=>"001011000",
  9867=>"011011101",
  9868=>"111000001",
  9869=>"011010001",
  9870=>"000001000",
  9871=>"101011001",
  9872=>"111110010",
  9873=>"001011011",
  9874=>"001111011",
  9875=>"000111110",
  9876=>"100010101",
  9877=>"001011000",
  9878=>"100010110",
  9879=>"011001000",
  9880=>"110101010",
  9881=>"111011101",
  9882=>"010000111",
  9883=>"100010100",
  9884=>"111101011",
  9885=>"001101111",
  9886=>"110101100",
  9887=>"111001101",
  9888=>"000111011",
  9889=>"010100010",
  9890=>"101010011",
  9891=>"111000110",
  9892=>"011011011",
  9893=>"001101010",
  9894=>"110010110",
  9895=>"011011001",
  9896=>"110001101",
  9897=>"100001000",
  9898=>"100001001",
  9899=>"101110001",
  9900=>"111010010",
  9901=>"000111101",
  9902=>"101110000",
  9903=>"000100001",
  9904=>"011110010",
  9905=>"100000000",
  9906=>"111111001",
  9907=>"011101001",
  9908=>"110101010",
  9909=>"010000111",
  9910=>"110111111",
  9911=>"101010111",
  9912=>"110100010",
  9913=>"010110000",
  9914=>"101100001",
  9915=>"101001111",
  9916=>"100000000",
  9917=>"011001011",
  9918=>"001010000",
  9919=>"110110011",
  9920=>"101001011",
  9921=>"000101111",
  9922=>"001001000",
  9923=>"011101111",
  9924=>"011101000",
  9925=>"101000011",
  9926=>"101010101",
  9927=>"111101011",
  9928=>"010010101",
  9929=>"010111110",
  9930=>"111011001",
  9931=>"110110110",
  9932=>"001110011",
  9933=>"011110001",
  9934=>"101010101",
  9935=>"001010111",
  9936=>"110101011",
  9937=>"001111001",
  9938=>"010001100",
  9939=>"100111100",
  9940=>"110110101",
  9941=>"010000000",
  9942=>"000001001",
  9943=>"010111100",
  9944=>"111100001",
  9945=>"110100010",
  9946=>"001001001",
  9947=>"011011001",
  9948=>"110111110",
  9949=>"100100101",
  9950=>"011011000",
  9951=>"110001011",
  9952=>"000011110",
  9953=>"011100100",
  9954=>"100011010",
  9955=>"111110100",
  9956=>"101111011",
  9957=>"111001111",
  9958=>"011010000",
  9959=>"001111010",
  9960=>"110000000",
  9961=>"011101000",
  9962=>"110000110",
  9963=>"000101111",
  9964=>"100000000",
  9965=>"111111011",
  9966=>"111100110",
  9967=>"010010101",
  9968=>"001001000",
  9969=>"111111011",
  9970=>"000100100",
  9971=>"100000010",
  9972=>"010100110",
  9973=>"100111011",
  9974=>"100101010",
  9975=>"111111011",
  9976=>"101000001",
  9977=>"110101110",
  9978=>"001111110",
  9979=>"011000111",
  9980=>"001111111",
  9981=>"001011101",
  9982=>"111100001",
  9983=>"000100100",
  9984=>"100011010",
  9985=>"110000110",
  9986=>"100110011",
  9987=>"011000110",
  9988=>"001001101",
  9989=>"001000111",
  9990=>"011001011",
  9991=>"001111111",
  9992=>"001011101",
  9993=>"111100101",
  9994=>"000010011",
  9995=>"111000100",
  9996=>"110110010",
  9997=>"111110100",
  9998=>"001111101",
  9999=>"001011011",
  10000=>"000101000",
  10001=>"001001001",
  10002=>"011111101",
  10003=>"110001111",
  10004=>"101101001",
  10005=>"010110101",
  10006=>"100111011",
  10007=>"100011001",
  10008=>"111101001",
  10009=>"001111001",
  10010=>"100001101",
  10011=>"100100010",
  10012=>"111111010",
  10013=>"101010100",
  10014=>"011000010",
  10015=>"001101001",
  10016=>"111001110",
  10017=>"110000111",
  10018=>"111110010",
  10019=>"110100101",
  10020=>"010111000",
  10021=>"101111100",
  10022=>"111010110",
  10023=>"010000100",
  10024=>"111111011",
  10025=>"100001100",
  10026=>"011101011",
  10027=>"100010100",
  10028=>"010011011",
  10029=>"111101111",
  10030=>"101101100",
  10031=>"111011100",
  10032=>"000001001",
  10033=>"111100000",
  10034=>"000100101",
  10035=>"110100111",
  10036=>"100100101",
  10037=>"110010100",
  10038=>"000110011",
  10039=>"101100000",
  10040=>"000110111",
  10041=>"011001001",
  10042=>"110110011",
  10043=>"011111011",
  10044=>"000100100",
  10045=>"011001000",
  10046=>"101000010",
  10047=>"001101011",
  10048=>"000010010",
  10049=>"101111101",
  10050=>"000000000",
  10051=>"100000100",
  10052=>"101010010",
  10053=>"100010110",
  10054=>"101000000",
  10055=>"101011100",
  10056=>"010001010",
  10057=>"100101111",
  10058=>"000100100",
  10059=>"001101011",
  10060=>"111101110",
  10061=>"011111101",
  10062=>"111001000",
  10063=>"000010011",
  10064=>"000011100",
  10065=>"001000010",
  10066=>"111111001",
  10067=>"111000010",
  10068=>"010100101",
  10069=>"000100100",
  10070=>"101000101",
  10071=>"000010010",
  10072=>"001010000",
  10073=>"001100010",
  10074=>"100010111",
  10075=>"010100100",
  10076=>"111011111",
  10077=>"010111010",
  10078=>"111001110",
  10079=>"000010100",
  10080=>"001101100",
  10081=>"111110111",
  10082=>"000111110",
  10083=>"011011100",
  10084=>"000011010",
  10085=>"001101010",
  10086=>"111010110",
  10087=>"110111000",
  10088=>"110001001",
  10089=>"001101110",
  10090=>"100111010",
  10091=>"001100000",
  10092=>"101110111",
  10093=>"011000110",
  10094=>"001100000",
  10095=>"001011011",
  10096=>"101101110",
  10097=>"110110111",
  10098=>"111011111",
  10099=>"111001000",
  10100=>"100011000",
  10101=>"000001100",
  10102=>"111001101",
  10103=>"000000011",
  10104=>"000011011",
  10105=>"011001111",
  10106=>"000101010",
  10107=>"000011101",
  10108=>"011000000",
  10109=>"111111110",
  10110=>"100001111",
  10111=>"110000110",
  10112=>"011011011",
  10113=>"101001100",
  10114=>"001010100",
  10115=>"000101111",
  10116=>"011011001",
  10117=>"111001101",
  10118=>"011100111",
  10119=>"100111001",
  10120=>"101000111",
  10121=>"101001001",
  10122=>"000101111",
  10123=>"110111011",
  10124=>"110001010",
  10125=>"111011110",
  10126=>"111001100",
  10127=>"010010110",
  10128=>"001011010",
  10129=>"010010101",
  10130=>"010000000",
  10131=>"111111001",
  10132=>"111011011",
  10133=>"000000011",
  10134=>"011001011",
  10135=>"101100111",
  10136=>"110101111",
  10137=>"011010001",
  10138=>"000111011",
  10139=>"100011110",
  10140=>"111111001",
  10141=>"111010001",
  10142=>"101111101",
  10143=>"101100110",
  10144=>"111010010",
  10145=>"111011101",
  10146=>"011010110",
  10147=>"100100001",
  10148=>"110111011",
  10149=>"101011001",
  10150=>"000100101",
  10151=>"111001110",
  10152=>"111010000",
  10153=>"010001000",
  10154=>"000100110",
  10155=>"101011110",
  10156=>"010001111",
  10157=>"111111000",
  10158=>"110111110",
  10159=>"111111101",
  10160=>"110001100",
  10161=>"100110011",
  10162=>"000011011",
  10163=>"101101010",
  10164=>"110010001",
  10165=>"010011101",
  10166=>"001000011",
  10167=>"111111010",
  10168=>"101111110",
  10169=>"100001001",
  10170=>"011110101",
  10171=>"111101011",
  10172=>"111000110",
  10173=>"011010101",
  10174=>"101011010",
  10175=>"111111001",
  10176=>"101101000",
  10177=>"100000010",
  10178=>"001011010",
  10179=>"111010011",
  10180=>"110011010",
  10181=>"100010111",
  10182=>"110110111",
  10183=>"000111000",
  10184=>"110100100",
  10185=>"111101000",
  10186=>"000100100",
  10187=>"100010000",
  10188=>"100100100",
  10189=>"001010001",
  10190=>"100110000",
  10191=>"001000101",
  10192=>"111011100",
  10193=>"010100100",
  10194=>"010101001",
  10195=>"010001111",
  10196=>"010011000",
  10197=>"101011110",
  10198=>"000010001",
  10199=>"010101111",
  10200=>"011110100",
  10201=>"110101010",
  10202=>"010000110",
  10203=>"110000010",
  10204=>"010110110",
  10205=>"001101010",
  10206=>"000011001",
  10207=>"101011001",
  10208=>"100011001",
  10209=>"001000000",
  10210=>"110111100",
  10211=>"011010011",
  10212=>"011001011",
  10213=>"110110001",
  10214=>"110101100",
  10215=>"110010000",
  10216=>"111111110",
  10217=>"110100111",
  10218=>"110011001",
  10219=>"001101010",
  10220=>"011011111",
  10221=>"001101100",
  10222=>"000010000",
  10223=>"000100111",
  10224=>"001001000",
  10225=>"111011101",
  10226=>"110010010",
  10227=>"100101011",
  10228=>"011011010",
  10229=>"011110110",
  10230=>"101010011",
  10231=>"100110111",
  10232=>"001111110",
  10233=>"110100100",
  10234=>"111010100",
  10235=>"000000101",
  10236=>"001100100",
  10237=>"010011001",
  10238=>"000000101",
  10239=>"001100010",
  10240=>"111010000",
  10241=>"110011100",
  10242=>"111010010",
  10243=>"001001110",
  10244=>"101111011",
  10245=>"000011101",
  10246=>"101000111",
  10247=>"100011010",
  10248=>"010110100",
  10249=>"110110110",
  10250=>"110010010",
  10251=>"111011011",
  10252=>"111111101",
  10253=>"110010011",
  10254=>"011100010",
  10255=>"000111000",
  10256=>"011111010",
  10257=>"000001000",
  10258=>"111011010",
  10259=>"101001111",
  10260=>"010100111",
  10261=>"111110110",
  10262=>"111011010",
  10263=>"111000011",
  10264=>"110110000",
  10265=>"101011011",
  10266=>"000010100",
  10267=>"010110001",
  10268=>"101110111",
  10269=>"011111011",
  10270=>"001110111",
  10271=>"111010011",
  10272=>"011010011",
  10273=>"101110001",
  10274=>"111000010",
  10275=>"010001001",
  10276=>"101001010",
  10277=>"100011110",
  10278=>"001000000",
  10279=>"011101000",
  10280=>"111111101",
  10281=>"111100001",
  10282=>"100000111",
  10283=>"111010101",
  10284=>"100001100",
  10285=>"011001110",
  10286=>"011111111",
  10287=>"010110111",
  10288=>"111000101",
  10289=>"100100101",
  10290=>"101000000",
  10291=>"100011111",
  10292=>"010111001",
  10293=>"000010100",
  10294=>"100001000",
  10295=>"100101010",
  10296=>"100001100",
  10297=>"110001001",
  10298=>"010011111",
  10299=>"111001110",
  10300=>"001100100",
  10301=>"110110001",
  10302=>"111110110",
  10303=>"100000101",
  10304=>"001011110",
  10305=>"010010110",
  10306=>"111001110",
  10307=>"001111100",
  10308=>"110100001",
  10309=>"111110011",
  10310=>"011111011",
  10311=>"100010001",
  10312=>"011001000",
  10313=>"010001101",
  10314=>"100001100",
  10315=>"001101110",
  10316=>"110001000",
  10317=>"000011001",
  10318=>"001101010",
  10319=>"101111011",
  10320=>"001010110",
  10321=>"000000111",
  10322=>"000010010",
  10323=>"100001010",
  10324=>"000000100",
  10325=>"010100000",
  10326=>"001100000",
  10327=>"111111100",
  10328=>"000101101",
  10329=>"100011111",
  10330=>"010011001",
  10331=>"010010001",
  10332=>"011010011",
  10333=>"010010000",
  10334=>"101100101",
  10335=>"110110011",
  10336=>"000000100",
  10337=>"011001010",
  10338=>"001000001",
  10339=>"011011111",
  10340=>"010101110",
  10341=>"000000000",
  10342=>"000011110",
  10343=>"010001010",
  10344=>"001010000",
  10345=>"111111011",
  10346=>"111110010",
  10347=>"100001011",
  10348=>"111010000",
  10349=>"110001001",
  10350=>"100001100",
  10351=>"011011010",
  10352=>"101110100",
  10353=>"000111011",
  10354=>"000011000",
  10355=>"000010100",
  10356=>"010001100",
  10357=>"111110100",
  10358=>"000100111",
  10359=>"000100110",
  10360=>"010111101",
  10361=>"111100010",
  10362=>"010001010",
  10363=>"010101001",
  10364=>"011110010",
  10365=>"010100101",
  10366=>"111111000",
  10367=>"110010110",
  10368=>"111001111",
  10369=>"110000011",
  10370=>"101100000",
  10371=>"011011011",
  10372=>"011101010",
  10373=>"111000000",
  10374=>"101111100",
  10375=>"000000001",
  10376=>"111100101",
  10377=>"010100101",
  10378=>"001010011",
  10379=>"100011111",
  10380=>"010000001",
  10381=>"011011001",
  10382=>"101101110",
  10383=>"101010110",
  10384=>"110000001",
  10385=>"011100010",
  10386=>"101010101",
  10387=>"100001001",
  10388=>"000011000",
  10389=>"101100000",
  10390=>"111011011",
  10391=>"000111000",
  10392=>"110001101",
  10393=>"011111011",
  10394=>"000100000",
  10395=>"111011111",
  10396=>"100110101",
  10397=>"000101001",
  10398=>"110001101",
  10399=>"010111010",
  10400=>"000101000",
  10401=>"001100001",
  10402=>"111110110",
  10403=>"011011110",
  10404=>"101100100",
  10405=>"001000110",
  10406=>"110001011",
  10407=>"011101001",
  10408=>"111011111",
  10409=>"011010111",
  10410=>"110000110",
  10411=>"101000000",
  10412=>"010110101",
  10413=>"111111101",
  10414=>"001011101",
  10415=>"000000000",
  10416=>"110110000",
  10417=>"000000000",
  10418=>"100111010",
  10419=>"000000110",
  10420=>"111011000",
  10421=>"101000110",
  10422=>"110100010",
  10423=>"011001100",
  10424=>"011010000",
  10425=>"110110100",
  10426=>"011110001",
  10427=>"111110100",
  10428=>"110100101",
  10429=>"110001111",
  10430=>"011101010",
  10431=>"000111110",
  10432=>"000100000",
  10433=>"100111000",
  10434=>"000001100",
  10435=>"101100000",
  10436=>"000000011",
  10437=>"001001010",
  10438=>"111101101",
  10439=>"101110011",
  10440=>"001000000",
  10441=>"000101011",
  10442=>"111110110",
  10443=>"111101011",
  10444=>"000111001",
  10445=>"111010001",
  10446=>"011010001",
  10447=>"011001010",
  10448=>"110100011",
  10449=>"001001010",
  10450=>"001010110",
  10451=>"100100010",
  10452=>"010001110",
  10453=>"010100100",
  10454=>"001110111",
  10455=>"100010110",
  10456=>"000001101",
  10457=>"010011001",
  10458=>"100001000",
  10459=>"101110000",
  10460=>"110101011",
  10461=>"100111011",
  10462=>"101111110",
  10463=>"000100100",
  10464=>"100100111",
  10465=>"001111110",
  10466=>"101110111",
  10467=>"110000001",
  10468=>"101101001",
  10469=>"100010110",
  10470=>"001000001",
  10471=>"011011100",
  10472=>"101000111",
  10473=>"111110110",
  10474=>"110000000",
  10475=>"100001110",
  10476=>"001110110",
  10477=>"001001010",
  10478=>"011110000",
  10479=>"001101101",
  10480=>"110100100",
  10481=>"010000101",
  10482=>"001001100",
  10483=>"110000010",
  10484=>"011110100",
  10485=>"100000010",
  10486=>"010001011",
  10487=>"011010100",
  10488=>"010000111",
  10489=>"000011110",
  10490=>"001010011",
  10491=>"010111100",
  10492=>"000100011",
  10493=>"000011010",
  10494=>"010011001",
  10495=>"000100101",
  10496=>"010010101",
  10497=>"001111100",
  10498=>"000010111",
  10499=>"110001001",
  10500=>"100111000",
  10501=>"010000010",
  10502=>"001001011",
  10503=>"100000111",
  10504=>"000101010",
  10505=>"010000101",
  10506=>"111011001",
  10507=>"101000011",
  10508=>"000001000",
  10509=>"011000101",
  10510=>"010000001",
  10511=>"000111100",
  10512=>"111110010",
  10513=>"101110110",
  10514=>"001100011",
  10515=>"111000110",
  10516=>"101110001",
  10517=>"011011111",
  10518=>"011111011",
  10519=>"101000101",
  10520=>"101111001",
  10521=>"000001001",
  10522=>"110001000",
  10523=>"100000100",
  10524=>"000011010",
  10525=>"110001100",
  10526=>"111100011",
  10527=>"111100001",
  10528=>"001000010",
  10529=>"100001000",
  10530=>"001010111",
  10531=>"101100110",
  10532=>"111110010",
  10533=>"010000000",
  10534=>"100000011",
  10535=>"000000101",
  10536=>"111011000",
  10537=>"100011101",
  10538=>"101000101",
  10539=>"100011010",
  10540=>"101101100",
  10541=>"011100000",
  10542=>"111001011",
  10543=>"110011111",
  10544=>"001100000",
  10545=>"011101100",
  10546=>"110010111",
  10547=>"001010000",
  10548=>"001110111",
  10549=>"001110011",
  10550=>"011010001",
  10551=>"000101110",
  10552=>"100010010",
  10553=>"110111111",
  10554=>"111001000",
  10555=>"110001001",
  10556=>"110001001",
  10557=>"011011101",
  10558=>"101100000",
  10559=>"010001010",
  10560=>"011101100",
  10561=>"000011010",
  10562=>"111111010",
  10563=>"101001101",
  10564=>"100110011",
  10565=>"100011010",
  10566=>"110100110",
  10567=>"011001010",
  10568=>"110010101",
  10569=>"001100100",
  10570=>"011100011",
  10571=>"000010000",
  10572=>"100111000",
  10573=>"100100111",
  10574=>"100001011",
  10575=>"101010001",
  10576=>"010100111",
  10577=>"101101100",
  10578=>"101011011",
  10579=>"011011001",
  10580=>"011110000",
  10581=>"010000011",
  10582=>"011100101",
  10583=>"000010110",
  10584=>"001000010",
  10585=>"111101011",
  10586=>"110000100",
  10587=>"101001110",
  10588=>"100011100",
  10589=>"110001111",
  10590=>"000000000",
  10591=>"001011010",
  10592=>"111111111",
  10593=>"111010010",
  10594=>"001001100",
  10595=>"101011100",
  10596=>"010001110",
  10597=>"110000011",
  10598=>"100100000",
  10599=>"001011000",
  10600=>"110110000",
  10601=>"001000010",
  10602=>"101001001",
  10603=>"111101001",
  10604=>"101011010",
  10605=>"100101011",
  10606=>"000100110",
  10607=>"100001001",
  10608=>"000010000",
  10609=>"000000010",
  10610=>"100101001",
  10611=>"100001110",
  10612=>"010001000",
  10613=>"000001111",
  10614=>"011010101",
  10615=>"010000100",
  10616=>"111100100",
  10617=>"011101110",
  10618=>"011010001",
  10619=>"110001101",
  10620=>"100010010",
  10621=>"100011110",
  10622=>"001110101",
  10623=>"110010001",
  10624=>"000001011",
  10625=>"000011101",
  10626=>"001111001",
  10627=>"001001001",
  10628=>"110011010",
  10629=>"011000000",
  10630=>"100000110",
  10631=>"101100001",
  10632=>"111010001",
  10633=>"111101010",
  10634=>"011101000",
  10635=>"001001001",
  10636=>"110000000",
  10637=>"000010001",
  10638=>"110000010",
  10639=>"110111000",
  10640=>"001111011",
  10641=>"010110111",
  10642=>"100000111",
  10643=>"011100011",
  10644=>"000010100",
  10645=>"110110110",
  10646=>"100011010",
  10647=>"000010110",
  10648=>"011001111",
  10649=>"101000001",
  10650=>"010011010",
  10651=>"010011001",
  10652=>"111000100",
  10653=>"011110010",
  10654=>"110101110",
  10655=>"011001100",
  10656=>"101010100",
  10657=>"110100100",
  10658=>"010100011",
  10659=>"010011010",
  10660=>"001101110",
  10661=>"110000111",
  10662=>"100001010",
  10663=>"010010101",
  10664=>"100100000",
  10665=>"010100101",
  10666=>"111110000",
  10667=>"011001001",
  10668=>"000111101",
  10669=>"010100000",
  10670=>"100111010",
  10671=>"101011000",
  10672=>"110110000",
  10673=>"011000100",
  10674=>"010011010",
  10675=>"100010011",
  10676=>"110000010",
  10677=>"001100010",
  10678=>"111010011",
  10679=>"101111011",
  10680=>"010100001",
  10681=>"101101111",
  10682=>"100010010",
  10683=>"110000111",
  10684=>"000011010",
  10685=>"101111011",
  10686=>"111000011",
  10687=>"110001001",
  10688=>"101101111",
  10689=>"110000111",
  10690=>"010100010",
  10691=>"011111010",
  10692=>"000110001",
  10693=>"010101000",
  10694=>"011111110",
  10695=>"100100101",
  10696=>"101011110",
  10697=>"000110111",
  10698=>"001101110",
  10699=>"011010100",
  10700=>"101010111",
  10701=>"101110110",
  10702=>"110111111",
  10703=>"110110111",
  10704=>"110101101",
  10705=>"000010001",
  10706=>"011011010",
  10707=>"000001000",
  10708=>"000101010",
  10709=>"001011010",
  10710=>"001010111",
  10711=>"110110011",
  10712=>"101010101",
  10713=>"000101110",
  10714=>"011111011",
  10715=>"010101100",
  10716=>"101001000",
  10717=>"110001101",
  10718=>"001011101",
  10719=>"110010100",
  10720=>"100100100",
  10721=>"100010111",
  10722=>"110000101",
  10723=>"010001001",
  10724=>"100010011",
  10725=>"111100100",
  10726=>"001111001",
  10727=>"110010111",
  10728=>"101111111",
  10729=>"110010000",
  10730=>"010000111",
  10731=>"111101010",
  10732=>"100001010",
  10733=>"101001110",
  10734=>"010011101",
  10735=>"011011010",
  10736=>"001000001",
  10737=>"010000111",
  10738=>"001001110",
  10739=>"110101011",
  10740=>"110001100",
  10741=>"101000010",
  10742=>"001001101",
  10743=>"110100110",
  10744=>"111011100",
  10745=>"011010001",
  10746=>"101110011",
  10747=>"000100100",
  10748=>"000101110",
  10749=>"011110011",
  10750=>"011000100",
  10751=>"011000111",
  10752=>"011110110",
  10753=>"000011110",
  10754=>"110011010",
  10755=>"100001111",
  10756=>"000110100",
  10757=>"100001001",
  10758=>"011011100",
  10759=>"001110000",
  10760=>"100000001",
  10761=>"011100010",
  10762=>"001011010",
  10763=>"011111010",
  10764=>"100000100",
  10765=>"110000001",
  10766=>"111000111",
  10767=>"101100111",
  10768=>"001011101",
  10769=>"100101001",
  10770=>"111111010",
  10771=>"001101111",
  10772=>"001010000",
  10773=>"011111100",
  10774=>"111111000",
  10775=>"101001010",
  10776=>"001100110",
  10777=>"111100011",
  10778=>"110111111",
  10779=>"000110111",
  10780=>"001000010",
  10781=>"011010011",
  10782=>"111001111",
  10783=>"001100010",
  10784=>"011000000",
  10785=>"111001111",
  10786=>"110111110",
  10787=>"111001101",
  10788=>"001010101",
  10789=>"001110111",
  10790=>"010010010",
  10791=>"111000000",
  10792=>"100100001",
  10793=>"011000001",
  10794=>"101001111",
  10795=>"101000011",
  10796=>"110111011",
  10797=>"000001000",
  10798=>"011010010",
  10799=>"000011001",
  10800=>"011011100",
  10801=>"100110111",
  10802=>"011001011",
  10803=>"001111101",
  10804=>"101111111",
  10805=>"111101011",
  10806=>"000100100",
  10807=>"010101010",
  10808=>"011100101",
  10809=>"000110001",
  10810=>"100111000",
  10811=>"110111010",
  10812=>"100011000",
  10813=>"101100101",
  10814=>"100011010",
  10815=>"010000011",
  10816=>"000010010",
  10817=>"000001000",
  10818=>"101111110",
  10819=>"101000110",
  10820=>"111000110",
  10821=>"010110101",
  10822=>"010101010",
  10823=>"110110000",
  10824=>"111001111",
  10825=>"001110001",
  10826=>"000100111",
  10827=>"101011011",
  10828=>"011110111",
  10829=>"011101011",
  10830=>"000000010",
  10831=>"010111111",
  10832=>"100100100",
  10833=>"000111101",
  10834=>"111110110",
  10835=>"101000010",
  10836=>"100011000",
  10837=>"110111000",
  10838=>"001010000",
  10839=>"111010111",
  10840=>"111010111",
  10841=>"111101111",
  10842=>"101000110",
  10843=>"101110111",
  10844=>"101101110",
  10845=>"011100010",
  10846=>"000011101",
  10847=>"101101111",
  10848=>"001010001",
  10849=>"011111111",
  10850=>"001101001",
  10851=>"011010001",
  10852=>"101101011",
  10853=>"010101000",
  10854=>"011110100",
  10855=>"111001010",
  10856=>"000000100",
  10857=>"100001001",
  10858=>"010011011",
  10859=>"001101010",
  10860=>"010001100",
  10861=>"100110101",
  10862=>"001010100",
  10863=>"100001110",
  10864=>"011000101",
  10865=>"101000000",
  10866=>"001100110",
  10867=>"100010101",
  10868=>"011111000",
  10869=>"001010001",
  10870=>"000000100",
  10871=>"100100111",
  10872=>"001110110",
  10873=>"011100110",
  10874=>"111111101",
  10875=>"111011010",
  10876=>"101101011",
  10877=>"011110001",
  10878=>"111110100",
  10879=>"011110100",
  10880=>"000000101",
  10881=>"101101001",
  10882=>"000110001",
  10883=>"000110001",
  10884=>"010011010",
  10885=>"000100001",
  10886=>"011100000",
  10887=>"001010110",
  10888=>"001101000",
  10889=>"101000010",
  10890=>"100011000",
  10891=>"100100111",
  10892=>"100110001",
  10893=>"010101000",
  10894=>"010011100",
  10895=>"001010001",
  10896=>"101010010",
  10897=>"101000011",
  10898=>"000010001",
  10899=>"000111100",
  10900=>"010100011",
  10901=>"101010110",
  10902=>"100100000",
  10903=>"101000111",
  10904=>"101111000",
  10905=>"111110111",
  10906=>"011000100",
  10907=>"010011110",
  10908=>"010010001",
  10909=>"010011100",
  10910=>"000000010",
  10911=>"011111000",
  10912=>"011100000",
  10913=>"001010101",
  10914=>"000110111",
  10915=>"111110111",
  10916=>"110010010",
  10917=>"010100010",
  10918=>"000000101",
  10919=>"110011001",
  10920=>"101100001",
  10921=>"001010000",
  10922=>"011000011",
  10923=>"001011110",
  10924=>"010001110",
  10925=>"001100001",
  10926=>"010011111",
  10927=>"110110011",
  10928=>"110010001",
  10929=>"001101000",
  10930=>"100011011",
  10931=>"101000011",
  10932=>"111000000",
  10933=>"101001101",
  10934=>"101010100",
  10935=>"011001001",
  10936=>"001100010",
  10937=>"001011001",
  10938=>"101100001",
  10939=>"101110001",
  10940=>"011110000",
  10941=>"100011000",
  10942=>"011010001",
  10943=>"010011100",
  10944=>"001000011",
  10945=>"011001100",
  10946=>"000011010",
  10947=>"011110001",
  10948=>"010110110",
  10949=>"010011000",
  10950=>"001100110",
  10951=>"000101000",
  10952=>"000111011",
  10953=>"111010111",
  10954=>"000011100",
  10955=>"010101111",
  10956=>"111011110",
  10957=>"011010001",
  10958=>"110101000",
  10959=>"111000010",
  10960=>"010111001",
  10961=>"101001110",
  10962=>"110110001",
  10963=>"100010010",
  10964=>"001111101",
  10965=>"111101000",
  10966=>"001000101",
  10967=>"011011111",
  10968=>"000001010",
  10969=>"010101000",
  10970=>"000100011",
  10971=>"010101010",
  10972=>"101011111",
  10973=>"010010101",
  10974=>"110110010",
  10975=>"010111100",
  10976=>"111101100",
  10977=>"000101111",
  10978=>"011110010",
  10979=>"100101111",
  10980=>"110010001",
  10981=>"001101000",
  10982=>"111110010",
  10983=>"110101100",
  10984=>"011110110",
  10985=>"001011111",
  10986=>"111011001",
  10987=>"000111000",
  10988=>"000100100",
  10989=>"000000001",
  10990=>"010011000",
  10991=>"100010111",
  10992=>"100010010",
  10993=>"100100111",
  10994=>"011010000",
  10995=>"110010110",
  10996=>"101011110",
  10997=>"101000110",
  10998=>"000000110",
  10999=>"101100100",
  11000=>"001100010",
  11001=>"101101011",
  11002=>"101101100",
  11003=>"011001010",
  11004=>"111110111",
  11005=>"001010110",
  11006=>"100110110",
  11007=>"000111001",
  11008=>"100100100",
  11009=>"001110011",
  11010=>"111011000",
  11011=>"011111110",
  11012=>"001011011",
  11013=>"000001100",
  11014=>"101100100",
  11015=>"011001101",
  11016=>"101000110",
  11017=>"010001101",
  11018=>"011111001",
  11019=>"010000011",
  11020=>"101110011",
  11021=>"111100110",
  11022=>"101001011",
  11023=>"101101010",
  11024=>"100000010",
  11025=>"001111000",
  11026=>"111110001",
  11027=>"111111001",
  11028=>"001111011",
  11029=>"000101001",
  11030=>"110001101",
  11031=>"101001110",
  11032=>"100110000",
  11033=>"110001010",
  11034=>"010100001",
  11035=>"001110011",
  11036=>"000111000",
  11037=>"000001000",
  11038=>"000010000",
  11039=>"011000011",
  11040=>"100000011",
  11041=>"100000101",
  11042=>"000001001",
  11043=>"011010010",
  11044=>"111010100",
  11045=>"101100111",
  11046=>"010000011",
  11047=>"011111011",
  11048=>"001100110",
  11049=>"101001111",
  11050=>"100100011",
  11051=>"101010001",
  11052=>"000010000",
  11053=>"110100010",
  11054=>"100111100",
  11055=>"001001010",
  11056=>"001000001",
  11057=>"101001101",
  11058=>"011101010",
  11059=>"000111011",
  11060=>"101100101",
  11061=>"011001111",
  11062=>"111011111",
  11063=>"001010110",
  11064=>"000110110",
  11065=>"111101011",
  11066=>"000110010",
  11067=>"100110001",
  11068=>"000111100",
  11069=>"010011100",
  11070=>"001100101",
  11071=>"000110000",
  11072=>"001010100",
  11073=>"101111111",
  11074=>"101001100",
  11075=>"101100010",
  11076=>"100011000",
  11077=>"001111000",
  11078=>"110001100",
  11079=>"011011101",
  11080=>"100100011",
  11081=>"010011110",
  11082=>"011011000",
  11083=>"000111101",
  11084=>"111011110",
  11085=>"111011101",
  11086=>"001101010",
  11087=>"111000110",
  11088=>"000101000",
  11089=>"101111100",
  11090=>"000111001",
  11091=>"100100100",
  11092=>"011101000",
  11093=>"011000001",
  11094=>"110100011",
  11095=>"010000010",
  11096=>"111011101",
  11097=>"110111100",
  11098=>"100111101",
  11099=>"101010110",
  11100=>"101000110",
  11101=>"111111100",
  11102=>"011001111",
  11103=>"010101000",
  11104=>"100101011",
  11105=>"001010011",
  11106=>"110011111",
  11107=>"100110011",
  11108=>"111000011",
  11109=>"011000010",
  11110=>"000010110",
  11111=>"111111011",
  11112=>"010000000",
  11113=>"010010111",
  11114=>"011000111",
  11115=>"101110101",
  11116=>"100011001",
  11117=>"101100011",
  11118=>"011001111",
  11119=>"001000010",
  11120=>"001011111",
  11121=>"011101101",
  11122=>"101001110",
  11123=>"000010110",
  11124=>"111100000",
  11125=>"101111010",
  11126=>"010110100",
  11127=>"001001011",
  11128=>"110111010",
  11129=>"001101101",
  11130=>"000001011",
  11131=>"100110100",
  11132=>"011100010",
  11133=>"111111000",
  11134=>"001011011",
  11135=>"111001000",
  11136=>"010101001",
  11137=>"001011011",
  11138=>"001100100",
  11139=>"100110111",
  11140=>"111001001",
  11141=>"011111110",
  11142=>"101100011",
  11143=>"010100110",
  11144=>"101000100",
  11145=>"110011101",
  11146=>"111100111",
  11147=>"011111010",
  11148=>"111111100",
  11149=>"010111001",
  11150=>"001101011",
  11151=>"110100010",
  11152=>"010010101",
  11153=>"111111110",
  11154=>"011010000",
  11155=>"111110000",
  11156=>"101000100",
  11157=>"011000001",
  11158=>"110001101",
  11159=>"111101110",
  11160=>"110011100",
  11161=>"111101001",
  11162=>"110001010",
  11163=>"000001000",
  11164=>"101101101",
  11165=>"001101011",
  11166=>"000111111",
  11167=>"000100111",
  11168=>"100100101",
  11169=>"010111010",
  11170=>"010011001",
  11171=>"100101100",
  11172=>"100101100",
  11173=>"000011011",
  11174=>"111000000",
  11175=>"111111000",
  11176=>"000111010",
  11177=>"101001010",
  11178=>"010110010",
  11179=>"010010110",
  11180=>"001100110",
  11181=>"000011001",
  11182=>"110111001",
  11183=>"100100111",
  11184=>"111011010",
  11185=>"010100101",
  11186=>"110011011",
  11187=>"001100101",
  11188=>"011110111",
  11189=>"110101011",
  11190=>"100101001",
  11191=>"110001001",
  11192=>"110110101",
  11193=>"101011001",
  11194=>"110110101",
  11195=>"000011100",
  11196=>"101011101",
  11197=>"010011111",
  11198=>"101110010",
  11199=>"001111001",
  11200=>"010001011",
  11201=>"001010001",
  11202=>"110101001",
  11203=>"011111000",
  11204=>"110001001",
  11205=>"000010100",
  11206=>"100001101",
  11207=>"101101011",
  11208=>"001000111",
  11209=>"110010111",
  11210=>"010011111",
  11211=>"101011010",
  11212=>"011010010",
  11213=>"100000001",
  11214=>"000100000",
  11215=>"010011000",
  11216=>"110000011",
  11217=>"000011101",
  11218=>"010001001",
  11219=>"010011010",
  11220=>"110101110",
  11221=>"111111001",
  11222=>"100100111",
  11223=>"110100010",
  11224=>"110101001",
  11225=>"100111110",
  11226=>"100111111",
  11227=>"011110111",
  11228=>"111111001",
  11229=>"100100110",
  11230=>"011011100",
  11231=>"100010011",
  11232=>"010100011",
  11233=>"000111101",
  11234=>"010000100",
  11235=>"001101101",
  11236=>"001010001",
  11237=>"011001010",
  11238=>"010111010",
  11239=>"000000010",
  11240=>"100110111",
  11241=>"010001100",
  11242=>"110110101",
  11243=>"001010011",
  11244=>"100000011",
  11245=>"011110101",
  11246=>"000001111",
  11247=>"100010001",
  11248=>"110001011",
  11249=>"110011010",
  11250=>"101001111",
  11251=>"010101011",
  11252=>"011011101",
  11253=>"000000100",
  11254=>"000001001",
  11255=>"111011110",
  11256=>"111011111",
  11257=>"110001100",
  11258=>"110100001",
  11259=>"101010101",
  11260=>"001000010",
  11261=>"011000011",
  11262=>"011011001",
  11263=>"111100110",
  11264=>"100101001",
  11265=>"110100111",
  11266=>"001011000",
  11267=>"011101101",
  11268=>"100001111",
  11269=>"101011010",
  11270=>"011001110",
  11271=>"111101111",
  11272=>"001011100",
  11273=>"001001011",
  11274=>"011010001",
  11275=>"011001111",
  11276=>"110111000",
  11277=>"000101010",
  11278=>"100100000",
  11279=>"000011011",
  11280=>"101001000",
  11281=>"011100000",
  11282=>"011010110",
  11283=>"000000101",
  11284=>"000110101",
  11285=>"101010100",
  11286=>"010000100",
  11287=>"011000100",
  11288=>"000011101",
  11289=>"001100101",
  11290=>"001111010",
  11291=>"011001001",
  11292=>"101111100",
  11293=>"101111100",
  11294=>"000100110",
  11295=>"010010001",
  11296=>"010010101",
  11297=>"100000011",
  11298=>"110101111",
  11299=>"010011101",
  11300=>"111101001",
  11301=>"011100000",
  11302=>"001100110",
  11303=>"100010011",
  11304=>"111001101",
  11305=>"100000100",
  11306=>"001101111",
  11307=>"111010011",
  11308=>"001101000",
  11309=>"100010100",
  11310=>"100101010",
  11311=>"011000101",
  11312=>"100101000",
  11313=>"101101110",
  11314=>"111101101",
  11315=>"001111011",
  11316=>"100101011",
  11317=>"010000010",
  11318=>"111101111",
  11319=>"110101101",
  11320=>"001010000",
  11321=>"101011111",
  11322=>"011011100",
  11323=>"010001101",
  11324=>"101000100",
  11325=>"110010010",
  11326=>"110111001",
  11327=>"101010011",
  11328=>"011001000",
  11329=>"100101101",
  11330=>"100100110",
  11331=>"000110001",
  11332=>"011100000",
  11333=>"010011001",
  11334=>"010110100",
  11335=>"010101100",
  11336=>"100010111",
  11337=>"000111010",
  11338=>"111111000",
  11339=>"000011100",
  11340=>"010000000",
  11341=>"111011001",
  11342=>"110010000",
  11343=>"000000100",
  11344=>"011110011",
  11345=>"111110000",
  11346=>"000111000",
  11347=>"110000110",
  11348=>"000110010",
  11349=>"010000101",
  11350=>"110100000",
  11351=>"100100110",
  11352=>"101111101",
  11353=>"001011111",
  11354=>"111101110",
  11355=>"010000100",
  11356=>"111011001",
  11357=>"111001001",
  11358=>"001000001",
  11359=>"100111010",
  11360=>"101110111",
  11361=>"111101000",
  11362=>"011100001",
  11363=>"101001100",
  11364=>"010110010",
  11365=>"001000000",
  11366=>"011101011",
  11367=>"010110000",
  11368=>"011111100",
  11369=>"101110011",
  11370=>"001100000",
  11371=>"000110011",
  11372=>"000101011",
  11373=>"000000101",
  11374=>"010001110",
  11375=>"001110110",
  11376=>"100000011",
  11377=>"101110110",
  11378=>"100111011",
  11379=>"111101000",
  11380=>"010111110",
  11381=>"101100011",
  11382=>"101111010",
  11383=>"101001000",
  11384=>"101101000",
  11385=>"000001110",
  11386=>"110110111",
  11387=>"011000001",
  11388=>"011001010",
  11389=>"011111101",
  11390=>"010000011",
  11391=>"010000000",
  11392=>"101001111",
  11393=>"110101000",
  11394=>"101011101",
  11395=>"100000001",
  11396=>"101000010",
  11397=>"011010000",
  11398=>"100011101",
  11399=>"000110100",
  11400=>"010100111",
  11401=>"111100001",
  11402=>"110000101",
  11403=>"111011111",
  11404=>"100011111",
  11405=>"000000010",
  11406=>"100011001",
  11407=>"000100110",
  11408=>"000111100",
  11409=>"101001011",
  11410=>"011010011",
  11411=>"100110001",
  11412=>"000000111",
  11413=>"110000100",
  11414=>"011100011",
  11415=>"010010011",
  11416=>"100001000",
  11417=>"100001101",
  11418=>"100101111",
  11419=>"000000010",
  11420=>"000000001",
  11421=>"001101100",
  11422=>"100010110",
  11423=>"100111011",
  11424=>"100001010",
  11425=>"110011011",
  11426=>"111001100",
  11427=>"010100011",
  11428=>"011010111",
  11429=>"001000101",
  11430=>"010111110",
  11431=>"000101111",
  11432=>"001001101",
  11433=>"000011111",
  11434=>"001101101",
  11435=>"111110000",
  11436=>"111100001",
  11437=>"110110010",
  11438=>"100100111",
  11439=>"111011010",
  11440=>"010110100",
  11441=>"001001111",
  11442=>"100110001",
  11443=>"000000101",
  11444=>"100100000",
  11445=>"100011001",
  11446=>"111001000",
  11447=>"101100011",
  11448=>"001101011",
  11449=>"000001011",
  11450=>"000001001",
  11451=>"111110111",
  11452=>"110111110",
  11453=>"010011101",
  11454=>"010001000",
  11455=>"010010111",
  11456=>"000000000",
  11457=>"100111011",
  11458=>"110001110",
  11459=>"100100101",
  11460=>"010110111",
  11461=>"100110011",
  11462=>"000100001",
  11463=>"111000111",
  11464=>"011101011",
  11465=>"100100101",
  11466=>"001110001",
  11467=>"000100000",
  11468=>"000100011",
  11469=>"111010010",
  11470=>"111111011",
  11471=>"111110111",
  11472=>"110100111",
  11473=>"110010001",
  11474=>"011110111",
  11475=>"000101010",
  11476=>"001001100",
  11477=>"111111011",
  11478=>"100001001",
  11479=>"011100001",
  11480=>"011011001",
  11481=>"010001100",
  11482=>"010001111",
  11483=>"000101111",
  11484=>"000001010",
  11485=>"001010011",
  11486=>"001101001",
  11487=>"110000101",
  11488=>"000101010",
  11489=>"010101000",
  11490=>"100000010",
  11491=>"100011100",
  11492=>"111111011",
  11493=>"111001110",
  11494=>"111110011",
  11495=>"100110010",
  11496=>"011111110",
  11497=>"111101110",
  11498=>"101110001",
  11499=>"000100100",
  11500=>"010110011",
  11501=>"101001110",
  11502=>"001001100",
  11503=>"010100110",
  11504=>"011010100",
  11505=>"110000101",
  11506=>"110101011",
  11507=>"000010010",
  11508=>"010100010",
  11509=>"101101101",
  11510=>"000011000",
  11511=>"110000110",
  11512=>"001110000",
  11513=>"111000100",
  11514=>"011010101",
  11515=>"010001100",
  11516=>"011111100",
  11517=>"110010110",
  11518=>"000100100",
  11519=>"011101101",
  11520=>"011000001",
  11521=>"000001100",
  11522=>"100010110",
  11523=>"100011000",
  11524=>"001111000",
  11525=>"010010010",
  11526=>"111111000",
  11527=>"001001000",
  11528=>"010000110",
  11529=>"011101000",
  11530=>"111011100",
  11531=>"111010100",
  11532=>"110101110",
  11533=>"011110001",
  11534=>"110011110",
  11535=>"001100101",
  11536=>"111000100",
  11537=>"000000000",
  11538=>"101010100",
  11539=>"000010111",
  11540=>"011011110",
  11541=>"010001000",
  11542=>"011111110",
  11543=>"000101011",
  11544=>"010001001",
  11545=>"000011100",
  11546=>"100101111",
  11547=>"101000110",
  11548=>"011000111",
  11549=>"100000010",
  11550=>"110111011",
  11551=>"000110110",
  11552=>"010001001",
  11553=>"001000111",
  11554=>"010001001",
  11555=>"100001000",
  11556=>"000111110",
  11557=>"111101000",
  11558=>"110000100",
  11559=>"111110011",
  11560=>"001001011",
  11561=>"011010101",
  11562=>"000111111",
  11563=>"100100010",
  11564=>"100001001",
  11565=>"111011001",
  11566=>"001101110",
  11567=>"001011101",
  11568=>"000111000",
  11569=>"000000110",
  11570=>"010010000",
  11571=>"110101111",
  11572=>"001110010",
  11573=>"000011000",
  11574=>"000001111",
  11575=>"101000001",
  11576=>"000001111",
  11577=>"100110111",
  11578=>"001000110",
  11579=>"001101000",
  11580=>"011000000",
  11581=>"111010011",
  11582=>"011001110",
  11583=>"100100101",
  11584=>"101010100",
  11585=>"011111011",
  11586=>"011001010",
  11587=>"111011011",
  11588=>"010011010",
  11589=>"010000100",
  11590=>"110101010",
  11591=>"010011000",
  11592=>"001101011",
  11593=>"110101100",
  11594=>"101010010",
  11595=>"110100111",
  11596=>"110100011",
  11597=>"001010001",
  11598=>"100010111",
  11599=>"100101001",
  11600=>"001101101",
  11601=>"011001111",
  11602=>"100001011",
  11603=>"011000000",
  11604=>"100110110",
  11605=>"101010000",
  11606=>"110100111",
  11607=>"111010101",
  11608=>"001010010",
  11609=>"100000001",
  11610=>"110010001",
  11611=>"010010001",
  11612=>"011010110",
  11613=>"001100010",
  11614=>"010010000",
  11615=>"000000010",
  11616=>"010100010",
  11617=>"100011111",
  11618=>"111001000",
  11619=>"011000001",
  11620=>"111001010",
  11621=>"001110011",
  11622=>"001000111",
  11623=>"101011101",
  11624=>"000100100",
  11625=>"010111010",
  11626=>"100111101",
  11627=>"101111111",
  11628=>"000001110",
  11629=>"001100010",
  11630=>"000100000",
  11631=>"101100111",
  11632=>"011001111",
  11633=>"011010011",
  11634=>"101100010",
  11635=>"110011101",
  11636=>"101000001",
  11637=>"110001001",
  11638=>"010101101",
  11639=>"101010111",
  11640=>"100110011",
  11641=>"011100011",
  11642=>"011111110",
  11643=>"110010100",
  11644=>"001011010",
  11645=>"101000111",
  11646=>"111001000",
  11647=>"101100111",
  11648=>"101111010",
  11649=>"011010011",
  11650=>"100111001",
  11651=>"001011000",
  11652=>"010000110",
  11653=>"010001011",
  11654=>"110010100",
  11655=>"000000100",
  11656=>"100100000",
  11657=>"111001001",
  11658=>"100110001",
  11659=>"111011010",
  11660=>"111001101",
  11661=>"010011111",
  11662=>"111001010",
  11663=>"000100000",
  11664=>"101101010",
  11665=>"000000011",
  11666=>"000101011",
  11667=>"100101001",
  11668=>"110111010",
  11669=>"111111100",
  11670=>"010100011",
  11671=>"101011110",
  11672=>"001011110",
  11673=>"111000010",
  11674=>"111101111",
  11675=>"110000000",
  11676=>"101011101",
  11677=>"010010000",
  11678=>"111001101",
  11679=>"011010000",
  11680=>"000101000",
  11681=>"001100111",
  11682=>"010010001",
  11683=>"011001001",
  11684=>"110111011",
  11685=>"000010001",
  11686=>"100011000",
  11687=>"010001011",
  11688=>"001101111",
  11689=>"100111101",
  11690=>"100010000",
  11691=>"011010110",
  11692=>"000010011",
  11693=>"110011111",
  11694=>"011011010",
  11695=>"001100101",
  11696=>"001000011",
  11697=>"011110111",
  11698=>"101001000",
  11699=>"001001101",
  11700=>"000111101",
  11701=>"111111110",
  11702=>"011111111",
  11703=>"110011110",
  11704=>"110010101",
  11705=>"010100010",
  11706=>"110100111",
  11707=>"001010010",
  11708=>"011111000",
  11709=>"110000101",
  11710=>"110011101",
  11711=>"000001001",
  11712=>"010000101",
  11713=>"111001110",
  11714=>"011111010",
  11715=>"110111100",
  11716=>"011110101",
  11717=>"111001011",
  11718=>"101011000",
  11719=>"010011111",
  11720=>"011110101",
  11721=>"000001000",
  11722=>"011001111",
  11723=>"001111100",
  11724=>"101001010",
  11725=>"101001010",
  11726=>"101110011",
  11727=>"100000110",
  11728=>"110011110",
  11729=>"111011010",
  11730=>"010110101",
  11731=>"100000101",
  11732=>"000010010",
  11733=>"011101111",
  11734=>"011111000",
  11735=>"010101010",
  11736=>"010111011",
  11737=>"011110100",
  11738=>"110111010",
  11739=>"111011001",
  11740=>"110111010",
  11741=>"111101010",
  11742=>"010000011",
  11743=>"011111110",
  11744=>"100101101",
  11745=>"000000011",
  11746=>"110000010",
  11747=>"111000100",
  11748=>"000110000",
  11749=>"001011001",
  11750=>"100100000",
  11751=>"110110011",
  11752=>"111101111",
  11753=>"001010110",
  11754=>"101100001",
  11755=>"111100001",
  11756=>"000111111",
  11757=>"110000101",
  11758=>"000101010",
  11759=>"100100000",
  11760=>"010010001",
  11761=>"100101101",
  11762=>"111111101",
  11763=>"111001011",
  11764=>"101101111",
  11765=>"101000110",
  11766=>"001001011",
  11767=>"100100000",
  11768=>"010011011",
  11769=>"111100000",
  11770=>"101000001",
  11771=>"111001010",
  11772=>"110011010",
  11773=>"000111100",
  11774=>"111100100",
  11775=>"001111101",
  11776=>"110100010",
  11777=>"000001011",
  11778=>"010110100",
  11779=>"010100000",
  11780=>"101100011",
  11781=>"001000000",
  11782=>"011101110",
  11783=>"000010010",
  11784=>"100000011",
  11785=>"011101111",
  11786=>"011011100",
  11787=>"010000000",
  11788=>"000110111",
  11789=>"111010100",
  11790=>"111111010",
  11791=>"011110110",
  11792=>"111010100",
  11793=>"000010111",
  11794=>"110110011",
  11795=>"111100110",
  11796=>"011101000",
  11797=>"000010010",
  11798=>"100110000",
  11799=>"111100010",
  11800=>"011101001",
  11801=>"011001110",
  11802=>"111000101",
  11803=>"010011011",
  11804=>"001000110",
  11805=>"110110001",
  11806=>"010100101",
  11807=>"110111011",
  11808=>"110100111",
  11809=>"111001101",
  11810=>"100101001",
  11811=>"111110000",
  11812=>"000000011",
  11813=>"110100100",
  11814=>"000000110",
  11815=>"010101000",
  11816=>"101000111",
  11817=>"101101010",
  11818=>"101110010",
  11819=>"011010000",
  11820=>"011100100",
  11821=>"010100000",
  11822=>"110011111",
  11823=>"101000000",
  11824=>"011000011",
  11825=>"011100110",
  11826=>"100100000",
  11827=>"000110110",
  11828=>"110000101",
  11829=>"100001001",
  11830=>"010111000",
  11831=>"010111101",
  11832=>"111010110",
  11833=>"111100110",
  11834=>"011000010",
  11835=>"010100111",
  11836=>"100100011",
  11837=>"100110011",
  11838=>"100111110",
  11839=>"101011011",
  11840=>"000111000",
  11841=>"010001000",
  11842=>"011010000",
  11843=>"101111010",
  11844=>"000011110",
  11845=>"000100110",
  11846=>"010011111",
  11847=>"010010000",
  11848=>"010100101",
  11849=>"001000000",
  11850=>"011100001",
  11851=>"111110101",
  11852=>"110100000",
  11853=>"000100001",
  11854=>"100010000",
  11855=>"111111110",
  11856=>"111001110",
  11857=>"000110101",
  11858=>"100011101",
  11859=>"000111100",
  11860=>"110110010",
  11861=>"101011011",
  11862=>"010100000",
  11863=>"000010001",
  11864=>"111001101",
  11865=>"111010110",
  11866=>"000001000",
  11867=>"010001010",
  11868=>"000100000",
  11869=>"001101000",
  11870=>"001011010",
  11871=>"001010101",
  11872=>"100111110",
  11873=>"100001110",
  11874=>"000000011",
  11875=>"110110100",
  11876=>"000000101",
  11877=>"000100111",
  11878=>"001000001",
  11879=>"100101100",
  11880=>"000100101",
  11881=>"001110011",
  11882=>"111011101",
  11883=>"100100001",
  11884=>"100001001",
  11885=>"111000000",
  11886=>"101100111",
  11887=>"000010101",
  11888=>"001001101",
  11889=>"011101001",
  11890=>"111101001",
  11891=>"111000000",
  11892=>"011000011",
  11893=>"001001110",
  11894=>"100000110",
  11895=>"000000110",
  11896=>"000001001",
  11897=>"110111010",
  11898=>"111011101",
  11899=>"011001100",
  11900=>"100000101",
  11901=>"111100010",
  11902=>"010010100",
  11903=>"111100010",
  11904=>"001000101",
  11905=>"010011000",
  11906=>"010010001",
  11907=>"000101001",
  11908=>"100101101",
  11909=>"111110000",
  11910=>"111011111",
  11911=>"011011000",
  11912=>"111100100",
  11913=>"000111101",
  11914=>"010010101",
  11915=>"100000111",
  11916=>"111100001",
  11917=>"010101000",
  11918=>"001001001",
  11919=>"011110100",
  11920=>"110110111",
  11921=>"001110010",
  11922=>"010011110",
  11923=>"111000100",
  11924=>"000110001",
  11925=>"011110111",
  11926=>"011101010",
  11927=>"000111100",
  11928=>"101010000",
  11929=>"011000011",
  11930=>"100111000",
  11931=>"110111101",
  11932=>"011011010",
  11933=>"110100010",
  11934=>"111000000",
  11935=>"100001000",
  11936=>"001111111",
  11937=>"011111010",
  11938=>"101100000",
  11939=>"101010001",
  11940=>"101110100",
  11941=>"001110000",
  11942=>"111011110",
  11943=>"000010111",
  11944=>"100110110",
  11945=>"001010001",
  11946=>"101001001",
  11947=>"100111111",
  11948=>"000010100",
  11949=>"010000101",
  11950=>"010011100",
  11951=>"011000100",
  11952=>"101000011",
  11953=>"100010101",
  11954=>"010000000",
  11955=>"100111000",
  11956=>"111010100",
  11957=>"000101010",
  11958=>"011011111",
  11959=>"011010001",
  11960=>"110110110",
  11961=>"110101000",
  11962=>"011111110",
  11963=>"010100100",
  11964=>"100011010",
  11965=>"000101011",
  11966=>"100101000",
  11967=>"010000010",
  11968=>"011010000",
  11969=>"000100000",
  11970=>"101000001",
  11971=>"111111110",
  11972=>"101000000",
  11973=>"100000000",
  11974=>"011000101",
  11975=>"010111011",
  11976=>"100110000",
  11977=>"001110110",
  11978=>"011011110",
  11979=>"101110100",
  11980=>"000010010",
  11981=>"011110110",
  11982=>"010000011",
  11983=>"000001101",
  11984=>"001000010",
  11985=>"010100100",
  11986=>"010001111",
  11987=>"000000011",
  11988=>"111011111",
  11989=>"110011101",
  11990=>"011101011",
  11991=>"010001001",
  11992=>"100000101",
  11993=>"010001111",
  11994=>"111100100",
  11995=>"111000100",
  11996=>"111101111",
  11997=>"011000110",
  11998=>"110001011",
  11999=>"100010011",
  12000=>"101100011",
  12001=>"110100101",
  12002=>"100010000",
  12003=>"110010101",
  12004=>"111000110",
  12005=>"011101111",
  12006=>"000111101",
  12007=>"011111101",
  12008=>"101000000",
  12009=>"011100001",
  12010=>"110110110",
  12011=>"000110001",
  12012=>"001101110",
  12013=>"100111111",
  12014=>"000000000",
  12015=>"100110110",
  12016=>"010010010",
  12017=>"001111110",
  12018=>"000001011",
  12019=>"001010100",
  12020=>"111010111",
  12021=>"110011011",
  12022=>"000101111",
  12023=>"110011111",
  12024=>"111000101",
  12025=>"011111010",
  12026=>"100101100",
  12027=>"100110001",
  12028=>"100010000",
  12029=>"100000011",
  12030=>"010110000",
  12031=>"011001010",
  12032=>"111111110",
  12033=>"001001010",
  12034=>"010100000",
  12035=>"101111111",
  12036=>"110110010",
  12037=>"010001101",
  12038=>"111010010",
  12039=>"101010011",
  12040=>"101000011",
  12041=>"111111111",
  12042=>"110100110",
  12043=>"101111110",
  12044=>"010111110",
  12045=>"000101100",
  12046=>"011011010",
  12047=>"000100100",
  12048=>"101100100",
  12049=>"010100010",
  12050=>"001000110",
  12051=>"011001010",
  12052=>"011111001",
  12053=>"000001011",
  12054=>"011110100",
  12055=>"100100000",
  12056=>"101110010",
  12057=>"100100001",
  12058=>"101000011",
  12059=>"101000111",
  12060=>"101011110",
  12061=>"101111101",
  12062=>"110100000",
  12063=>"110000110",
  12064=>"010100000",
  12065=>"100001101",
  12066=>"101001110",
  12067=>"000001000",
  12068=>"100101110",
  12069=>"101101010",
  12070=>"101101010",
  12071=>"100111111",
  12072=>"010100001",
  12073=>"010001101",
  12074=>"100111011",
  12075=>"100011011",
  12076=>"110111100",
  12077=>"100001101",
  12078=>"110001001",
  12079=>"101110000",
  12080=>"000011100",
  12081=>"111010110",
  12082=>"011110111",
  12083=>"110010100",
  12084=>"000110101",
  12085=>"000110001",
  12086=>"101010100",
  12087=>"010101100",
  12088=>"001111001",
  12089=>"010010100",
  12090=>"010010101",
  12091=>"011111111",
  12092=>"110011001",
  12093=>"010111001",
  12094=>"001101001",
  12095=>"000110110",
  12096=>"010000010",
  12097=>"001001010",
  12098=>"001011010",
  12099=>"100001010",
  12100=>"101011100",
  12101=>"110011110",
  12102=>"111101100",
  12103=>"011000010",
  12104=>"100100101",
  12105=>"010111101",
  12106=>"001011000",
  12107=>"111100000",
  12108=>"010000010",
  12109=>"011111111",
  12110=>"011111100",
  12111=>"110000100",
  12112=>"110011101",
  12113=>"000000001",
  12114=>"010001111",
  12115=>"010111110",
  12116=>"111101010",
  12117=>"000000001",
  12118=>"001010001",
  12119=>"110000010",
  12120=>"000100011",
  12121=>"110011110",
  12122=>"010111010",
  12123=>"100010010",
  12124=>"001110110",
  12125=>"110111111",
  12126=>"100110010",
  12127=>"001100101",
  12128=>"001010111",
  12129=>"000110111",
  12130=>"011100011",
  12131=>"001001101",
  12132=>"011110011",
  12133=>"001011101",
  12134=>"100111001",
  12135=>"000010101",
  12136=>"111111111",
  12137=>"111010100",
  12138=>"010011110",
  12139=>"111110010",
  12140=>"100011000",
  12141=>"001100010",
  12142=>"001101111",
  12143=>"010011001",
  12144=>"000110111",
  12145=>"000001000",
  12146=>"101101010",
  12147=>"100001010",
  12148=>"000010110",
  12149=>"010010001",
  12150=>"111111011",
  12151=>"000001111",
  12152=>"000010000",
  12153=>"010101000",
  12154=>"100101111",
  12155=>"110111010",
  12156=>"101101001",
  12157=>"011110101",
  12158=>"001000011",
  12159=>"110000111",
  12160=>"101100110",
  12161=>"101011011",
  12162=>"010110011",
  12163=>"010101010",
  12164=>"001100101",
  12165=>"010110001",
  12166=>"101010101",
  12167=>"001010000",
  12168=>"000101001",
  12169=>"110001111",
  12170=>"101010010",
  12171=>"010000111",
  12172=>"101001001",
  12173=>"100000011",
  12174=>"010110110",
  12175=>"011101001",
  12176=>"000100001",
  12177=>"001011001",
  12178=>"101000110",
  12179=>"000000000",
  12180=>"111100000",
  12181=>"011111000",
  12182=>"000001001",
  12183=>"011111111",
  12184=>"100100101",
  12185=>"111111111",
  12186=>"010001101",
  12187=>"001010011",
  12188=>"100011101",
  12189=>"000101111",
  12190=>"000011000",
  12191=>"100011100",
  12192=>"000001010",
  12193=>"111010101",
  12194=>"100100010",
  12195=>"000101111",
  12196=>"011000010",
  12197=>"011000100",
  12198=>"101011000",
  12199=>"010011100",
  12200=>"001111011",
  12201=>"011111000",
  12202=>"011101101",
  12203=>"100010000",
  12204=>"110101010",
  12205=>"000100101",
  12206=>"100000000",
  12207=>"111000010",
  12208=>"100010101",
  12209=>"000010011",
  12210=>"100101000",
  12211=>"001000001",
  12212=>"100110111",
  12213=>"000011001",
  12214=>"010011010",
  12215=>"001110101",
  12216=>"001111000",
  12217=>"001001010",
  12218=>"110010111",
  12219=>"111110001",
  12220=>"011110101",
  12221=>"000100101",
  12222=>"101100111",
  12223=>"000000001",
  12224=>"000010101",
  12225=>"100100000",
  12226=>"100001111",
  12227=>"111101100",
  12228=>"001010010",
  12229=>"010100000",
  12230=>"011110011",
  12231=>"010100000",
  12232=>"111100011",
  12233=>"001101111",
  12234=>"100101110",
  12235=>"000011111",
  12236=>"011000110",
  12237=>"101001101",
  12238=>"000001111",
  12239=>"111111111",
  12240=>"111000111",
  12241=>"010101000",
  12242=>"011000110",
  12243=>"110001010",
  12244=>"111000101",
  12245=>"100110101",
  12246=>"100010000",
  12247=>"000100101",
  12248=>"101000010",
  12249=>"100000100",
  12250=>"110011011",
  12251=>"000000101",
  12252=>"000001100",
  12253=>"001000001",
  12254=>"001100001",
  12255=>"001010010",
  12256=>"010101101",
  12257=>"010111111",
  12258=>"111010111",
  12259=>"100110010",
  12260=>"001100110",
  12261=>"110010111",
  12262=>"000100011",
  12263=>"110011110",
  12264=>"010111001",
  12265=>"010010000",
  12266=>"001011101",
  12267=>"111100100",
  12268=>"010000100",
  12269=>"101011000",
  12270=>"001111010",
  12271=>"100100100",
  12272=>"100110110",
  12273=>"101101111",
  12274=>"000010111",
  12275=>"000100101",
  12276=>"011000100",
  12277=>"111010010",
  12278=>"101011001",
  12279=>"100000010",
  12280=>"111001000",
  12281=>"010001001",
  12282=>"100110101",
  12283=>"100011001",
  12284=>"110000110",
  12285=>"111111001",
  12286=>"100001000",
  12287=>"001100000",
  12288=>"000100001",
  12289=>"000011011",
  12290=>"101000100",
  12291=>"001111010",
  12292=>"010000100",
  12293=>"001101101",
  12294=>"110000110",
  12295=>"111101010",
  12296=>"110111011",
  12297=>"001001001",
  12298=>"001101101",
  12299=>"111100010",
  12300=>"111100001",
  12301=>"101111111",
  12302=>"000001111",
  12303=>"001011101",
  12304=>"001101110",
  12305=>"101010010",
  12306=>"010000110",
  12307=>"010111101",
  12308=>"011100110",
  12309=>"100111110",
  12310=>"000011010",
  12311=>"001111110",
  12312=>"110000011",
  12313=>"110011000",
  12314=>"000111111",
  12315=>"000111100",
  12316=>"010111111",
  12317=>"111010001",
  12318=>"001101011",
  12319=>"110011100",
  12320=>"000011110",
  12321=>"100100010",
  12322=>"001110001",
  12323=>"110010010",
  12324=>"000100101",
  12325=>"111011111",
  12326=>"011001011",
  12327=>"111010001",
  12328=>"101011100",
  12329=>"001011001",
  12330=>"100000000",
  12331=>"000001101",
  12332=>"001110100",
  12333=>"000011100",
  12334=>"100111111",
  12335=>"010101110",
  12336=>"111011001",
  12337=>"011010111",
  12338=>"000101001",
  12339=>"111110110",
  12340=>"101001111",
  12341=>"100101100",
  12342=>"100110000",
  12343=>"001110011",
  12344=>"000100001",
  12345=>"101101101",
  12346=>"100010100",
  12347=>"011111110",
  12348=>"001100010",
  12349=>"001011011",
  12350=>"110100111",
  12351=>"010100111",
  12352=>"110110010",
  12353=>"000100000",
  12354=>"000010100",
  12355=>"000010110",
  12356=>"000101000",
  12357=>"111011100",
  12358=>"001000011",
  12359=>"001011100",
  12360=>"010101011",
  12361=>"000101000",
  12362=>"101000010",
  12363=>"001011110",
  12364=>"010100010",
  12365=>"001001010",
  12366=>"111000101",
  12367=>"110100010",
  12368=>"000100110",
  12369=>"001001001",
  12370=>"000010010",
  12371=>"011100001",
  12372=>"001110000",
  12373=>"011010010",
  12374=>"001011010",
  12375=>"100000000",
  12376=>"011111111",
  12377=>"110101110",
  12378=>"000000111",
  12379=>"011000110",
  12380=>"001001100",
  12381=>"000100110",
  12382=>"001111101",
  12383=>"011100001",
  12384=>"001000001",
  12385=>"111010011",
  12386=>"001011001",
  12387=>"000011100",
  12388=>"010111101",
  12389=>"100101110",
  12390=>"011010110",
  12391=>"000010000",
  12392=>"011111001",
  12393=>"110010101",
  12394=>"010011101",
  12395=>"000001101",
  12396=>"011000010",
  12397=>"110101101",
  12398=>"111100101",
  12399=>"000001110",
  12400=>"000001100",
  12401=>"000010000",
  12402=>"001011000",
  12403=>"110001110",
  12404=>"011011000",
  12405=>"111100111",
  12406=>"011111111",
  12407=>"100001111",
  12408=>"111011001",
  12409=>"000000100",
  12410=>"000100100",
  12411=>"101011001",
  12412=>"000000011",
  12413=>"110100001",
  12414=>"001110111",
  12415=>"001000001",
  12416=>"111100100",
  12417=>"001011101",
  12418=>"100100110",
  12419=>"001011000",
  12420=>"100000101",
  12421=>"010110111",
  12422=>"001110110",
  12423=>"011000100",
  12424=>"010000010",
  12425=>"110111100",
  12426=>"110100101",
  12427=>"101111001",
  12428=>"101000000",
  12429=>"111001101",
  12430=>"011101101",
  12431=>"001000100",
  12432=>"011010101",
  12433=>"011110100",
  12434=>"110000101",
  12435=>"000101101",
  12436=>"101100001",
  12437=>"110101010",
  12438=>"001111110",
  12439=>"100000101",
  12440=>"001100111",
  12441=>"101110000",
  12442=>"001010101",
  12443=>"001000000",
  12444=>"110110011",
  12445=>"000000000",
  12446=>"100010110",
  12447=>"110010000",
  12448=>"111011100",
  12449=>"011001111",
  12450=>"100000110",
  12451=>"101110100",
  12452=>"111101101",
  12453=>"110011110",
  12454=>"001001001",
  12455=>"111111111",
  12456=>"000010011",
  12457=>"000111101",
  12458=>"100010011",
  12459=>"100011110",
  12460=>"100111001",
  12461=>"101111001",
  12462=>"000101011",
  12463=>"111001101",
  12464=>"000001101",
  12465=>"000001010",
  12466=>"111010111",
  12467=>"101011110",
  12468=>"010000010",
  12469=>"010010101",
  12470=>"011100011",
  12471=>"001000000",
  12472=>"010110100",
  12473=>"101000110",
  12474=>"101001000",
  12475=>"011100010",
  12476=>"011111011",
  12477=>"011101011",
  12478=>"010001011",
  12479=>"101111001",
  12480=>"100110111",
  12481=>"010000010",
  12482=>"011000101",
  12483=>"100100111",
  12484=>"010110010",
  12485=>"000011011",
  12486=>"111000101",
  12487=>"110100001",
  12488=>"001100111",
  12489=>"001011010",
  12490=>"000000100",
  12491=>"001001100",
  12492=>"110100000",
  12493=>"010101001",
  12494=>"100100111",
  12495=>"001000010",
  12496=>"100100111",
  12497=>"111001000",
  12498=>"111110110",
  12499=>"010011110",
  12500=>"010000011",
  12501=>"101010110",
  12502=>"101001011",
  12503=>"010001001",
  12504=>"101001101",
  12505=>"000000010",
  12506=>"001101111",
  12507=>"001001100",
  12508=>"000101010",
  12509=>"001001100",
  12510=>"011001110",
  12511=>"110111001",
  12512=>"101000110",
  12513=>"011101001",
  12514=>"111011000",
  12515=>"111100111",
  12516=>"110001011",
  12517=>"001011011",
  12518=>"001001110",
  12519=>"101011010",
  12520=>"001111110",
  12521=>"110011001",
  12522=>"110011010",
  12523=>"101100100",
  12524=>"011111001",
  12525=>"011000110",
  12526=>"001110110",
  12527=>"000000000",
  12528=>"111111010",
  12529=>"111110111",
  12530=>"000111101",
  12531=>"011000100",
  12532=>"101100000",
  12533=>"101001001",
  12534=>"000101000",
  12535=>"100000100",
  12536=>"001101110",
  12537=>"101001001",
  12538=>"110010010",
  12539=>"000111000",
  12540=>"011001001",
  12541=>"011011100",
  12542=>"001010001",
  12543=>"000000110",
  12544=>"010111110",
  12545=>"001111011",
  12546=>"101000101",
  12547=>"011100011",
  12548=>"110000111",
  12549=>"101011001",
  12550=>"010001111",
  12551=>"101001001",
  12552=>"001100000",
  12553=>"010000001",
  12554=>"000101111",
  12555=>"110111011",
  12556=>"001110001",
  12557=>"101000100",
  12558=>"001011111",
  12559=>"000111101",
  12560=>"101111100",
  12561=>"001111010",
  12562=>"100110011",
  12563=>"111010001",
  12564=>"000110001",
  12565=>"100011110",
  12566=>"110011001",
  12567=>"101001111",
  12568=>"111110101",
  12569=>"000100010",
  12570=>"000111011",
  12571=>"001110000",
  12572=>"110001100",
  12573=>"011110100",
  12574=>"110010010",
  12575=>"000100111",
  12576=>"100111101",
  12577=>"111111111",
  12578=>"110000100",
  12579=>"101110110",
  12580=>"110110100",
  12581=>"000110101",
  12582=>"111011011",
  12583=>"010001100",
  12584=>"110001000",
  12585=>"100011110",
  12586=>"011101011",
  12587=>"100010000",
  12588=>"110100111",
  12589=>"000000000",
  12590=>"010000000",
  12591=>"011110111",
  12592=>"000010101",
  12593=>"011110110",
  12594=>"100101110",
  12595=>"111011110",
  12596=>"010001000",
  12597=>"100000001",
  12598=>"111010100",
  12599=>"110001001",
  12600=>"000000101",
  12601=>"100000111",
  12602=>"001101100",
  12603=>"111010010",
  12604=>"000011111",
  12605=>"000111101",
  12606=>"111001010",
  12607=>"111110101",
  12608=>"110111010",
  12609=>"100101110",
  12610=>"011101010",
  12611=>"110010100",
  12612=>"101001011",
  12613=>"000010000",
  12614=>"000001000",
  12615=>"111110011",
  12616=>"110000100",
  12617=>"010011010",
  12618=>"011100111",
  12619=>"101001000",
  12620=>"011011111",
  12621=>"100111010",
  12622=>"110110010",
  12623=>"100011000",
  12624=>"110001000",
  12625=>"110001010",
  12626=>"010011110",
  12627=>"100100111",
  12628=>"100111000",
  12629=>"111011000",
  12630=>"100010001",
  12631=>"000101000",
  12632=>"100100100",
  12633=>"000101001",
  12634=>"100011111",
  12635=>"110110010",
  12636=>"100111000",
  12637=>"011101101",
  12638=>"101111110",
  12639=>"111000101",
  12640=>"001101111",
  12641=>"110000010",
  12642=>"111011011",
  12643=>"000000101",
  12644=>"000010000",
  12645=>"111010101",
  12646=>"001011000",
  12647=>"011001111",
  12648=>"100100000",
  12649=>"010001000",
  12650=>"011100111",
  12651=>"000011111",
  12652=>"111101001",
  12653=>"111100001",
  12654=>"010001100",
  12655=>"010110000",
  12656=>"000110001",
  12657=>"101111011",
  12658=>"100001010",
  12659=>"001101000",
  12660=>"110111000",
  12661=>"100110101",
  12662=>"110001111",
  12663=>"100101110",
  12664=>"011111111",
  12665=>"001100000",
  12666=>"100111011",
  12667=>"101001111",
  12668=>"110111111",
  12669=>"111011100",
  12670=>"000100011",
  12671=>"111010011",
  12672=>"000101000",
  12673=>"001010000",
  12674=>"100000101",
  12675=>"001000010",
  12676=>"011111011",
  12677=>"001100000",
  12678=>"001010010",
  12679=>"011001110",
  12680=>"110000000",
  12681=>"001010100",
  12682=>"000001100",
  12683=>"001111101",
  12684=>"000111011",
  12685=>"011011000",
  12686=>"110000110",
  12687=>"010011101",
  12688=>"011000111",
  12689=>"000101010",
  12690=>"100011101",
  12691=>"110101000",
  12692=>"011011000",
  12693=>"001000011",
  12694=>"000100110",
  12695=>"111001000",
  12696=>"110110000",
  12697=>"100111111",
  12698=>"101001001",
  12699=>"010001101",
  12700=>"111000000",
  12701=>"101110100",
  12702=>"011000010",
  12703=>"011000101",
  12704=>"110110010",
  12705=>"000001011",
  12706=>"110001101",
  12707=>"000001010",
  12708=>"101111010",
  12709=>"001111001",
  12710=>"100100010",
  12711=>"101011111",
  12712=>"110100000",
  12713=>"101000001",
  12714=>"100100100",
  12715=>"001001111",
  12716=>"010000100",
  12717=>"110011110",
  12718=>"001010100",
  12719=>"001011000",
  12720=>"111111000",
  12721=>"001000101",
  12722=>"110001110",
  12723=>"100010011",
  12724=>"100000010",
  12725=>"011111011",
  12726=>"000000111",
  12727=>"011111010",
  12728=>"101100011",
  12729=>"111110000",
  12730=>"011011110",
  12731=>"111111100",
  12732=>"110100000",
  12733=>"110001001",
  12734=>"001111101",
  12735=>"110111001",
  12736=>"010001101",
  12737=>"100000101",
  12738=>"011000101",
  12739=>"010001110",
  12740=>"001000010",
  12741=>"011100011",
  12742=>"101100111",
  12743=>"110001101",
  12744=>"101000000",
  12745=>"100000011",
  12746=>"111000000",
  12747=>"001001100",
  12748=>"000101010",
  12749=>"110001000",
  12750=>"010100001",
  12751=>"000100010",
  12752=>"011101110",
  12753=>"001011011",
  12754=>"000111011",
  12755=>"111111110",
  12756=>"011011010",
  12757=>"100110111",
  12758=>"010100000",
  12759=>"010000100",
  12760=>"100001010",
  12761=>"011010100",
  12762=>"110010010",
  12763=>"111000110",
  12764=>"010001010",
  12765=>"001000100",
  12766=>"000111100",
  12767=>"110010100",
  12768=>"000001110",
  12769=>"001011100",
  12770=>"101000000",
  12771=>"110010111",
  12772=>"110101011",
  12773=>"001111101",
  12774=>"110101101",
  12775=>"001100001",
  12776=>"010011001",
  12777=>"011111010",
  12778=>"000110011",
  12779=>"110100000",
  12780=>"111111011",
  12781=>"101000010",
  12782=>"101001111",
  12783=>"111010110",
  12784=>"011110110",
  12785=>"101111101",
  12786=>"111010100",
  12787=>"111101100",
  12788=>"110011010",
  12789=>"111111000",
  12790=>"110010111",
  12791=>"010001111",
  12792=>"100000110",
  12793=>"001110111",
  12794=>"011100101",
  12795=>"100000010",
  12796=>"010010101",
  12797=>"100100001",
  12798=>"001010000",
  12799=>"100011001",
  12800=>"001000010",
  12801=>"001011010",
  12802=>"101110010",
  12803=>"101001011",
  12804=>"111100111",
  12805=>"011000001",
  12806=>"101001100",
  12807=>"110001000",
  12808=>"010000010",
  12809=>"000011001",
  12810=>"000010001",
  12811=>"000010100",
  12812=>"100010101",
  12813=>"100100011",
  12814=>"111110011",
  12815=>"001100100",
  12816=>"100110101",
  12817=>"111100011",
  12818=>"111100100",
  12819=>"111111011",
  12820=>"001001011",
  12821=>"101000010",
  12822=>"111110100",
  12823=>"111001010",
  12824=>"110000101",
  12825=>"110001110",
  12826=>"011001111",
  12827=>"111110101",
  12828=>"000100100",
  12829=>"111100001",
  12830=>"110010110",
  12831=>"000110001",
  12832=>"100001110",
  12833=>"000100011",
  12834=>"000001100",
  12835=>"101101110",
  12836=>"111110111",
  12837=>"010101010",
  12838=>"001000110",
  12839=>"110011101",
  12840=>"000000001",
  12841=>"101100011",
  12842=>"111110011",
  12843=>"111011111",
  12844=>"010001101",
  12845=>"001100100",
  12846=>"101010000",
  12847=>"001001001",
  12848=>"101011001",
  12849=>"111111011",
  12850=>"001001000",
  12851=>"100101100",
  12852=>"001101110",
  12853=>"010010000",
  12854=>"011011101",
  12855=>"111011111",
  12856=>"010100110",
  12857=>"011100101",
  12858=>"010111011",
  12859=>"100010000",
  12860=>"101111101",
  12861=>"010010000",
  12862=>"010111001",
  12863=>"010110111",
  12864=>"111001101",
  12865=>"011011011",
  12866=>"000010011",
  12867=>"101010001",
  12868=>"111001001",
  12869=>"110101101",
  12870=>"000100100",
  12871=>"000100100",
  12872=>"001100011",
  12873=>"011111111",
  12874=>"000001101",
  12875=>"111111010",
  12876=>"100001111",
  12877=>"111111101",
  12878=>"001111010",
  12879=>"101111100",
  12880=>"010101010",
  12881=>"011111011",
  12882=>"111001011",
  12883=>"001001010",
  12884=>"101000010",
  12885=>"000100001",
  12886=>"001000000",
  12887=>"000110010",
  12888=>"000000110",
  12889=>"010001101",
  12890=>"101100011",
  12891=>"000001110",
  12892=>"000110011",
  12893=>"100000001",
  12894=>"101110111",
  12895=>"111011001",
  12896=>"001100011",
  12897=>"100000010",
  12898=>"100001100",
  12899=>"000011010",
  12900=>"011000001",
  12901=>"100000000",
  12902=>"110100000",
  12903=>"001111110",
  12904=>"100000000",
  12905=>"101010111",
  12906=>"100110101",
  12907=>"010111011",
  12908=>"001001111",
  12909=>"100110111",
  12910=>"011111000",
  12911=>"000111110",
  12912=>"001001001",
  12913=>"101110110",
  12914=>"010010101",
  12915=>"001001010",
  12916=>"101101111",
  12917=>"000001000",
  12918=>"010000111",
  12919=>"110111011",
  12920=>"011000101",
  12921=>"101001100",
  12922=>"101011100",
  12923=>"010010100",
  12924=>"101101010",
  12925=>"001010001",
  12926=>"100111111",
  12927=>"110011001",
  12928=>"110010010",
  12929=>"011111100",
  12930=>"011011000",
  12931=>"000111101",
  12932=>"000100001",
  12933=>"100111111",
  12934=>"101101101",
  12935=>"111101011",
  12936=>"001110011",
  12937=>"110000001",
  12938=>"101111011",
  12939=>"011110010",
  12940=>"011011000",
  12941=>"011100011",
  12942=>"001001011",
  12943=>"000000010",
  12944=>"111010001",
  12945=>"011011110",
  12946=>"011011101",
  12947=>"111101110",
  12948=>"101111110",
  12949=>"010001001",
  12950=>"001100110",
  12951=>"101001100",
  12952=>"010001010",
  12953=>"000000011",
  12954=>"011110010",
  12955=>"111000100",
  12956=>"000000111",
  12957=>"011011000",
  12958=>"010111011",
  12959=>"100010001",
  12960=>"010111001",
  12961=>"100011010",
  12962=>"100111001",
  12963=>"010011111",
  12964=>"001010000",
  12965=>"001001011",
  12966=>"011001001",
  12967=>"010000010",
  12968=>"010010101",
  12969=>"111001000",
  12970=>"001101000",
  12971=>"101011111",
  12972=>"111111001",
  12973=>"000001001",
  12974=>"110100100",
  12975=>"001101100",
  12976=>"000110100",
  12977=>"000000000",
  12978=>"111110111",
  12979=>"111000010",
  12980=>"000000001",
  12981=>"111100100",
  12982=>"100111000",
  12983=>"101100010",
  12984=>"101010101",
  12985=>"000100110",
  12986=>"101111110",
  12987=>"010000001",
  12988=>"100000000",
  12989=>"110110001",
  12990=>"011010101",
  12991=>"000101110",
  12992=>"111001011",
  12993=>"000001001",
  12994=>"000011001",
  12995=>"010101000",
  12996=>"111110110",
  12997=>"110110111",
  12998=>"110010110",
  12999=>"000001101",
  13000=>"100000010",
  13001=>"010001011",
  13002=>"001000010",
  13003=>"000001111",
  13004=>"100010010",
  13005=>"100111011",
  13006=>"010101010",
  13007=>"100101000",
  13008=>"010110100",
  13009=>"001001101",
  13010=>"100101011",
  13011=>"110001000",
  13012=>"110001100",
  13013=>"100010110",
  13014=>"010110000",
  13015=>"001000101",
  13016=>"000000110",
  13017=>"100101101",
  13018=>"011100010",
  13019=>"111111110",
  13020=>"100101111",
  13021=>"110001010",
  13022=>"100011100",
  13023=>"000101101",
  13024=>"001011101",
  13025=>"111000111",
  13026=>"011001000",
  13027=>"101100110",
  13028=>"000100110",
  13029=>"011100111",
  13030=>"101001100",
  13031=>"010110111",
  13032=>"001001000",
  13033=>"101110000",
  13034=>"010100001",
  13035=>"000001111",
  13036=>"110000010",
  13037=>"000010000",
  13038=>"110111000",
  13039=>"110111110",
  13040=>"001000111",
  13041=>"101011010",
  13042=>"010110100",
  13043=>"111110100",
  13044=>"110110010",
  13045=>"001001100",
  13046=>"100110110",
  13047=>"100000101",
  13048=>"111111111",
  13049=>"111000000",
  13050=>"111111001",
  13051=>"001000100",
  13052=>"110010001",
  13053=>"011001010",
  13054=>"110101001",
  13055=>"100111101",
  13056=>"111010000",
  13057=>"000000110",
  13058=>"001110011",
  13059=>"110100011",
  13060=>"111110100",
  13061=>"010110010",
  13062=>"010011110",
  13063=>"111111110",
  13064=>"000100101",
  13065=>"011101111",
  13066=>"101001101",
  13067=>"010001011",
  13068=>"011001011",
  13069=>"110010011",
  13070=>"011111011",
  13071=>"001111100",
  13072=>"111000101",
  13073=>"111110011",
  13074=>"101101000",
  13075=>"100011001",
  13076=>"110110001",
  13077=>"111011101",
  13078=>"111100001",
  13079=>"010001010",
  13080=>"110111010",
  13081=>"001010010",
  13082=>"110100100",
  13083=>"000011000",
  13084=>"001001110",
  13085=>"000010110",
  13086=>"000011000",
  13087=>"100101010",
  13088=>"001110010",
  13089=>"001001100",
  13090=>"101001110",
  13091=>"001100111",
  13092=>"000010010",
  13093=>"000001010",
  13094=>"010000001",
  13095=>"010011000",
  13096=>"000000100",
  13097=>"101100101",
  13098=>"111100100",
  13099=>"011011100",
  13100=>"000000001",
  13101=>"110010001",
  13102=>"111000110",
  13103=>"100111110",
  13104=>"000001010",
  13105=>"010110010",
  13106=>"000110101",
  13107=>"010000101",
  13108=>"111000111",
  13109=>"000000111",
  13110=>"100100010",
  13111=>"011100010",
  13112=>"000101010",
  13113=>"000000111",
  13114=>"101000000",
  13115=>"100110111",
  13116=>"111101110",
  13117=>"000110010",
  13118=>"101000011",
  13119=>"110111101",
  13120=>"110101101",
  13121=>"011101101",
  13122=>"111001111",
  13123=>"101001100",
  13124=>"100001111",
  13125=>"000011000",
  13126=>"110101110",
  13127=>"000100101",
  13128=>"111111110",
  13129=>"100011110",
  13130=>"001111111",
  13131=>"100001110",
  13132=>"010010010",
  13133=>"111100101",
  13134=>"000001010",
  13135=>"001010010",
  13136=>"110100010",
  13137=>"000011110",
  13138=>"111100101",
  13139=>"111100000",
  13140=>"010000110",
  13141=>"101101001",
  13142=>"000010111",
  13143=>"011111111",
  13144=>"010001001",
  13145=>"010010000",
  13146=>"100011000",
  13147=>"110000101",
  13148=>"111001100",
  13149=>"110000011",
  13150=>"010111001",
  13151=>"011001011",
  13152=>"111110011",
  13153=>"000000010",
  13154=>"000010101",
  13155=>"111101011",
  13156=>"101110010",
  13157=>"100010010",
  13158=>"111100111",
  13159=>"011001101",
  13160=>"011001101",
  13161=>"000000010",
  13162=>"100001100",
  13163=>"100000100",
  13164=>"110000010",
  13165=>"010101100",
  13166=>"100101110",
  13167=>"011100111",
  13168=>"010001111",
  13169=>"110100010",
  13170=>"010011100",
  13171=>"001011001",
  13172=>"000011000",
  13173=>"110010001",
  13174=>"000001010",
  13175=>"111101100",
  13176=>"110001000",
  13177=>"010001101",
  13178=>"101000001",
  13179=>"011010110",
  13180=>"011011110",
  13181=>"111001011",
  13182=>"100011111",
  13183=>"011111111",
  13184=>"000111000",
  13185=>"001110000",
  13186=>"001100110",
  13187=>"000100100",
  13188=>"111101101",
  13189=>"111011100",
  13190=>"010101011",
  13191=>"010000111",
  13192=>"101000101",
  13193=>"110101101",
  13194=>"010000111",
  13195=>"000110110",
  13196=>"010000000",
  13197=>"100111000",
  13198=>"010011010",
  13199=>"100110000",
  13200=>"011001010",
  13201=>"001111010",
  13202=>"000110001",
  13203=>"000011000",
  13204=>"101010101",
  13205=>"100000001",
  13206=>"101100011",
  13207=>"111010110",
  13208=>"100100011",
  13209=>"100010110",
  13210=>"110111011",
  13211=>"100101011",
  13212=>"110100110",
  13213=>"101010010",
  13214=>"000100011",
  13215=>"000110101",
  13216=>"001001101",
  13217=>"110110111",
  13218=>"000111101",
  13219=>"000000111",
  13220=>"110101010",
  13221=>"000000001",
  13222=>"000101101",
  13223=>"001000000",
  13224=>"100000001",
  13225=>"110010110",
  13226=>"111111100",
  13227=>"000001111",
  13228=>"001111100",
  13229=>"000000000",
  13230=>"001100111",
  13231=>"100001000",
  13232=>"101000011",
  13233=>"101001100",
  13234=>"101011110",
  13235=>"010100010",
  13236=>"000010010",
  13237=>"011001110",
  13238=>"110100100",
  13239=>"011101101",
  13240=>"100000011",
  13241=>"001010101",
  13242=>"001000010",
  13243=>"111110011",
  13244=>"110100011",
  13245=>"110010011",
  13246=>"011110011",
  13247=>"111011011",
  13248=>"010111111",
  13249=>"110000010",
  13250=>"111100101",
  13251=>"100000110",
  13252=>"110001011",
  13253=>"111100110",
  13254=>"000101010",
  13255=>"010101100",
  13256=>"000010001",
  13257=>"000011111",
  13258=>"111100100",
  13259=>"000110100",
  13260=>"000111110",
  13261=>"100111110",
  13262=>"000011100",
  13263=>"011010110",
  13264=>"011100110",
  13265=>"101001110",
  13266=>"011011001",
  13267=>"110101010",
  13268=>"011000011",
  13269=>"110000100",
  13270=>"000110000",
  13271=>"000001111",
  13272=>"110100000",
  13273=>"001111001",
  13274=>"011010110",
  13275=>"111110101",
  13276=>"110010111",
  13277=>"100011000",
  13278=>"110100110",
  13279=>"011000011",
  13280=>"111110111",
  13281=>"011000101",
  13282=>"101011111",
  13283=>"111110001",
  13284=>"010001010",
  13285=>"110010110",
  13286=>"111101110",
  13287=>"010010001",
  13288=>"000010001",
  13289=>"111110000",
  13290=>"001000110",
  13291=>"011101011",
  13292=>"011010110",
  13293=>"000000000",
  13294=>"000001101",
  13295=>"001100110",
  13296=>"011011101",
  13297=>"100000001",
  13298=>"001011111",
  13299=>"010010100",
  13300=>"010101011",
  13301=>"011100100",
  13302=>"011111001",
  13303=>"011000101",
  13304=>"000000111",
  13305=>"011000000",
  13306=>"101111111",
  13307=>"111100001",
  13308=>"000001000",
  13309=>"110011101",
  13310=>"010010010",
  13311=>"011111001",
  13312=>"010000101",
  13313=>"111101100",
  13314=>"100001001",
  13315=>"110111011",
  13316=>"001111101",
  13317=>"111010010",
  13318=>"011110010",
  13319=>"111000000",
  13320=>"101011011",
  13321=>"010000000",
  13322=>"101111100",
  13323=>"000010000",
  13324=>"100000100",
  13325=>"000000000",
  13326=>"111111111",
  13327=>"001100111",
  13328=>"101010101",
  13329=>"101001111",
  13330=>"111011101",
  13331=>"100111101",
  13332=>"000000000",
  13333=>"101010011",
  13334=>"110110010",
  13335=>"010011000",
  13336=>"001000110",
  13337=>"001101011",
  13338=>"101101101",
  13339=>"101111110",
  13340=>"011001010",
  13341=>"101001001",
  13342=>"010111000",
  13343=>"111110110",
  13344=>"010010101",
  13345=>"001011111",
  13346=>"000011000",
  13347=>"111001010",
  13348=>"100110111",
  13349=>"111101000",
  13350=>"101001010",
  13351=>"110110010",
  13352=>"000011011",
  13353=>"101000010",
  13354=>"110111001",
  13355=>"000110101",
  13356=>"000000101",
  13357=>"000100101",
  13358=>"000011111",
  13359=>"000001101",
  13360=>"000000111",
  13361=>"001011001",
  13362=>"100110101",
  13363=>"010000011",
  13364=>"110001100",
  13365=>"111111001",
  13366=>"111000001",
  13367=>"100010001",
  13368=>"011111000",
  13369=>"111110001",
  13370=>"000100110",
  13371=>"010110110",
  13372=>"011011000",
  13373=>"111110100",
  13374=>"001100010",
  13375=>"001111100",
  13376=>"001100001",
  13377=>"000000010",
  13378=>"000101100",
  13379=>"001100001",
  13380=>"110010101",
  13381=>"101011010",
  13382=>"111101110",
  13383=>"100010101",
  13384=>"010011001",
  13385=>"101000010",
  13386=>"010110001",
  13387=>"010000001",
  13388=>"001100011",
  13389=>"111110111",
  13390=>"111111001",
  13391=>"000110100",
  13392=>"010101011",
  13393=>"010010100",
  13394=>"010011010",
  13395=>"001000001",
  13396=>"100110101",
  13397=>"110001001",
  13398=>"111000101",
  13399=>"000101011",
  13400=>"011011011",
  13401=>"101010010",
  13402=>"011011001",
  13403=>"000110110",
  13404=>"111010110",
  13405=>"100011010",
  13406=>"000011010",
  13407=>"000110011",
  13408=>"011000010",
  13409=>"001010101",
  13410=>"000111011",
  13411=>"000011001",
  13412=>"000001010",
  13413=>"011110011",
  13414=>"111101111",
  13415=>"101000100",
  13416=>"000111111",
  13417=>"110000010",
  13418=>"001000011",
  13419=>"101110001",
  13420=>"010001001",
  13421=>"101100110",
  13422=>"100000010",
  13423=>"001111111",
  13424=>"110100000",
  13425=>"110011000",
  13426=>"101010111",
  13427=>"110110101",
  13428=>"011101011",
  13429=>"111110010",
  13430=>"001100011",
  13431=>"000011000",
  13432=>"111101101",
  13433=>"011000100",
  13434=>"011100101",
  13435=>"000000110",
  13436=>"101101010",
  13437=>"000000100",
  13438=>"010011011",
  13439=>"110011101",
  13440=>"110001100",
  13441=>"000000101",
  13442=>"111000100",
  13443=>"001000110",
  13444=>"001001110",
  13445=>"001000111",
  13446=>"000111010",
  13447=>"111010100",
  13448=>"110111111",
  13449=>"100011000",
  13450=>"010001111",
  13451=>"001110111",
  13452=>"111010100",
  13453=>"011101110",
  13454=>"111100101",
  13455=>"001001110",
  13456=>"101111111",
  13457=>"000111010",
  13458=>"001011110",
  13459=>"111100101",
  13460=>"111010001",
  13461=>"010001100",
  13462=>"000011011",
  13463=>"000101101",
  13464=>"100001001",
  13465=>"010000010",
  13466=>"100100100",
  13467=>"101011101",
  13468=>"101001110",
  13469=>"111011010",
  13470=>"000000010",
  13471=>"001111110",
  13472=>"000000100",
  13473=>"110101110",
  13474=>"100000111",
  13475=>"101100100",
  13476=>"000101100",
  13477=>"101001011",
  13478=>"101001000",
  13479=>"010001111",
  13480=>"010011000",
  13481=>"011100010",
  13482=>"000010101",
  13483=>"001011101",
  13484=>"011010111",
  13485=>"101111111",
  13486=>"000011100",
  13487=>"111000011",
  13488=>"010110011",
  13489=>"010000000",
  13490=>"001000101",
  13491=>"000101000",
  13492=>"010100000",
  13493=>"111000100",
  13494=>"011101000",
  13495=>"000111010",
  13496=>"010110010",
  13497=>"001100001",
  13498=>"001010000",
  13499=>"011011100",
  13500=>"010100011",
  13501=>"010011001",
  13502=>"011000011",
  13503=>"110010000",
  13504=>"111111111",
  13505=>"110100110",
  13506=>"110101000",
  13507=>"011010011",
  13508=>"011100101",
  13509=>"010011110",
  13510=>"000111000",
  13511=>"000000000",
  13512=>"101000010",
  13513=>"001100100",
  13514=>"101100001",
  13515=>"010100001",
  13516=>"111111110",
  13517=>"010111011",
  13518=>"011001010",
  13519=>"110010100",
  13520=>"011111001",
  13521=>"100110010",
  13522=>"111001100",
  13523=>"100100111",
  13524=>"000000111",
  13525=>"001100011",
  13526=>"010011000",
  13527=>"100111110",
  13528=>"100101000",
  13529=>"111011000",
  13530=>"111011100",
  13531=>"010110000",
  13532=>"110011010",
  13533=>"100110101",
  13534=>"010101001",
  13535=>"000000001",
  13536=>"111101110",
  13537=>"011011111",
  13538=>"111010011",
  13539=>"100010100",
  13540=>"100111001",
  13541=>"010101111",
  13542=>"001011001",
  13543=>"100011110",
  13544=>"100000100",
  13545=>"101101101",
  13546=>"001001011",
  13547=>"100001100",
  13548=>"000000010",
  13549=>"101010010",
  13550=>"001100000",
  13551=>"011000000",
  13552=>"110110101",
  13553=>"101001101",
  13554=>"010010111",
  13555=>"100011011",
  13556=>"101000000",
  13557=>"001000000",
  13558=>"001100001",
  13559=>"010101111",
  13560=>"110111111",
  13561=>"000011011",
  13562=>"111100011",
  13563=>"100010110",
  13564=>"010010000",
  13565=>"101111011",
  13566=>"111010111",
  13567=>"101001111",
  13568=>"111110111",
  13569=>"010111110",
  13570=>"000001000",
  13571=>"011101001",
  13572=>"110110011",
  13573=>"101101011",
  13574=>"100101111",
  13575=>"000111011",
  13576=>"010111001",
  13577=>"001100000",
  13578=>"111101101",
  13579=>"001100001",
  13580=>"001000000",
  13581=>"111001010",
  13582=>"100110010",
  13583=>"111110010",
  13584=>"111100100",
  13585=>"010010110",
  13586=>"111011000",
  13587=>"000111111",
  13588=>"100011011",
  13589=>"101101110",
  13590=>"100101100",
  13591=>"010100000",
  13592=>"110000000",
  13593=>"000000110",
  13594=>"111100111",
  13595=>"110111100",
  13596=>"000001111",
  13597=>"011000000",
  13598=>"100010110",
  13599=>"000111010",
  13600=>"000010011",
  13601=>"110011101",
  13602=>"010111001",
  13603=>"000001100",
  13604=>"111001100",
  13605=>"001111100",
  13606=>"100101011",
  13607=>"100001001",
  13608=>"000101010",
  13609=>"110110001",
  13610=>"000100010",
  13611=>"110100010",
  13612=>"010010111",
  13613=>"111000110",
  13614=>"000001111",
  13615=>"100001100",
  13616=>"110010000",
  13617=>"100100110",
  13618=>"110101111",
  13619=>"000100110",
  13620=>"010000001",
  13621=>"101010011",
  13622=>"101100110",
  13623=>"111110000",
  13624=>"101001001",
  13625=>"111111000",
  13626=>"010111011",
  13627=>"101100010",
  13628=>"000100001",
  13629=>"011111101",
  13630=>"110000011",
  13631=>"011000111",
  13632=>"010111100",
  13633=>"001000100",
  13634=>"000000010",
  13635=>"110111110",
  13636=>"001110011",
  13637=>"111000000",
  13638=>"110101110",
  13639=>"001001001",
  13640=>"011010110",
  13641=>"001010000",
  13642=>"000011010",
  13643=>"010000000",
  13644=>"001001000",
  13645=>"111001001",
  13646=>"011001101",
  13647=>"011110000",
  13648=>"001111001",
  13649=>"110011110",
  13650=>"100010001",
  13651=>"000011001",
  13652=>"101000111",
  13653=>"110101111",
  13654=>"111101000",
  13655=>"100000110",
  13656=>"100011111",
  13657=>"000000000",
  13658=>"101001001",
  13659=>"010000100",
  13660=>"110111010",
  13661=>"011110110",
  13662=>"000100010",
  13663=>"110000001",
  13664=>"100010110",
  13665=>"010110111",
  13666=>"010100101",
  13667=>"111100011",
  13668=>"110111001",
  13669=>"000011100",
  13670=>"101000011",
  13671=>"011010110",
  13672=>"011111001",
  13673=>"010010101",
  13674=>"010010111",
  13675=>"000011011",
  13676=>"011111001",
  13677=>"100101000",
  13678=>"001101010",
  13679=>"011110010",
  13680=>"010100101",
  13681=>"100000101",
  13682=>"111111101",
  13683=>"010110010",
  13684=>"111011110",
  13685=>"011000011",
  13686=>"111000010",
  13687=>"111110001",
  13688=>"011000001",
  13689=>"000100100",
  13690=>"011001000",
  13691=>"101110000",
  13692=>"111010010",
  13693=>"110100100",
  13694=>"010001101",
  13695=>"011100100",
  13696=>"000111101",
  13697=>"010011110",
  13698=>"111010001",
  13699=>"100110111",
  13700=>"110011100",
  13701=>"010100000",
  13702=>"101010110",
  13703=>"100111101",
  13704=>"111000011",
  13705=>"101110100",
  13706=>"111011011",
  13707=>"010101001",
  13708=>"011101000",
  13709=>"111101000",
  13710=>"111010000",
  13711=>"111110001",
  13712=>"111010101",
  13713=>"001011100",
  13714=>"101000001",
  13715=>"010100001",
  13716=>"110111111",
  13717=>"001100010",
  13718=>"111001110",
  13719=>"100011011",
  13720=>"000101110",
  13721=>"001001001",
  13722=>"001010011",
  13723=>"000110000",
  13724=>"111000111",
  13725=>"000000000",
  13726=>"011010011",
  13727=>"100101000",
  13728=>"100010000",
  13729=>"010000010",
  13730=>"000000110",
  13731=>"001001101",
  13732=>"011101000",
  13733=>"101110100",
  13734=>"001110000",
  13735=>"001111001",
  13736=>"000111111",
  13737=>"111010011",
  13738=>"000100101",
  13739=>"010001000",
  13740=>"110111101",
  13741=>"001111110",
  13742=>"000001010",
  13743=>"110000110",
  13744=>"000010100",
  13745=>"011010001",
  13746=>"000100101",
  13747=>"011001000",
  13748=>"110101111",
  13749=>"111110110",
  13750=>"001111011",
  13751=>"000111100",
  13752=>"100001011",
  13753=>"010011100",
  13754=>"010010001",
  13755=>"001011101",
  13756=>"101011111",
  13757=>"010101111",
  13758=>"000001100",
  13759=>"010001011",
  13760=>"000110100",
  13761=>"100010111",
  13762=>"001010100",
  13763=>"111110111",
  13764=>"110000011",
  13765=>"000001111",
  13766=>"000010011",
  13767=>"000001001",
  13768=>"001011111",
  13769=>"010011100",
  13770=>"100100000",
  13771=>"000001110",
  13772=>"110001011",
  13773=>"111001010",
  13774=>"100000011",
  13775=>"110010010",
  13776=>"100011000",
  13777=>"001000110",
  13778=>"000011101",
  13779=>"100101011",
  13780=>"101010001",
  13781=>"010100110",
  13782=>"100011101",
  13783=>"100001100",
  13784=>"011110111",
  13785=>"010000010",
  13786=>"010101000",
  13787=>"101001110",
  13788=>"010011011",
  13789=>"111111011",
  13790=>"011010000",
  13791=>"100011011",
  13792=>"110111010",
  13793=>"100001011",
  13794=>"011000000",
  13795=>"010110100",
  13796=>"111101111",
  13797=>"111000011",
  13798=>"000000010",
  13799=>"011010001",
  13800=>"101110001",
  13801=>"110100001",
  13802=>"001110000",
  13803=>"010111000",
  13804=>"101100010",
  13805=>"101010100",
  13806=>"001100000",
  13807=>"100000010",
  13808=>"111001010",
  13809=>"111001011",
  13810=>"111010011",
  13811=>"010010100",
  13812=>"001101001",
  13813=>"100101101",
  13814=>"000100000",
  13815=>"110001111",
  13816=>"010000000",
  13817=>"001100000",
  13818=>"011010010",
  13819=>"011001000",
  13820=>"101010011",
  13821=>"011111000",
  13822=>"010001100",
  13823=>"000001000",
  13824=>"111101111",
  13825=>"010110101",
  13826=>"101100010",
  13827=>"001000001",
  13828=>"000000000",
  13829=>"100000111",
  13830=>"011100000",
  13831=>"111011000",
  13832=>"100101011",
  13833=>"101110100",
  13834=>"100001111",
  13835=>"101100011",
  13836=>"000111000",
  13837=>"100111011",
  13838=>"011100101",
  13839=>"011111011",
  13840=>"101111010",
  13841=>"111110011",
  13842=>"101111000",
  13843=>"000000100",
  13844=>"001001001",
  13845=>"101000011",
  13846=>"101000000",
  13847=>"110101011",
  13848=>"000010101",
  13849=>"101101110",
  13850=>"101011101",
  13851=>"010000000",
  13852=>"101101010",
  13853=>"011000101",
  13854=>"000111010",
  13855=>"101000110",
  13856=>"100101111",
  13857=>"101011100",
  13858=>"000101001",
  13859=>"011100010",
  13860=>"101100011",
  13861=>"001010101",
  13862=>"110001001",
  13863=>"101110000",
  13864=>"111011000",
  13865=>"101011101",
  13866=>"111000001",
  13867=>"010001011",
  13868=>"011101001",
  13869=>"100110100",
  13870=>"111001101",
  13871=>"111010000",
  13872=>"011000001",
  13873=>"010101111",
  13874=>"010000111",
  13875=>"110001100",
  13876=>"010110010",
  13877=>"100111000",
  13878=>"011111101",
  13879=>"100101101",
  13880=>"111010100",
  13881=>"000111011",
  13882=>"101100011",
  13883=>"110101010",
  13884=>"000100111",
  13885=>"100000010",
  13886=>"100001110",
  13887=>"111101000",
  13888=>"010100010",
  13889=>"000010000",
  13890=>"011101010",
  13891=>"000111100",
  13892=>"101101101",
  13893=>"101111101",
  13894=>"011101010",
  13895=>"001010000",
  13896=>"001100100",
  13897=>"010000100",
  13898=>"000111101",
  13899=>"110110011",
  13900=>"101111010",
  13901=>"101000110",
  13902=>"010101101",
  13903=>"010011110",
  13904=>"000111001",
  13905=>"111110001",
  13906=>"010101000",
  13907=>"110000001",
  13908=>"011000000",
  13909=>"110011000",
  13910=>"111011010",
  13911=>"111110101",
  13912=>"010100101",
  13913=>"111011110",
  13914=>"100101010",
  13915=>"101000101",
  13916=>"101101010",
  13917=>"110010011",
  13918=>"100111000",
  13919=>"011000001",
  13920=>"111011010",
  13921=>"100000101",
  13922=>"110001110",
  13923=>"100000010",
  13924=>"000100111",
  13925=>"101100101",
  13926=>"100001001",
  13927=>"000110101",
  13928=>"000000000",
  13929=>"101010101",
  13930=>"101010101",
  13931=>"000100011",
  13932=>"011110111",
  13933=>"110000100",
  13934=>"110110111",
  13935=>"110000011",
  13936=>"001010000",
  13937=>"100100000",
  13938=>"111101110",
  13939=>"011100011",
  13940=>"100111110",
  13941=>"100110100",
  13942=>"100100101",
  13943=>"110100110",
  13944=>"001001101",
  13945=>"000111111",
  13946=>"000011101",
  13947=>"111100111",
  13948=>"111010001",
  13949=>"001000010",
  13950=>"010100010",
  13951=>"110000011",
  13952=>"100001100",
  13953=>"011110110",
  13954=>"000101111",
  13955=>"100111000",
  13956=>"001010101",
  13957=>"010001000",
  13958=>"001001100",
  13959=>"011011110",
  13960=>"001111001",
  13961=>"010011101",
  13962=>"110011100",
  13963=>"010010111",
  13964=>"001001011",
  13965=>"111110111",
  13966=>"100011011",
  13967=>"111000101",
  13968=>"011111000",
  13969=>"011010010",
  13970=>"000011001",
  13971=>"010010001",
  13972=>"101001010",
  13973=>"100100100",
  13974=>"001010010",
  13975=>"101111001",
  13976=>"001111100",
  13977=>"101101001",
  13978=>"111101101",
  13979=>"111010110",
  13980=>"101011110",
  13981=>"101110011",
  13982=>"010011110",
  13983=>"010001011",
  13984=>"110000101",
  13985=>"011011011",
  13986=>"111000110",
  13987=>"101001101",
  13988=>"010111001",
  13989=>"101111000",
  13990=>"011100100",
  13991=>"000001011",
  13992=>"010010110",
  13993=>"100100101",
  13994=>"100100000",
  13995=>"011010010",
  13996=>"011011101",
  13997=>"100001101",
  13998=>"000100101",
  13999=>"001101110",
  14000=>"010001111",
  14001=>"001001100",
  14002=>"110101010",
  14003=>"010000101",
  14004=>"000011110",
  14005=>"110000101",
  14006=>"011110101",
  14007=>"001111011",
  14008=>"010111110",
  14009=>"001111101",
  14010=>"111011011",
  14011=>"110011000",
  14012=>"000100100",
  14013=>"001110101",
  14014=>"000111111",
  14015=>"110011110",
  14016=>"111001111",
  14017=>"101111101",
  14018=>"100111000",
  14019=>"111111011",
  14020=>"001101010",
  14021=>"110010110",
  14022=>"111000001",
  14023=>"100101011",
  14024=>"001011001",
  14025=>"101000101",
  14026=>"101100011",
  14027=>"101101110",
  14028=>"011011111",
  14029=>"100111000",
  14030=>"100010111",
  14031=>"100001111",
  14032=>"100101011",
  14033=>"101000000",
  14034=>"011110011",
  14035=>"001101110",
  14036=>"000001011",
  14037=>"000000000",
  14038=>"101000100",
  14039=>"110100101",
  14040=>"000100111",
  14041=>"001010001",
  14042=>"001111011",
  14043=>"100011000",
  14044=>"101100010",
  14045=>"101011010",
  14046=>"011100001",
  14047=>"100010001",
  14048=>"010001101",
  14049=>"001101100",
  14050=>"001101001",
  14051=>"001000111",
  14052=>"010000010",
  14053=>"100001101",
  14054=>"001011100",
  14055=>"000000001",
  14056=>"010111010",
  14057=>"100011110",
  14058=>"110001101",
  14059=>"001110010",
  14060=>"110000000",
  14061=>"111001011",
  14062=>"010011111",
  14063=>"000010111",
  14064=>"000001000",
  14065=>"101010110",
  14066=>"011111011",
  14067=>"111010000",
  14068=>"100011100",
  14069=>"000001001",
  14070=>"001010100",
  14071=>"011001111",
  14072=>"000100001",
  14073=>"001010110",
  14074=>"010011110",
  14075=>"111001100",
  14076=>"001111110",
  14077=>"110001101",
  14078=>"010110000",
  14079=>"000111100",
  14080=>"011110000",
  14081=>"010001010",
  14082=>"000011001",
  14083=>"100101101",
  14084=>"011110001",
  14085=>"101001001",
  14086=>"100100100",
  14087=>"011000111",
  14088=>"001101000",
  14089=>"000101100",
  14090=>"010100110",
  14091=>"101100100",
  14092=>"010101111",
  14093=>"111001011",
  14094=>"000001010",
  14095=>"000010000",
  14096=>"000100100",
  14097=>"010010000",
  14098=>"010001110",
  14099=>"010001111",
  14100=>"010101101",
  14101=>"110001011",
  14102=>"100100000",
  14103=>"010000000",
  14104=>"100001100",
  14105=>"110010101",
  14106=>"001101101",
  14107=>"111101011",
  14108=>"100010001",
  14109=>"110010100",
  14110=>"001010111",
  14111=>"001111011",
  14112=>"011110000",
  14113=>"000011100",
  14114=>"000110010",
  14115=>"001101100",
  14116=>"000010111",
  14117=>"000011000",
  14118=>"010001001",
  14119=>"001110011",
  14120=>"011011010",
  14121=>"111001001",
  14122=>"011101010",
  14123=>"110101001",
  14124=>"101000111",
  14125=>"100000010",
  14126=>"000101011",
  14127=>"100110010",
  14128=>"011000010",
  14129=>"001101110",
  14130=>"001011001",
  14131=>"111000001",
  14132=>"011111101",
  14133=>"101111001",
  14134=>"010111000",
  14135=>"100011000",
  14136=>"000010101",
  14137=>"110101011",
  14138=>"010000010",
  14139=>"011101101",
  14140=>"010111110",
  14141=>"111101101",
  14142=>"011001111",
  14143=>"111111111",
  14144=>"001101101",
  14145=>"011011001",
  14146=>"101101111",
  14147=>"110001100",
  14148=>"010101101",
  14149=>"111110110",
  14150=>"101011011",
  14151=>"011011111",
  14152=>"011100100",
  14153=>"111011111",
  14154=>"110011011",
  14155=>"100101000",
  14156=>"101101001",
  14157=>"101110011",
  14158=>"101010111",
  14159=>"110010111",
  14160=>"101000101",
  14161=>"101111111",
  14162=>"110000011",
  14163=>"111000000",
  14164=>"101000011",
  14165=>"001011001",
  14166=>"101100000",
  14167=>"111100010",
  14168=>"001000111",
  14169=>"010010100",
  14170=>"001000011",
  14171=>"000001000",
  14172=>"000011010",
  14173=>"100101011",
  14174=>"111101110",
  14175=>"101110010",
  14176=>"011000000",
  14177=>"010010100",
  14178=>"001000001",
  14179=>"011111110",
  14180=>"110011010",
  14181=>"011110000",
  14182=>"001000010",
  14183=>"010001101",
  14184=>"110010101",
  14185=>"110001011",
  14186=>"001100100",
  14187=>"011000110",
  14188=>"101101101",
  14189=>"001001110",
  14190=>"000010000",
  14191=>"011100010",
  14192=>"111101001",
  14193=>"100101111",
  14194=>"111000011",
  14195=>"111110100",
  14196=>"100000111",
  14197=>"010111100",
  14198=>"011111011",
  14199=>"001011010",
  14200=>"000110001",
  14201=>"000001011",
  14202=>"100011001",
  14203=>"100001100",
  14204=>"101100110",
  14205=>"110010011",
  14206=>"011010000",
  14207=>"001110111",
  14208=>"111101000",
  14209=>"011011101",
  14210=>"000110100",
  14211=>"111101101",
  14212=>"101010110",
  14213=>"111110101",
  14214=>"110011110",
  14215=>"010111110",
  14216=>"110111111",
  14217=>"101111100",
  14218=>"111101111",
  14219=>"111010001",
  14220=>"000110110",
  14221=>"110110110",
  14222=>"000001101",
  14223=>"010010010",
  14224=>"011101101",
  14225=>"010101100",
  14226=>"011000000",
  14227=>"011101111",
  14228=>"011010011",
  14229=>"001011111",
  14230=>"000010001",
  14231=>"110110001",
  14232=>"111110101",
  14233=>"001000000",
  14234=>"110001101",
  14235=>"110101001",
  14236=>"111001101",
  14237=>"111110101",
  14238=>"101100111",
  14239=>"100011111",
  14240=>"110110001",
  14241=>"000110001",
  14242=>"000111000",
  14243=>"001000100",
  14244=>"100110010",
  14245=>"101111111",
  14246=>"001101110",
  14247=>"011010000",
  14248=>"111101110",
  14249=>"001000010",
  14250=>"001101100",
  14251=>"111100001",
  14252=>"011100010",
  14253=>"001001010",
  14254=>"101010111",
  14255=>"011001110",
  14256=>"001011111",
  14257=>"101001001",
  14258=>"100011010",
  14259=>"111110000",
  14260=>"000011001",
  14261=>"110101100",
  14262=>"110101101",
  14263=>"101011111",
  14264=>"000001111",
  14265=>"000101100",
  14266=>"100000000",
  14267=>"100000010",
  14268=>"011111101",
  14269=>"000110001",
  14270=>"111001010",
  14271=>"000101101",
  14272=>"000000010",
  14273=>"101001000",
  14274=>"010111110",
  14275=>"101101100",
  14276=>"001000000",
  14277=>"010011001",
  14278=>"000110010",
  14279=>"001010001",
  14280=>"000000011",
  14281=>"000010001",
  14282=>"000100010",
  14283=>"100111000",
  14284=>"010101100",
  14285=>"000101000",
  14286=>"001101011",
  14287=>"010110110",
  14288=>"011010110",
  14289=>"111101101",
  14290=>"001100010",
  14291=>"011110000",
  14292=>"101111010",
  14293=>"010101011",
  14294=>"001000000",
  14295=>"111000010",
  14296=>"101000100",
  14297=>"000010001",
  14298=>"100001000",
  14299=>"010000001",
  14300=>"110000110",
  14301=>"101111010",
  14302=>"000001011",
  14303=>"111101101",
  14304=>"001001101",
  14305=>"101001100",
  14306=>"011010001",
  14307=>"100100111",
  14308=>"001011000",
  14309=>"001010100",
  14310=>"000000001",
  14311=>"110001000",
  14312=>"110100000",
  14313=>"100111001",
  14314=>"100110100",
  14315=>"001001101",
  14316=>"100101001",
  14317=>"111100010",
  14318=>"010101011",
  14319=>"101010111",
  14320=>"111010010",
  14321=>"010111010",
  14322=>"101001001",
  14323=>"111001010",
  14324=>"010101111",
  14325=>"100011000",
  14326=>"010000111",
  14327=>"000100101",
  14328=>"101111000",
  14329=>"011100001",
  14330=>"101111100",
  14331=>"001101000",
  14332=>"001110001",
  14333=>"111010101",
  14334=>"010001111",
  14335=>"011110111",
  14336=>"101111101",
  14337=>"011011101",
  14338=>"011100101",
  14339=>"001001111",
  14340=>"101110100",
  14341=>"010010111",
  14342=>"111010110",
  14343=>"000001111",
  14344=>"001111011",
  14345=>"000001100",
  14346=>"100011111",
  14347=>"101011000",
  14348=>"101010010",
  14349=>"010110000",
  14350=>"001110110",
  14351=>"110100110",
  14352=>"001100100",
  14353=>"101001100",
  14354=>"010000101",
  14355=>"110110100",
  14356=>"001111000",
  14357=>"000100111",
  14358=>"101001101",
  14359=>"001101001",
  14360=>"000110011",
  14361=>"010111110",
  14362=>"010110111",
  14363=>"101101111",
  14364=>"110001100",
  14365=>"100111101",
  14366=>"000100111",
  14367=>"000000001",
  14368=>"110000011",
  14369=>"111110010",
  14370=>"000011100",
  14371=>"000000000",
  14372=>"010001001",
  14373=>"000001011",
  14374=>"001010101",
  14375=>"110101000",
  14376=>"100100011",
  14377=>"100100101",
  14378=>"110100111",
  14379=>"101110001",
  14380=>"100000110",
  14381=>"101101110",
  14382=>"111010011",
  14383=>"011101101",
  14384=>"000101000",
  14385=>"110110111",
  14386=>"110010110",
  14387=>"101010000",
  14388=>"010000101",
  14389=>"110110010",
  14390=>"001000000",
  14391=>"010001100",
  14392=>"100000011",
  14393=>"010101111",
  14394=>"000110100",
  14395=>"110010100",
  14396=>"010000110",
  14397=>"110000111",
  14398=>"011101110",
  14399=>"111010100",
  14400=>"110000011",
  14401=>"010110110",
  14402=>"000101011",
  14403=>"111001100",
  14404=>"011111111",
  14405=>"000111001",
  14406=>"001110100",
  14407=>"001000011",
  14408=>"111010111",
  14409=>"111011111",
  14410=>"011011000",
  14411=>"111010000",
  14412=>"110010101",
  14413=>"100001011",
  14414=>"000010101",
  14415=>"011101011",
  14416=>"011000110",
  14417=>"010111101",
  14418=>"100101100",
  14419=>"001010111",
  14420=>"110101101",
  14421=>"001101100",
  14422=>"110101000",
  14423=>"000001011",
  14424=>"100011101",
  14425=>"101010001",
  14426=>"010111011",
  14427=>"100010101",
  14428=>"000011110",
  14429=>"001011000",
  14430=>"111000011",
  14431=>"111100101",
  14432=>"011100101",
  14433=>"000011101",
  14434=>"001001011",
  14435=>"111101010",
  14436=>"000011111",
  14437=>"011000001",
  14438=>"000010010",
  14439=>"101110000",
  14440=>"011000010",
  14441=>"010000111",
  14442=>"110100110",
  14443=>"111001100",
  14444=>"000110011",
  14445=>"001000100",
  14446=>"111011011",
  14447=>"111000001",
  14448=>"000011111",
  14449=>"111111101",
  14450=>"000000001",
  14451=>"011110010",
  14452=>"001101111",
  14453=>"001001000",
  14454=>"100111111",
  14455=>"111110111",
  14456=>"000110001",
  14457=>"010011101",
  14458=>"111101011",
  14459=>"110001101",
  14460=>"101110000",
  14461=>"000111100",
  14462=>"111101111",
  14463=>"001000100",
  14464=>"001100100",
  14465=>"111010001",
  14466=>"010101100",
  14467=>"011111000",
  14468=>"100011010",
  14469=>"001101000",
  14470=>"111001010",
  14471=>"001011000",
  14472=>"000111110",
  14473=>"010010110",
  14474=>"100010110",
  14475=>"111001111",
  14476=>"110101011",
  14477=>"101001001",
  14478=>"110101011",
  14479=>"011101101",
  14480=>"110000000",
  14481=>"011111110",
  14482=>"101101001",
  14483=>"001101111",
  14484=>"010100111",
  14485=>"011001011",
  14486=>"000000000",
  14487=>"011111011",
  14488=>"011010000",
  14489=>"010001011",
  14490=>"011001000",
  14491=>"100101001",
  14492=>"100001000",
  14493=>"101110111",
  14494=>"001011010",
  14495=>"001011010",
  14496=>"101101111",
  14497=>"110100010",
  14498=>"011101000",
  14499=>"010001111",
  14500=>"100100011",
  14501=>"100100010",
  14502=>"000110001",
  14503=>"110001000",
  14504=>"111101110",
  14505=>"100010110",
  14506=>"000100001",
  14507=>"110111101",
  14508=>"001100100",
  14509=>"001000110",
  14510=>"011111001",
  14511=>"100110100",
  14512=>"111011111",
  14513=>"111011010",
  14514=>"001101101",
  14515=>"010110111",
  14516=>"001001010",
  14517=>"011100111",
  14518=>"011101010",
  14519=>"000010001",
  14520=>"100000100",
  14521=>"000110010",
  14522=>"101010001",
  14523=>"110111110",
  14524=>"010111111",
  14525=>"110011110",
  14526=>"101111000",
  14527=>"001011000",
  14528=>"001000100",
  14529=>"011011010",
  14530=>"101100101",
  14531=>"000110000",
  14532=>"100110110",
  14533=>"011010000",
  14534=>"010000110",
  14535=>"001111110",
  14536=>"101111101",
  14537=>"100010000",
  14538=>"100010101",
  14539=>"001000000",
  14540=>"110110110",
  14541=>"101111011",
  14542=>"001010010",
  14543=>"000010011",
  14544=>"111011010",
  14545=>"000111000",
  14546=>"101101011",
  14547=>"001011110",
  14548=>"000000010",
  14549=>"100100111",
  14550=>"100101111",
  14551=>"000011111",
  14552=>"010010000",
  14553=>"000100010",
  14554=>"101101010",
  14555=>"001001010",
  14556=>"001010000",
  14557=>"001010010",
  14558=>"111101110",
  14559=>"011110100",
  14560=>"000010000",
  14561=>"001110111",
  14562=>"101110010",
  14563=>"110110000",
  14564=>"110100110",
  14565=>"011000100",
  14566=>"011000000",
  14567=>"010001001",
  14568=>"001000001",
  14569=>"000000001",
  14570=>"100101100",
  14571=>"101000001",
  14572=>"101111011",
  14573=>"000110100",
  14574=>"111101011",
  14575=>"010011010",
  14576=>"110010111",
  14577=>"000110000",
  14578=>"010111001",
  14579=>"000011001",
  14580=>"100011101",
  14581=>"010110011",
  14582=>"000101110",
  14583=>"111000111",
  14584=>"100111111",
  14585=>"010011011",
  14586=>"110000110",
  14587=>"110011100",
  14588=>"010000101",
  14589=>"111000101",
  14590=>"101100011",
  14591=>"101011101",
  14592=>"100111000",
  14593=>"000101001",
  14594=>"100001011",
  14595=>"101101010",
  14596=>"001010110",
  14597=>"010100001",
  14598=>"100001101",
  14599=>"101001000",
  14600=>"011001111",
  14601=>"000111010",
  14602=>"111111101",
  14603=>"100000100",
  14604=>"000000001",
  14605=>"001010100",
  14606=>"000010010",
  14607=>"010010001",
  14608=>"101011000",
  14609=>"110101000",
  14610=>"100001011",
  14611=>"101010101",
  14612=>"111101001",
  14613=>"110000001",
  14614=>"111001001",
  14615=>"000111010",
  14616=>"011010011",
  14617=>"100110001",
  14618=>"000110010",
  14619=>"111001101",
  14620=>"000110000",
  14621=>"011110011",
  14622=>"111011011",
  14623=>"111000110",
  14624=>"011000000",
  14625=>"000001100",
  14626=>"000101010",
  14627=>"110101000",
  14628=>"110010000",
  14629=>"001100001",
  14630=>"010110101",
  14631=>"110101111",
  14632=>"110001010",
  14633=>"000100010",
  14634=>"000000011",
  14635=>"100001101",
  14636=>"011111111",
  14637=>"000011000",
  14638=>"111001110",
  14639=>"011000110",
  14640=>"110011101",
  14641=>"110111001",
  14642=>"111010101",
  14643=>"010011111",
  14644=>"110110101",
  14645=>"000001001",
  14646=>"011001100",
  14647=>"111110101",
  14648=>"110100000",
  14649=>"011101101",
  14650=>"001001111",
  14651=>"111101101",
  14652=>"010100000",
  14653=>"001010001",
  14654=>"100001000",
  14655=>"001110001",
  14656=>"000111010",
  14657=>"111010111",
  14658=>"000011010",
  14659=>"101110101",
  14660=>"010010100",
  14661=>"111010010",
  14662=>"111000001",
  14663=>"111001100",
  14664=>"110111011",
  14665=>"100110101",
  14666=>"111001000",
  14667=>"111010010",
  14668=>"001011101",
  14669=>"000111110",
  14670=>"000000101",
  14671=>"010000001",
  14672=>"010011111",
  14673=>"010011110",
  14674=>"100010100",
  14675=>"001010110",
  14676=>"001110100",
  14677=>"001100010",
  14678=>"010111010",
  14679=>"000111101",
  14680=>"001010001",
  14681=>"101010000",
  14682=>"010001011",
  14683=>"111010000",
  14684=>"111011111",
  14685=>"000101111",
  14686=>"010010001",
  14687=>"010000111",
  14688=>"110001111",
  14689=>"010000100",
  14690=>"000110001",
  14691=>"001110011",
  14692=>"001110011",
  14693=>"100101101",
  14694=>"011111011",
  14695=>"000100001",
  14696=>"101000101",
  14697=>"111011100",
  14698=>"100000101",
  14699=>"001000011",
  14700=>"000110101",
  14701=>"111111000",
  14702=>"100001010",
  14703=>"111000110",
  14704=>"110100001",
  14705=>"000000111",
  14706=>"011001011",
  14707=>"101000001",
  14708=>"111110100",
  14709=>"010100111",
  14710=>"000010111",
  14711=>"000101001",
  14712=>"011101000",
  14713=>"011001001",
  14714=>"111100110",
  14715=>"011110101",
  14716=>"100110110",
  14717=>"000000110",
  14718=>"001001110",
  14719=>"010101100",
  14720=>"110100010",
  14721=>"010110001",
  14722=>"100101010",
  14723=>"100000000",
  14724=>"111101111",
  14725=>"010001001",
  14726=>"001110001",
  14727=>"001110110",
  14728=>"000000110",
  14729=>"001011001",
  14730=>"001101111",
  14731=>"010001110",
  14732=>"111010101",
  14733=>"000000101",
  14734=>"101011110",
  14735=>"001100100",
  14736=>"011101100",
  14737=>"001101000",
  14738=>"010010000",
  14739=>"000100011",
  14740=>"010101001",
  14741=>"000101101",
  14742=>"000000010",
  14743=>"101111011",
  14744=>"100111111",
  14745=>"110011001",
  14746=>"001101110",
  14747=>"010011110",
  14748=>"000011011",
  14749=>"001100100",
  14750=>"011110101",
  14751=>"000100101",
  14752=>"111011010",
  14753=>"000010010",
  14754=>"001011100",
  14755=>"100100001",
  14756=>"110100010",
  14757=>"111100000",
  14758=>"001100100",
  14759=>"011101000",
  14760=>"111101000",
  14761=>"100010101",
  14762=>"101101110",
  14763=>"111101000",
  14764=>"010011110",
  14765=>"000101101",
  14766=>"101110111",
  14767=>"000101000",
  14768=>"000011101",
  14769=>"000010001",
  14770=>"001111101",
  14771=>"110001111",
  14772=>"010100001",
  14773=>"110011111",
  14774=>"110000110",
  14775=>"101111101",
  14776=>"111101011",
  14777=>"110111100",
  14778=>"111101110",
  14779=>"000101011",
  14780=>"110011001",
  14781=>"011110111",
  14782=>"000001101",
  14783=>"000001100",
  14784=>"010110101",
  14785=>"001101010",
  14786=>"100111001",
  14787=>"110001100",
  14788=>"111101111",
  14789=>"100000110",
  14790=>"111110101",
  14791=>"011111011",
  14792=>"110100110",
  14793=>"000110101",
  14794=>"001101010",
  14795=>"100011101",
  14796=>"101111111",
  14797=>"100100011",
  14798=>"001011001",
  14799=>"010011100",
  14800=>"110010101",
  14801=>"011111001",
  14802=>"011011110",
  14803=>"010010001",
  14804=>"110110110",
  14805=>"000011011",
  14806=>"100011011",
  14807=>"100100100",
  14808=>"001000010",
  14809=>"010110001",
  14810=>"001000011",
  14811=>"111110110",
  14812=>"111101100",
  14813=>"010001001",
  14814=>"011000101",
  14815=>"110010000",
  14816=>"011001111",
  14817=>"111110011",
  14818=>"001001000",
  14819=>"111000101",
  14820=>"000110001",
  14821=>"110101101",
  14822=>"010001011",
  14823=>"110011110",
  14824=>"000111011",
  14825=>"101111111",
  14826=>"101110011",
  14827=>"101000100",
  14828=>"000000101",
  14829=>"111011100",
  14830=>"111110011",
  14831=>"000001000",
  14832=>"100110001",
  14833=>"110011011",
  14834=>"010100111",
  14835=>"101100011",
  14836=>"000000111",
  14837=>"010100001",
  14838=>"010100100",
  14839=>"100111001",
  14840=>"010001010",
  14841=>"101000001",
  14842=>"100010010",
  14843=>"101101101",
  14844=>"111101000",
  14845=>"111101100",
  14846=>"010011011",
  14847=>"111000001",
  14848=>"111100000",
  14849=>"111010101",
  14850=>"011100010",
  14851=>"110011110",
  14852=>"010010101",
  14853=>"010111110",
  14854=>"101011000",
  14855=>"001101111",
  14856=>"101100000",
  14857=>"010010010",
  14858=>"000010000",
  14859=>"101000101",
  14860=>"000100010",
  14861=>"001100011",
  14862=>"100010011",
  14863=>"111101110",
  14864=>"000010011",
  14865=>"001000001",
  14866=>"111001111",
  14867=>"010111101",
  14868=>"000110010",
  14869=>"101111011",
  14870=>"101001011",
  14871=>"111000001",
  14872=>"010111101",
  14873=>"001000100",
  14874=>"101011011",
  14875=>"010101000",
  14876=>"000101000",
  14877=>"010000011",
  14878=>"001010010",
  14879=>"110111011",
  14880=>"110101010",
  14881=>"010000101",
  14882=>"001010110",
  14883=>"110011110",
  14884=>"001001101",
  14885=>"010000100",
  14886=>"101010001",
  14887=>"010011000",
  14888=>"000000000",
  14889=>"011010100",
  14890=>"000011101",
  14891=>"101101010",
  14892=>"111010100",
  14893=>"010001100",
  14894=>"101110011",
  14895=>"000101000",
  14896=>"100100011",
  14897=>"010110000",
  14898=>"000101111",
  14899=>"110011101",
  14900=>"011010011",
  14901=>"111001001",
  14902=>"100110111",
  14903=>"010011111",
  14904=>"000000000",
  14905=>"110001110",
  14906=>"110010101",
  14907=>"111100100",
  14908=>"001111000",
  14909=>"010111001",
  14910=>"001011001",
  14911=>"001110010",
  14912=>"110000000",
  14913=>"000011011",
  14914=>"100100111",
  14915=>"111111010",
  14916=>"100100111",
  14917=>"011011010",
  14918=>"001101111",
  14919=>"000101000",
  14920=>"011000100",
  14921=>"111100110",
  14922=>"010100010",
  14923=>"111100101",
  14924=>"010001001",
  14925=>"011101101",
  14926=>"101011001",
  14927=>"001001000",
  14928=>"011011000",
  14929=>"100110000",
  14930=>"001110110",
  14931=>"000101110",
  14932=>"010111100",
  14933=>"101001001",
  14934=>"011001000",
  14935=>"111101010",
  14936=>"001101110",
  14937=>"010001110",
  14938=>"111010001",
  14939=>"110100101",
  14940=>"000010000",
  14941=>"001000001",
  14942=>"101010110",
  14943=>"110100010",
  14944=>"010001011",
  14945=>"101000000",
  14946=>"111111111",
  14947=>"011100010",
  14948=>"100101001",
  14949=>"000000010",
  14950=>"011001111",
  14951=>"010100001",
  14952=>"000000101",
  14953=>"010010010",
  14954=>"110001111",
  14955=>"000001000",
  14956=>"101101000",
  14957=>"110100111",
  14958=>"100011110",
  14959=>"100101001",
  14960=>"110100101",
  14961=>"001110100",
  14962=>"001101100",
  14963=>"011010100",
  14964=>"101001010",
  14965=>"011100110",
  14966=>"011101000",
  14967=>"101000100",
  14968=>"000011100",
  14969=>"001010101",
  14970=>"010110101",
  14971=>"101010010",
  14972=>"001011010",
  14973=>"111001001",
  14974=>"011111100",
  14975=>"101101000",
  14976=>"010101000",
  14977=>"110001101",
  14978=>"101110010",
  14979=>"001001101",
  14980=>"100100111",
  14981=>"110000110",
  14982=>"001100001",
  14983=>"101100001",
  14984=>"111000111",
  14985=>"100110100",
  14986=>"110000100",
  14987=>"010001110",
  14988=>"001100111",
  14989=>"110001110",
  14990=>"000010111",
  14991=>"110111110",
  14992=>"010011010",
  14993=>"110011101",
  14994=>"100010110",
  14995=>"101011110",
  14996=>"001110010",
  14997=>"101001111",
  14998=>"101101111",
  14999=>"000011010",
  15000=>"000001010",
  15001=>"011010110",
  15002=>"100011010",
  15003=>"001100101",
  15004=>"101110001",
  15005=>"111101000",
  15006=>"010000100",
  15007=>"000000010",
  15008=>"101100101",
  15009=>"100110110",
  15010=>"001101111",
  15011=>"011100010",
  15012=>"110000011",
  15013=>"111000101",
  15014=>"111000011",
  15015=>"001001001",
  15016=>"111111010",
  15017=>"010101011",
  15018=>"001010100",
  15019=>"001000100",
  15020=>"001100111",
  15021=>"001001000",
  15022=>"101110111",
  15023=>"011001010",
  15024=>"101110001",
  15025=>"010111000",
  15026=>"001100000",
  15027=>"010010000",
  15028=>"010000110",
  15029=>"001011010",
  15030=>"101000001",
  15031=>"110100000",
  15032=>"101000011",
  15033=>"100010111",
  15034=>"101110010",
  15035=>"001001000",
  15036=>"100000101",
  15037=>"101001000",
  15038=>"100011011",
  15039=>"001110101",
  15040=>"110010001",
  15041=>"011101100",
  15042=>"000101110",
  15043=>"001110100",
  15044=>"110110101",
  15045=>"001000100",
  15046=>"000001110",
  15047=>"011001000",
  15048=>"000001100",
  15049=>"110000101",
  15050=>"001100110",
  15051=>"010011100",
  15052=>"000100110",
  15053=>"001111000",
  15054=>"011110100",
  15055=>"111100110",
  15056=>"010001000",
  15057=>"100001111",
  15058=>"110000111",
  15059=>"111011111",
  15060=>"101110011",
  15061=>"001110010",
  15062=>"010010010",
  15063=>"101000011",
  15064=>"000101010",
  15065=>"110111011",
  15066=>"100101101",
  15067=>"101111000",
  15068=>"111101100",
  15069=>"100010111",
  15070=>"101110011",
  15071=>"011011001",
  15072=>"101000010",
  15073=>"000010000",
  15074=>"011011001",
  15075=>"100110010",
  15076=>"101110100",
  15077=>"010000000",
  15078=>"011111101",
  15079=>"000001000",
  15080=>"001100011",
  15081=>"000101000",
  15082=>"100001000",
  15083=>"110010100",
  15084=>"111000011",
  15085=>"010100000",
  15086=>"011010010",
  15087=>"011111001",
  15088=>"010100101",
  15089=>"100011011",
  15090=>"011100110",
  15091=>"010110000",
  15092=>"011111101",
  15093=>"100110001",
  15094=>"010100111",
  15095=>"111011111",
  15096=>"110001000",
  15097=>"101000010",
  15098=>"110101101",
  15099=>"100000101",
  15100=>"011010011",
  15101=>"101000101",
  15102=>"010010111",
  15103=>"111001011",
  15104=>"000110011",
  15105=>"011111010",
  15106=>"011100101",
  15107=>"001101100",
  15108=>"000110110",
  15109=>"010100000",
  15110=>"000000101",
  15111=>"010001011",
  15112=>"100111010",
  15113=>"001011110",
  15114=>"010010010",
  15115=>"000011010",
  15116=>"010100000",
  15117=>"110011010",
  15118=>"100010010",
  15119=>"100000010",
  15120=>"110110111",
  15121=>"001101001",
  15122=>"001101100",
  15123=>"111001011",
  15124=>"010001011",
  15125=>"010100100",
  15126=>"101100101",
  15127=>"011010000",
  15128=>"010110110",
  15129=>"100000000",
  15130=>"101011110",
  15131=>"001000110",
  15132=>"101101101",
  15133=>"100010001",
  15134=>"010110001",
  15135=>"010111001",
  15136=>"110011100",
  15137=>"100000100",
  15138=>"101010000",
  15139=>"000000010",
  15140=>"100000111",
  15141=>"001101001",
  15142=>"101110100",
  15143=>"110111000",
  15144=>"101001011",
  15145=>"001110011",
  15146=>"011101000",
  15147=>"100110101",
  15148=>"011010010",
  15149=>"011010001",
  15150=>"101011111",
  15151=>"010101101",
  15152=>"110010000",
  15153=>"101011001",
  15154=>"111110110",
  15155=>"101010111",
  15156=>"100001101",
  15157=>"111010000",
  15158=>"111101101",
  15159=>"011111000",
  15160=>"001110000",
  15161=>"111101100",
  15162=>"010000110",
  15163=>"000100011",
  15164=>"110101010",
  15165=>"001011111",
  15166=>"100100110",
  15167=>"110111100",
  15168=>"010100010",
  15169=>"000011111",
  15170=>"010100101",
  15171=>"010001100",
  15172=>"011011001",
  15173=>"000101000",
  15174=>"000010000",
  15175=>"010010100",
  15176=>"100000101",
  15177=>"101110011",
  15178=>"010001111",
  15179=>"001000010",
  15180=>"101011110",
  15181=>"010111000",
  15182=>"001100100",
  15183=>"111000100",
  15184=>"011111011",
  15185=>"100100001",
  15186=>"110001000",
  15187=>"011001010",
  15188=>"011110111",
  15189=>"001101100",
  15190=>"000000011",
  15191=>"011011110",
  15192=>"111010010",
  15193=>"011000100",
  15194=>"000100011",
  15195=>"000011011",
  15196=>"001100001",
  15197=>"001100100",
  15198=>"100011010",
  15199=>"000110111",
  15200=>"100100111",
  15201=>"000100011",
  15202=>"110110111",
  15203=>"000101001",
  15204=>"001000101",
  15205=>"101010010",
  15206=>"100111010",
  15207=>"110101001",
  15208=>"101111010",
  15209=>"000101110",
  15210=>"011111101",
  15211=>"010000100",
  15212=>"010011001",
  15213=>"110011000",
  15214=>"011100000",
  15215=>"111100101",
  15216=>"010110000",
  15217=>"100000000",
  15218=>"011001100",
  15219=>"111100100",
  15220=>"000000011",
  15221=>"100001000",
  15222=>"110010100",
  15223=>"001111000",
  15224=>"000010000",
  15225=>"100100101",
  15226=>"110001110",
  15227=>"100110110",
  15228=>"000101001",
  15229=>"000000010",
  15230=>"100000001",
  15231=>"010100000",
  15232=>"111011100",
  15233=>"000001100",
  15234=>"000010011",
  15235=>"000101101",
  15236=>"111111000",
  15237=>"000001001",
  15238=>"000001000",
  15239=>"110100010",
  15240=>"001001110",
  15241=>"110101100",
  15242=>"000111100",
  15243=>"011100011",
  15244=>"001001010",
  15245=>"000100111",
  15246=>"110111001",
  15247=>"111110011",
  15248=>"100010101",
  15249=>"100111011",
  15250=>"110101011",
  15251=>"000101101",
  15252=>"110010000",
  15253=>"000100001",
  15254=>"111001011",
  15255=>"010100001",
  15256=>"110111110",
  15257=>"111010100",
  15258=>"100000100",
  15259=>"101110011",
  15260=>"110000111",
  15261=>"000000111",
  15262=>"110000000",
  15263=>"100101000",
  15264=>"011010011",
  15265=>"100001000",
  15266=>"000111101",
  15267=>"001111101",
  15268=>"110101111",
  15269=>"101100010",
  15270=>"011101101",
  15271=>"111110100",
  15272=>"111011111",
  15273=>"111100000",
  15274=>"110110001",
  15275=>"010000001",
  15276=>"010000100",
  15277=>"110000111",
  15278=>"101101101",
  15279=>"000111000",
  15280=>"111100110",
  15281=>"000101101",
  15282=>"110101111",
  15283=>"111000010",
  15284=>"011000101",
  15285=>"011011001",
  15286=>"101101011",
  15287=>"111111101",
  15288=>"111101001",
  15289=>"101000111",
  15290=>"000011111",
  15291=>"101001011",
  15292=>"111110101",
  15293=>"101000011",
  15294=>"010001110",
  15295=>"000011010",
  15296=>"101011010",
  15297=>"000011111",
  15298=>"111000011",
  15299=>"100011000",
  15300=>"000110110",
  15301=>"011010111",
  15302=>"010110100",
  15303=>"010111111",
  15304=>"000010101",
  15305=>"000001011",
  15306=>"111000010",
  15307=>"001010111",
  15308=>"011100100",
  15309=>"111100011",
  15310=>"010110101",
  15311=>"101100100",
  15312=>"110110101",
  15313=>"000111011",
  15314=>"010101000",
  15315=>"100001100",
  15316=>"011110011",
  15317=>"011110011",
  15318=>"101100001",
  15319=>"001101101",
  15320=>"100101001",
  15321=>"111011001",
  15322=>"110110101",
  15323=>"010111001",
  15324=>"010101111",
  15325=>"010101000",
  15326=>"110101100",
  15327=>"000001001",
  15328=>"111100100",
  15329=>"101111101",
  15330=>"101100111",
  15331=>"110110000",
  15332=>"100010110",
  15333=>"000110111",
  15334=>"000100011",
  15335=>"000010010",
  15336=>"010010110",
  15337=>"011010111",
  15338=>"100100000",
  15339=>"010011001",
  15340=>"000101100",
  15341=>"010011110",
  15342=>"011000000",
  15343=>"111111110",
  15344=>"011010100",
  15345=>"011111101",
  15346=>"100001111",
  15347=>"110111000",
  15348=>"000110110",
  15349=>"100011100",
  15350=>"001011010",
  15351=>"000000010",
  15352=>"010001110",
  15353=>"011111010",
  15354=>"101010101",
  15355=>"101100011",
  15356=>"100011101",
  15357=>"011111110",
  15358=>"001011010",
  15359=>"001100000",
  15360=>"001110100",
  15361=>"001101111",
  15362=>"011100100",
  15363=>"101011011",
  15364=>"100110110",
  15365=>"111101011",
  15366=>"001100010",
  15367=>"011101011",
  15368=>"001111010",
  15369=>"001110111",
  15370=>"000001101",
  15371=>"101011100",
  15372=>"100110101",
  15373=>"001101100",
  15374=>"001011110",
  15375=>"110001000",
  15376=>"101100010",
  15377=>"011000000",
  15378=>"100001100",
  15379=>"111000101",
  15380=>"111010000",
  15381=>"001001011",
  15382=>"010101100",
  15383=>"110010001",
  15384=>"000110001",
  15385=>"000010000",
  15386=>"000110000",
  15387=>"000111100",
  15388=>"010001101",
  15389=>"100101010",
  15390=>"011011010",
  15391=>"111101001",
  15392=>"100010111",
  15393=>"111001111",
  15394=>"010110000",
  15395=>"111011101",
  15396=>"001111111",
  15397=>"011101110",
  15398=>"010011000",
  15399=>"111111010",
  15400=>"000100010",
  15401=>"111011001",
  15402=>"001001001",
  15403=>"100000011",
  15404=>"010010011",
  15405=>"100101011",
  15406=>"110011010",
  15407=>"111000010",
  15408=>"100101111",
  15409=>"010000011",
  15410=>"110010111",
  15411=>"000110101",
  15412=>"010000001",
  15413=>"100000001",
  15414=>"101111010",
  15415=>"110100100",
  15416=>"010001110",
  15417=>"111111110",
  15418=>"000100110",
  15419=>"111111010",
  15420=>"000011001",
  15421=>"001011101",
  15422=>"101001110",
  15423=>"001101011",
  15424=>"000011010",
  15425=>"000001001",
  15426=>"111000010",
  15427=>"111101101",
  15428=>"011100010",
  15429=>"110111101",
  15430=>"100010101",
  15431=>"001011101",
  15432=>"011101100",
  15433=>"011001001",
  15434=>"111000001",
  15435=>"101110100",
  15436=>"011100000",
  15437=>"111011001",
  15438=>"100000000",
  15439=>"110000111",
  15440=>"011101010",
  15441=>"000110001",
  15442=>"111101101",
  15443=>"001100010",
  15444=>"110010010",
  15445=>"110011110",
  15446=>"101011101",
  15447=>"100010010",
  15448=>"110101011",
  15449=>"011001100",
  15450=>"000100101",
  15451=>"010001000",
  15452=>"011110010",
  15453=>"000111001",
  15454=>"010010010",
  15455=>"001010001",
  15456=>"111000100",
  15457=>"110100101",
  15458=>"101010001",
  15459=>"000101000",
  15460=>"111000010",
  15461=>"110101010",
  15462=>"010001000",
  15463=>"011110010",
  15464=>"010001110",
  15465=>"000110110",
  15466=>"010000010",
  15467=>"111100111",
  15468=>"000111110",
  15469=>"111001011",
  15470=>"101110001",
  15471=>"100111011",
  15472=>"000101000",
  15473=>"010001110",
  15474=>"001001011",
  15475=>"010100001",
  15476=>"000010110",
  15477=>"010110011",
  15478=>"001101001",
  15479=>"001110010",
  15480=>"111100110",
  15481=>"010100001",
  15482=>"101110111",
  15483=>"101001011",
  15484=>"110110000",
  15485=>"111011001",
  15486=>"010010111",
  15487=>"001110100",
  15488=>"001010000",
  15489=>"100110010",
  15490=>"110110011",
  15491=>"110111000",
  15492=>"101001110",
  15493=>"000011100",
  15494=>"111101100",
  15495=>"010010110",
  15496=>"111011011",
  15497=>"100101110",
  15498=>"000011100",
  15499=>"110001000",
  15500=>"101100100",
  15501=>"100111001",
  15502=>"111110101",
  15503=>"110101001",
  15504=>"111010011",
  15505=>"111000110",
  15506=>"010100001",
  15507=>"111011010",
  15508=>"100110000",
  15509=>"110100101",
  15510=>"001011100",
  15511=>"100010110",
  15512=>"000010100",
  15513=>"101111011",
  15514=>"101000000",
  15515=>"011110111",
  15516=>"011101010",
  15517=>"111010010",
  15518=>"011111100",
  15519=>"100101011",
  15520=>"110101011",
  15521=>"110110001",
  15522=>"111011001",
  15523=>"011110001",
  15524=>"011100111",
  15525=>"000100101",
  15526=>"111100101",
  15527=>"000111101",
  15528=>"111111111",
  15529=>"000010100",
  15530=>"100001100",
  15531=>"100001001",
  15532=>"011001001",
  15533=>"111011101",
  15534=>"001010100",
  15535=>"101001101",
  15536=>"111000000",
  15537=>"001101111",
  15538=>"101011111",
  15539=>"001111010",
  15540=>"111111000",
  15541=>"011111011",
  15542=>"001000000",
  15543=>"011001101",
  15544=>"110101110",
  15545=>"010010001",
  15546=>"011000001",
  15547=>"101110100",
  15548=>"111001000",
  15549=>"111111101",
  15550=>"000000011",
  15551=>"111111110",
  15552=>"001100110",
  15553=>"000011010",
  15554=>"010010001",
  15555=>"011010100",
  15556=>"110110001",
  15557=>"000110111",
  15558=>"110111101",
  15559=>"011100100",
  15560=>"010001110",
  15561=>"010010000",
  15562=>"010101000",
  15563=>"011101000",
  15564=>"101011110",
  15565=>"111110100",
  15566=>"111000101",
  15567=>"000100111",
  15568=>"010100000",
  15569=>"111010111",
  15570=>"000001010",
  15571=>"111101110",
  15572=>"100110101",
  15573=>"100111010",
  15574=>"000101011",
  15575=>"111011001",
  15576=>"011010011",
  15577=>"011000110",
  15578=>"010011100",
  15579=>"001010100",
  15580=>"011101110",
  15581=>"101011011",
  15582=>"001011111",
  15583=>"011111111",
  15584=>"100111010",
  15585=>"000101000",
  15586=>"001011000",
  15587=>"111001101",
  15588=>"111011011",
  15589=>"110101100",
  15590=>"101110101",
  15591=>"100011011",
  15592=>"110110010",
  15593=>"100010111",
  15594=>"001000001",
  15595=>"001001100",
  15596=>"101100000",
  15597=>"100010001",
  15598=>"001110001",
  15599=>"101001110",
  15600=>"011011011",
  15601=>"111111011",
  15602=>"000010010",
  15603=>"011011101",
  15604=>"000000010",
  15605=>"111010111",
  15606=>"111011100",
  15607=>"111000110",
  15608=>"001011001",
  15609=>"000010010",
  15610=>"110011100",
  15611=>"101001011",
  15612=>"011001101",
  15613=>"111001011",
  15614=>"011001010",
  15615=>"001100110",
  15616=>"111110111",
  15617=>"110011101",
  15618=>"101111111",
  15619=>"001000011",
  15620=>"111001000",
  15621=>"010001000",
  15622=>"001000010",
  15623=>"100111011",
  15624=>"110001111",
  15625=>"110110100",
  15626=>"010100011",
  15627=>"001011010",
  15628=>"100000101",
  15629=>"100000011",
  15630=>"111111011",
  15631=>"001010000",
  15632=>"001101111",
  15633=>"101011011",
  15634=>"001000100",
  15635=>"000110110",
  15636=>"001101111",
  15637=>"011101001",
  15638=>"101000001",
  15639=>"010111111",
  15640=>"101001110",
  15641=>"010011110",
  15642=>"000000000",
  15643=>"011011111",
  15644=>"011001110",
  15645=>"100110011",
  15646=>"111100111",
  15647=>"001001010",
  15648=>"111010001",
  15649=>"010100000",
  15650=>"010001100",
  15651=>"110100011",
  15652=>"011111011",
  15653=>"001100001",
  15654=>"100111110",
  15655=>"111000000",
  15656=>"000010010",
  15657=>"011000001",
  15658=>"110010101",
  15659=>"000110100",
  15660=>"000110100",
  15661=>"101101000",
  15662=>"101001001",
  15663=>"000100100",
  15664=>"101011001",
  15665=>"110000111",
  15666=>"100100111",
  15667=>"000100010",
  15668=>"111000010",
  15669=>"110000000",
  15670=>"101110101",
  15671=>"011001110",
  15672=>"001110100",
  15673=>"110101101",
  15674=>"011000001",
  15675=>"100010000",
  15676=>"110100001",
  15677=>"111010001",
  15678=>"101000101",
  15679=>"000010111",
  15680=>"011110000",
  15681=>"100011001",
  15682=>"110000110",
  15683=>"101101000",
  15684=>"101101101",
  15685=>"110100110",
  15686=>"101110111",
  15687=>"111100010",
  15688=>"011000110",
  15689=>"001101001",
  15690=>"010000011",
  15691=>"001100011",
  15692=>"001110010",
  15693=>"111010110",
  15694=>"010111110",
  15695=>"010011111",
  15696=>"010011100",
  15697=>"110011011",
  15698=>"000000100",
  15699=>"100100011",
  15700=>"111011011",
  15701=>"001110001",
  15702=>"000110000",
  15703=>"000001000",
  15704=>"100101000",
  15705=>"000110011",
  15706=>"100100110",
  15707=>"011100001",
  15708=>"110111111",
  15709=>"110111101",
  15710=>"100010111",
  15711=>"011100101",
  15712=>"111100010",
  15713=>"101001100",
  15714=>"000000001",
  15715=>"011100001",
  15716=>"100011001",
  15717=>"110011001",
  15718=>"001001101",
  15719=>"111100010",
  15720=>"010011010",
  15721=>"000001111",
  15722=>"010011011",
  15723=>"001000101",
  15724=>"111001100",
  15725=>"010001011",
  15726=>"100100001",
  15727=>"010011111",
  15728=>"100000010",
  15729=>"111111110",
  15730=>"010000011",
  15731=>"110001001",
  15732=>"000101110",
  15733=>"010001000",
  15734=>"110001001",
  15735=>"111100010",
  15736=>"100111011",
  15737=>"100110100",
  15738=>"011001101",
  15739=>"011110101",
  15740=>"011000000",
  15741=>"100111111",
  15742=>"111100111",
  15743=>"101110011",
  15744=>"000110010",
  15745=>"000001101",
  15746=>"000111000",
  15747=>"110111101",
  15748=>"010011000",
  15749=>"001001100",
  15750=>"111011000",
  15751=>"001100010",
  15752=>"111101000",
  15753=>"010101000",
  15754=>"000110111",
  15755=>"110010110",
  15756=>"101100010",
  15757=>"001010101",
  15758=>"000000101",
  15759=>"100010110",
  15760=>"000100000",
  15761=>"010111001",
  15762=>"110110000",
  15763=>"011100010",
  15764=>"010110010",
  15765=>"110100110",
  15766=>"000000000",
  15767=>"001111000",
  15768=>"110010000",
  15769=>"100100011",
  15770=>"000101100",
  15771=>"001100101",
  15772=>"000011110",
  15773=>"111000111",
  15774=>"101000110",
  15775=>"010011001",
  15776=>"100000010",
  15777=>"011111111",
  15778=>"111111010",
  15779=>"101100000",
  15780=>"011110010",
  15781=>"000011101",
  15782=>"011001000",
  15783=>"101011000",
  15784=>"001001100",
  15785=>"110011110",
  15786=>"100101010",
  15787=>"110011000",
  15788=>"010101111",
  15789=>"011010101",
  15790=>"110101111",
  15791=>"100100001",
  15792=>"101010101",
  15793=>"100011100",
  15794=>"101011111",
  15795=>"100010110",
  15796=>"110101001",
  15797=>"110010100",
  15798=>"111100001",
  15799=>"001000110",
  15800=>"011011001",
  15801=>"111110100",
  15802=>"011101111",
  15803=>"101011110",
  15804=>"101000010",
  15805=>"111010111",
  15806=>"101000100",
  15807=>"100010100",
  15808=>"010010010",
  15809=>"011100110",
  15810=>"011001001",
  15811=>"101101010",
  15812=>"110101100",
  15813=>"011110101",
  15814=>"101011110",
  15815=>"101100001",
  15816=>"111101111",
  15817=>"011100101",
  15818=>"001001000",
  15819=>"101111111",
  15820=>"000110100",
  15821=>"101110000",
  15822=>"010110100",
  15823=>"011000111",
  15824=>"111000100",
  15825=>"101110111",
  15826=>"001011001",
  15827=>"111010011",
  15828=>"001000100",
  15829=>"001100100",
  15830=>"000100010",
  15831=>"101001011",
  15832=>"010110010",
  15833=>"001010100",
  15834=>"111000110",
  15835=>"110101110",
  15836=>"101111100",
  15837=>"111110110",
  15838=>"011101011",
  15839=>"000111011",
  15840=>"001001100",
  15841=>"110001010",
  15842=>"101101101",
  15843=>"111111110",
  15844=>"010100010",
  15845=>"111001110",
  15846=>"101000101",
  15847=>"101100000",
  15848=>"001000001",
  15849=>"010001111",
  15850=>"100100111",
  15851=>"001001011",
  15852=>"101101110",
  15853=>"101101000",
  15854=>"011000100",
  15855=>"110110111",
  15856=>"000101011",
  15857=>"111000001",
  15858=>"000001111",
  15859=>"101110110",
  15860=>"000101000",
  15861=>"000001111",
  15862=>"100001011",
  15863=>"000100111",
  15864=>"100111011",
  15865=>"001110000",
  15866=>"000010010",
  15867=>"101000110",
  15868=>"000000100",
  15869=>"000111111",
  15870=>"010001011",
  15871=>"111001110",
  15872=>"010011000",
  15873=>"011100001",
  15874=>"011100111",
  15875=>"111110001",
  15876=>"110111010",
  15877=>"100100000",
  15878=>"001010011",
  15879=>"110001010",
  15880=>"000001101",
  15881=>"100010100",
  15882=>"111100111",
  15883=>"010111000",
  15884=>"010111011",
  15885=>"101100000",
  15886=>"110001100",
  15887=>"111111110",
  15888=>"100011010",
  15889=>"000000001",
  15890=>"101111111",
  15891=>"110001110",
  15892=>"011000100",
  15893=>"110001010",
  15894=>"001100111",
  15895=>"000001010",
  15896=>"010001110",
  15897=>"010111111",
  15898=>"000100011",
  15899=>"000011111",
  15900=>"110010011",
  15901=>"100001000",
  15902=>"110110001",
  15903=>"111110000",
  15904=>"011000010",
  15905=>"101000000",
  15906=>"110010111",
  15907=>"010111010",
  15908=>"000101100",
  15909=>"001111011",
  15910=>"010001010",
  15911=>"001110000",
  15912=>"000101101",
  15913=>"001111111",
  15914=>"101100101",
  15915=>"100010111",
  15916=>"001010111",
  15917=>"011000111",
  15918=>"101100110",
  15919=>"101110010",
  15920=>"111010001",
  15921=>"110011000",
  15922=>"101111110",
  15923=>"010000111",
  15924=>"001111011",
  15925=>"010000000",
  15926=>"111011010",
  15927=>"110101001",
  15928=>"001110011",
  15929=>"001111000",
  15930=>"000000010",
  15931=>"001100100",
  15932=>"100110000",
  15933=>"010001111",
  15934=>"010100001",
  15935=>"111111001",
  15936=>"111010101",
  15937=>"101010001",
  15938=>"100001111",
  15939=>"110011011",
  15940=>"010000100",
  15941=>"010011011",
  15942=>"011101010",
  15943=>"110101011",
  15944=>"000011110",
  15945=>"000001100",
  15946=>"000101110",
  15947=>"111000000",
  15948=>"011101100",
  15949=>"101011111",
  15950=>"111101110",
  15951=>"000010110",
  15952=>"101010110",
  15953=>"111011011",
  15954=>"111010010",
  15955=>"111111110",
  15956=>"100010110",
  15957=>"100011010",
  15958=>"101111011",
  15959=>"100101000",
  15960=>"100010000",
  15961=>"010111100",
  15962=>"001100000",
  15963=>"001100000",
  15964=>"101001000",
  15965=>"001000010",
  15966=>"000110010",
  15967=>"010010010",
  15968=>"010011011",
  15969=>"100111010",
  15970=>"001001010",
  15971=>"000001000",
  15972=>"010101011",
  15973=>"000101110",
  15974=>"001111111",
  15975=>"100100000",
  15976=>"100011111",
  15977=>"101100000",
  15978=>"010000101",
  15979=>"111001011",
  15980=>"110101100",
  15981=>"111010001",
  15982=>"110000100",
  15983=>"100011110",
  15984=>"110100001",
  15985=>"000011000",
  15986=>"101011011",
  15987=>"111010111",
  15988=>"101110011",
  15989=>"100000001",
  15990=>"001000100",
  15991=>"001101101",
  15992=>"100101101",
  15993=>"111101000",
  15994=>"001111100",
  15995=>"100011101",
  15996=>"000000111",
  15997=>"100011100",
  15998=>"111111011",
  15999=>"101110010",
  16000=>"011010011",
  16001=>"100110011",
  16002=>"110011001",
  16003=>"001011010",
  16004=>"000011101",
  16005=>"110000111",
  16006=>"110111000",
  16007=>"110101100",
  16008=>"011010110",
  16009=>"111110001",
  16010=>"111011101",
  16011=>"010101011",
  16012=>"100100000",
  16013=>"000110101",
  16014=>"011100111",
  16015=>"110010101",
  16016=>"011011101",
  16017=>"101101000",
  16018=>"111011100",
  16019=>"011110100",
  16020=>"011011000",
  16021=>"100000111",
  16022=>"001111010",
  16023=>"111101100",
  16024=>"110101101",
  16025=>"110101100",
  16026=>"001100001",
  16027=>"111110000",
  16028=>"010010111",
  16029=>"001000000",
  16030=>"110000000",
  16031=>"001011000",
  16032=>"010010000",
  16033=>"100100011",
  16034=>"011011101",
  16035=>"011101010",
  16036=>"111110101",
  16037=>"110001111",
  16038=>"100001101",
  16039=>"000110001",
  16040=>"110001010",
  16041=>"111100111",
  16042=>"011000010",
  16043=>"101010010",
  16044=>"000101010",
  16045=>"000011001",
  16046=>"000101101",
  16047=>"101011111",
  16048=>"000111111",
  16049=>"111100000",
  16050=>"010100010",
  16051=>"111001111",
  16052=>"010010110",
  16053=>"100010000",
  16054=>"110101010",
  16055=>"001011001",
  16056=>"110011110",
  16057=>"101110110",
  16058=>"100111011",
  16059=>"001111010",
  16060=>"111001101",
  16061=>"111001100",
  16062=>"110100100",
  16063=>"010111000",
  16064=>"000001011",
  16065=>"011111101",
  16066=>"111010001",
  16067=>"010010010",
  16068=>"000001010",
  16069=>"110000010",
  16070=>"111010100",
  16071=>"111010011",
  16072=>"001010101",
  16073=>"000010100",
  16074=>"010011111",
  16075=>"000000010",
  16076=>"011110100",
  16077=>"110111011",
  16078=>"110111111",
  16079=>"011101010",
  16080=>"010100100",
  16081=>"110001011",
  16082=>"010011111",
  16083=>"001110001",
  16084=>"000101100",
  16085=>"011110010",
  16086=>"110101110",
  16087=>"101000110",
  16088=>"101101111",
  16089=>"011010010",
  16090=>"100010001",
  16091=>"111000101",
  16092=>"000100101",
  16093=>"000110000",
  16094=>"110011101",
  16095=>"100010100",
  16096=>"111101011",
  16097=>"100011010",
  16098=>"111100101",
  16099=>"011010010",
  16100=>"110100100",
  16101=>"101101110",
  16102=>"110000001",
  16103=>"101000011",
  16104=>"101110111",
  16105=>"101110101",
  16106=>"111100000",
  16107=>"111000000",
  16108=>"010001111",
  16109=>"001010000",
  16110=>"011101000",
  16111=>"100110010",
  16112=>"000111100",
  16113=>"001110000",
  16114=>"100100010",
  16115=>"011100110",
  16116=>"010111000",
  16117=>"111000110",
  16118=>"110110000",
  16119=>"100111001",
  16120=>"110001010",
  16121=>"011110110",
  16122=>"110011010",
  16123=>"110011100",
  16124=>"000010110",
  16125=>"111110010",
  16126=>"111000010",
  16127=>"000101110",
  16128=>"000011010",
  16129=>"111111000",
  16130=>"000111010",
  16131=>"101001010",
  16132=>"000010010",
  16133=>"000011101",
  16134=>"010100011",
  16135=>"001101011",
  16136=>"000101110",
  16137=>"100010101",
  16138=>"011011000",
  16139=>"000010101",
  16140=>"110111110",
  16141=>"011100111",
  16142=>"110000001",
  16143=>"111101000",
  16144=>"110001000",
  16145=>"101001100",
  16146=>"110111100",
  16147=>"001011001",
  16148=>"011110101",
  16149=>"010001101",
  16150=>"110110100",
  16151=>"010000110",
  16152=>"011110001",
  16153=>"011100100",
  16154=>"011001100",
  16155=>"111000110",
  16156=>"000100111",
  16157=>"011111101",
  16158=>"000100100",
  16159=>"010010101",
  16160=>"100101101",
  16161=>"011000110",
  16162=>"101000000",
  16163=>"100010110",
  16164=>"100110000",
  16165=>"010101010",
  16166=>"001110101",
  16167=>"110011110",
  16168=>"101011010",
  16169=>"011001011",
  16170=>"010010101",
  16171=>"111001111",
  16172=>"010110000",
  16173=>"010001001",
  16174=>"011101110",
  16175=>"001010100",
  16176=>"011010100",
  16177=>"101011010",
  16178=>"101010000",
  16179=>"010110000",
  16180=>"110111111",
  16181=>"000100100",
  16182=>"010110001",
  16183=>"011011100",
  16184=>"011111100",
  16185=>"110100000",
  16186=>"101000010",
  16187=>"000101011",
  16188=>"010000000",
  16189=>"110101001",
  16190=>"110011000",
  16191=>"100001110",
  16192=>"101010111",
  16193=>"001001100",
  16194=>"110100111",
  16195=>"100110100",
  16196=>"111011001",
  16197=>"110001110",
  16198=>"111000100",
  16199=>"000011011",
  16200=>"001010001",
  16201=>"011001010",
  16202=>"011011011",
  16203=>"010100000",
  16204=>"001100011",
  16205=>"011010001",
  16206=>"001111001",
  16207=>"111010011",
  16208=>"100001101",
  16209=>"101100101",
  16210=>"010001011",
  16211=>"000001011",
  16212=>"001100111",
  16213=>"100010011",
  16214=>"001000101",
  16215=>"010110110",
  16216=>"010011001",
  16217=>"111101100",
  16218=>"100110100",
  16219=>"100011100",
  16220=>"100001101",
  16221=>"100000111",
  16222=>"000101101",
  16223=>"111100011",
  16224=>"001000010",
  16225=>"110100110",
  16226=>"101010110",
  16227=>"111001100",
  16228=>"100000010",
  16229=>"101100000",
  16230=>"010101110",
  16231=>"110111100",
  16232=>"111000000",
  16233=>"011101100",
  16234=>"111100111",
  16235=>"011111011",
  16236=>"100000001",
  16237=>"001010011",
  16238=>"100010001",
  16239=>"111010101",
  16240=>"110010100",
  16241=>"111111000",
  16242=>"010000011",
  16243=>"001010010",
  16244=>"111100101",
  16245=>"001000111",
  16246=>"110101000",
  16247=>"110101000",
  16248=>"110100011",
  16249=>"000100010",
  16250=>"101101111",
  16251=>"011001111",
  16252=>"111111100",
  16253=>"100010001",
  16254=>"101111101",
  16255=>"011011001",
  16256=>"011111100",
  16257=>"011100011",
  16258=>"001001100",
  16259=>"010100111",
  16260=>"011010100",
  16261=>"010110110",
  16262=>"000110011",
  16263=>"011000101",
  16264=>"000100000",
  16265=>"110101010",
  16266=>"001000100",
  16267=>"001111000",
  16268=>"010000000",
  16269=>"010100000",
  16270=>"001100001",
  16271=>"110111000",
  16272=>"111101101",
  16273=>"111110010",
  16274=>"001011000",
  16275=>"011110101",
  16276=>"010011000",
  16277=>"111001100",
  16278=>"101110101",
  16279=>"100101101",
  16280=>"000011011",
  16281=>"111000101",
  16282=>"111110101",
  16283=>"100000110",
  16284=>"011011111",
  16285=>"010001111",
  16286=>"001100001",
  16287=>"011000001",
  16288=>"000001011",
  16289=>"001110100",
  16290=>"101011100",
  16291=>"010011110",
  16292=>"111010011",
  16293=>"100101111",
  16294=>"111110001",
  16295=>"111000110",
  16296=>"000011111",
  16297=>"000100010",
  16298=>"110110111",
  16299=>"010101101",
  16300=>"001100000",
  16301=>"100100010",
  16302=>"111111101",
  16303=>"010010011",
  16304=>"000110010",
  16305=>"100111000",
  16306=>"110111100",
  16307=>"000110100",
  16308=>"111101110",
  16309=>"101100111",
  16310=>"111010001",
  16311=>"000101010",
  16312=>"010100010",
  16313=>"010101100",
  16314=>"100110100",
  16315=>"110010001",
  16316=>"010110100",
  16317=>"111010110",
  16318=>"000000110",
  16319=>"110000111",
  16320=>"010110001",
  16321=>"110101000",
  16322=>"001111001",
  16323=>"101001000",
  16324=>"100101110",
  16325=>"010001010",
  16326=>"101011000",
  16327=>"000101011",
  16328=>"100110001",
  16329=>"011010001",
  16330=>"001110111",
  16331=>"001000100",
  16332=>"011011000",
  16333=>"000100100",
  16334=>"011110110",
  16335=>"111000111",
  16336=>"110111010",
  16337=>"110110111",
  16338=>"101001100",
  16339=>"101100100",
  16340=>"111101100",
  16341=>"011011110",
  16342=>"010101000",
  16343=>"000110111",
  16344=>"100000101",
  16345=>"100010100",
  16346=>"110000000",
  16347=>"011110001",
  16348=>"001010100",
  16349=>"001111101",
  16350=>"000011000",
  16351=>"111100001",
  16352=>"001100001",
  16353=>"111001111",
  16354=>"000111101",
  16355=>"111100111",
  16356=>"001011101",
  16357=>"000000000",
  16358=>"110000011",
  16359=>"111011010",
  16360=>"011101000",
  16361=>"110110000",
  16362=>"110001011",
  16363=>"101100100",
  16364=>"001011010",
  16365=>"100111000",
  16366=>"001100110",
  16367=>"110111111",
  16368=>"100110010",
  16369=>"101100100",
  16370=>"110001100",
  16371=>"010101110",
  16372=>"010100001",
  16373=>"100101100",
  16374=>"010001110",
  16375=>"011000011",
  16376=>"111000110",
  16377=>"000110101",
  16378=>"110010001",
  16379=>"010010011",
  16380=>"000011100",
  16381=>"101010000",
  16382=>"001010010",
  16383=>"000001110",
  16384=>"000000110",
  16385=>"010100000",
  16386=>"100010111",
  16387=>"000010010",
  16388=>"011101000",
  16389=>"101101111",
  16390=>"000111001",
  16391=>"101110100",
  16392=>"110101100",
  16393=>"100100100",
  16394=>"100001010",
  16395=>"010101000",
  16396=>"001101111",
  16397=>"001000110",
  16398=>"010001010",
  16399=>"000100010",
  16400=>"111111101",
  16401=>"011000011",
  16402=>"011001010",
  16403=>"100001010",
  16404=>"110010101",
  16405=>"000110110",
  16406=>"100100100",
  16407=>"011100000",
  16408=>"000011010",
  16409=>"001110100",
  16410=>"101000101",
  16411=>"101100101",
  16412=>"010000000",
  16413=>"001101001",
  16414=>"011110100",
  16415=>"100011101",
  16416=>"000011001",
  16417=>"101111111",
  16418=>"000010000",
  16419=>"010001000",
  16420=>"011101100",
  16421=>"111000011",
  16422=>"100100000",
  16423=>"111010011",
  16424=>"111001001",
  16425=>"001001001",
  16426=>"000111101",
  16427=>"100000000",
  16428=>"100100000",
  16429=>"011101010",
  16430=>"000111111",
  16431=>"011011010",
  16432=>"001000100",
  16433=>"001001101",
  16434=>"010000011",
  16435=>"111111001",
  16436=>"000100110",
  16437=>"011110000",
  16438=>"001001100",
  16439=>"000001010",
  16440=>"001000100",
  16441=>"010011001",
  16442=>"010000110",
  16443=>"100101100",
  16444=>"101011101",
  16445=>"011110101",
  16446=>"001110101",
  16447=>"001111010",
  16448=>"011110011",
  16449=>"000010000",
  16450=>"001011000",
  16451=>"010101011",
  16452=>"010001010",
  16453=>"001111010",
  16454=>"111001111",
  16455=>"111000101",
  16456=>"010101110",
  16457=>"010011010",
  16458=>"010001101",
  16459=>"011100001",
  16460=>"111001010",
  16461=>"001000000",
  16462=>"101100011",
  16463=>"101000100",
  16464=>"011010001",
  16465=>"111001111",
  16466=>"010111111",
  16467=>"011100110",
  16468=>"011110010",
  16469=>"100000001",
  16470=>"111100011",
  16471=>"101100001",
  16472=>"101111010",
  16473=>"001101001",
  16474=>"100001100",
  16475=>"100100000",
  16476=>"101001110",
  16477=>"001011101",
  16478=>"010011001",
  16479=>"001001100",
  16480=>"101111111",
  16481=>"111000000",
  16482=>"000001111",
  16483=>"100101100",
  16484=>"111000000",
  16485=>"110110011",
  16486=>"011100001",
  16487=>"101111101",
  16488=>"011100100",
  16489=>"011110111",
  16490=>"110100100",
  16491=>"111010011",
  16492=>"100101101",
  16493=>"011011000",
  16494=>"100001111",
  16495=>"000000000",
  16496=>"111000101",
  16497=>"010011010",
  16498=>"011111001",
  16499=>"110100001",
  16500=>"001001110",
  16501=>"000101000",
  16502=>"001010010",
  16503=>"101001110",
  16504=>"111100110",
  16505=>"011011111",
  16506=>"001111010",
  16507=>"011001011",
  16508=>"111100101",
  16509=>"000100010",
  16510=>"001000000",
  16511=>"110100001",
  16512=>"001001000",
  16513=>"111111100",
  16514=>"101011001",
  16515=>"101010110",
  16516=>"100001101",
  16517=>"110010110",
  16518=>"001010111",
  16519=>"011111011",
  16520=>"011111110",
  16521=>"011010001",
  16522=>"011001100",
  16523=>"001001000",
  16524=>"100101111",
  16525=>"111101001",
  16526=>"010000011",
  16527=>"101000000",
  16528=>"010110000",
  16529=>"110110100",
  16530=>"010000110",
  16531=>"100000011",
  16532=>"100001001",
  16533=>"000111010",
  16534=>"101000110",
  16535=>"110101101",
  16536=>"100100100",
  16537=>"001100101",
  16538=>"111110000",
  16539=>"101111111",
  16540=>"100111001",
  16541=>"101011111",
  16542=>"111001100",
  16543=>"100010001",
  16544=>"100000000",
  16545=>"101000111",
  16546=>"001010101",
  16547=>"001110000",
  16548=>"111101000",
  16549=>"111100010",
  16550=>"000001101",
  16551=>"011000000",
  16552=>"001011001",
  16553=>"111100001",
  16554=>"101011111",
  16555=>"001100100",
  16556=>"111100010",
  16557=>"001010001",
  16558=>"110011001",
  16559=>"101011101",
  16560=>"000101111",
  16561=>"001010000",
  16562=>"001001000",
  16563=>"000101011",
  16564=>"001111010",
  16565=>"000110101",
  16566=>"010100010",
  16567=>"100000011",
  16568=>"101010111",
  16569=>"001111111",
  16570=>"001011100",
  16571=>"100100000",
  16572=>"100001110",
  16573=>"000010100",
  16574=>"110001001",
  16575=>"110100100",
  16576=>"110011000",
  16577=>"101101000",
  16578=>"001000000",
  16579=>"000111110",
  16580=>"100011001",
  16581=>"110110011",
  16582=>"001000001",
  16583=>"100011100",
  16584=>"101011010",
  16585=>"110100101",
  16586=>"101000101",
  16587=>"010000010",
  16588=>"101111001",
  16589=>"110011011",
  16590=>"011011001",
  16591=>"101100100",
  16592=>"111001110",
  16593=>"010011111",
  16594=>"100010101",
  16595=>"000101110",
  16596=>"010101001",
  16597=>"011101100",
  16598=>"001011000",
  16599=>"000110110",
  16600=>"010011000",
  16601=>"111111010",
  16602=>"001010001",
  16603=>"000010001",
  16604=>"100100011",
  16605=>"010110100",
  16606=>"001001110",
  16607=>"110100011",
  16608=>"000101111",
  16609=>"101110101",
  16610=>"011110110",
  16611=>"000100010",
  16612=>"100000110",
  16613=>"110110001",
  16614=>"001101101",
  16615=>"101100000",
  16616=>"010110000",
  16617=>"000100111",
  16618=>"000101101",
  16619=>"101111101",
  16620=>"111110011",
  16621=>"101001101",
  16622=>"000110111",
  16623=>"110000100",
  16624=>"101010100",
  16625=>"111111111",
  16626=>"101000101",
  16627=>"011111100",
  16628=>"111110101",
  16629=>"010110000",
  16630=>"000000001",
  16631=>"111011110",
  16632=>"111111000",
  16633=>"111101110",
  16634=>"110111001",
  16635=>"011010111",
  16636=>"000101010",
  16637=>"111001000",
  16638=>"011110100",
  16639=>"101101100",
  16640=>"100101110",
  16641=>"000101000",
  16642=>"111111000",
  16643=>"000011110",
  16644=>"001101100",
  16645=>"101011100",
  16646=>"011111000",
  16647=>"001111000",
  16648=>"000111001",
  16649=>"111010110",
  16650=>"010101011",
  16651=>"110000010",
  16652=>"110011010",
  16653=>"101111001",
  16654=>"011111111",
  16655=>"000001110",
  16656=>"010111011",
  16657=>"110111011",
  16658=>"011111011",
  16659=>"000000111",
  16660=>"010111111",
  16661=>"101100001",
  16662=>"001011101",
  16663=>"111000010",
  16664=>"110011010",
  16665=>"110001011",
  16666=>"101100011",
  16667=>"011111000",
  16668=>"101110001",
  16669=>"000101010",
  16670=>"001110000",
  16671=>"100001011",
  16672=>"010010011",
  16673=>"101101100",
  16674=>"100101010",
  16675=>"011000000",
  16676=>"010000001",
  16677=>"011110011",
  16678=>"000000100",
  16679=>"010001001",
  16680=>"111001111",
  16681=>"010111110",
  16682=>"011100100",
  16683=>"110000110",
  16684=>"011011000",
  16685=>"001010111",
  16686=>"011010101",
  16687=>"001110010",
  16688=>"000001011",
  16689=>"111011111",
  16690=>"011101011",
  16691=>"101100101",
  16692=>"110101100",
  16693=>"101100110",
  16694=>"101011010",
  16695=>"000101111",
  16696=>"101001001",
  16697=>"110000110",
  16698=>"111110000",
  16699=>"000000000",
  16700=>"100101000",
  16701=>"101101001",
  16702=>"100101111",
  16703=>"101001110",
  16704=>"010000010",
  16705=>"001100101",
  16706=>"001011000",
  16707=>"011011111",
  16708=>"111111000",
  16709=>"111101111",
  16710=>"011110010",
  16711=>"101100010",
  16712=>"100010100",
  16713=>"110001000",
  16714=>"110011101",
  16715=>"000101110",
  16716=>"010100110",
  16717=>"101001000",
  16718=>"101111100",
  16719=>"100001100",
  16720=>"101100101",
  16721=>"011101000",
  16722=>"101111110",
  16723=>"010001000",
  16724=>"010101000",
  16725=>"011010100",
  16726=>"111111101",
  16727=>"100110010",
  16728=>"000100010",
  16729=>"110000110",
  16730=>"110011110",
  16731=>"011010101",
  16732=>"111110011",
  16733=>"000001111",
  16734=>"000001011",
  16735=>"000000100",
  16736=>"000101010",
  16737=>"011110100",
  16738=>"111101100",
  16739=>"000001011",
  16740=>"001101000",
  16741=>"011100010",
  16742=>"000010010",
  16743=>"100100011",
  16744=>"101011110",
  16745=>"111001101",
  16746=>"111011000",
  16747=>"100111011",
  16748=>"101100001",
  16749=>"011011110",
  16750=>"011010001",
  16751=>"100010100",
  16752=>"001100111",
  16753=>"010100001",
  16754=>"111000111",
  16755=>"010010011",
  16756=>"000110010",
  16757=>"001010000",
  16758=>"011010111",
  16759=>"000011010",
  16760=>"010100000",
  16761=>"101110110",
  16762=>"100101100",
  16763=>"010000000",
  16764=>"101100000",
  16765=>"011110100",
  16766=>"010000001",
  16767=>"101100010",
  16768=>"010100110",
  16769=>"111001011",
  16770=>"000010100",
  16771=>"111110111",
  16772=>"010101010",
  16773=>"111101000",
  16774=>"001110010",
  16775=>"110010100",
  16776=>"101101111",
  16777=>"011101111",
  16778=>"110000001",
  16779=>"110001111",
  16780=>"101010110",
  16781=>"110011110",
  16782=>"101110010",
  16783=>"011110111",
  16784=>"111000011",
  16785=>"001001000",
  16786=>"000000001",
  16787=>"011010001",
  16788=>"000001101",
  16789=>"111000111",
  16790=>"101111010",
  16791=>"110010010",
  16792=>"101001010",
  16793=>"101101010",
  16794=>"111000100",
  16795=>"110001010",
  16796=>"001000000",
  16797=>"100011100",
  16798=>"011100111",
  16799=>"110111100",
  16800=>"100010001",
  16801=>"111000000",
  16802=>"001000110",
  16803=>"100000000",
  16804=>"110110100",
  16805=>"001010000",
  16806=>"111111111",
  16807=>"100010001",
  16808=>"011011001",
  16809=>"001011000",
  16810=>"010110010",
  16811=>"011101101",
  16812=>"111111101",
  16813=>"011111110",
  16814=>"010110111",
  16815=>"001110010",
  16816=>"000100010",
  16817=>"011101101",
  16818=>"100010000",
  16819=>"101111010",
  16820=>"001001010",
  16821=>"110011010",
  16822=>"110101001",
  16823=>"000010011",
  16824=>"011010011",
  16825=>"110111000",
  16826=>"010001111",
  16827=>"111111000",
  16828=>"110100001",
  16829=>"110010010",
  16830=>"101101011",
  16831=>"001000110",
  16832=>"010010101",
  16833=>"101110101",
  16834=>"011111101",
  16835=>"111001111",
  16836=>"110011111",
  16837=>"101000100",
  16838=>"100111011",
  16839=>"111011101",
  16840=>"010011100",
  16841=>"111111011",
  16842=>"110101010",
  16843=>"100011111",
  16844=>"110100000",
  16845=>"001110011",
  16846=>"101000000",
  16847=>"100010110",
  16848=>"111111101",
  16849=>"100100100",
  16850=>"100111011",
  16851=>"010111110",
  16852=>"000001101",
  16853=>"010010111",
  16854=>"111010100",
  16855=>"001010100",
  16856=>"000100011",
  16857=>"111001100",
  16858=>"011000000",
  16859=>"000001100",
  16860=>"010001101",
  16861=>"000111111",
  16862=>"110100010",
  16863=>"110011111",
  16864=>"110011000",
  16865=>"011011110",
  16866=>"001010111",
  16867=>"000011011",
  16868=>"000100101",
  16869=>"010011000",
  16870=>"110011100",
  16871=>"111001011",
  16872=>"000111001",
  16873=>"100000100",
  16874=>"010100000",
  16875=>"110111111",
  16876=>"010011101",
  16877=>"010010100",
  16878=>"111010100",
  16879=>"100001011",
  16880=>"011110000",
  16881=>"011010000",
  16882=>"101101100",
  16883=>"111011111",
  16884=>"001001110",
  16885=>"001110011",
  16886=>"101100101",
  16887=>"000101110",
  16888=>"100010100",
  16889=>"001001011",
  16890=>"000011010",
  16891=>"001110011",
  16892=>"010001011",
  16893=>"010011011",
  16894=>"000011101",
  16895=>"011011011",
  16896=>"010101001",
  16897=>"011110101",
  16898=>"100001001",
  16899=>"110110010",
  16900=>"010100100",
  16901=>"010100001",
  16902=>"010101001",
  16903=>"001001101",
  16904=>"001101100",
  16905=>"001011000",
  16906=>"000011101",
  16907=>"010000010",
  16908=>"010101100",
  16909=>"011111101",
  16910=>"111000000",
  16911=>"101100000",
  16912=>"111111110",
  16913=>"110010110",
  16914=>"001011111",
  16915=>"010100001",
  16916=>"111000101",
  16917=>"101000111",
  16918=>"000001100",
  16919=>"110010110",
  16920=>"101101000",
  16921=>"001010000",
  16922=>"001010001",
  16923=>"100111100",
  16924=>"111000100",
  16925=>"010101001",
  16926=>"111000101",
  16927=>"010010011",
  16928=>"010010100",
  16929=>"010011000",
  16930=>"010100001",
  16931=>"111010000",
  16932=>"010000100",
  16933=>"100101101",
  16934=>"111100000",
  16935=>"101101110",
  16936=>"100000011",
  16937=>"010111101",
  16938=>"101101010",
  16939=>"010010010",
  16940=>"100100101",
  16941=>"001101000",
  16942=>"000110011",
  16943=>"001110000",
  16944=>"010111110",
  16945=>"001010011",
  16946=>"001001101",
  16947=>"110101111",
  16948=>"101011100",
  16949=>"010000111",
  16950=>"000011011",
  16951=>"011010010",
  16952=>"110111110",
  16953=>"111100010",
  16954=>"011001100",
  16955=>"011000110",
  16956=>"011010011",
  16957=>"100100100",
  16958=>"000010000",
  16959=>"111101111",
  16960=>"111001001",
  16961=>"110100001",
  16962=>"010001001",
  16963=>"100000010",
  16964=>"101111111",
  16965=>"010000011",
  16966=>"100100011",
  16967=>"010011000",
  16968=>"101001000",
  16969=>"101000001",
  16970=>"100000100",
  16971=>"011101000",
  16972=>"001110001",
  16973=>"001111000",
  16974=>"110101110",
  16975=>"001110100",
  16976=>"100001001",
  16977=>"001001101",
  16978=>"011101000",
  16979=>"100000011",
  16980=>"010000101",
  16981=>"000111001",
  16982=>"100000101",
  16983=>"010000000",
  16984=>"001011111",
  16985=>"010111011",
  16986=>"000110011",
  16987=>"011100000",
  16988=>"001101010",
  16989=>"111101000",
  16990=>"000010101",
  16991=>"001011101",
  16992=>"011011101",
  16993=>"111000001",
  16994=>"001100101",
  16995=>"010000111",
  16996=>"000011111",
  16997=>"001111101",
  16998=>"011001111",
  16999=>"100111110",
  17000=>"010110111",
  17001=>"010010100",
  17002=>"111110101",
  17003=>"101000100",
  17004=>"101101000",
  17005=>"000100111",
  17006=>"110110101",
  17007=>"111011010",
  17008=>"011000111",
  17009=>"100100000",
  17010=>"011000110",
  17011=>"110001000",
  17012=>"101000110",
  17013=>"101010100",
  17014=>"111111110",
  17015=>"111101011",
  17016=>"111001100",
  17017=>"100111101",
  17018=>"101010110",
  17019=>"111010011",
  17020=>"011100001",
  17021=>"000010110",
  17022=>"011001011",
  17023=>"110011011",
  17024=>"001001101",
  17025=>"001111111",
  17026=>"000111111",
  17027=>"110000110",
  17028=>"111110101",
  17029=>"010111000",
  17030=>"111111111",
  17031=>"111011001",
  17032=>"000101000",
  17033=>"100100110",
  17034=>"001111100",
  17035=>"101000001",
  17036=>"101011111",
  17037=>"111011111",
  17038=>"101010001",
  17039=>"001100001",
  17040=>"011010111",
  17041=>"111111111",
  17042=>"111101000",
  17043=>"010010101",
  17044=>"001001000",
  17045=>"000100010",
  17046=>"011010100",
  17047=>"100100001",
  17048=>"010110100",
  17049=>"011111000",
  17050=>"011001100",
  17051=>"001100100",
  17052=>"111100000",
  17053=>"110000010",
  17054=>"000110001",
  17055=>"100011100",
  17056=>"001101011",
  17057=>"001110001",
  17058=>"010011010",
  17059=>"011100010",
  17060=>"111101010",
  17061=>"111110110",
  17062=>"100000110",
  17063=>"101000100",
  17064=>"010101011",
  17065=>"111111110",
  17066=>"110011011",
  17067=>"110001011",
  17068=>"000111110",
  17069=>"110110011",
  17070=>"111110100",
  17071=>"010110000",
  17072=>"011100001",
  17073=>"001111101",
  17074=>"001000111",
  17075=>"000001010",
  17076=>"011011111",
  17077=>"010010000",
  17078=>"010010010",
  17079=>"010100010",
  17080=>"011100000",
  17081=>"000111101",
  17082=>"000110111",
  17083=>"110101111",
  17084=>"010001000",
  17085=>"001100010",
  17086=>"001011111",
  17087=>"011010100",
  17088=>"011100111",
  17089=>"110000110",
  17090=>"011100010",
  17091=>"111010011",
  17092=>"000100101",
  17093=>"000010111",
  17094=>"010010110",
  17095=>"010101001",
  17096=>"010010011",
  17097=>"011111000",
  17098=>"110111011",
  17099=>"111101100",
  17100=>"000000100",
  17101=>"100111101",
  17102=>"100011001",
  17103=>"000011000",
  17104=>"010000101",
  17105=>"111101111",
  17106=>"100101000",
  17107=>"001011001",
  17108=>"000011100",
  17109=>"000001110",
  17110=>"000100000",
  17111=>"000010000",
  17112=>"011111110",
  17113=>"010010100",
  17114=>"001010001",
  17115=>"111111000",
  17116=>"000011101",
  17117=>"111110111",
  17118=>"000011001",
  17119=>"010100011",
  17120=>"101010010",
  17121=>"001010001",
  17122=>"100110100",
  17123=>"101001011",
  17124=>"100011010",
  17125=>"001101111",
  17126=>"000100011",
  17127=>"001000001",
  17128=>"000101000",
  17129=>"011100110",
  17130=>"000010010",
  17131=>"000010100",
  17132=>"001100000",
  17133=>"101000011",
  17134=>"100000010",
  17135=>"100101001",
  17136=>"000110101",
  17137=>"100111100",
  17138=>"001000110",
  17139=>"011000000",
  17140=>"000011101",
  17141=>"011110100",
  17142=>"111011110",
  17143=>"101011011",
  17144=>"011011101",
  17145=>"101101101",
  17146=>"100111110",
  17147=>"000111111",
  17148=>"111011110",
  17149=>"000111011",
  17150=>"100111000",
  17151=>"100011010",
  17152=>"011011111",
  17153=>"011101000",
  17154=>"001110101",
  17155=>"000101011",
  17156=>"011101000",
  17157=>"100010000",
  17158=>"000111001",
  17159=>"011100010",
  17160=>"000101101",
  17161=>"011011101",
  17162=>"001111111",
  17163=>"101001101",
  17164=>"110011100",
  17165=>"111010011",
  17166=>"100001100",
  17167=>"010011011",
  17168=>"001100000",
  17169=>"000111001",
  17170=>"000011010",
  17171=>"101011000",
  17172=>"000111110",
  17173=>"011011010",
  17174=>"100010100",
  17175=>"100101100",
  17176=>"011101001",
  17177=>"001000100",
  17178=>"101011111",
  17179=>"011101011",
  17180=>"100000110",
  17181=>"100000110",
  17182=>"101000110",
  17183=>"100011000",
  17184=>"001010110",
  17185=>"110000101",
  17186=>"001010001",
  17187=>"000011001",
  17188=>"010010111",
  17189=>"011110100",
  17190=>"100110010",
  17191=>"110001110",
  17192=>"000101100",
  17193=>"100111100",
  17194=>"010000000",
  17195=>"010111101",
  17196=>"011111111",
  17197=>"000100010",
  17198=>"000100100",
  17199=>"101001010",
  17200=>"111110011",
  17201=>"011000011",
  17202=>"010000100",
  17203=>"100001111",
  17204=>"001011011",
  17205=>"110001011",
  17206=>"000101101",
  17207=>"110100011",
  17208=>"111001001",
  17209=>"111011001",
  17210=>"001101010",
  17211=>"111110100",
  17212=>"111110101",
  17213=>"101010010",
  17214=>"010001110",
  17215=>"011101001",
  17216=>"011010001",
  17217=>"000010000",
  17218=>"010010000",
  17219=>"111011010",
  17220=>"111000101",
  17221=>"101101111",
  17222=>"001101011",
  17223=>"110100000",
  17224=>"011001010",
  17225=>"110110110",
  17226=>"010101100",
  17227=>"111000100",
  17228=>"101101011",
  17229=>"110101110",
  17230=>"111001100",
  17231=>"110101100",
  17232=>"110111111",
  17233=>"111100001",
  17234=>"001000111",
  17235=>"110000000",
  17236=>"010011100",
  17237=>"101001111",
  17238=>"101111100",
  17239=>"111101000",
  17240=>"110001000",
  17241=>"111010011",
  17242=>"011111010",
  17243=>"100111010",
  17244=>"011001001",
  17245=>"000011001",
  17246=>"101001000",
  17247=>"000001000",
  17248=>"000111111",
  17249=>"111010111",
  17250=>"000100000",
  17251=>"010011000",
  17252=>"001111101",
  17253=>"110010000",
  17254=>"001110011",
  17255=>"000100000",
  17256=>"110111111",
  17257=>"100110011",
  17258=>"011111100",
  17259=>"001010101",
  17260=>"101001111",
  17261=>"111110010",
  17262=>"011010101",
  17263=>"110100100",
  17264=>"111000000",
  17265=>"111110110",
  17266=>"010110111",
  17267=>"101001111",
  17268=>"011001100",
  17269=>"000001100",
  17270=>"001001000",
  17271=>"100000001",
  17272=>"101101110",
  17273=>"111110111",
  17274=>"110110010",
  17275=>"111101000",
  17276=>"100011001",
  17277=>"101011010",
  17278=>"010101110",
  17279=>"110010000",
  17280=>"001010111",
  17281=>"000100100",
  17282=>"010100001",
  17283=>"111000100",
  17284=>"101101000",
  17285=>"011100001",
  17286=>"000000101",
  17287=>"001001010",
  17288=>"101010100",
  17289=>"000010010",
  17290=>"111010000",
  17291=>"100100011",
  17292=>"001111011",
  17293=>"111000000",
  17294=>"000100110",
  17295=>"111100111",
  17296=>"100110010",
  17297=>"000001111",
  17298=>"101000000",
  17299=>"100100010",
  17300=>"010000111",
  17301=>"110011001",
  17302=>"111110101",
  17303=>"000110000",
  17304=>"111001110",
  17305=>"011101110",
  17306=>"010111000",
  17307=>"010000000",
  17308=>"101000100",
  17309=>"101100000",
  17310=>"101011001",
  17311=>"100100100",
  17312=>"001111010",
  17313=>"111110111",
  17314=>"000010010",
  17315=>"101001111",
  17316=>"000110011",
  17317=>"010010011",
  17318=>"100000101",
  17319=>"011001111",
  17320=>"110001111",
  17321=>"111101111",
  17322=>"100111110",
  17323=>"111011001",
  17324=>"000100000",
  17325=>"011010001",
  17326=>"011000100",
  17327=>"110100001",
  17328=>"001111010",
  17329=>"110010000",
  17330=>"111111001",
  17331=>"001100111",
  17332=>"100111101",
  17333=>"011001000",
  17334=>"100111101",
  17335=>"101011100",
  17336=>"101001011",
  17337=>"111001101",
  17338=>"010010100",
  17339=>"111101010",
  17340=>"111011110",
  17341=>"000010001",
  17342=>"101101010",
  17343=>"000011001",
  17344=>"101010001",
  17345=>"100100110",
  17346=>"001101101",
  17347=>"110010110",
  17348=>"000111001",
  17349=>"011001000",
  17350=>"011001010",
  17351=>"111111011",
  17352=>"011101000",
  17353=>"000010011",
  17354=>"101010110",
  17355=>"000101110",
  17356=>"111010101",
  17357=>"111111011",
  17358=>"100111111",
  17359=>"111100110",
  17360=>"100100010",
  17361=>"101111010",
  17362=>"110001000",
  17363=>"000000110",
  17364=>"010110111",
  17365=>"111010010",
  17366=>"001110111",
  17367=>"110000010",
  17368=>"100100111",
  17369=>"110111111",
  17370=>"010110000",
  17371=>"010000110",
  17372=>"101110010",
  17373=>"111001010",
  17374=>"011100110",
  17375=>"100001010",
  17376=>"001111101",
  17377=>"111111110",
  17378=>"101000111",
  17379=>"111001011",
  17380=>"110100011",
  17381=>"000001001",
  17382=>"000111111",
  17383=>"011110100",
  17384=>"110100001",
  17385=>"101010111",
  17386=>"000000101",
  17387=>"100010010",
  17388=>"110010111",
  17389=>"011111000",
  17390=>"011001110",
  17391=>"110111000",
  17392=>"000001101",
  17393=>"001110001",
  17394=>"001111100",
  17395=>"100110011",
  17396=>"111000000",
  17397=>"110110000",
  17398=>"101011111",
  17399=>"010010001",
  17400=>"001000110",
  17401=>"000001011",
  17402=>"000110101",
  17403=>"000101011",
  17404=>"101000010",
  17405=>"110011100",
  17406=>"001101010",
  17407=>"100110111",
  17408=>"101001000",
  17409=>"111010111",
  17410=>"111011001",
  17411=>"110111010",
  17412=>"011110100",
  17413=>"101010101",
  17414=>"100101111",
  17415=>"000100000",
  17416=>"100110001",
  17417=>"110000111",
  17418=>"000000011",
  17419=>"100110111",
  17420=>"101101010",
  17421=>"000011001",
  17422=>"111001011",
  17423=>"010011011",
  17424=>"110001001",
  17425=>"111000100",
  17426=>"100000001",
  17427=>"111000110",
  17428=>"100011001",
  17429=>"000110010",
  17430=>"101111111",
  17431=>"001000110",
  17432=>"111111100",
  17433=>"010000000",
  17434=>"101100011",
  17435=>"110111011",
  17436=>"100000010",
  17437=>"100101010",
  17438=>"001011110",
  17439=>"111011100",
  17440=>"110000010",
  17441=>"011110010",
  17442=>"111001100",
  17443=>"101100100",
  17444=>"011101110",
  17445=>"111101111",
  17446=>"000110111",
  17447=>"010100000",
  17448=>"011110011",
  17449=>"110100110",
  17450=>"010010000",
  17451=>"111100010",
  17452=>"100110111",
  17453=>"000111101",
  17454=>"100001110",
  17455=>"000010111",
  17456=>"100101011",
  17457=>"011110011",
  17458=>"000000010",
  17459=>"001001100",
  17460=>"100001000",
  17461=>"100001010",
  17462=>"110011101",
  17463=>"111111100",
  17464=>"001001000",
  17465=>"000100100",
  17466=>"110010000",
  17467=>"000011111",
  17468=>"011000010",
  17469=>"011001110",
  17470=>"011011000",
  17471=>"111111111",
  17472=>"111000000",
  17473=>"000000111",
  17474=>"001001010",
  17475=>"101101000",
  17476=>"111001100",
  17477=>"111101111",
  17478=>"011001110",
  17479=>"100110000",
  17480=>"011100010",
  17481=>"110000000",
  17482=>"001010110",
  17483=>"100011110",
  17484=>"001111101",
  17485=>"111011011",
  17486=>"111101100",
  17487=>"100101101",
  17488=>"100011000",
  17489=>"011000101",
  17490=>"100010010",
  17491=>"010001000",
  17492=>"111110101",
  17493=>"010110010",
  17494=>"000001111",
  17495=>"000001101",
  17496=>"001101100",
  17497=>"000011100",
  17498=>"001111110",
  17499=>"100000000",
  17500=>"000100000",
  17501=>"101111001",
  17502=>"101000111",
  17503=>"010010111",
  17504=>"001000001",
  17505=>"100001101",
  17506=>"011100000",
  17507=>"001010000",
  17508=>"010000110",
  17509=>"010010010",
  17510=>"001011001",
  17511=>"000101010",
  17512=>"000111111",
  17513=>"011000110",
  17514=>"100010101",
  17515=>"110110100",
  17516=>"101101100",
  17517=>"100010001",
  17518=>"010101100",
  17519=>"001000001",
  17520=>"010010000",
  17521=>"111001110",
  17522=>"010111001",
  17523=>"100111101",
  17524=>"010110111",
  17525=>"000000010",
  17526=>"010011000",
  17527=>"010101010",
  17528=>"100001000",
  17529=>"000001010",
  17530=>"010000000",
  17531=>"000101011",
  17532=>"101101101",
  17533=>"001001111",
  17534=>"101010001",
  17535=>"010001101",
  17536=>"010000101",
  17537=>"000011110",
  17538=>"000001110",
  17539=>"010001001",
  17540=>"001001101",
  17541=>"000110111",
  17542=>"000010010",
  17543=>"011011111",
  17544=>"100111000",
  17545=>"110001110",
  17546=>"111001100",
  17547=>"110111110",
  17548=>"101011001",
  17549=>"100110101",
  17550=>"100111100",
  17551=>"100110111",
  17552=>"100010110",
  17553=>"110101110",
  17554=>"010000010",
  17555=>"111000110",
  17556=>"110111001",
  17557=>"111110000",
  17558=>"110101101",
  17559=>"011001010",
  17560=>"110110001",
  17561=>"010101101",
  17562=>"001001001",
  17563=>"101101010",
  17564=>"001000001",
  17565=>"101010000",
  17566=>"011000000",
  17567=>"100101100",
  17568=>"110001011",
  17569=>"001101001",
  17570=>"111001100",
  17571=>"010001110",
  17572=>"111001010",
  17573=>"111100001",
  17574=>"111001000",
  17575=>"001000001",
  17576=>"011000000",
  17577=>"111010010",
  17578=>"101111111",
  17579=>"100001010",
  17580=>"001110111",
  17581=>"000100101",
  17582=>"111001011",
  17583=>"001011110",
  17584=>"000110001",
  17585=>"000000001",
  17586=>"111111011",
  17587=>"010011110",
  17588=>"011100010",
  17589=>"010110111",
  17590=>"111000110",
  17591=>"100111100",
  17592=>"000000101",
  17593=>"110100110",
  17594=>"000110110",
  17595=>"111111101",
  17596=>"111111001",
  17597=>"111101011",
  17598=>"111100110",
  17599=>"010011010",
  17600=>"111101101",
  17601=>"000011111",
  17602=>"000010000",
  17603=>"011001111",
  17604=>"000010010",
  17605=>"000101111",
  17606=>"011011001",
  17607=>"101100101",
  17608=>"011111111",
  17609=>"010110011",
  17610=>"101101100",
  17611=>"110101101",
  17612=>"001000001",
  17613=>"101011010",
  17614=>"000110110",
  17615=>"001011010",
  17616=>"000011101",
  17617=>"101101101",
  17618=>"011101010",
  17619=>"001110111",
  17620=>"011000001",
  17621=>"101101010",
  17622=>"100100101",
  17623=>"011000011",
  17624=>"000000001",
  17625=>"011001110",
  17626=>"101110101",
  17627=>"100011000",
  17628=>"101110010",
  17629=>"001001101",
  17630=>"011000001",
  17631=>"010111000",
  17632=>"000011010",
  17633=>"011111000",
  17634=>"111110111",
  17635=>"011010101",
  17636=>"101100110",
  17637=>"000110000",
  17638=>"000100110",
  17639=>"010101001",
  17640=>"010100011",
  17641=>"010000101",
  17642=>"101001011",
  17643=>"101001011",
  17644=>"010000001",
  17645=>"111011011",
  17646=>"101000110",
  17647=>"010011110",
  17648=>"010100110",
  17649=>"010010000",
  17650=>"010101101",
  17651=>"111110000",
  17652=>"111111110",
  17653=>"001001101",
  17654=>"001011110",
  17655=>"000000110",
  17656=>"110010001",
  17657=>"111100000",
  17658=>"001100001",
  17659=>"000000001",
  17660=>"101001011",
  17661=>"000100111",
  17662=>"101010110",
  17663=>"101000011",
  17664=>"100110111",
  17665=>"100110010",
  17666=>"111100011",
  17667=>"100010010",
  17668=>"101001010",
  17669=>"100101111",
  17670=>"011110110",
  17671=>"100110011",
  17672=>"000111011",
  17673=>"110010001",
  17674=>"111010100",
  17675=>"101000100",
  17676=>"001010100",
  17677=>"100100101",
  17678=>"111100110",
  17679=>"010000010",
  17680=>"100001111",
  17681=>"111111010",
  17682=>"110110101",
  17683=>"000001101",
  17684=>"111000000",
  17685=>"111000010",
  17686=>"010100101",
  17687=>"000010100",
  17688=>"011000001",
  17689=>"111111101",
  17690=>"101110100",
  17691=>"110001010",
  17692=>"001010110",
  17693=>"111001101",
  17694=>"001001010",
  17695=>"011101100",
  17696=>"000011100",
  17697=>"101100000",
  17698=>"011011111",
  17699=>"110101111",
  17700=>"101100111",
  17701=>"100101100",
  17702=>"000000110",
  17703=>"000001001",
  17704=>"011001001",
  17705=>"100010110",
  17706=>"100111110",
  17707=>"000000100",
  17708=>"111000110",
  17709=>"100001010",
  17710=>"000010001",
  17711=>"111110111",
  17712=>"001001100",
  17713=>"111011100",
  17714=>"000110010",
  17715=>"110110000",
  17716=>"001000010",
  17717=>"111111011",
  17718=>"001111100",
  17719=>"001111010",
  17720=>"000011010",
  17721=>"010000111",
  17722=>"010000101",
  17723=>"111011000",
  17724=>"000110110",
  17725=>"100110110",
  17726=>"110100101",
  17727=>"110001001",
  17728=>"110111111",
  17729=>"111001111",
  17730=>"000000000",
  17731=>"000110000",
  17732=>"101101011",
  17733=>"100111111",
  17734=>"010001101",
  17735=>"000011011",
  17736=>"110011100",
  17737=>"001101111",
  17738=>"111010000",
  17739=>"101000100",
  17740=>"111111110",
  17741=>"010011001",
  17742=>"001100010",
  17743=>"111001100",
  17744=>"110101100",
  17745=>"101011000",
  17746=>"111101010",
  17747=>"100010000",
  17748=>"101000010",
  17749=>"111000111",
  17750=>"101110101",
  17751=>"110011100",
  17752=>"101101001",
  17753=>"000111101",
  17754=>"101010001",
  17755=>"110010100",
  17756=>"010100010",
  17757=>"110100110",
  17758=>"011010011",
  17759=>"010000100",
  17760=>"000011010",
  17761=>"101011111",
  17762=>"011100011",
  17763=>"000010100",
  17764=>"010000000",
  17765=>"011010111",
  17766=>"001010000",
  17767=>"110100111",
  17768=>"000111101",
  17769=>"010001100",
  17770=>"000010110",
  17771=>"110101101",
  17772=>"110000101",
  17773=>"101100100",
  17774=>"101010111",
  17775=>"010111101",
  17776=>"000010000",
  17777=>"001000000",
  17778=>"101111111",
  17779=>"101101110",
  17780=>"101110100",
  17781=>"111010101",
  17782=>"100010101",
  17783=>"001111110",
  17784=>"100111110",
  17785=>"111001100",
  17786=>"000010100",
  17787=>"001111110",
  17788=>"100011101",
  17789=>"100111110",
  17790=>"000100110",
  17791=>"010111110",
  17792=>"001000101",
  17793=>"000000001",
  17794=>"111011111",
  17795=>"001100010",
  17796=>"000010011",
  17797=>"101111100",
  17798=>"111000111",
  17799=>"100011000",
  17800=>"110010010",
  17801=>"101010111",
  17802=>"000100001",
  17803=>"010110100",
  17804=>"101011011",
  17805=>"111000100",
  17806=>"000011001",
  17807=>"101110100",
  17808=>"010101010",
  17809=>"000001111",
  17810=>"100000000",
  17811=>"000011001",
  17812=>"011010111",
  17813=>"000000111",
  17814=>"001010111",
  17815=>"010010100",
  17816=>"111000110",
  17817=>"011000110",
  17818=>"001111110",
  17819=>"001101111",
  17820=>"110010001",
  17821=>"100101101",
  17822=>"010101101",
  17823=>"011100000",
  17824=>"100000110",
  17825=>"101001101",
  17826=>"110011010",
  17827=>"000001101",
  17828=>"011110000",
  17829=>"001100000",
  17830=>"101001101",
  17831=>"111101010",
  17832=>"111001110",
  17833=>"000101010",
  17834=>"000100100",
  17835=>"010101100",
  17836=>"111111001",
  17837=>"011000001",
  17838=>"110111110",
  17839=>"001110001",
  17840=>"010100110",
  17841=>"010101001",
  17842=>"101010100",
  17843=>"001001101",
  17844=>"111010110",
  17845=>"111110010",
  17846=>"111101110",
  17847=>"010110110",
  17848=>"100110000",
  17849=>"110101011",
  17850=>"001000000",
  17851=>"000111111",
  17852=>"101011001",
  17853=>"111100001",
  17854=>"100001010",
  17855=>"111011011",
  17856=>"110110010",
  17857=>"101000011",
  17858=>"110100111",
  17859=>"110000110",
  17860=>"100011100",
  17861=>"111000101",
  17862=>"110010000",
  17863=>"011011011",
  17864=>"100101010",
  17865=>"100100110",
  17866=>"110010110",
  17867=>"111110101",
  17868=>"010111001",
  17869=>"110010100",
  17870=>"101100111",
  17871=>"000110001",
  17872=>"111101011",
  17873=>"001100000",
  17874=>"011100011",
  17875=>"001001011",
  17876=>"101011001",
  17877=>"011011011",
  17878=>"111101101",
  17879=>"001001110",
  17880=>"010010001",
  17881=>"101110001",
  17882=>"011010111",
  17883=>"000111000",
  17884=>"001000111",
  17885=>"101000001",
  17886=>"101010010",
  17887=>"110100001",
  17888=>"000100011",
  17889=>"000011110",
  17890=>"000100110",
  17891=>"000111100",
  17892=>"000110011",
  17893=>"111000010",
  17894=>"000010101",
  17895=>"000100011",
  17896=>"011011011",
  17897=>"000111111",
  17898=>"000000100",
  17899=>"101110001",
  17900=>"010100111",
  17901=>"101000001",
  17902=>"000101000",
  17903=>"011111001",
  17904=>"000011111",
  17905=>"010000010",
  17906=>"101000101",
  17907=>"100010111",
  17908=>"111010111",
  17909=>"001100000",
  17910=>"100011100",
  17911=>"110111000",
  17912=>"110011111",
  17913=>"111101110",
  17914=>"100100110",
  17915=>"110100011",
  17916=>"010100110",
  17917=>"010100101",
  17918=>"011111100",
  17919=>"001010110",
  17920=>"101110111",
  17921=>"001011100",
  17922=>"101101001",
  17923=>"111000101",
  17924=>"000111000",
  17925=>"010001100",
  17926=>"110100011",
  17927=>"110000110",
  17928=>"000100011",
  17929=>"001001110",
  17930=>"100111111",
  17931=>"011110100",
  17932=>"010111101",
  17933=>"010011000",
  17934=>"001000100",
  17935=>"001001011",
  17936=>"101110111",
  17937=>"000100111",
  17938=>"100000110",
  17939=>"100101110",
  17940=>"110100111",
  17941=>"001000001",
  17942=>"110000000",
  17943=>"011110001",
  17944=>"100100001",
  17945=>"001111111",
  17946=>"001001101",
  17947=>"000110010",
  17948=>"110101011",
  17949=>"011100001",
  17950=>"101110010",
  17951=>"001111111",
  17952=>"101000010",
  17953=>"011100100",
  17954=>"001011001",
  17955=>"101010101",
  17956=>"000011000",
  17957=>"100111110",
  17958=>"001011001",
  17959=>"100000110",
  17960=>"000011100",
  17961=>"100000100",
  17962=>"110011001",
  17963=>"111101010",
  17964=>"011000001",
  17965=>"010100011",
  17966=>"010110100",
  17967=>"010111101",
  17968=>"110001110",
  17969=>"100001101",
  17970=>"110101011",
  17971=>"101101110",
  17972=>"101010000",
  17973=>"011101001",
  17974=>"101110001",
  17975=>"000001000",
  17976=>"000110100",
  17977=>"110000110",
  17978=>"010111111",
  17979=>"000101000",
  17980=>"011000110",
  17981=>"100100001",
  17982=>"001011100",
  17983=>"001110011",
  17984=>"000101100",
  17985=>"101111101",
  17986=>"000100011",
  17987=>"011100011",
  17988=>"100001101",
  17989=>"100010011",
  17990=>"100100100",
  17991=>"100001000",
  17992=>"001001111",
  17993=>"001101010",
  17994=>"010111111",
  17995=>"100110101",
  17996=>"110100010",
  17997=>"010001110",
  17998=>"110100110",
  17999=>"110000010",
  18000=>"000100000",
  18001=>"000101111",
  18002=>"111100011",
  18003=>"011100000",
  18004=>"001000110",
  18005=>"011001111",
  18006=>"010000000",
  18007=>"000011101",
  18008=>"111010000",
  18009=>"110000011",
  18010=>"011010101",
  18011=>"101001101",
  18012=>"100010010",
  18013=>"001011001",
  18014=>"001011011",
  18015=>"110000100",
  18016=>"111000010",
  18017=>"110100000",
  18018=>"000100000",
  18019=>"010111111",
  18020=>"001001101",
  18021=>"011111011",
  18022=>"011000101",
  18023=>"011111101",
  18024=>"010111100",
  18025=>"010110001",
  18026=>"111001101",
  18027=>"010001101",
  18028=>"000010001",
  18029=>"010000010",
  18030=>"001001011",
  18031=>"101010001",
  18032=>"000011100",
  18033=>"101010110",
  18034=>"010011001",
  18035=>"001000010",
  18036=>"000111000",
  18037=>"111000001",
  18038=>"001000111",
  18039=>"010010000",
  18040=>"000011110",
  18041=>"000101110",
  18042=>"101010010",
  18043=>"010010011",
  18044=>"001001100",
  18045=>"001101010",
  18046=>"100000000",
  18047=>"011000111",
  18048=>"100110100",
  18049=>"110101001",
  18050=>"010100000",
  18051=>"111001001",
  18052=>"101010110",
  18053=>"101100011",
  18054=>"001110111",
  18055=>"100010110",
  18056=>"001100110",
  18057=>"010100011",
  18058=>"111101101",
  18059=>"111111001",
  18060=>"001001000",
  18061=>"100100000",
  18062=>"001000001",
  18063=>"100110001",
  18064=>"111010101",
  18065=>"111101101",
  18066=>"011001110",
  18067=>"111110111",
  18068=>"101001011",
  18069=>"011111011",
  18070=>"000100011",
  18071=>"001110101",
  18072=>"100000001",
  18073=>"101111001",
  18074=>"001010000",
  18075=>"100101100",
  18076=>"100101000",
  18077=>"001011110",
  18078=>"011000010",
  18079=>"011010101",
  18080=>"110000100",
  18081=>"001101100",
  18082=>"111001010",
  18083=>"011000000",
  18084=>"111101100",
  18085=>"111110101",
  18086=>"000011011",
  18087=>"001001100",
  18088=>"101111011",
  18089=>"000001000",
  18090=>"100111110",
  18091=>"110100000",
  18092=>"100001100",
  18093=>"011110000",
  18094=>"000011100",
  18095=>"110011110",
  18096=>"110000000",
  18097=>"000011001",
  18098=>"011011010",
  18099=>"011000011",
  18100=>"010101001",
  18101=>"010101101",
  18102=>"101000010",
  18103=>"010100000",
  18104=>"101111101",
  18105=>"100110011",
  18106=>"111011111",
  18107=>"011111110",
  18108=>"001001111",
  18109=>"001110100",
  18110=>"000001001",
  18111=>"110101110",
  18112=>"100000100",
  18113=>"011001001",
  18114=>"100010110",
  18115=>"100010011",
  18116=>"111011001",
  18117=>"010100010",
  18118=>"110000000",
  18119=>"000001001",
  18120=>"100100000",
  18121=>"000111010",
  18122=>"011000111",
  18123=>"111000100",
  18124=>"101011111",
  18125=>"111101011",
  18126=>"000011000",
  18127=>"010101010",
  18128=>"000011000",
  18129=>"010000100",
  18130=>"000101000",
  18131=>"111010010",
  18132=>"101000100",
  18133=>"110101010",
  18134=>"110111101",
  18135=>"000001110",
  18136=>"001001100",
  18137=>"100111010",
  18138=>"011010111",
  18139=>"110010000",
  18140=>"001011011",
  18141=>"000111110",
  18142=>"101100100",
  18143=>"000101010",
  18144=>"110000111",
  18145=>"100001101",
  18146=>"110110001",
  18147=>"000100101",
  18148=>"000111010",
  18149=>"110110110",
  18150=>"010101101",
  18151=>"000100101",
  18152=>"101000110",
  18153=>"111111011",
  18154=>"110101111",
  18155=>"111000010",
  18156=>"110101001",
  18157=>"100101000",
  18158=>"110111101",
  18159=>"101011000",
  18160=>"001110011",
  18161=>"101001010",
  18162=>"010111010",
  18163=>"010100000",
  18164=>"000100100",
  18165=>"010000101",
  18166=>"000100110",
  18167=>"110011011",
  18168=>"010111000",
  18169=>"000111101",
  18170=>"101001101",
  18171=>"000001001",
  18172=>"001111110",
  18173=>"011010110",
  18174=>"111010101",
  18175=>"011110001",
  18176=>"011110011",
  18177=>"011101101",
  18178=>"111011010",
  18179=>"101000100",
  18180=>"100111110",
  18181=>"011100110",
  18182=>"001110001",
  18183=>"111111111",
  18184=>"101100001",
  18185=>"101101111",
  18186=>"101010111",
  18187=>"000000000",
  18188=>"001001010",
  18189=>"010111011",
  18190=>"000011000",
  18191=>"011100110",
  18192=>"000101000",
  18193=>"101111011",
  18194=>"110011111",
  18195=>"100010011",
  18196=>"011000101",
  18197=>"000000010",
  18198=>"001000000",
  18199=>"111111100",
  18200=>"010111110",
  18201=>"101000100",
  18202=>"111110110",
  18203=>"110110101",
  18204=>"111111110",
  18205=>"011001000",
  18206=>"000010001",
  18207=>"001010000",
  18208=>"100111100",
  18209=>"101110011",
  18210=>"000110110",
  18211=>"000000100",
  18212=>"110000000",
  18213=>"001000101",
  18214=>"111100101",
  18215=>"010011010",
  18216=>"100101110",
  18217=>"010101100",
  18218=>"000000000",
  18219=>"010010101",
  18220=>"101110101",
  18221=>"101111011",
  18222=>"010110000",
  18223=>"000011110",
  18224=>"000000101",
  18225=>"001010101",
  18226=>"100111110",
  18227=>"011010111",
  18228=>"001010010",
  18229=>"101100111",
  18230=>"001000000",
  18231=>"000000110",
  18232=>"100111001",
  18233=>"110111000",
  18234=>"101111010",
  18235=>"011101111",
  18236=>"001000010",
  18237=>"001000001",
  18238=>"101010001",
  18239=>"101010010",
  18240=>"110011001",
  18241=>"000000101",
  18242=>"010101110",
  18243=>"100111001",
  18244=>"101110110",
  18245=>"010011010",
  18246=>"000010010",
  18247=>"100110111",
  18248=>"101000000",
  18249=>"111010000",
  18250=>"001000111",
  18251=>"000011111",
  18252=>"000010011",
  18253=>"001010001",
  18254=>"010011011",
  18255=>"011011001",
  18256=>"000000011",
  18257=>"000111101",
  18258=>"001010111",
  18259=>"000011110",
  18260=>"110101011",
  18261=>"100110111",
  18262=>"011001000",
  18263=>"111011011",
  18264=>"110010110",
  18265=>"101001011",
  18266=>"110010010",
  18267=>"111001011",
  18268=>"010001001",
  18269=>"011001010",
  18270=>"110110111",
  18271=>"001000111",
  18272=>"100011010",
  18273=>"010001111",
  18274=>"000101110",
  18275=>"001110100",
  18276=>"101000011",
  18277=>"001100011",
  18278=>"000011000",
  18279=>"001110010",
  18280=>"110111011",
  18281=>"111110100",
  18282=>"100001100",
  18283=>"000101111",
  18284=>"101101010",
  18285=>"011011110",
  18286=>"110111101",
  18287=>"101111000",
  18288=>"111001100",
  18289=>"101111000",
  18290=>"001011101",
  18291=>"110100101",
  18292=>"110110101",
  18293=>"010110000",
  18294=>"011110011",
  18295=>"001011000",
  18296=>"101000100",
  18297=>"011110010",
  18298=>"111000000",
  18299=>"111001101",
  18300=>"010100000",
  18301=>"111101110",
  18302=>"111000010",
  18303=>"110110110",
  18304=>"111111111",
  18305=>"001000000",
  18306=>"101010001",
  18307=>"010100101",
  18308=>"110100100",
  18309=>"111110110",
  18310=>"110101010",
  18311=>"000000010",
  18312=>"001101000",
  18313=>"111111011",
  18314=>"110101111",
  18315=>"010111011",
  18316=>"000011001",
  18317=>"100100010",
  18318=>"111011000",
  18319=>"100110111",
  18320=>"100000100",
  18321=>"111101000",
  18322=>"101010001",
  18323=>"001001000",
  18324=>"100010001",
  18325=>"111000011",
  18326=>"000000010",
  18327=>"011011101",
  18328=>"000110111",
  18329=>"111111011",
  18330=>"001110110",
  18331=>"110111110",
  18332=>"100110001",
  18333=>"111101011",
  18334=>"110110000",
  18335=>"101001111",
  18336=>"110011100",
  18337=>"110001100",
  18338=>"111111111",
  18339=>"000000111",
  18340=>"110101101",
  18341=>"100101010",
  18342=>"110100111",
  18343=>"001100111",
  18344=>"010001001",
  18345=>"010010000",
  18346=>"111011111",
  18347=>"001110111",
  18348=>"000100010",
  18349=>"111000011",
  18350=>"111010110",
  18351=>"110101110",
  18352=>"001011100",
  18353=>"111111010",
  18354=>"100100010",
  18355=>"111010110",
  18356=>"110110000",
  18357=>"001100110",
  18358=>"101110100",
  18359=>"101111010",
  18360=>"100101111",
  18361=>"111101101",
  18362=>"101111111",
  18363=>"110110101",
  18364=>"011000111",
  18365=>"100000000",
  18366=>"100010100",
  18367=>"001110001",
  18368=>"100011100",
  18369=>"001111100",
  18370=>"101000110",
  18371=>"010111000",
  18372=>"011111001",
  18373=>"010110111",
  18374=>"110110011",
  18375=>"001111000",
  18376=>"101101000",
  18377=>"011101100",
  18378=>"010110101",
  18379=>"000000001",
  18380=>"101011001",
  18381=>"100001001",
  18382=>"111100101",
  18383=>"010110101",
  18384=>"000011100",
  18385=>"000001010",
  18386=>"011011011",
  18387=>"011111001",
  18388=>"001000111",
  18389=>"011100111",
  18390=>"000001101",
  18391=>"011011001",
  18392=>"010000110",
  18393=>"010001100",
  18394=>"101111010",
  18395=>"001011111",
  18396=>"111010001",
  18397=>"111110001",
  18398=>"101000110",
  18399=>"001001100",
  18400=>"001110101",
  18401=>"100101010",
  18402=>"100111111",
  18403=>"001110000",
  18404=>"100001110",
  18405=>"011000001",
  18406=>"100111101",
  18407=>"100000111",
  18408=>"100000110",
  18409=>"110011100",
  18410=>"110001110",
  18411=>"110111011",
  18412=>"100000000",
  18413=>"010001110",
  18414=>"000000011",
  18415=>"000101101",
  18416=>"111110100",
  18417=>"111001111",
  18418=>"101011001",
  18419=>"011111100",
  18420=>"001100101",
  18421=>"011000001",
  18422=>"111110110",
  18423=>"011110010",
  18424=>"101111101",
  18425=>"000000110",
  18426=>"110011100",
  18427=>"110110001",
  18428=>"001001110",
  18429=>"001000100",
  18430=>"011100100",
  18431=>"111100101",
  18432=>"010110001",
  18433=>"111001100",
  18434=>"010010010",
  18435=>"001010001",
  18436=>"110110110",
  18437=>"010000100",
  18438=>"111011111",
  18439=>"101100110",
  18440=>"110011010",
  18441=>"000000010",
  18442=>"001100011",
  18443=>"111010011",
  18444=>"010011100",
  18445=>"001000000",
  18446=>"000101000",
  18447=>"111001110",
  18448=>"100101100",
  18449=>"000011010",
  18450=>"001011101",
  18451=>"010001101",
  18452=>"000100010",
  18453=>"001100001",
  18454=>"010101110",
  18455=>"011000000",
  18456=>"100010010",
  18457=>"010010011",
  18458=>"011000101",
  18459=>"111010010",
  18460=>"111101000",
  18461=>"010011010",
  18462=>"110010001",
  18463=>"110100000",
  18464=>"101000011",
  18465=>"001010100",
  18466=>"111100111",
  18467=>"001101010",
  18468=>"100000110",
  18469=>"000001011",
  18470=>"011000110",
  18471=>"111001000",
  18472=>"101100001",
  18473=>"000100111",
  18474=>"100111110",
  18475=>"000011000",
  18476=>"110110011",
  18477=>"100111111",
  18478=>"101111010",
  18479=>"111110100",
  18480=>"001010111",
  18481=>"011000100",
  18482=>"101000000",
  18483=>"000111010",
  18484=>"110111001",
  18485=>"001010000",
  18486=>"101110001",
  18487=>"110001111",
  18488=>"011100011",
  18489=>"110110011",
  18490=>"110010101",
  18491=>"110011011",
  18492=>"001011001",
  18493=>"110001100",
  18494=>"101110011",
  18495=>"001011111",
  18496=>"101010001",
  18497=>"101001101",
  18498=>"110111000",
  18499=>"011000011",
  18500=>"111011111",
  18501=>"110010010",
  18502=>"110100100",
  18503=>"110010011",
  18504=>"000100010",
  18505=>"011001001",
  18506=>"111100111",
  18507=>"100000001",
  18508=>"000011000",
  18509=>"010010101",
  18510=>"101100110",
  18511=>"011110000",
  18512=>"011110100",
  18513=>"010000101",
  18514=>"110000011",
  18515=>"001110010",
  18516=>"110100000",
  18517=>"000000000",
  18518=>"000011111",
  18519=>"011111001",
  18520=>"010100000",
  18521=>"011011111",
  18522=>"010000010",
  18523=>"111110000",
  18524=>"000011001",
  18525=>"101000111",
  18526=>"010111111",
  18527=>"010100010",
  18528=>"101101100",
  18529=>"010100100",
  18530=>"111001011",
  18531=>"011110011",
  18532=>"001001001",
  18533=>"101101000",
  18534=>"011111100",
  18535=>"110010000",
  18536=>"111100010",
  18537=>"101101010",
  18538=>"011111111",
  18539=>"101010011",
  18540=>"000000000",
  18541=>"100000111",
  18542=>"001111101",
  18543=>"010110000",
  18544=>"010111000",
  18545=>"001010110",
  18546=>"001000100",
  18547=>"101110001",
  18548=>"111111111",
  18549=>"110000111",
  18550=>"011110011",
  18551=>"011100000",
  18552=>"110011001",
  18553=>"110100111",
  18554=>"101010001",
  18555=>"000001110",
  18556=>"001000001",
  18557=>"101111011",
  18558=>"110001010",
  18559=>"010111100",
  18560=>"010001110",
  18561=>"110110110",
  18562=>"100011011",
  18563=>"111010100",
  18564=>"000100111",
  18565=>"101000000",
  18566=>"010010111",
  18567=>"001110000",
  18568=>"110110010",
  18569=>"101100101",
  18570=>"001010111",
  18571=>"101011100",
  18572=>"011000001",
  18573=>"100111001",
  18574=>"010011110",
  18575=>"011010001",
  18576=>"010101011",
  18577=>"101011100",
  18578=>"000011011",
  18579=>"101111111",
  18580=>"101001000",
  18581=>"110001010",
  18582=>"010100011",
  18583=>"110101101",
  18584=>"010101010",
  18585=>"111110100",
  18586=>"000101010",
  18587=>"000000011",
  18588=>"010010100",
  18589=>"001000100",
  18590=>"101111001",
  18591=>"011110000",
  18592=>"000100111",
  18593=>"001110011",
  18594=>"111010010",
  18595=>"111101101",
  18596=>"011010000",
  18597=>"001000010",
  18598=>"111011111",
  18599=>"010000110",
  18600=>"010000101",
  18601=>"000010011",
  18602=>"011111101",
  18603=>"000000000",
  18604=>"100001111",
  18605=>"001010101",
  18606=>"010000001",
  18607=>"011111010",
  18608=>"110001001",
  18609=>"000010000",
  18610=>"001100111",
  18611=>"001111011",
  18612=>"101101111",
  18613=>"111001111",
  18614=>"011000101",
  18615=>"000111100",
  18616=>"101000100",
  18617=>"000010001",
  18618=>"001001001",
  18619=>"000010010",
  18620=>"111110011",
  18621=>"110010000",
  18622=>"011010001",
  18623=>"001010101",
  18624=>"001000010",
  18625=>"000011010",
  18626=>"000101010",
  18627=>"011101101",
  18628=>"011100001",
  18629=>"001001000",
  18630=>"100001010",
  18631=>"110110010",
  18632=>"110110101",
  18633=>"001101001",
  18634=>"111011100",
  18635=>"111100011",
  18636=>"001011101",
  18637=>"100101010",
  18638=>"001010100",
  18639=>"011110011",
  18640=>"010011100",
  18641=>"011100001",
  18642=>"101100110",
  18643=>"101011111",
  18644=>"101111101",
  18645=>"100110001",
  18646=>"011011001",
  18647=>"010101100",
  18648=>"110010111",
  18649=>"001111010",
  18650=>"000100001",
  18651=>"000011000",
  18652=>"100011001",
  18653=>"100001100",
  18654=>"101111001",
  18655=>"110111111",
  18656=>"000101011",
  18657=>"000000010",
  18658=>"110011100",
  18659=>"000100011",
  18660=>"000001011",
  18661=>"110100101",
  18662=>"011010110",
  18663=>"010100001",
  18664=>"110111000",
  18665=>"101000110",
  18666=>"010010010",
  18667=>"000000000",
  18668=>"011101001",
  18669=>"101000000",
  18670=>"010010010",
  18671=>"010001000",
  18672=>"110101001",
  18673=>"010110010",
  18674=>"001001100",
  18675=>"110011000",
  18676=>"001110011",
  18677=>"001111010",
  18678=>"111110110",
  18679=>"000100100",
  18680=>"100110001",
  18681=>"001011100",
  18682=>"010111011",
  18683=>"000011010",
  18684=>"110110011",
  18685=>"111111000",
  18686=>"111101110",
  18687=>"110001011",
  18688=>"000000100",
  18689=>"001001111",
  18690=>"010101001",
  18691=>"111011000",
  18692=>"010111001",
  18693=>"101010000",
  18694=>"111110000",
  18695=>"000001001",
  18696=>"000100011",
  18697=>"110111010",
  18698=>"010110101",
  18699=>"010011110",
  18700=>"101101100",
  18701=>"000010010",
  18702=>"100011101",
  18703=>"111110100",
  18704=>"100011111",
  18705=>"100111011",
  18706=>"111111111",
  18707=>"000000111",
  18708=>"001011111",
  18709=>"010110101",
  18710=>"010010000",
  18711=>"111000110",
  18712=>"101011110",
  18713=>"111001000",
  18714=>"100010110",
  18715=>"011000010",
  18716=>"101111101",
  18717=>"001100101",
  18718=>"001001010",
  18719=>"011001001",
  18720=>"111010000",
  18721=>"001001010",
  18722=>"010001110",
  18723=>"100110001",
  18724=>"110001110",
  18725=>"111101000",
  18726=>"101101001",
  18727=>"011010010",
  18728=>"101101101",
  18729=>"000110011",
  18730=>"010001001",
  18731=>"000100101",
  18732=>"101111101",
  18733=>"110100110",
  18734=>"110101000",
  18735=>"100010001",
  18736=>"110010111",
  18737=>"100110011",
  18738=>"001011000",
  18739=>"111001110",
  18740=>"010011110",
  18741=>"110010010",
  18742=>"001110001",
  18743=>"011111111",
  18744=>"000000000",
  18745=>"011110010",
  18746=>"001000110",
  18747=>"000001111",
  18748=>"111010010",
  18749=>"011010011",
  18750=>"011100111",
  18751=>"100001100",
  18752=>"000010001",
  18753=>"010010101",
  18754=>"010001011",
  18755=>"011010001",
  18756=>"100011110",
  18757=>"000010011",
  18758=>"001101111",
  18759=>"001110101",
  18760=>"100110011",
  18761=>"111011100",
  18762=>"001000100",
  18763=>"100110011",
  18764=>"011000111",
  18765=>"110100101",
  18766=>"111010011",
  18767=>"111100001",
  18768=>"000001111",
  18769=>"110010011",
  18770=>"001011101",
  18771=>"111100110",
  18772=>"000001100",
  18773=>"111111010",
  18774=>"100000010",
  18775=>"011001011",
  18776=>"010001100",
  18777=>"010001111",
  18778=>"000010101",
  18779=>"001010000",
  18780=>"111010010",
  18781=>"111111111",
  18782=>"101110010",
  18783=>"100011010",
  18784=>"001100100",
  18785=>"011111001",
  18786=>"111001100",
  18787=>"000100011",
  18788=>"011010101",
  18789=>"111010101",
  18790=>"111100111",
  18791=>"010100011",
  18792=>"100001001",
  18793=>"001110100",
  18794=>"100010100",
  18795=>"110000011",
  18796=>"111000001",
  18797=>"100011011",
  18798=>"100101101",
  18799=>"001001011",
  18800=>"000010000",
  18801=>"101110111",
  18802=>"111100000",
  18803=>"110111110",
  18804=>"000000000",
  18805=>"110011000",
  18806=>"000101111",
  18807=>"111010000",
  18808=>"100110101",
  18809=>"100111001",
  18810=>"011110010",
  18811=>"100101111",
  18812=>"111100101",
  18813=>"001010010",
  18814=>"101110110",
  18815=>"100001110",
  18816=>"010101011",
  18817=>"110001001",
  18818=>"001011110",
  18819=>"011010101",
  18820=>"111011110",
  18821=>"010001100",
  18822=>"100100101",
  18823=>"010110100",
  18824=>"010000100",
  18825=>"011011100",
  18826=>"111110010",
  18827=>"100111110",
  18828=>"100000111",
  18829=>"101011000",
  18830=>"100100011",
  18831=>"111111010",
  18832=>"000010110",
  18833=>"101010010",
  18834=>"010011100",
  18835=>"110101100",
  18836=>"000010101",
  18837=>"011010010",
  18838=>"011100101",
  18839=>"011101100",
  18840=>"111110010",
  18841=>"100101011",
  18842=>"111011000",
  18843=>"101110011",
  18844=>"111011000",
  18845=>"010110100",
  18846=>"101100010",
  18847=>"001011100",
  18848=>"111110100",
  18849=>"000100101",
  18850=>"111001111",
  18851=>"011100001",
  18852=>"101111100",
  18853=>"000000001",
  18854=>"100111101",
  18855=>"000010001",
  18856=>"111101110",
  18857=>"111010101",
  18858=>"001000100",
  18859=>"010000100",
  18860=>"110000111",
  18861=>"000110101",
  18862=>"111111100",
  18863=>"011100001",
  18864=>"000010001",
  18865=>"111010011",
  18866=>"000011100",
  18867=>"000011100",
  18868=>"111100010",
  18869=>"100100100",
  18870=>"101000010",
  18871=>"100001111",
  18872=>"111111111",
  18873=>"100000101",
  18874=>"010111111",
  18875=>"001100010",
  18876=>"011111110",
  18877=>"000100001",
  18878=>"111101101",
  18879=>"000000001",
  18880=>"001000000",
  18881=>"000000011",
  18882=>"101010100",
  18883=>"001001101",
  18884=>"111110100",
  18885=>"010110110",
  18886=>"101011110",
  18887=>"001001000",
  18888=>"000000001",
  18889=>"110011111",
  18890=>"010110011",
  18891=>"010011001",
  18892=>"111001100",
  18893=>"011000110",
  18894=>"000100001",
  18895=>"010001010",
  18896=>"100000001",
  18897=>"010111000",
  18898=>"001001000",
  18899=>"011001000",
  18900=>"100010110",
  18901=>"101110110",
  18902=>"000001000",
  18903=>"011010010",
  18904=>"000010111",
  18905=>"111011011",
  18906=>"100100111",
  18907=>"110100000",
  18908=>"001000000",
  18909=>"111001100",
  18910=>"111101000",
  18911=>"000011000",
  18912=>"001110001",
  18913=>"111000101",
  18914=>"100101010",
  18915=>"010011100",
  18916=>"011100110",
  18917=>"010100001",
  18918=>"100110001",
  18919=>"100000001",
  18920=>"110110011",
  18921=>"111000000",
  18922=>"110100011",
  18923=>"011011101",
  18924=>"000100100",
  18925=>"101010000",
  18926=>"110001000",
  18927=>"001100011",
  18928=>"110011110",
  18929=>"110001011",
  18930=>"100000100",
  18931=>"011101000",
  18932=>"100110011",
  18933=>"111111011",
  18934=>"011110011",
  18935=>"010101100",
  18936=>"100101101",
  18937=>"101100100",
  18938=>"111111011",
  18939=>"100001011",
  18940=>"011110111",
  18941=>"101100010",
  18942=>"001000000",
  18943=>"110111100",
  18944=>"110100001",
  18945=>"100111111",
  18946=>"110011011",
  18947=>"000000110",
  18948=>"011100001",
  18949=>"111111010",
  18950=>"101110100",
  18951=>"100001110",
  18952=>"111111001",
  18953=>"101101111",
  18954=>"000010100",
  18955=>"110011100",
  18956=>"100011111",
  18957=>"000010010",
  18958=>"001000101",
  18959=>"000110010",
  18960=>"111000101",
  18961=>"011101111",
  18962=>"101111101",
  18963=>"011000011",
  18964=>"101111111",
  18965=>"010110100",
  18966=>"100010101",
  18967=>"011101111",
  18968=>"011101100",
  18969=>"010101011",
  18970=>"101011100",
  18971=>"111110101",
  18972=>"000000100",
  18973=>"000011000",
  18974=>"010001011",
  18975=>"111111111",
  18976=>"100111111",
  18977=>"001110101",
  18978=>"100000011",
  18979=>"000101010",
  18980=>"101010001",
  18981=>"100000000",
  18982=>"101000000",
  18983=>"101010000",
  18984=>"001001011",
  18985=>"001011000",
  18986=>"010010010",
  18987=>"110100010",
  18988=>"000100110",
  18989=>"011000111",
  18990=>"101011110",
  18991=>"111110011",
  18992=>"101010111",
  18993=>"000000000",
  18994=>"101101111",
  18995=>"011010111",
  18996=>"111100100",
  18997=>"001001001",
  18998=>"000000101",
  18999=>"011111011",
  19000=>"110010100",
  19001=>"101011111",
  19002=>"010010010",
  19003=>"101011110",
  19004=>"111101010",
  19005=>"111100010",
  19006=>"010100110",
  19007=>"000101110",
  19008=>"011111111",
  19009=>"011011100",
  19010=>"101100100",
  19011=>"010101001",
  19012=>"110100111",
  19013=>"101011111",
  19014=>"001110100",
  19015=>"000000010",
  19016=>"001100101",
  19017=>"100000110",
  19018=>"101000000",
  19019=>"110111111",
  19020=>"100100001",
  19021=>"010110111",
  19022=>"110000000",
  19023=>"010010000",
  19024=>"101011010",
  19025=>"000000010",
  19026=>"000100100",
  19027=>"000001001",
  19028=>"110100100",
  19029=>"010110111",
  19030=>"011000111",
  19031=>"011001111",
  19032=>"111000000",
  19033=>"110011001",
  19034=>"110000000",
  19035=>"110100110",
  19036=>"000010011",
  19037=>"000010000",
  19038=>"011111000",
  19039=>"001101111",
  19040=>"111101001",
  19041=>"011111010",
  19042=>"110001011",
  19043=>"111110000",
  19044=>"001110100",
  19045=>"111101001",
  19046=>"000001110",
  19047=>"111111110",
  19048=>"100011001",
  19049=>"110101101",
  19050=>"101010111",
  19051=>"100001101",
  19052=>"110001101",
  19053=>"010000111",
  19054=>"111111110",
  19055=>"111001011",
  19056=>"001010011",
  19057=>"000000111",
  19058=>"111100001",
  19059=>"010011111",
  19060=>"100101000",
  19061=>"101100101",
  19062=>"000111010",
  19063=>"000100001",
  19064=>"110101101",
  19065=>"111000001",
  19066=>"011111010",
  19067=>"001000101",
  19068=>"000101010",
  19069=>"100001110",
  19070=>"101000101",
  19071=>"001001010",
  19072=>"010000010",
  19073=>"100001010",
  19074=>"011111101",
  19075=>"101000100",
  19076=>"111000011",
  19077=>"010001001",
  19078=>"011010110",
  19079=>"100010101",
  19080=>"001100100",
  19081=>"100100101",
  19082=>"110110110",
  19083=>"010011001",
  19084=>"100110011",
  19085=>"001111011",
  19086=>"101010111",
  19087=>"000010110",
  19088=>"101011001",
  19089=>"011001101",
  19090=>"110010101",
  19091=>"110101010",
  19092=>"011110111",
  19093=>"000101111",
  19094=>"001000011",
  19095=>"001100001",
  19096=>"111000110",
  19097=>"111000000",
  19098=>"011000110",
  19099=>"001100110",
  19100=>"100100010",
  19101=>"100100100",
  19102=>"101000000",
  19103=>"011000001",
  19104=>"100111010",
  19105=>"000101110",
  19106=>"100100110",
  19107=>"001111001",
  19108=>"100111000",
  19109=>"100110111",
  19110=>"010011010",
  19111=>"100000111",
  19112=>"100110000",
  19113=>"001111001",
  19114=>"101101011",
  19115=>"011100101",
  19116=>"001000001",
  19117=>"110010101",
  19118=>"010011011",
  19119=>"110110001",
  19120=>"100101110",
  19121=>"011111111",
  19122=>"010001011",
  19123=>"001001000",
  19124=>"010011000",
  19125=>"101110101",
  19126=>"100100001",
  19127=>"110111101",
  19128=>"000000110",
  19129=>"010100110",
  19130=>"011111110",
  19131=>"100111111",
  19132=>"010010101",
  19133=>"001111111",
  19134=>"000101110",
  19135=>"011111001",
  19136=>"110001110",
  19137=>"011010100",
  19138=>"010001011",
  19139=>"100010010",
  19140=>"000001010",
  19141=>"001000111",
  19142=>"010011100",
  19143=>"111000011",
  19144=>"000111000",
  19145=>"111000100",
  19146=>"010111111",
  19147=>"110011101",
  19148=>"110101111",
  19149=>"000000011",
  19150=>"100101011",
  19151=>"010100101",
  19152=>"110111010",
  19153=>"000111011",
  19154=>"110111100",
  19155=>"000000110",
  19156=>"010010110",
  19157=>"011110001",
  19158=>"100101011",
  19159=>"000010100",
  19160=>"111111011",
  19161=>"110110010",
  19162=>"111110010",
  19163=>"110101111",
  19164=>"100010001",
  19165=>"111110101",
  19166=>"101010000",
  19167=>"010100000",
  19168=>"001000111",
  19169=>"010011010",
  19170=>"010100111",
  19171=>"000011001",
  19172=>"101100110",
  19173=>"011101011",
  19174=>"111101001",
  19175=>"111100100",
  19176=>"010000011",
  19177=>"101010111",
  19178=>"110011100",
  19179=>"000110011",
  19180=>"000000110",
  19181=>"000111100",
  19182=>"101101010",
  19183=>"010100000",
  19184=>"110111011",
  19185=>"101011111",
  19186=>"111000000",
  19187=>"011100000",
  19188=>"101010000",
  19189=>"101101000",
  19190=>"011010110",
  19191=>"010010100",
  19192=>"111001101",
  19193=>"100011000",
  19194=>"100100000",
  19195=>"101000100",
  19196=>"101100000",
  19197=>"010111010",
  19198=>"011100000",
  19199=>"001010000",
  19200=>"101010000",
  19201=>"111011101",
  19202=>"100000010",
  19203=>"100111001",
  19204=>"001000001",
  19205=>"000011101",
  19206=>"000001101",
  19207=>"111010001",
  19208=>"101011101",
  19209=>"010101101",
  19210=>"101000010",
  19211=>"000011100",
  19212=>"100000000",
  19213=>"001110110",
  19214=>"000010110",
  19215=>"010111111",
  19216=>"100000001",
  19217=>"011010001",
  19218=>"111101011",
  19219=>"111111111",
  19220=>"010101111",
  19221=>"101110111",
  19222=>"001000010",
  19223=>"111111110",
  19224=>"011011000",
  19225=>"010001001",
  19226=>"111111100",
  19227=>"000001010",
  19228=>"110000001",
  19229=>"000011100",
  19230=>"010010001",
  19231=>"001001001",
  19232=>"010101101",
  19233=>"111110010",
  19234=>"011011010",
  19235=>"011100010",
  19236=>"111001110",
  19237=>"011000110",
  19238=>"101001101",
  19239=>"000100100",
  19240=>"010001000",
  19241=>"100000100",
  19242=>"110001100",
  19243=>"111111101",
  19244=>"100101101",
  19245=>"001011110",
  19246=>"000011001",
  19247=>"001110111",
  19248=>"011111100",
  19249=>"111100011",
  19250=>"000101101",
  19251=>"011101001",
  19252=>"111011000",
  19253=>"011010100",
  19254=>"110100010",
  19255=>"101111110",
  19256=>"111111000",
  19257=>"011110000",
  19258=>"000001001",
  19259=>"110101011",
  19260=>"101111111",
  19261=>"111000111",
  19262=>"000110000",
  19263=>"110100101",
  19264=>"000111010",
  19265=>"000100001",
  19266=>"100001010",
  19267=>"000100000",
  19268=>"000001000",
  19269=>"010111111",
  19270=>"111111010",
  19271=>"110001000",
  19272=>"011000011",
  19273=>"100111000",
  19274=>"010000110",
  19275=>"000100010",
  19276=>"011011011",
  19277=>"000101010",
  19278=>"000011100",
  19279=>"101011110",
  19280=>"110010000",
  19281=>"000000010",
  19282=>"011010110",
  19283=>"010100111",
  19284=>"001010011",
  19285=>"001010010",
  19286=>"010001110",
  19287=>"111010001",
  19288=>"111000111",
  19289=>"011111111",
  19290=>"101101010",
  19291=>"101101011",
  19292=>"111111001",
  19293=>"100110001",
  19294=>"110101001",
  19295=>"000001110",
  19296=>"111111111",
  19297=>"000101001",
  19298=>"111100111",
  19299=>"000110110",
  19300=>"101011011",
  19301=>"010010001",
  19302=>"110101101",
  19303=>"010000000",
  19304=>"010010011",
  19305=>"100100010",
  19306=>"110011010",
  19307=>"100000001",
  19308=>"011010001",
  19309=>"100101001",
  19310=>"011011111",
  19311=>"110101110",
  19312=>"111000000",
  19313=>"000000111",
  19314=>"101101101",
  19315=>"110100101",
  19316=>"001100000",
  19317=>"110111011",
  19318=>"100110111",
  19319=>"001110011",
  19320=>"100001010",
  19321=>"010110100",
  19322=>"111100111",
  19323=>"101010100",
  19324=>"001001100",
  19325=>"011010000",
  19326=>"010100100",
  19327=>"101100101",
  19328=>"010110000",
  19329=>"101001101",
  19330=>"111011111",
  19331=>"001111010",
  19332=>"001100000",
  19333=>"011011000",
  19334=>"011010010",
  19335=>"100110011",
  19336=>"001101101",
  19337=>"111001001",
  19338=>"100101000",
  19339=>"000100110",
  19340=>"000000001",
  19341=>"011100101",
  19342=>"001010010",
  19343=>"000100001",
  19344=>"100111000",
  19345=>"101110110",
  19346=>"000000100",
  19347=>"011110011",
  19348=>"010110010",
  19349=>"101011010",
  19350=>"101111111",
  19351=>"111111101",
  19352=>"010001010",
  19353=>"111011011",
  19354=>"111100011",
  19355=>"011000101",
  19356=>"000001011",
  19357=>"111100001",
  19358=>"001111101",
  19359=>"011100000",
  19360=>"101101001",
  19361=>"101110110",
  19362=>"010110110",
  19363=>"010110000",
  19364=>"110110001",
  19365=>"101000000",
  19366=>"100100001",
  19367=>"011110110",
  19368=>"001001101",
  19369=>"000010000",
  19370=>"011011100",
  19371=>"000010110",
  19372=>"111011001",
  19373=>"110110000",
  19374=>"110100101",
  19375=>"101010100",
  19376=>"110101110",
  19377=>"011011101",
  19378=>"111100010",
  19379=>"000101111",
  19380=>"011110011",
  19381=>"010001100",
  19382=>"010001011",
  19383=>"000111001",
  19384=>"011000100",
  19385=>"100100010",
  19386=>"111000111",
  19387=>"100011100",
  19388=>"001110110",
  19389=>"101101111",
  19390=>"101010110",
  19391=>"110000100",
  19392=>"101000000",
  19393=>"011011100",
  19394=>"000001100",
  19395=>"000001110",
  19396=>"100000101",
  19397=>"100000001",
  19398=>"100101000",
  19399=>"101111010",
  19400=>"010100111",
  19401=>"000000000",
  19402=>"011101001",
  19403=>"001001100",
  19404=>"000111111",
  19405=>"000011000",
  19406=>"000111000",
  19407=>"010011110",
  19408=>"011011001",
  19409=>"011010010",
  19410=>"000000100",
  19411=>"111101101",
  19412=>"111010010",
  19413=>"000110001",
  19414=>"010001011",
  19415=>"111000110",
  19416=>"001010000",
  19417=>"110110100",
  19418=>"100011011",
  19419=>"010011101",
  19420=>"110011111",
  19421=>"101010000",
  19422=>"000111001",
  19423=>"001101100",
  19424=>"111010010",
  19425=>"100101101",
  19426=>"000001001",
  19427=>"100011001",
  19428=>"110100000",
  19429=>"011000111",
  19430=>"011010001",
  19431=>"001100001",
  19432=>"111101100",
  19433=>"101001010",
  19434=>"011000010",
  19435=>"101110110",
  19436=>"010101110",
  19437=>"011101111",
  19438=>"101000111",
  19439=>"100010110",
  19440=>"100101100",
  19441=>"011010010",
  19442=>"110001110",
  19443=>"101001000",
  19444=>"010000011",
  19445=>"001000111",
  19446=>"101001100",
  19447=>"111000111",
  19448=>"010101010",
  19449=>"011111011",
  19450=>"010011110",
  19451=>"011011111",
  19452=>"110000101",
  19453=>"111000100",
  19454=>"101000001",
  19455=>"000110001",
  19456=>"001011101",
  19457=>"000011110",
  19458=>"011001000",
  19459=>"101111111",
  19460=>"000010011",
  19461=>"110110010",
  19462=>"010101100",
  19463=>"111100101",
  19464=>"100101111",
  19465=>"100000100",
  19466=>"001111100",
  19467=>"100011101",
  19468=>"101011100",
  19469=>"100001001",
  19470=>"000110100",
  19471=>"100111110",
  19472=>"011101110",
  19473=>"101001011",
  19474=>"010110010",
  19475=>"000110101",
  19476=>"000110000",
  19477=>"000001011",
  19478=>"111101100",
  19479=>"010000110",
  19480=>"110011001",
  19481=>"010010110",
  19482=>"000111101",
  19483=>"010101111",
  19484=>"100010101",
  19485=>"110011001",
  19486=>"001011010",
  19487=>"001100110",
  19488=>"000101111",
  19489=>"100011011",
  19490=>"110011111",
  19491=>"110001001",
  19492=>"000110101",
  19493=>"001101101",
  19494=>"100101110",
  19495=>"110011111",
  19496=>"100111101",
  19497=>"000011001",
  19498=>"100010100",
  19499=>"111011101",
  19500=>"001111101",
  19501=>"011001111",
  19502=>"011001000",
  19503=>"000011111",
  19504=>"000101110",
  19505=>"001000111",
  19506=>"010010100",
  19507=>"101001001",
  19508=>"010010111",
  19509=>"010101011",
  19510=>"011100000",
  19511=>"111110010",
  19512=>"001011111",
  19513=>"111000010",
  19514=>"001100001",
  19515=>"000000010",
  19516=>"101101011",
  19517=>"101100100",
  19518=>"000001111",
  19519=>"010011111",
  19520=>"001011010",
  19521=>"010010001",
  19522=>"100101111",
  19523=>"000000010",
  19524=>"110011011",
  19525=>"100000101",
  19526=>"000001000",
  19527=>"101000110",
  19528=>"110011101",
  19529=>"110100010",
  19530=>"111111111",
  19531=>"100010001",
  19532=>"100001100",
  19533=>"101011000",
  19534=>"111010111",
  19535=>"101000111",
  19536=>"001100001",
  19537=>"000101000",
  19538=>"111001011",
  19539=>"100001010",
  19540=>"101111111",
  19541=>"001101011",
  19542=>"001001110",
  19543=>"111101011",
  19544=>"100010010",
  19545=>"000001110",
  19546=>"001001001",
  19547=>"010011000",
  19548=>"010011111",
  19549=>"000011101",
  19550=>"100011111",
  19551=>"001101010",
  19552=>"011010101",
  19553=>"000000110",
  19554=>"001010111",
  19555=>"011000011",
  19556=>"100011000",
  19557=>"100110100",
  19558=>"100011100",
  19559=>"101010101",
  19560=>"001100100",
  19561=>"000100111",
  19562=>"001110100",
  19563=>"100010101",
  19564=>"010001110",
  19565=>"100101010",
  19566=>"111101100",
  19567=>"001111111",
  19568=>"001100010",
  19569=>"110011001",
  19570=>"000110111",
  19571=>"001000111",
  19572=>"110011011",
  19573=>"101101101",
  19574=>"111111000",
  19575=>"100101000",
  19576=>"000110001",
  19577=>"001000010",
  19578=>"000011111",
  19579=>"010101001",
  19580=>"101000100",
  19581=>"000101001",
  19582=>"111000011",
  19583=>"111000000",
  19584=>"000110000",
  19585=>"010111010",
  19586=>"111011100",
  19587=>"100011011",
  19588=>"100001000",
  19589=>"000010010",
  19590=>"100101001",
  19591=>"010010001",
  19592=>"010111100",
  19593=>"000001100",
  19594=>"011000000",
  19595=>"001011011",
  19596=>"110111001",
  19597=>"110101001",
  19598=>"111010011",
  19599=>"100010011",
  19600=>"110011100",
  19601=>"111111110",
  19602=>"100011100",
  19603=>"100101111",
  19604=>"110011110",
  19605=>"000101010",
  19606=>"100000011",
  19607=>"011100111",
  19608=>"101000001",
  19609=>"100000000",
  19610=>"110111000",
  19611=>"000011100",
  19612=>"011101111",
  19613=>"110011101",
  19614=>"011001101",
  19615=>"001100111",
  19616=>"101101000",
  19617=>"110011111",
  19618=>"110101111",
  19619=>"110001011",
  19620=>"100101000",
  19621=>"110110100",
  19622=>"011010101",
  19623=>"000000000",
  19624=>"001101010",
  19625=>"010000000",
  19626=>"101011001",
  19627=>"100011000",
  19628=>"110111000",
  19629=>"101111010",
  19630=>"000001110",
  19631=>"110101001",
  19632=>"101100000",
  19633=>"000000001",
  19634=>"011101000",
  19635=>"101100101",
  19636=>"100001010",
  19637=>"100110111",
  19638=>"010011101",
  19639=>"111010111",
  19640=>"101010001",
  19641=>"110110101",
  19642=>"010110111",
  19643=>"101101001",
  19644=>"110110010",
  19645=>"000010111",
  19646=>"100101000",
  19647=>"011111000",
  19648=>"011000110",
  19649=>"101010100",
  19650=>"001010111",
  19651=>"010011101",
  19652=>"010000000",
  19653=>"000111010",
  19654=>"110101011",
  19655=>"001010001",
  19656=>"110000000",
  19657=>"000100111",
  19658=>"100110000",
  19659=>"100111111",
  19660=>"011110101",
  19661=>"011111110",
  19662=>"100000010",
  19663=>"010101110",
  19664=>"110110001",
  19665=>"001110100",
  19666=>"000101101",
  19667=>"011010110",
  19668=>"110111011",
  19669=>"000010010",
  19670=>"011010110",
  19671=>"001010100",
  19672=>"011000101",
  19673=>"101001111",
  19674=>"100000100",
  19675=>"011000110",
  19676=>"100100011",
  19677=>"110010111",
  19678=>"011111111",
  19679=>"000011000",
  19680=>"111000011",
  19681=>"100010000",
  19682=>"000101001",
  19683=>"001110100",
  19684=>"010001100",
  19685=>"011010010",
  19686=>"010000010",
  19687=>"010111110",
  19688=>"010000101",
  19689=>"110000001",
  19690=>"101110000",
  19691=>"101101001",
  19692=>"000000000",
  19693=>"000111010",
  19694=>"011010010",
  19695=>"011111001",
  19696=>"010001110",
  19697=>"100000011",
  19698=>"001000101",
  19699=>"110010110",
  19700=>"010110000",
  19701=>"000011101",
  19702=>"000111100",
  19703=>"101101101",
  19704=>"001011011",
  19705=>"111111111",
  19706=>"001001000",
  19707=>"001000011",
  19708=>"011101110",
  19709=>"011011100",
  19710=>"100100110",
  19711=>"100101000",
  19712=>"111101100",
  19713=>"100110111",
  19714=>"001001010",
  19715=>"000010011",
  19716=>"101110111",
  19717=>"000110010",
  19718=>"100100000",
  19719=>"001101101",
  19720=>"110111000",
  19721=>"110000000",
  19722=>"100101101",
  19723=>"001001011",
  19724=>"000001110",
  19725=>"101001111",
  19726=>"000010100",
  19727=>"000011000",
  19728=>"101111001",
  19729=>"111100100",
  19730=>"000011111",
  19731=>"000010100",
  19732=>"110001000",
  19733=>"101101111",
  19734=>"110111100",
  19735=>"110011000",
  19736=>"011001101",
  19737=>"010110001",
  19738=>"111011111",
  19739=>"011100001",
  19740=>"001111000",
  19741=>"011100100",
  19742=>"111001001",
  19743=>"100001000",
  19744=>"001110110",
  19745=>"100100110",
  19746=>"001010001",
  19747=>"101100101",
  19748=>"010101000",
  19749=>"100000110",
  19750=>"011101101",
  19751=>"000001110",
  19752=>"100111110",
  19753=>"010000111",
  19754=>"010010010",
  19755=>"010000010",
  19756=>"010010100",
  19757=>"010101111",
  19758=>"000000100",
  19759=>"110100000",
  19760=>"110100011",
  19761=>"011111000",
  19762=>"101010010",
  19763=>"001111111",
  19764=>"011100011",
  19765=>"000100010",
  19766=>"111001010",
  19767=>"110011011",
  19768=>"101101111",
  19769=>"110111011",
  19770=>"010110100",
  19771=>"111111110",
  19772=>"000000011",
  19773=>"101111100",
  19774=>"000101010",
  19775=>"010111111",
  19776=>"010010110",
  19777=>"001100110",
  19778=>"101000110",
  19779=>"010001101",
  19780=>"000101001",
  19781=>"001101001",
  19782=>"100000011",
  19783=>"000110011",
  19784=>"011100011",
  19785=>"100100000",
  19786=>"011010011",
  19787=>"010000001",
  19788=>"000101101",
  19789=>"000011001",
  19790=>"000010001",
  19791=>"101011110",
  19792=>"001111011",
  19793=>"010001000",
  19794=>"111001110",
  19795=>"101000000",
  19796=>"000011011",
  19797=>"100001100",
  19798=>"111111110",
  19799=>"100011011",
  19800=>"011000010",
  19801=>"111000101",
  19802=>"100101000",
  19803=>"011110110",
  19804=>"111011011",
  19805=>"111110011",
  19806=>"000001001",
  19807=>"100110110",
  19808=>"000111101",
  19809=>"010111101",
  19810=>"100010110",
  19811=>"101110110",
  19812=>"101100110",
  19813=>"110001000",
  19814=>"100100100",
  19815=>"111111001",
  19816=>"100010100",
  19817=>"000100000",
  19818=>"111001100",
  19819=>"001001100",
  19820=>"000010010",
  19821=>"011100110",
  19822=>"011100000",
  19823=>"101100011",
  19824=>"000010111",
  19825=>"010111010",
  19826=>"000101110",
  19827=>"111100010",
  19828=>"100011001",
  19829=>"111101111",
  19830=>"000100010",
  19831=>"001110000",
  19832=>"010100000",
  19833=>"101110110",
  19834=>"111001000",
  19835=>"011111111",
  19836=>"101110100",
  19837=>"111010001",
  19838=>"000100101",
  19839=>"011111110",
  19840=>"101001100",
  19841=>"010011110",
  19842=>"110110011",
  19843=>"101101010",
  19844=>"100101011",
  19845=>"101000010",
  19846=>"101000111",
  19847=>"111000000",
  19848=>"110101011",
  19849=>"011101001",
  19850=>"101010111",
  19851=>"110011100",
  19852=>"000001111",
  19853=>"001011010",
  19854=>"000000000",
  19855=>"111000000",
  19856=>"011011100",
  19857=>"000101000",
  19858=>"010010110",
  19859=>"111011100",
  19860=>"000110100",
  19861=>"110000111",
  19862=>"000110111",
  19863=>"100110000",
  19864=>"000011100",
  19865=>"111110111",
  19866=>"010011111",
  19867=>"010001000",
  19868=>"111110101",
  19869=>"011011000",
  19870=>"010001100",
  19871=>"110110110",
  19872=>"110001001",
  19873=>"101000010",
  19874=>"000010110",
  19875=>"001001000",
  19876=>"000110000",
  19877=>"101010100",
  19878=>"111110000",
  19879=>"000001101",
  19880=>"101000110",
  19881=>"000011011",
  19882=>"111101001",
  19883=>"111111110",
  19884=>"110000000",
  19885=>"011111101",
  19886=>"110000111",
  19887=>"001101101",
  19888=>"010011011",
  19889=>"101100100",
  19890=>"010010100",
  19891=>"110011001",
  19892=>"011101000",
  19893=>"100000001",
  19894=>"000111100",
  19895=>"111100011",
  19896=>"101110001",
  19897=>"001110000",
  19898=>"101011001",
  19899=>"000001000",
  19900=>"000100100",
  19901=>"011010001",
  19902=>"100111011",
  19903=>"110101010",
  19904=>"010101111",
  19905=>"111110101",
  19906=>"101111111",
  19907=>"111000001",
  19908=>"011110110",
  19909=>"100111000",
  19910=>"011111101",
  19911=>"000001001",
  19912=>"000001101",
  19913=>"110011111",
  19914=>"001000011",
  19915=>"000010101",
  19916=>"101110110",
  19917=>"111000000",
  19918=>"000111011",
  19919=>"011101011",
  19920=>"100110101",
  19921=>"100110111",
  19922=>"111000100",
  19923=>"111000100",
  19924=>"000101100",
  19925=>"000111010",
  19926=>"111011011",
  19927=>"000010100",
  19928=>"001100101",
  19929=>"110101001",
  19930=>"000011100",
  19931=>"111000010",
  19932=>"000000001",
  19933=>"100101011",
  19934=>"101000001",
  19935=>"000010111",
  19936=>"001100011",
  19937=>"110011101",
  19938=>"000101011",
  19939=>"010001111",
  19940=>"111011111",
  19941=>"011111010",
  19942=>"001111001",
  19943=>"101100100",
  19944=>"110010111",
  19945=>"100100110",
  19946=>"100001011",
  19947=>"110100000",
  19948=>"010011111",
  19949=>"100100010",
  19950=>"110100000",
  19951=>"011001110",
  19952=>"000111011",
  19953=>"111110011",
  19954=>"011001011",
  19955=>"000010000",
  19956=>"001111011",
  19957=>"011010000",
  19958=>"110111000",
  19959=>"111110111",
  19960=>"111000110",
  19961=>"001111001",
  19962=>"100010111",
  19963=>"011001111",
  19964=>"101011011",
  19965=>"100011001",
  19966=>"000000001",
  19967=>"010011000",
  19968=>"001111000",
  19969=>"111111000",
  19970=>"001110100",
  19971=>"110011101",
  19972=>"101000110",
  19973=>"000111011",
  19974=>"110000101",
  19975=>"011110110",
  19976=>"011001101",
  19977=>"100101000",
  19978=>"011110111",
  19979=>"000000010",
  19980=>"011111100",
  19981=>"110110111",
  19982=>"100011000",
  19983=>"011111101",
  19984=>"101111010",
  19985=>"000110100",
  19986=>"111101100",
  19987=>"111111111",
  19988=>"010111011",
  19989=>"001110000",
  19990=>"101010100",
  19991=>"110000110",
  19992=>"000000000",
  19993=>"011101000",
  19994=>"001000111",
  19995=>"011011011",
  19996=>"101100111",
  19997=>"010110111",
  19998=>"111110010",
  19999=>"101011111",
  20000=>"000101101",
  20001=>"010011001",
  20002=>"000100010",
  20003=>"100100111",
  20004=>"101000110",
  20005=>"110001111",
  20006=>"010111100",
  20007=>"111010101",
  20008=>"000000100",
  20009=>"101011110",
  20010=>"111011110",
  20011=>"110101111",
  20012=>"010011010",
  20013=>"010011011",
  20014=>"000000111",
  20015=>"011010001",
  20016=>"001001110",
  20017=>"001100111",
  20018=>"100110001",
  20019=>"111100100",
  20020=>"010100100",
  20021=>"011110000",
  20022=>"000001001",
  20023=>"011100010",
  20024=>"011110110",
  20025=>"110101011",
  20026=>"011100001",
  20027=>"101011100",
  20028=>"001001101",
  20029=>"110010000",
  20030=>"011101000",
  20031=>"100111101",
  20032=>"001000010",
  20033=>"100001001",
  20034=>"000000010",
  20035=>"100110111",
  20036=>"101100011",
  20037=>"101101001",
  20038=>"000000101",
  20039=>"100010011",
  20040=>"001111011",
  20041=>"010001111",
  20042=>"111001001",
  20043=>"111111010",
  20044=>"000000001",
  20045=>"100100100",
  20046=>"001000100",
  20047=>"010100000",
  20048=>"111110010",
  20049=>"101100010",
  20050=>"100011011",
  20051=>"010010000",
  20052=>"001110101",
  20053=>"000101000",
  20054=>"011001101",
  20055=>"101100111",
  20056=>"001010111",
  20057=>"011111101",
  20058=>"101111110",
  20059=>"110011011",
  20060=>"100011001",
  20061=>"000000100",
  20062=>"011101111",
  20063=>"010101101",
  20064=>"111011001",
  20065=>"110100110",
  20066=>"111011010",
  20067=>"001011101",
  20068=>"111111110",
  20069=>"001111111",
  20070=>"000011101",
  20071=>"111001000",
  20072=>"011000001",
  20073=>"110011100",
  20074=>"010100111",
  20075=>"000100101",
  20076=>"110011101",
  20077=>"111111010",
  20078=>"011000100",
  20079=>"010111100",
  20080=>"100110110",
  20081=>"100111011",
  20082=>"001111111",
  20083=>"000100110",
  20084=>"111101100",
  20085=>"001010001",
  20086=>"000101110",
  20087=>"000111001",
  20088=>"100101111",
  20089=>"011110011",
  20090=>"010000011",
  20091=>"100100100",
  20092=>"100000001",
  20093=>"001100010",
  20094=>"011011000",
  20095=>"111001101",
  20096=>"111111111",
  20097=>"000110110",
  20098=>"101010110",
  20099=>"100011010",
  20100=>"101010111",
  20101=>"001011111",
  20102=>"010001100",
  20103=>"111001101",
  20104=>"000001110",
  20105=>"000000110",
  20106=>"111101000",
  20107=>"001001010",
  20108=>"001101010",
  20109=>"110111000",
  20110=>"111000111",
  20111=>"100101111",
  20112=>"001110101",
  20113=>"100000101",
  20114=>"010100110",
  20115=>"010010100",
  20116=>"000010101",
  20117=>"011000011",
  20118=>"100010011",
  20119=>"010001001",
  20120=>"101001011",
  20121=>"100111111",
  20122=>"010010111",
  20123=>"001111100",
  20124=>"000111010",
  20125=>"100101110",
  20126=>"010100000",
  20127=>"100111011",
  20128=>"000110111",
  20129=>"101011111",
  20130=>"111010110",
  20131=>"100000010",
  20132=>"110001010",
  20133=>"111001101",
  20134=>"111000000",
  20135=>"111000111",
  20136=>"110000100",
  20137=>"011111010",
  20138=>"111010111",
  20139=>"110100000",
  20140=>"111101101",
  20141=>"011000100",
  20142=>"000111011",
  20143=>"000111110",
  20144=>"010011100",
  20145=>"001100000",
  20146=>"001100101",
  20147=>"111000000",
  20148=>"111111000",
  20149=>"111101100",
  20150=>"111111111",
  20151=>"100111101",
  20152=>"010110001",
  20153=>"110001100",
  20154=>"111001000",
  20155=>"011011010",
  20156=>"011011110",
  20157=>"010001001",
  20158=>"001110000",
  20159=>"101111110",
  20160=>"000001100",
  20161=>"010001111",
  20162=>"001011000",
  20163=>"100111011",
  20164=>"010000000",
  20165=>"101100011",
  20166=>"110000001",
  20167=>"111110110",
  20168=>"111111001",
  20169=>"000000000",
  20170=>"010000101",
  20171=>"010110001",
  20172=>"011010111",
  20173=>"001111010",
  20174=>"010110011",
  20175=>"011111010",
  20176=>"110010001",
  20177=>"100010111",
  20178=>"011110111",
  20179=>"111100110",
  20180=>"110111001",
  20181=>"010001101",
  20182=>"011110000",
  20183=>"000000110",
  20184=>"100101101",
  20185=>"001001100",
  20186=>"101010000",
  20187=>"000010111",
  20188=>"001110110",
  20189=>"000011111",
  20190=>"101001001",
  20191=>"010000011",
  20192=>"010100010",
  20193=>"001101100",
  20194=>"011110010",
  20195=>"000110111",
  20196=>"010001101",
  20197=>"110011111",
  20198=>"111101111",
  20199=>"101011010",
  20200=>"100101111",
  20201=>"101011111",
  20202=>"110000000",
  20203=>"100011010",
  20204=>"101110001",
  20205=>"001110001",
  20206=>"001100100",
  20207=>"101100100",
  20208=>"010110000",
  20209=>"110011011",
  20210=>"111100001",
  20211=>"011011010",
  20212=>"100110101",
  20213=>"010101100",
  20214=>"000100010",
  20215=>"111110111",
  20216=>"001001010",
  20217=>"110011100",
  20218=>"101101111",
  20219=>"110010010",
  20220=>"010001011",
  20221=>"000100000",
  20222=>"000111111",
  20223=>"101001111",
  20224=>"010000011",
  20225=>"110010000",
  20226=>"111001001",
  20227=>"010100100",
  20228=>"010001001",
  20229=>"110101001",
  20230=>"100111010",
  20231=>"011100111",
  20232=>"100110110",
  20233=>"010010010",
  20234=>"011001000",
  20235=>"111000101",
  20236=>"110000110",
  20237=>"110001010",
  20238=>"110110101",
  20239=>"110110011",
  20240=>"110011011",
  20241=>"110010001",
  20242=>"111101110",
  20243=>"100010011",
  20244=>"111111010",
  20245=>"101010001",
  20246=>"110011110",
  20247=>"110111011",
  20248=>"011001111",
  20249=>"110010111",
  20250=>"000100110",
  20251=>"101101010",
  20252=>"100001110",
  20253=>"010001101",
  20254=>"000101011",
  20255=>"111010000",
  20256=>"001110111",
  20257=>"111000110",
  20258=>"011100110",
  20259=>"111011111",
  20260=>"000100101",
  20261=>"110011110",
  20262=>"110001111",
  20263=>"110111011",
  20264=>"110110111",
  20265=>"111000000",
  20266=>"010101101",
  20267=>"100111111",
  20268=>"110111011",
  20269=>"110010111",
  20270=>"001000010",
  20271=>"110001101",
  20272=>"001101001",
  20273=>"010011110",
  20274=>"100111010",
  20275=>"000101001",
  20276=>"001110100",
  20277=>"110001011",
  20278=>"101111011",
  20279=>"110011010",
  20280=>"111000111",
  20281=>"110001101",
  20282=>"000100110",
  20283=>"000011110",
  20284=>"111110011",
  20285=>"000001111",
  20286=>"000000000",
  20287=>"000111011",
  20288=>"001001001",
  20289=>"000001111",
  20290=>"000101010",
  20291=>"010101001",
  20292=>"001111000",
  20293=>"011000110",
  20294=>"000100010",
  20295=>"101100000",
  20296=>"010010010",
  20297=>"000010110",
  20298=>"100010011",
  20299=>"011010101",
  20300=>"101000010",
  20301=>"111100001",
  20302=>"101110001",
  20303=>"000011001",
  20304=>"001100101",
  20305=>"001000000",
  20306=>"000110000",
  20307=>"000101100",
  20308=>"111101111",
  20309=>"010001101",
  20310=>"011111010",
  20311=>"100001100",
  20312=>"001001010",
  20313=>"001101000",
  20314=>"010101001",
  20315=>"100000100",
  20316=>"111110111",
  20317=>"000111101",
  20318=>"000001001",
  20319=>"000010010",
  20320=>"001001011",
  20321=>"101111011",
  20322=>"111010101",
  20323=>"001011111",
  20324=>"101000111",
  20325=>"111000101",
  20326=>"100100010",
  20327=>"111100110",
  20328=>"101111001",
  20329=>"001001001",
  20330=>"100100000",
  20331=>"110110000",
  20332=>"100111011",
  20333=>"000110111",
  20334=>"011100111",
  20335=>"001000000",
  20336=>"000000010",
  20337=>"100000101",
  20338=>"100000000",
  20339=>"000000011",
  20340=>"000111100",
  20341=>"111111001",
  20342=>"110110001",
  20343=>"100111101",
  20344=>"111101100",
  20345=>"110100010",
  20346=>"101011001",
  20347=>"111101011",
  20348=>"101101101",
  20349=>"111101001",
  20350=>"110111101",
  20351=>"000011001",
  20352=>"110000000",
  20353=>"110110111",
  20354=>"010001000",
  20355=>"011111101",
  20356=>"101101101",
  20357=>"100110110",
  20358=>"001111010",
  20359=>"111111110",
  20360=>"000000110",
  20361=>"101010100",
  20362=>"011111111",
  20363=>"101100000",
  20364=>"111111110",
  20365=>"000010000",
  20366=>"110111110",
  20367=>"110100100",
  20368=>"000001110",
  20369=>"111011100",
  20370=>"101001010",
  20371=>"001001111",
  20372=>"010100010",
  20373=>"001001001",
  20374=>"011111100",
  20375=>"010001101",
  20376=>"111111110",
  20377=>"000101000",
  20378=>"100010000",
  20379=>"010101011",
  20380=>"010000001",
  20381=>"001010010",
  20382=>"000110001",
  20383=>"000001100",
  20384=>"001010001",
  20385=>"101101000",
  20386=>"110010101",
  20387=>"010101110",
  20388=>"100111110",
  20389=>"000111011",
  20390=>"101101100",
  20391=>"011111101",
  20392=>"010001100",
  20393=>"101000111",
  20394=>"111100111",
  20395=>"011101001",
  20396=>"100101101",
  20397=>"101010100",
  20398=>"010101011",
  20399=>"000100011",
  20400=>"111010001",
  20401=>"000100110",
  20402=>"100000100",
  20403=>"000010000",
  20404=>"001011111",
  20405=>"111100011",
  20406=>"001110010",
  20407=>"110101000",
  20408=>"110000001",
  20409=>"000110111",
  20410=>"011111101",
  20411=>"000111100",
  20412=>"000000100",
  20413=>"101010000",
  20414=>"111100100",
  20415=>"110001100",
  20416=>"010001001",
  20417=>"101001000",
  20418=>"100011100",
  20419=>"110000101",
  20420=>"100010000",
  20421=>"000000110",
  20422=>"110100110",
  20423=>"011110000",
  20424=>"000010000",
  20425=>"101010011",
  20426=>"010110001",
  20427=>"010100000",
  20428=>"011101001",
  20429=>"010100010",
  20430=>"000110111",
  20431=>"110101010",
  20432=>"011110010",
  20433=>"010000101",
  20434=>"111000101",
  20435=>"110110010",
  20436=>"000101111",
  20437=>"001011111",
  20438=>"001111000",
  20439=>"000000011",
  20440=>"110110111",
  20441=>"011011000",
  20442=>"111110110",
  20443=>"001110010",
  20444=>"000001100",
  20445=>"111000100",
  20446=>"000100000",
  20447=>"001011010",
  20448=>"111001001",
  20449=>"100001101",
  20450=>"000000001",
  20451=>"111010010",
  20452=>"101101100",
  20453=>"000010011",
  20454=>"110011000",
  20455=>"000111000",
  20456=>"111110101",
  20457=>"011111001",
  20458=>"100011000",
  20459=>"000011001",
  20460=>"001011100",
  20461=>"111101111",
  20462=>"100101110",
  20463=>"011111111",
  20464=>"010101110",
  20465=>"000101010",
  20466=>"111111000",
  20467=>"010100100",
  20468=>"100100101",
  20469=>"100110101",
  20470=>"010101000",
  20471=>"011001000",
  20472=>"111101101",
  20473=>"010101000",
  20474=>"000100011",
  20475=>"001001000",
  20476=>"100100101",
  20477=>"001001110",
  20478=>"011110000",
  20479=>"011111111",
  20480=>"010111011",
  20481=>"110010000",
  20482=>"011000011",
  20483=>"101111101",
  20484=>"000101000",
  20485=>"010001010",
  20486=>"011010110",
  20487=>"110101001",
  20488=>"010100110",
  20489=>"101101101",
  20490=>"000011100",
  20491=>"011000111",
  20492=>"111001000",
  20493=>"001101111",
  20494=>"011000000",
  20495=>"001111111",
  20496=>"100010101",
  20497=>"001111101",
  20498=>"010110010",
  20499=>"100101001",
  20500=>"111101110",
  20501=>"011010111",
  20502=>"100011111",
  20503=>"110001000",
  20504=>"100011110",
  20505=>"001001111",
  20506=>"111100111",
  20507=>"010100101",
  20508=>"101110101",
  20509=>"111000010",
  20510=>"110011000",
  20511=>"100110110",
  20512=>"010101111",
  20513=>"101011001",
  20514=>"000100010",
  20515=>"100111010",
  20516=>"100100000",
  20517=>"000111101",
  20518=>"011101100",
  20519=>"110010000",
  20520=>"011100001",
  20521=>"111111101",
  20522=>"011110110",
  20523=>"111101101",
  20524=>"111111010",
  20525=>"100010010",
  20526=>"111001110",
  20527=>"001000011",
  20528=>"001010101",
  20529=>"100100110",
  20530=>"000100010",
  20531=>"010110100",
  20532=>"100100000",
  20533=>"101110100",
  20534=>"110100001",
  20535=>"001101010",
  20536=>"001100111",
  20537=>"010100001",
  20538=>"001011101",
  20539=>"101100110",
  20540=>"100111110",
  20541=>"011101000",
  20542=>"001110011",
  20543=>"011101111",
  20544=>"111000101",
  20545=>"000000000",
  20546=>"010000101",
  20547=>"100001100",
  20548=>"010000001",
  20549=>"000111101",
  20550=>"011111011",
  20551=>"010110110",
  20552=>"101011101",
  20553=>"100000101",
  20554=>"111111100",
  20555=>"100010101",
  20556=>"000100001",
  20557=>"111111001",
  20558=>"011011011",
  20559=>"011000010",
  20560=>"001111100",
  20561=>"000100110",
  20562=>"101011111",
  20563=>"001101000",
  20564=>"001010111",
  20565=>"101111011",
  20566=>"110110011",
  20567=>"010110101",
  20568=>"100110011",
  20569=>"001101011",
  20570=>"100000010",
  20571=>"001101000",
  20572=>"000010101",
  20573=>"110010101",
  20574=>"000011110",
  20575=>"110001000",
  20576=>"100111001",
  20577=>"001100010",
  20578=>"010000000",
  20579=>"100000110",
  20580=>"000000000",
  20581=>"011111011",
  20582=>"010001101",
  20583=>"111011010",
  20584=>"101011111",
  20585=>"111010000",
  20586=>"110010010",
  20587=>"100110011",
  20588=>"010101100",
  20589=>"111010110",
  20590=>"111011001",
  20591=>"010110100",
  20592=>"011100000",
  20593=>"011000000",
  20594=>"000110010",
  20595=>"011000110",
  20596=>"001110011",
  20597=>"001110000",
  20598=>"101001111",
  20599=>"011011011",
  20600=>"010111100",
  20601=>"010101001",
  20602=>"001101111",
  20603=>"010000001",
  20604=>"010101110",
  20605=>"010001011",
  20606=>"100000000",
  20607=>"101000111",
  20608=>"010010000",
  20609=>"100111000",
  20610=>"111111100",
  20611=>"011000010",
  20612=>"110011000",
  20613=>"001111011",
  20614=>"101101110",
  20615=>"001111101",
  20616=>"101011110",
  20617=>"001010011",
  20618=>"110111100",
  20619=>"101011110",
  20620=>"110010000",
  20621=>"000011111",
  20622=>"010101010",
  20623=>"000100000",
  20624=>"000110100",
  20625=>"110010111",
  20626=>"010101011",
  20627=>"000001101",
  20628=>"100011000",
  20629=>"111011110",
  20630=>"111000100",
  20631=>"101101100",
  20632=>"000100110",
  20633=>"011000000",
  20634=>"101100110",
  20635=>"000111001",
  20636=>"011000010",
  20637=>"110110111",
  20638=>"000100100",
  20639=>"010010011",
  20640=>"010111000",
  20641=>"001011000",
  20642=>"100111000",
  20643=>"001111000",
  20644=>"111100000",
  20645=>"101111010",
  20646=>"110000011",
  20647=>"100111001",
  20648=>"011000100",
  20649=>"101100000",
  20650=>"010110100",
  20651=>"100110010",
  20652=>"111100111",
  20653=>"100011111",
  20654=>"101000010",
  20655=>"000111111",
  20656=>"011111100",
  20657=>"010010110",
  20658=>"001110111",
  20659=>"101000000",
  20660=>"100010010",
  20661=>"011010001",
  20662=>"100111000",
  20663=>"001111000",
  20664=>"100100000",
  20665=>"111111011",
  20666=>"001110000",
  20667=>"110000111",
  20668=>"111001101",
  20669=>"101001001",
  20670=>"111101110",
  20671=>"001000001",
  20672=>"101100000",
  20673=>"011111000",
  20674=>"001010000",
  20675=>"001000010",
  20676=>"011101010",
  20677=>"010000000",
  20678=>"000101111",
  20679=>"100010100",
  20680=>"000011100",
  20681=>"001010110",
  20682=>"011000111",
  20683=>"000111110",
  20684=>"110111100",
  20685=>"101100011",
  20686=>"100100111",
  20687=>"011100000",
  20688=>"111011010",
  20689=>"011001010",
  20690=>"110011000",
  20691=>"110101111",
  20692=>"110100001",
  20693=>"000000001",
  20694=>"000000000",
  20695=>"010000111",
  20696=>"100101011",
  20697=>"010111011",
  20698=>"001010011",
  20699=>"111011001",
  20700=>"100110111",
  20701=>"111000101",
  20702=>"010100100",
  20703=>"010001000",
  20704=>"110101100",
  20705=>"110010110",
  20706=>"001000001",
  20707=>"011100101",
  20708=>"110101011",
  20709=>"000111110",
  20710=>"100100001",
  20711=>"111111101",
  20712=>"101001110",
  20713=>"101100010",
  20714=>"111111000",
  20715=>"101110100",
  20716=>"000000011",
  20717=>"000110001",
  20718=>"101100000",
  20719=>"011011100",
  20720=>"001101011",
  20721=>"111000001",
  20722=>"010011101",
  20723=>"101101101",
  20724=>"110000001",
  20725=>"000110100",
  20726=>"110011010",
  20727=>"101001111",
  20728=>"111010010",
  20729=>"010100010",
  20730=>"001100010",
  20731=>"101111101",
  20732=>"100011000",
  20733=>"110000010",
  20734=>"011111111",
  20735=>"011000101",
  20736=>"010100010",
  20737=>"100111000",
  20738=>"010111111",
  20739=>"000011110",
  20740=>"101101010",
  20741=>"100000010",
  20742=>"100111000",
  20743=>"110101101",
  20744=>"101001101",
  20745=>"111100110",
  20746=>"010011110",
  20747=>"110101000",
  20748=>"101111110",
  20749=>"100001011",
  20750=>"011010001",
  20751=>"100000110",
  20752=>"111110111",
  20753=>"100001011",
  20754=>"000100101",
  20755=>"001110010",
  20756=>"001010000",
  20757=>"010101101",
  20758=>"011001111",
  20759=>"000110010",
  20760=>"011100001",
  20761=>"101111010",
  20762=>"011000011",
  20763=>"111100100",
  20764=>"001101110",
  20765=>"000001001",
  20766=>"110000110",
  20767=>"000111110",
  20768=>"000000000",
  20769=>"011101010",
  20770=>"001000100",
  20771=>"111010101",
  20772=>"110011011",
  20773=>"110110101",
  20774=>"100011101",
  20775=>"010101101",
  20776=>"010001001",
  20777=>"111011111",
  20778=>"111011111",
  20779=>"010101001",
  20780=>"001101000",
  20781=>"101010001",
  20782=>"100000101",
  20783=>"100001001",
  20784=>"110101010",
  20785=>"001011111",
  20786=>"001010111",
  20787=>"000000010",
  20788=>"110010100",
  20789=>"000011000",
  20790=>"010110110",
  20791=>"111011011",
  20792=>"111001111",
  20793=>"110000001",
  20794=>"010111110",
  20795=>"000101010",
  20796=>"111011010",
  20797=>"101011100",
  20798=>"010111100",
  20799=>"101001000",
  20800=>"110011110",
  20801=>"010101011",
  20802=>"101100000",
  20803=>"011111111",
  20804=>"001110110",
  20805=>"010011100",
  20806=>"011100000",
  20807=>"100100000",
  20808=>"101010010",
  20809=>"110110100",
  20810=>"111010010",
  20811=>"001000000",
  20812=>"101111001",
  20813=>"101011101",
  20814=>"010110000",
  20815=>"111111111",
  20816=>"111111111",
  20817=>"110011101",
  20818=>"100011010",
  20819=>"011111111",
  20820=>"110111110",
  20821=>"101100110",
  20822=>"111001001",
  20823=>"000010100",
  20824=>"101110100",
  20825=>"001001001",
  20826=>"101011101",
  20827=>"100000000",
  20828=>"001001101",
  20829=>"000101100",
  20830=>"101111110",
  20831=>"000101000",
  20832=>"010010010",
  20833=>"001000111",
  20834=>"111101010",
  20835=>"110100000",
  20836=>"001000011",
  20837=>"011000000",
  20838=>"000010010",
  20839=>"110101010",
  20840=>"101011110",
  20841=>"100110100",
  20842=>"011001100",
  20843=>"001000010",
  20844=>"110010011",
  20845=>"010010001",
  20846=>"011010001",
  20847=>"000100001",
  20848=>"001101011",
  20849=>"101000010",
  20850=>"100111110",
  20851=>"111110010",
  20852=>"001110101",
  20853=>"000001010",
  20854=>"011111011",
  20855=>"111111100",
  20856=>"101000101",
  20857=>"010100101",
  20858=>"000000110",
  20859=>"010110111",
  20860=>"110001100",
  20861=>"010100100",
  20862=>"110101100",
  20863=>"110100111",
  20864=>"111111011",
  20865=>"101101001",
  20866=>"000101000",
  20867=>"000011111",
  20868=>"110001000",
  20869=>"100100111",
  20870=>"001101111",
  20871=>"111000100",
  20872=>"100001110",
  20873=>"010000111",
  20874=>"110111000",
  20875=>"111000111",
  20876=>"100010010",
  20877=>"110011000",
  20878=>"101101001",
  20879=>"111000101",
  20880=>"010010011",
  20881=>"100010000",
  20882=>"101100000",
  20883=>"001000110",
  20884=>"001001001",
  20885=>"011000000",
  20886=>"001110011",
  20887=>"100110001",
  20888=>"110011000",
  20889=>"110111101",
  20890=>"010000111",
  20891=>"000111111",
  20892=>"011100101",
  20893=>"101000010",
  20894=>"110100001",
  20895=>"011101110",
  20896=>"111101110",
  20897=>"000111000",
  20898=>"011100001",
  20899=>"101000111",
  20900=>"111111000",
  20901=>"111110011",
  20902=>"110110010",
  20903=>"000010111",
  20904=>"110011001",
  20905=>"111011000",
  20906=>"101010011",
  20907=>"101100100",
  20908=>"111110000",
  20909=>"010011010",
  20910=>"001011100",
  20911=>"100111001",
  20912=>"010011101",
  20913=>"000011110",
  20914=>"111101000",
  20915=>"010000000",
  20916=>"010100000",
  20917=>"101001100",
  20918=>"100110110",
  20919=>"010000010",
  20920=>"101101101",
  20921=>"011000001",
  20922=>"110110011",
  20923=>"101111000",
  20924=>"001000010",
  20925=>"000010001",
  20926=>"101011000",
  20927=>"011010000",
  20928=>"010011100",
  20929=>"101110011",
  20930=>"010110110",
  20931=>"110010000",
  20932=>"000110000",
  20933=>"110001111",
  20934=>"110101001",
  20935=>"110100100",
  20936=>"010000000",
  20937=>"000110010",
  20938=>"111100110",
  20939=>"100100010",
  20940=>"101110100",
  20941=>"011111111",
  20942=>"110111010",
  20943=>"111110111",
  20944=>"100100111",
  20945=>"000000001",
  20946=>"000010110",
  20947=>"001100011",
  20948=>"000101001",
  20949=>"000101000",
  20950=>"100001100",
  20951=>"101011100",
  20952=>"110110010",
  20953=>"110010111",
  20954=>"001000011",
  20955=>"111110010",
  20956=>"100100111",
  20957=>"101010000",
  20958=>"001000111",
  20959=>"111111100",
  20960=>"111000101",
  20961=>"101010100",
  20962=>"011111000",
  20963=>"000000101",
  20964=>"001100110",
  20965=>"100010100",
  20966=>"111111001",
  20967=>"100001111",
  20968=>"000001000",
  20969=>"001111011",
  20970=>"111111011",
  20971=>"101110010",
  20972=>"000110100",
  20973=>"000000100",
  20974=>"100100011",
  20975=>"011111010",
  20976=>"101110111",
  20977=>"101101110",
  20978=>"101111000",
  20979=>"000101000",
  20980=>"001100000",
  20981=>"010010011",
  20982=>"100001111",
  20983=>"000010100",
  20984=>"101011001",
  20985=>"000000001",
  20986=>"110110001",
  20987=>"000101111",
  20988=>"111000100",
  20989=>"000100000",
  20990=>"100111111",
  20991=>"000001111",
  20992=>"100110001",
  20993=>"101100010",
  20994=>"011100100",
  20995=>"111110110",
  20996=>"001111111",
  20997=>"111010110",
  20998=>"000100101",
  20999=>"101101011",
  21000=>"100100100",
  21001=>"101110011",
  21002=>"001001010",
  21003=>"010111010",
  21004=>"101000001",
  21005=>"100111011",
  21006=>"011000010",
  21007=>"000010100",
  21008=>"100011100",
  21009=>"000011011",
  21010=>"101001001",
  21011=>"000110000",
  21012=>"100001000",
  21013=>"000001100",
  21014=>"111111111",
  21015=>"001011110",
  21016=>"000101100",
  21017=>"010111000",
  21018=>"100000000",
  21019=>"000100000",
  21020=>"001011100",
  21021=>"111001000",
  21022=>"101111100",
  21023=>"011001110",
  21024=>"010011100",
  21025=>"110101100",
  21026=>"000100011",
  21027=>"110100011",
  21028=>"010001100",
  21029=>"010001000",
  21030=>"111111111",
  21031=>"010111100",
  21032=>"110100001",
  21033=>"110111101",
  21034=>"000001101",
  21035=>"100010010",
  21036=>"110000101",
  21037=>"011100101",
  21038=>"101110110",
  21039=>"001000011",
  21040=>"101011001",
  21041=>"100100110",
  21042=>"110011101",
  21043=>"001001011",
  21044=>"111100100",
  21045=>"000010100",
  21046=>"110001001",
  21047=>"000100111",
  21048=>"111001011",
  21049=>"101101111",
  21050=>"110111001",
  21051=>"011111011",
  21052=>"010111101",
  21053=>"010101101",
  21054=>"101011000",
  21055=>"110010110",
  21056=>"001101000",
  21057=>"010100110",
  21058=>"110010010",
  21059=>"001100000",
  21060=>"111111101",
  21061=>"001110111",
  21062=>"010001010",
  21063=>"000110001",
  21064=>"100110011",
  21065=>"011010100",
  21066=>"110111001",
  21067=>"001000110",
  21068=>"111100010",
  21069=>"100010111",
  21070=>"000111110",
  21071=>"101101010",
  21072=>"001110010",
  21073=>"001011000",
  21074=>"000101000",
  21075=>"010010110",
  21076=>"110100101",
  21077=>"111110000",
  21078=>"111101111",
  21079=>"000001001",
  21080=>"110001001",
  21081=>"000101111",
  21082=>"100011001",
  21083=>"001011111",
  21084=>"100100111",
  21085=>"001000110",
  21086=>"010001000",
  21087=>"110111000",
  21088=>"010101111",
  21089=>"000010011",
  21090=>"010011000",
  21091=>"110011110",
  21092=>"111100001",
  21093=>"001001110",
  21094=>"001000011",
  21095=>"010100011",
  21096=>"010011101",
  21097=>"000111010",
  21098=>"001111001",
  21099=>"001011100",
  21100=>"011101110",
  21101=>"111100011",
  21102=>"011110110",
  21103=>"000100011",
  21104=>"000100110",
  21105=>"100000101",
  21106=>"111101011",
  21107=>"000101010",
  21108=>"011001000",
  21109=>"110011110",
  21110=>"110100111",
  21111=>"100110010",
  21112=>"111010110",
  21113=>"111100111",
  21114=>"111011010",
  21115=>"101011000",
  21116=>"110101110",
  21117=>"110001111",
  21118=>"000101100",
  21119=>"001111011",
  21120=>"011000010",
  21121=>"001011101",
  21122=>"011100001",
  21123=>"011100111",
  21124=>"001001011",
  21125=>"101000001",
  21126=>"010011110",
  21127=>"110010011",
  21128=>"001111010",
  21129=>"110100000",
  21130=>"110011100",
  21131=>"100110000",
  21132=>"010000000",
  21133=>"100100000",
  21134=>"111011110",
  21135=>"001100111",
  21136=>"010000100",
  21137=>"000001111",
  21138=>"111111110",
  21139=>"101101011",
  21140=>"111010000",
  21141=>"111000100",
  21142=>"111100000",
  21143=>"110111101",
  21144=>"110000111",
  21145=>"011000101",
  21146=>"110011100",
  21147=>"011110011",
  21148=>"110010011",
  21149=>"111000011",
  21150=>"001011101",
  21151=>"010111110",
  21152=>"111000011",
  21153=>"101000011",
  21154=>"000100100",
  21155=>"111111101",
  21156=>"001011010",
  21157=>"001000111",
  21158=>"111101000",
  21159=>"100101111",
  21160=>"110111001",
  21161=>"011101111",
  21162=>"100110111",
  21163=>"000100001",
  21164=>"000011001",
  21165=>"101110000",
  21166=>"111001110",
  21167=>"110011100",
  21168=>"011011010",
  21169=>"011001000",
  21170=>"111101101",
  21171=>"001001010",
  21172=>"101111101",
  21173=>"000011000",
  21174=>"001111100",
  21175=>"010010010",
  21176=>"010110011",
  21177=>"000001110",
  21178=>"001000011",
  21179=>"101101001",
  21180=>"001111110",
  21181=>"010110010",
  21182=>"011110010",
  21183=>"011000111",
  21184=>"111101111",
  21185=>"001001001",
  21186=>"011101001",
  21187=>"000000100",
  21188=>"010011111",
  21189=>"111001101",
  21190=>"110000101",
  21191=>"011101000",
  21192=>"100010010",
  21193=>"111101101",
  21194=>"000111100",
  21195=>"000110110",
  21196=>"000010000",
  21197=>"110111101",
  21198=>"111100011",
  21199=>"110110100",
  21200=>"111010000",
  21201=>"101101111",
  21202=>"111001111",
  21203=>"110101110",
  21204=>"010111011",
  21205=>"000000111",
  21206=>"111110111",
  21207=>"010100001",
  21208=>"100001001",
  21209=>"110100010",
  21210=>"101111001",
  21211=>"001000110",
  21212=>"001010101",
  21213=>"110111110",
  21214=>"011010110",
  21215=>"000100001",
  21216=>"000100010",
  21217=>"101010111",
  21218=>"011001000",
  21219=>"011011111",
  21220=>"101100011",
  21221=>"111110010",
  21222=>"001110010",
  21223=>"001000101",
  21224=>"011010101",
  21225=>"111011100",
  21226=>"111110001",
  21227=>"100001111",
  21228=>"101101111",
  21229=>"101010100",
  21230=>"101010001",
  21231=>"010111110",
  21232=>"000010001",
  21233=>"111010111",
  21234=>"001101001",
  21235=>"000011111",
  21236=>"101111010",
  21237=>"100000101",
  21238=>"010110011",
  21239=>"011111101",
  21240=>"110101010",
  21241=>"000011001",
  21242=>"110111010",
  21243=>"011100001",
  21244=>"101111010",
  21245=>"100010101",
  21246=>"010100010",
  21247=>"100101110",
  21248=>"000100000",
  21249=>"010100100",
  21250=>"111111001",
  21251=>"011001111",
  21252=>"110010011",
  21253=>"101000100",
  21254=>"011011101",
  21255=>"101101000",
  21256=>"110111010",
  21257=>"100110001",
  21258=>"100100010",
  21259=>"100111100",
  21260=>"001101001",
  21261=>"011111001",
  21262=>"011101110",
  21263=>"111101110",
  21264=>"010111010",
  21265=>"101100001",
  21266=>"011111101",
  21267=>"000000010",
  21268=>"010110001",
  21269=>"111001010",
  21270=>"100000111",
  21271=>"000000010",
  21272=>"100000110",
  21273=>"010000010",
  21274=>"110001100",
  21275=>"110110011",
  21276=>"111001010",
  21277=>"110011110",
  21278=>"000000100",
  21279=>"111111110",
  21280=>"000010001",
  21281=>"010001111",
  21282=>"010001010",
  21283=>"001011010",
  21284=>"110000100",
  21285=>"000001010",
  21286=>"100101101",
  21287=>"010110010",
  21288=>"000110001",
  21289=>"000000001",
  21290=>"110100001",
  21291=>"101010011",
  21292=>"001100000",
  21293=>"000000000",
  21294=>"000011110",
  21295=>"010100101",
  21296=>"110001111",
  21297=>"110001110",
  21298=>"010111010",
  21299=>"110001001",
  21300=>"011010111",
  21301=>"100111110",
  21302=>"100101101",
  21303=>"001011110",
  21304=>"011100111",
  21305=>"110001001",
  21306=>"101000101",
  21307=>"111100110",
  21308=>"111000101",
  21309=>"011110101",
  21310=>"001111101",
  21311=>"111010101",
  21312=>"110110111",
  21313=>"000001010",
  21314=>"011001110",
  21315=>"111011111",
  21316=>"110100010",
  21317=>"100011110",
  21318=>"110110001",
  21319=>"000100101",
  21320=>"001010100",
  21321=>"110111001",
  21322=>"001011111",
  21323=>"000100110",
  21324=>"110000001",
  21325=>"010111100",
  21326=>"111100111",
  21327=>"111100001",
  21328=>"011010010",
  21329=>"100010010",
  21330=>"000011000",
  21331=>"111010001",
  21332=>"111111010",
  21333=>"110101010",
  21334=>"001010101",
  21335=>"111000111",
  21336=>"010001010",
  21337=>"100000001",
  21338=>"110101011",
  21339=>"110000000",
  21340=>"000000110",
  21341=>"101101110",
  21342=>"011100001",
  21343=>"001110101",
  21344=>"011101000",
  21345=>"000010001",
  21346=>"000000010",
  21347=>"100110001",
  21348=>"011011100",
  21349=>"000011010",
  21350=>"111100001",
  21351=>"111011100",
  21352=>"100000000",
  21353=>"111001011",
  21354=>"011100101",
  21355=>"100000101",
  21356=>"110101110",
  21357=>"111010110",
  21358=>"101101111",
  21359=>"010110111",
  21360=>"101000100",
  21361=>"110010100",
  21362=>"101001000",
  21363=>"100011101",
  21364=>"101001111",
  21365=>"001110011",
  21366=>"011001101",
  21367=>"011111100",
  21368=>"111001011",
  21369=>"000010100",
  21370=>"111011010",
  21371=>"011000000",
  21372=>"110101000",
  21373=>"110010100",
  21374=>"110111110",
  21375=>"111010011",
  21376=>"100011100",
  21377=>"110001000",
  21378=>"011111010",
  21379=>"100100000",
  21380=>"110111000",
  21381=>"111110100",
  21382=>"000101010",
  21383=>"001011111",
  21384=>"001110010",
  21385=>"111110110",
  21386=>"010100100",
  21387=>"010000110",
  21388=>"011001010",
  21389=>"010100100",
  21390=>"011100000",
  21391=>"000101011",
  21392=>"011011100",
  21393=>"100000101",
  21394=>"100111100",
  21395=>"111111000",
  21396=>"100110001",
  21397=>"100000100",
  21398=>"100010001",
  21399=>"000110100",
  21400=>"000010001",
  21401=>"010100011",
  21402=>"001011010",
  21403=>"110101000",
  21404=>"111011000",
  21405=>"001100100",
  21406=>"000100010",
  21407=>"111001010",
  21408=>"111001010",
  21409=>"010100000",
  21410=>"100010100",
  21411=>"111101010",
  21412=>"110001110",
  21413=>"100111011",
  21414=>"011000001",
  21415=>"000000000",
  21416=>"011011111",
  21417=>"011111100",
  21418=>"010011010",
  21419=>"101001111",
  21420=>"110011111",
  21421=>"100101011",
  21422=>"000100000",
  21423=>"100110000",
  21424=>"101110101",
  21425=>"001011001",
  21426=>"110001101",
  21427=>"111001100",
  21428=>"111100001",
  21429=>"110110101",
  21430=>"001100001",
  21431=>"101001100",
  21432=>"001101001",
  21433=>"001110001",
  21434=>"110011011",
  21435=>"011110110",
  21436=>"101100111",
  21437=>"000001100",
  21438=>"010110101",
  21439=>"011101000",
  21440=>"110101100",
  21441=>"101000100",
  21442=>"110100010",
  21443=>"010011101",
  21444=>"101011011",
  21445=>"101111000",
  21446=>"010100011",
  21447=>"111111001",
  21448=>"100010010",
  21449=>"110000010",
  21450=>"111011111",
  21451=>"111011101",
  21452=>"100110100",
  21453=>"110001010",
  21454=>"100011011",
  21455=>"101101110",
  21456=>"100011010",
  21457=>"010110100",
  21458=>"001100010",
  21459=>"010000111",
  21460=>"101011000",
  21461=>"101111001",
  21462=>"001000101",
  21463=>"100111011",
  21464=>"100010001",
  21465=>"010010101",
  21466=>"111010000",
  21467=>"101000010",
  21468=>"111010111",
  21469=>"010100011",
  21470=>"110100001",
  21471=>"111000001",
  21472=>"000000111",
  21473=>"110100100",
  21474=>"011011110",
  21475=>"011101101",
  21476=>"011011101",
  21477=>"010101000",
  21478=>"000100001",
  21479=>"011011010",
  21480=>"111100101",
  21481=>"110000101",
  21482=>"010100100",
  21483=>"000101000",
  21484=>"100101111",
  21485=>"110110100",
  21486=>"111000101",
  21487=>"110101001",
  21488=>"100111110",
  21489=>"100010001",
  21490=>"011000100",
  21491=>"010000100",
  21492=>"011010100",
  21493=>"000110101",
  21494=>"010001100",
  21495=>"110111000",
  21496=>"011111110",
  21497=>"011010011",
  21498=>"001111111",
  21499=>"101111001",
  21500=>"000011010",
  21501=>"000001000",
  21502=>"100101110",
  21503=>"000100011",
  21504=>"011100111",
  21505=>"101000010",
  21506=>"100100101",
  21507=>"100000100",
  21508=>"011010110",
  21509=>"010111100",
  21510=>"000111000",
  21511=>"000100001",
  21512=>"100100001",
  21513=>"010010101",
  21514=>"010010000",
  21515=>"011000001",
  21516=>"101000010",
  21517=>"011000101",
  21518=>"110011111",
  21519=>"001110011",
  21520=>"100010100",
  21521=>"100100111",
  21522=>"101010000",
  21523=>"000100101",
  21524=>"000100111",
  21525=>"111111110",
  21526=>"010011011",
  21527=>"011011000",
  21528=>"000100011",
  21529=>"011111111",
  21530=>"000110101",
  21531=>"000110110",
  21532=>"010001100",
  21533=>"101011000",
  21534=>"000001100",
  21535=>"110010000",
  21536=>"011100001",
  21537=>"110000011",
  21538=>"101011011",
  21539=>"101111100",
  21540=>"110110110",
  21541=>"101001001",
  21542=>"011011001",
  21543=>"111100011",
  21544=>"001101011",
  21545=>"001111111",
  21546=>"110110101",
  21547=>"011000111",
  21548=>"000000100",
  21549=>"011011010",
  21550=>"101100001",
  21551=>"000101000",
  21552=>"100000001",
  21553=>"110010101",
  21554=>"000010111",
  21555=>"111000010",
  21556=>"110001100",
  21557=>"011101101",
  21558=>"010111100",
  21559=>"110011000",
  21560=>"001101101",
  21561=>"101100111",
  21562=>"100010100",
  21563=>"110111100",
  21564=>"000100110",
  21565=>"010000110",
  21566=>"001010101",
  21567=>"101100100",
  21568=>"011010110",
  21569=>"001011010",
  21570=>"111001011",
  21571=>"000111011",
  21572=>"101100101",
  21573=>"010000010",
  21574=>"100110100",
  21575=>"111111111",
  21576=>"101000111",
  21577=>"101000001",
  21578=>"111111101",
  21579=>"000111001",
  21580=>"100111000",
  21581=>"000100111",
  21582=>"011010100",
  21583=>"011111111",
  21584=>"101110010",
  21585=>"110001001",
  21586=>"001100010",
  21587=>"110010110",
  21588=>"011000111",
  21589=>"110001111",
  21590=>"001010000",
  21591=>"101101101",
  21592=>"000100000",
  21593=>"100001101",
  21594=>"011011111",
  21595=>"011001100",
  21596=>"100011001",
  21597=>"110000101",
  21598=>"000010110",
  21599=>"100100100",
  21600=>"110010010",
  21601=>"111011111",
  21602=>"110101010",
  21603=>"010100001",
  21604=>"001000000",
  21605=>"011111101",
  21606=>"101100111",
  21607=>"010011110",
  21608=>"000010101",
  21609=>"111000111",
  21610=>"010001001",
  21611=>"011011111",
  21612=>"110100101",
  21613=>"101010110",
  21614=>"101100110",
  21615=>"100000111",
  21616=>"000101010",
  21617=>"000000010",
  21618=>"111000110",
  21619=>"010100001",
  21620=>"110001001",
  21621=>"100111100",
  21622=>"110001000",
  21623=>"000001110",
  21624=>"010000100",
  21625=>"101001000",
  21626=>"010000011",
  21627=>"100100011",
  21628=>"100001001",
  21629=>"000000001",
  21630=>"110110111",
  21631=>"100101000",
  21632=>"100000111",
  21633=>"100110101",
  21634=>"010011111",
  21635=>"110110111",
  21636=>"001001010",
  21637=>"011000100",
  21638=>"010011000",
  21639=>"111100000",
  21640=>"110000000",
  21641=>"110000001",
  21642=>"101001110",
  21643=>"000001011",
  21644=>"110100000",
  21645=>"111000001",
  21646=>"101101010",
  21647=>"001011011",
  21648=>"010101110",
  21649=>"010011110",
  21650=>"100111111",
  21651=>"010110111",
  21652=>"101111110",
  21653=>"001100000",
  21654=>"111001101",
  21655=>"101001100",
  21656=>"000011011",
  21657=>"111101101",
  21658=>"110011101",
  21659=>"000001001",
  21660=>"100001000",
  21661=>"010010010",
  21662=>"110000101",
  21663=>"001010111",
  21664=>"110110000",
  21665=>"110101101",
  21666=>"010100100",
  21667=>"011111100",
  21668=>"001110100",
  21669=>"000010000",
  21670=>"101001111",
  21671=>"111110101",
  21672=>"100001110",
  21673=>"011101011",
  21674=>"010101101",
  21675=>"110010110",
  21676=>"101101100",
  21677=>"011011111",
  21678=>"100111101",
  21679=>"100011011",
  21680=>"100001001",
  21681=>"100100110",
  21682=>"100001000",
  21683=>"011001001",
  21684=>"010101001",
  21685=>"011111101",
  21686=>"100001010",
  21687=>"001010111",
  21688=>"011001110",
  21689=>"011101100",
  21690=>"100110011",
  21691=>"100001000",
  21692=>"111000010",
  21693=>"110001000",
  21694=>"100110111",
  21695=>"110100001",
  21696=>"010110111",
  21697=>"101011001",
  21698=>"100111100",
  21699=>"111001110",
  21700=>"010110110",
  21701=>"010011010",
  21702=>"101001100",
  21703=>"101111100",
  21704=>"011001101",
  21705=>"011100010",
  21706=>"011000010",
  21707=>"111001111",
  21708=>"100011000",
  21709=>"011110010",
  21710=>"100100110",
  21711=>"000010100",
  21712=>"101100111",
  21713=>"001110010",
  21714=>"101110110",
  21715=>"000111111",
  21716=>"111011011",
  21717=>"110101101",
  21718=>"100111001",
  21719=>"110001011",
  21720=>"010111010",
  21721=>"000000100",
  21722=>"010110100",
  21723=>"010010001",
  21724=>"110001001",
  21725=>"111100010",
  21726=>"101010010",
  21727=>"110110011",
  21728=>"101111111",
  21729=>"100011100",
  21730=>"011001111",
  21731=>"001001011",
  21732=>"111011011",
  21733=>"101110111",
  21734=>"111011001",
  21735=>"101100001",
  21736=>"001110011",
  21737=>"101000011",
  21738=>"100001001",
  21739=>"101110011",
  21740=>"011010100",
  21741=>"101010001",
  21742=>"100110011",
  21743=>"001011111",
  21744=>"110010000",
  21745=>"111010100",
  21746=>"000110110",
  21747=>"111010110",
  21748=>"101010000",
  21749=>"000100010",
  21750=>"101110100",
  21751=>"111011111",
  21752=>"001111100",
  21753=>"011010000",
  21754=>"111110101",
  21755=>"001110101",
  21756=>"010110101",
  21757=>"100010110",
  21758=>"110101101",
  21759=>"111010100",
  21760=>"000011000",
  21761=>"010110000",
  21762=>"000010001",
  21763=>"100100000",
  21764=>"100000011",
  21765=>"100100010",
  21766=>"010000000",
  21767=>"100101011",
  21768=>"000011011",
  21769=>"010001110",
  21770=>"100011001",
  21771=>"110100100",
  21772=>"001111100",
  21773=>"101011000",
  21774=>"011011101",
  21775=>"001110101",
  21776=>"000010000",
  21777=>"101010011",
  21778=>"110100110",
  21779=>"110011001",
  21780=>"001100000",
  21781=>"010011001",
  21782=>"111000100",
  21783=>"111100110",
  21784=>"010011001",
  21785=>"010101000",
  21786=>"001101011",
  21787=>"000100110",
  21788=>"100100110",
  21789=>"111110100",
  21790=>"111110010",
  21791=>"000000101",
  21792=>"110010100",
  21793=>"001010010",
  21794=>"011110111",
  21795=>"001001000",
  21796=>"101000010",
  21797=>"111100110",
  21798=>"110111101",
  21799=>"001100110",
  21800=>"101111101",
  21801=>"101100110",
  21802=>"000010001",
  21803=>"010001000",
  21804=>"000110111",
  21805=>"010101010",
  21806=>"011000101",
  21807=>"111101101",
  21808=>"010110011",
  21809=>"111001011",
  21810=>"100111111",
  21811=>"001100000",
  21812=>"001011100",
  21813=>"111011011",
  21814=>"000110101",
  21815=>"011100001",
  21816=>"100111110",
  21817=>"101000011",
  21818=>"111110100",
  21819=>"001010001",
  21820=>"011001001",
  21821=>"000010101",
  21822=>"110001010",
  21823=>"000101001",
  21824=>"111000101",
  21825=>"100111001",
  21826=>"100111111",
  21827=>"110111111",
  21828=>"010110001",
  21829=>"000001110",
  21830=>"111010000",
  21831=>"000010111",
  21832=>"011010010",
  21833=>"100001111",
  21834=>"000111010",
  21835=>"111010100",
  21836=>"011000101",
  21837=>"100001001",
  21838=>"010000000",
  21839=>"000001001",
  21840=>"100010101",
  21841=>"110011100",
  21842=>"100010000",
  21843=>"011110011",
  21844=>"011011000",
  21845=>"011011111",
  21846=>"101000100",
  21847=>"001011010",
  21848=>"101100010",
  21849=>"010101000",
  21850=>"101100100",
  21851=>"000110000",
  21852=>"101100010",
  21853=>"101101000",
  21854=>"001011011",
  21855=>"101101011",
  21856=>"101010110",
  21857=>"101011101",
  21858=>"100111011",
  21859=>"101111111",
  21860=>"110001111",
  21861=>"101110010",
  21862=>"011100101",
  21863=>"111000001",
  21864=>"100101011",
  21865=>"000101101",
  21866=>"000001010",
  21867=>"111110101",
  21868=>"000100110",
  21869=>"000000100",
  21870=>"111010110",
  21871=>"101001010",
  21872=>"010101011",
  21873=>"000000001",
  21874=>"111011011",
  21875=>"101010000",
  21876=>"001000110",
  21877=>"111111101",
  21878=>"000101110",
  21879=>"111001010",
  21880=>"101001111",
  21881=>"001101000",
  21882=>"100000100",
  21883=>"110000000",
  21884=>"100011010",
  21885=>"010011101",
  21886=>"000111110",
  21887=>"111011100",
  21888=>"001001111",
  21889=>"000000010",
  21890=>"001001101",
  21891=>"100110111",
  21892=>"110100110",
  21893=>"010001001",
  21894=>"100100101",
  21895=>"011101001",
  21896=>"000000001",
  21897=>"001101110",
  21898=>"011010011",
  21899=>"101111011",
  21900=>"100010001",
  21901=>"000011001",
  21902=>"000101111",
  21903=>"101111100",
  21904=>"001001111",
  21905=>"100001110",
  21906=>"111101001",
  21907=>"011011010",
  21908=>"011100011",
  21909=>"111101000",
  21910=>"101000111",
  21911=>"111000111",
  21912=>"001111110",
  21913=>"111001001",
  21914=>"100000000",
  21915=>"001000000",
  21916=>"011011011",
  21917=>"100001101",
  21918=>"001111000",
  21919=>"010010011",
  21920=>"100101111",
  21921=>"001010000",
  21922=>"001001101",
  21923=>"110101111",
  21924=>"010010011",
  21925=>"000110000",
  21926=>"011100011",
  21927=>"111001000",
  21928=>"100111110",
  21929=>"000100101",
  21930=>"001111101",
  21931=>"011100011",
  21932=>"111111000",
  21933=>"010110010",
  21934=>"100111000",
  21935=>"000001100",
  21936=>"100110101",
  21937=>"000011100",
  21938=>"011101101",
  21939=>"100100011",
  21940=>"011011000",
  21941=>"101010000",
  21942=>"101111101",
  21943=>"000111011",
  21944=>"011110010",
  21945=>"100011000",
  21946=>"000101100",
  21947=>"110000001",
  21948=>"111000100",
  21949=>"100111010",
  21950=>"101001010",
  21951=>"010001001",
  21952=>"000011001",
  21953=>"110101010",
  21954=>"000010000",
  21955=>"101110011",
  21956=>"100111100",
  21957=>"111010001",
  21958=>"010110100",
  21959=>"111100101",
  21960=>"110100000",
  21961=>"100101110",
  21962=>"001100011",
  21963=>"011001100",
  21964=>"111110010",
  21965=>"100001111",
  21966=>"100110001",
  21967=>"011101000",
  21968=>"100101001",
  21969=>"011111000",
  21970=>"110010011",
  21971=>"111111111",
  21972=>"010011100",
  21973=>"100010100",
  21974=>"101010010",
  21975=>"101111001",
  21976=>"101011001",
  21977=>"111111001",
  21978=>"100101101",
  21979=>"001001101",
  21980=>"111111001",
  21981=>"010000101",
  21982=>"010000101",
  21983=>"001111010",
  21984=>"010110110",
  21985=>"000010011",
  21986=>"111100111",
  21987=>"010000110",
  21988=>"111101000",
  21989=>"000101111",
  21990=>"100100000",
  21991=>"011101011",
  21992=>"011101001",
  21993=>"010111100",
  21994=>"110110110",
  21995=>"100000000",
  21996=>"100010001",
  21997=>"000011111",
  21998=>"110000001",
  21999=>"010111001",
  22000=>"010010010",
  22001=>"000001100",
  22002=>"001011000",
  22003=>"001111010",
  22004=>"110101101",
  22005=>"100100100",
  22006=>"010011110",
  22007=>"110100110",
  22008=>"111111101",
  22009=>"111100010",
  22010=>"111111101",
  22011=>"001010100",
  22012=>"011111111",
  22013=>"000001110",
  22014=>"111011100",
  22015=>"110000001",
  22016=>"111011101",
  22017=>"101011111",
  22018=>"111011111",
  22019=>"001111110",
  22020=>"001001100",
  22021=>"000101101",
  22022=>"000100001",
  22023=>"111000100",
  22024=>"001000110",
  22025=>"010101011",
  22026=>"000011010",
  22027=>"000110100",
  22028=>"110000000",
  22029=>"001010011",
  22030=>"011001111",
  22031=>"101001000",
  22032=>"010010001",
  22033=>"101101000",
  22034=>"011011010",
  22035=>"100011001",
  22036=>"011000111",
  22037=>"101101011",
  22038=>"010011011",
  22039=>"011101111",
  22040=>"100000111",
  22041=>"110100001",
  22042=>"001101110",
  22043=>"001111011",
  22044=>"110110100",
  22045=>"001001100",
  22046=>"011000011",
  22047=>"000100010",
  22048=>"010111010",
  22049=>"110010000",
  22050=>"110011111",
  22051=>"000000010",
  22052=>"010011001",
  22053=>"001110100",
  22054=>"000000110",
  22055=>"100000000",
  22056=>"011100100",
  22057=>"010000011",
  22058=>"100000101",
  22059=>"011011100",
  22060=>"100100011",
  22061=>"010000010",
  22062=>"100000010",
  22063=>"101101001",
  22064=>"000110111",
  22065=>"101001100",
  22066=>"101110110",
  22067=>"000111001",
  22068=>"111110010",
  22069=>"001001000",
  22070=>"011110010",
  22071=>"100010011",
  22072=>"010000001",
  22073=>"100101011",
  22074=>"110011001",
  22075=>"100100110",
  22076=>"011001000",
  22077=>"010110110",
  22078=>"000110001",
  22079=>"010100000",
  22080=>"011111011",
  22081=>"000000110",
  22082=>"000000000",
  22083=>"001011111",
  22084=>"010000000",
  22085=>"100111111",
  22086=>"000101111",
  22087=>"011110011",
  22088=>"010101010",
  22089=>"100111101",
  22090=>"100110111",
  22091=>"111001011",
  22092=>"100011000",
  22093=>"000010010",
  22094=>"101000000",
  22095=>"110010100",
  22096=>"111111010",
  22097=>"010010010",
  22098=>"001011101",
  22099=>"011000110",
  22100=>"000000011",
  22101=>"111001000",
  22102=>"110110000",
  22103=>"110011001",
  22104=>"000100011",
  22105=>"010011111",
  22106=>"010100100",
  22107=>"010010111",
  22108=>"010011010",
  22109=>"010010111",
  22110=>"111110100",
  22111=>"010101000",
  22112=>"001110110",
  22113=>"101010100",
  22114=>"000000100",
  22115=>"010000011",
  22116=>"111000100",
  22117=>"010011100",
  22118=>"111000101",
  22119=>"101111110",
  22120=>"011000111",
  22121=>"111111011",
  22122=>"100100100",
  22123=>"100101100",
  22124=>"111110111",
  22125=>"010011001",
  22126=>"100110110",
  22127=>"110111101",
  22128=>"010100010",
  22129=>"110101110",
  22130=>"010000001",
  22131=>"010011110",
  22132=>"011010100",
  22133=>"000100111",
  22134=>"101111111",
  22135=>"010111000",
  22136=>"011100001",
  22137=>"000100100",
  22138=>"010101111",
  22139=>"011100101",
  22140=>"001100111",
  22141=>"011111101",
  22142=>"010000100",
  22143=>"000101110",
  22144=>"000110100",
  22145=>"011101001",
  22146=>"000010100",
  22147=>"001000000",
  22148=>"010101110",
  22149=>"000100010",
  22150=>"011000011",
  22151=>"111100101",
  22152=>"111111011",
  22153=>"011101111",
  22154=>"111010110",
  22155=>"011100000",
  22156=>"110110000",
  22157=>"001000110",
  22158=>"101010101",
  22159=>"011011001",
  22160=>"101111011",
  22161=>"110011010",
  22162=>"011111100",
  22163=>"011111100",
  22164=>"011010000",
  22165=>"000101000",
  22166=>"010001011",
  22167=>"001000010",
  22168=>"000100110",
  22169=>"110010101",
  22170=>"000000011",
  22171=>"111101001",
  22172=>"000010111",
  22173=>"101010101",
  22174=>"111111111",
  22175=>"101101000",
  22176=>"010111110",
  22177=>"111000000",
  22178=>"111100100",
  22179=>"100010001",
  22180=>"001100111",
  22181=>"011100111",
  22182=>"111110011",
  22183=>"000100001",
  22184=>"000110110",
  22185=>"100111111",
  22186=>"100110110",
  22187=>"010101101",
  22188=>"110110100",
  22189=>"001000111",
  22190=>"010011110",
  22191=>"110000001",
  22192=>"110110101",
  22193=>"001010011",
  22194=>"001001111",
  22195=>"101101100",
  22196=>"111001100",
  22197=>"110101100",
  22198=>"001010001",
  22199=>"110001100",
  22200=>"101101001",
  22201=>"111101101",
  22202=>"000011011",
  22203=>"110001100",
  22204=>"000100111",
  22205=>"101111101",
  22206=>"101101111",
  22207=>"100110101",
  22208=>"011110001",
  22209=>"011000101",
  22210=>"010011000",
  22211=>"000000011",
  22212=>"001101100",
  22213=>"000000001",
  22214=>"100110101",
  22215=>"101101101",
  22216=>"010100000",
  22217=>"111100110",
  22218=>"010011100",
  22219=>"010000010",
  22220=>"110111111",
  22221=>"010001100",
  22222=>"111100111",
  22223=>"011010001",
  22224=>"101001101",
  22225=>"101010011",
  22226=>"110010011",
  22227=>"001000111",
  22228=>"011100110",
  22229=>"010101010",
  22230=>"011100100",
  22231=>"011110011",
  22232=>"100000001",
  22233=>"101110101",
  22234=>"100001111",
  22235=>"001110001",
  22236=>"101101001",
  22237=>"101100101",
  22238=>"100100010",
  22239=>"111001110",
  22240=>"100000010",
  22241=>"111011111",
  22242=>"000110010",
  22243=>"010000010",
  22244=>"110110011",
  22245=>"110010111",
  22246=>"011100101",
  22247=>"010100101",
  22248=>"110110100",
  22249=>"011000110",
  22250=>"011000101",
  22251=>"000111100",
  22252=>"101101111",
  22253=>"011001001",
  22254=>"000000101",
  22255=>"110001100",
  22256=>"001100011",
  22257=>"011000010",
  22258=>"000010101",
  22259=>"011100000",
  22260=>"010010011",
  22261=>"011111111",
  22262=>"111011001",
  22263=>"001010110",
  22264=>"011110000",
  22265=>"000011000",
  22266=>"111111101",
  22267=>"100100100",
  22268=>"011001100",
  22269=>"001100010",
  22270=>"001101010",
  22271=>"011111001",
  22272=>"110000000",
  22273=>"100010111",
  22274=>"010001011",
  22275=>"111010101",
  22276=>"101000010",
  22277=>"101111011",
  22278=>"011110101",
  22279=>"011010001",
  22280=>"110101111",
  22281=>"001111000",
  22282=>"001000100",
  22283=>"010101010",
  22284=>"101111010",
  22285=>"011001000",
  22286=>"100111011",
  22287=>"111000100",
  22288=>"100001100",
  22289=>"100101011",
  22290=>"000010101",
  22291=>"100011000",
  22292=>"000010110",
  22293=>"101001100",
  22294=>"001001011",
  22295=>"101100111",
  22296=>"010101011",
  22297=>"010111010",
  22298=>"101011100",
  22299=>"100111110",
  22300=>"010011101",
  22301=>"001001010",
  22302=>"011001100",
  22303=>"110100101",
  22304=>"000100000",
  22305=>"011010001",
  22306=>"011001011",
  22307=>"110010011",
  22308=>"100100110",
  22309=>"010110101",
  22310=>"010000011",
  22311=>"111011110",
  22312=>"100101101",
  22313=>"110111010",
  22314=>"001001111",
  22315=>"101010010",
  22316=>"001000111",
  22317=>"011101111",
  22318=>"000110111",
  22319=>"000001011",
  22320=>"101110101",
  22321=>"110101010",
  22322=>"001000110",
  22323=>"100101000",
  22324=>"111000000",
  22325=>"010010111",
  22326=>"100010100",
  22327=>"000101111",
  22328=>"110100100",
  22329=>"100111101",
  22330=>"110101100",
  22331=>"100100110",
  22332=>"011011010",
  22333=>"001111010",
  22334=>"000000000",
  22335=>"111000100",
  22336=>"000011110",
  22337=>"010110010",
  22338=>"001000000",
  22339=>"100110111",
  22340=>"011100100",
  22341=>"010001011",
  22342=>"100001101",
  22343=>"100110101",
  22344=>"100000111",
  22345=>"011000010",
  22346=>"000011010",
  22347=>"101001101",
  22348=>"011010110",
  22349=>"111011011",
  22350=>"001101001",
  22351=>"011011111",
  22352=>"010011111",
  22353=>"101000110",
  22354=>"000111011",
  22355=>"101010101",
  22356=>"111011010",
  22357=>"010111110",
  22358=>"111000110",
  22359=>"010100111",
  22360=>"111011110",
  22361=>"111000010",
  22362=>"001100101",
  22363=>"100110010",
  22364=>"101100101",
  22365=>"010010010",
  22366=>"111011001",
  22367=>"000000111",
  22368=>"101010010",
  22369=>"101011110",
  22370=>"100011011",
  22371=>"001110111",
  22372=>"101001000",
  22373=>"010000101",
  22374=>"111110111",
  22375=>"101000000",
  22376=>"000010000",
  22377=>"001110100",
  22378=>"101111111",
  22379=>"110010000",
  22380=>"001101001",
  22381=>"111101000",
  22382=>"011010010",
  22383=>"101011101",
  22384=>"111111110",
  22385=>"111010110",
  22386=>"100000101",
  22387=>"001100110",
  22388=>"001100100",
  22389=>"010111010",
  22390=>"111011011",
  22391=>"001001011",
  22392=>"010111100",
  22393=>"110111100",
  22394=>"001011101",
  22395=>"101100101",
  22396=>"110110111",
  22397=>"001110001",
  22398=>"100111111",
  22399=>"110110110",
  22400=>"111110011",
  22401=>"011010110",
  22402=>"101011000",
  22403=>"101010000",
  22404=>"011001000",
  22405=>"000010000",
  22406=>"111111110",
  22407=>"111001110",
  22408=>"110010100",
  22409=>"100000011",
  22410=>"111001001",
  22411=>"001011011",
  22412=>"101000111",
  22413=>"011001001",
  22414=>"110110010",
  22415=>"001110111",
  22416=>"010110011",
  22417=>"000101011",
  22418=>"001111111",
  22419=>"100010111",
  22420=>"111110110",
  22421=>"100111111",
  22422=>"001010101",
  22423=>"000100010",
  22424=>"100010000",
  22425=>"010101101",
  22426=>"010110100",
  22427=>"110100100",
  22428=>"111010100",
  22429=>"101111100",
  22430=>"110101111",
  22431=>"011100100",
  22432=>"001100000",
  22433=>"110111001",
  22434=>"101001000",
  22435=>"110000111",
  22436=>"100110111",
  22437=>"010010001",
  22438=>"111111011",
  22439=>"001011100",
  22440=>"010000111",
  22441=>"110100101",
  22442=>"001010111",
  22443=>"001110110",
  22444=>"011000011",
  22445=>"101110011",
  22446=>"000111000",
  22447=>"100001011",
  22448=>"101010101",
  22449=>"111101000",
  22450=>"111111000",
  22451=>"101111101",
  22452=>"110111100",
  22453=>"100000101",
  22454=>"101100000",
  22455=>"010000100",
  22456=>"101110000",
  22457=>"010100101",
  22458=>"010111000",
  22459=>"001111001",
  22460=>"000000101",
  22461=>"110111101",
  22462=>"001111000",
  22463=>"011111101",
  22464=>"110111110",
  22465=>"000111110",
  22466=>"101000101",
  22467=>"011111101",
  22468=>"011001000",
  22469=>"010101100",
  22470=>"101000001",
  22471=>"000110010",
  22472=>"101010111",
  22473=>"001010111",
  22474=>"001011000",
  22475=>"000101010",
  22476=>"001100111",
  22477=>"001111100",
  22478=>"101000000",
  22479=>"101000001",
  22480=>"001110010",
  22481=>"000110001",
  22482=>"001001110",
  22483=>"001010100",
  22484=>"110110000",
  22485=>"010001011",
  22486=>"000111010",
  22487=>"000100001",
  22488=>"000111110",
  22489=>"101000110",
  22490=>"000001000",
  22491=>"100101100",
  22492=>"100010101",
  22493=>"010010001",
  22494=>"100111010",
  22495=>"111100000",
  22496=>"100001001",
  22497=>"111000111",
  22498=>"110010000",
  22499=>"010111101",
  22500=>"100011000",
  22501=>"110000101",
  22502=>"110000011",
  22503=>"110110000",
  22504=>"011010010",
  22505=>"100000100",
  22506=>"110110000",
  22507=>"000100111",
  22508=>"000111000",
  22509=>"101000111",
  22510=>"100100001",
  22511=>"111010111",
  22512=>"110101000",
  22513=>"010010011",
  22514=>"111111110",
  22515=>"101011111",
  22516=>"010101011",
  22517=>"110011000",
  22518=>"101010100",
  22519=>"101101110",
  22520=>"001101011",
  22521=>"011011011",
  22522=>"111101100",
  22523=>"100110001",
  22524=>"010110101",
  22525=>"100000010",
  22526=>"010000001",
  22527=>"010001000",
  22528=>"100101001",
  22529=>"011110111",
  22530=>"100010010",
  22531=>"001011101",
  22532=>"000010101",
  22533=>"001111000",
  22534=>"010010000",
  22535=>"010001010",
  22536=>"101011100",
  22537=>"101011100",
  22538=>"101111011",
  22539=>"100011110",
  22540=>"011100011",
  22541=>"101110111",
  22542=>"000110001",
  22543=>"111010111",
  22544=>"110100000",
  22545=>"000000010",
  22546=>"100001101",
  22547=>"010110101",
  22548=>"100010010",
  22549=>"000110101",
  22550=>"101101010",
  22551=>"000001001",
  22552=>"110101010",
  22553=>"111000000",
  22554=>"100111011",
  22555=>"101010100",
  22556=>"110001111",
  22557=>"101000010",
  22558=>"000010101",
  22559=>"100111010",
  22560=>"010111101",
  22561=>"101011011",
  22562=>"000000100",
  22563=>"000101010",
  22564=>"111100100",
  22565=>"110001011",
  22566=>"101011000",
  22567=>"000101000",
  22568=>"101001010",
  22569=>"111000000",
  22570=>"110010000",
  22571=>"011011010",
  22572=>"110111110",
  22573=>"111011101",
  22574=>"111011101",
  22575=>"100100001",
  22576=>"011111111",
  22577=>"001100100",
  22578=>"011101010",
  22579=>"011000010",
  22580=>"100001011",
  22581=>"101011110",
  22582=>"111001101",
  22583=>"011001011",
  22584=>"001100110",
  22585=>"101101111",
  22586=>"100101000",
  22587=>"110000010",
  22588=>"110101001",
  22589=>"010100010",
  22590=>"001111101",
  22591=>"011100010",
  22592=>"100110001",
  22593=>"111011100",
  22594=>"101000001",
  22595=>"101000111",
  22596=>"011100100",
  22597=>"001111100",
  22598=>"011000100",
  22599=>"100001000",
  22600=>"010101001",
  22601=>"000001000",
  22602=>"001111100",
  22603=>"100100000",
  22604=>"010111000",
  22605=>"100010101",
  22606=>"101111001",
  22607=>"010111011",
  22608=>"010011110",
  22609=>"011101101",
  22610=>"101000010",
  22611=>"011111100",
  22612=>"011101111",
  22613=>"111101101",
  22614=>"001000000",
  22615=>"111100101",
  22616=>"010101101",
  22617=>"110010101",
  22618=>"101111000",
  22619=>"110010111",
  22620=>"100010100",
  22621=>"101101100",
  22622=>"011000000",
  22623=>"011100011",
  22624=>"001101010",
  22625=>"011010001",
  22626=>"000110111",
  22627=>"000111101",
  22628=>"101000110",
  22629=>"010001101",
  22630=>"110111111",
  22631=>"111100000",
  22632=>"100111010",
  22633=>"100011001",
  22634=>"001000010",
  22635=>"001100101",
  22636=>"100111101",
  22637=>"110111011",
  22638=>"110011101",
  22639=>"100100010",
  22640=>"111010101",
  22641=>"111100101",
  22642=>"000101110",
  22643=>"011111001",
  22644=>"011011101",
  22645=>"110010100",
  22646=>"110101110",
  22647=>"010101011",
  22648=>"101111110",
  22649=>"010111000",
  22650=>"111101110",
  22651=>"101111000",
  22652=>"100000111",
  22653=>"010110110",
  22654=>"010010000",
  22655=>"111011110",
  22656=>"111111111",
  22657=>"111111000",
  22658=>"100101000",
  22659=>"001001011",
  22660=>"001111011",
  22661=>"111100010",
  22662=>"000110111",
  22663=>"000110100",
  22664=>"000110010",
  22665=>"111001010",
  22666=>"100001100",
  22667=>"111011111",
  22668=>"101011111",
  22669=>"110100001",
  22670=>"101001101",
  22671=>"100110000",
  22672=>"110001100",
  22673=>"111111111",
  22674=>"000100010",
  22675=>"110111110",
  22676=>"000101010",
  22677=>"000111011",
  22678=>"010010111",
  22679=>"010101001",
  22680=>"111111010",
  22681=>"010111001",
  22682=>"010101100",
  22683=>"100010111",
  22684=>"111000010",
  22685=>"111100111",
  22686=>"111101001",
  22687=>"010010010",
  22688=>"010111101",
  22689=>"001011111",
  22690=>"111101100",
  22691=>"000110101",
  22692=>"110110110",
  22693=>"011100111",
  22694=>"010100010",
  22695=>"011110001",
  22696=>"101101010",
  22697=>"101011111",
  22698=>"111111010",
  22699=>"111111100",
  22700=>"001000001",
  22701=>"001110111",
  22702=>"001101110",
  22703=>"000011011",
  22704=>"001001101",
  22705=>"111100010",
  22706=>"100111001",
  22707=>"100010100",
  22708=>"111010001",
  22709=>"001100000",
  22710=>"000001110",
  22711=>"000110001",
  22712=>"101100011",
  22713=>"100101010",
  22714=>"100001100",
  22715=>"011100110",
  22716=>"000001011",
  22717=>"101011000",
  22718=>"111000011",
  22719=>"110101001",
  22720=>"111101001",
  22721=>"011101001",
  22722=>"001100011",
  22723=>"000001000",
  22724=>"011110101",
  22725=>"110001101",
  22726=>"111011110",
  22727=>"100101100",
  22728=>"111100101",
  22729=>"001110100",
  22730=>"010000101",
  22731=>"011110001",
  22732=>"100111000",
  22733=>"111001011",
  22734=>"100010111",
  22735=>"010110001",
  22736=>"001101001",
  22737=>"111101001",
  22738=>"110000101",
  22739=>"100011001",
  22740=>"010101000",
  22741=>"000100111",
  22742=>"001110001",
  22743=>"110011110",
  22744=>"100101010",
  22745=>"011011110",
  22746=>"111101111",
  22747=>"010010101",
  22748=>"000110001",
  22749=>"111010001",
  22750=>"001101000",
  22751=>"110001010",
  22752=>"111011001",
  22753=>"000000101",
  22754=>"000011110",
  22755=>"000111101",
  22756=>"101010011",
  22757=>"111100101",
  22758=>"100011010",
  22759=>"010110100",
  22760=>"001100110",
  22761=>"111000111",
  22762=>"000100001",
  22763=>"111110111",
  22764=>"100000011",
  22765=>"000100011",
  22766=>"001011111",
  22767=>"100000100",
  22768=>"101100001",
  22769=>"111011011",
  22770=>"011101011",
  22771=>"111100001",
  22772=>"101010111",
  22773=>"101100101",
  22774=>"100000011",
  22775=>"111000101",
  22776=>"011101111",
  22777=>"101100110",
  22778=>"010101111",
  22779=>"100101001",
  22780=>"110111100",
  22781=>"100000101",
  22782=>"000111010",
  22783=>"111110000",
  22784=>"010010101",
  22785=>"011001101",
  22786=>"110101111",
  22787=>"001001111",
  22788=>"011111100",
  22789=>"101011000",
  22790=>"000010100",
  22791=>"110111000",
  22792=>"011000001",
  22793=>"100011011",
  22794=>"001101110",
  22795=>"001011000",
  22796=>"011001000",
  22797=>"101010011",
  22798=>"010111000",
  22799=>"101000100",
  22800=>"001110111",
  22801=>"100001111",
  22802=>"011110110",
  22803=>"111101011",
  22804=>"010010110",
  22805=>"110000010",
  22806=>"001110001",
  22807=>"011100011",
  22808=>"000010000",
  22809=>"011000111",
  22810=>"010010110",
  22811=>"000110110",
  22812=>"110100110",
  22813=>"010010010",
  22814=>"110010010",
  22815=>"000110011",
  22816=>"011110011",
  22817=>"100111111",
  22818=>"011101000",
  22819=>"000011100",
  22820=>"111000011",
  22821=>"110100101",
  22822=>"000110111",
  22823=>"110001111",
  22824=>"111111000",
  22825=>"100110110",
  22826=>"111100000",
  22827=>"100101100",
  22828=>"101110111",
  22829=>"001000101",
  22830=>"000010011",
  22831=>"001100110",
  22832=>"111111100",
  22833=>"111100110",
  22834=>"000111101",
  22835=>"111100000",
  22836=>"011110000",
  22837=>"010110111",
  22838=>"110000010",
  22839=>"101010111",
  22840=>"000011111",
  22841=>"010001111",
  22842=>"101100010",
  22843=>"000001011",
  22844=>"001010010",
  22845=>"000000110",
  22846=>"001010110",
  22847=>"100011010",
  22848=>"000000110",
  22849=>"100000111",
  22850=>"011100110",
  22851=>"111110011",
  22852=>"100001000",
  22853=>"000001011",
  22854=>"000100111",
  22855=>"101110110",
  22856=>"011011110",
  22857=>"001000101",
  22858=>"110000110",
  22859=>"101011111",
  22860=>"010110001",
  22861=>"111010111",
  22862=>"000111110",
  22863=>"000011011",
  22864=>"001001100",
  22865=>"001110001",
  22866=>"011011000",
  22867=>"010100100",
  22868=>"011110011",
  22869=>"111010000",
  22870=>"110010010",
  22871=>"111000010",
  22872=>"001011110",
  22873=>"111110111",
  22874=>"101110100",
  22875=>"111110001",
  22876=>"111110001",
  22877=>"011001101",
  22878=>"110001111",
  22879=>"001101010",
  22880=>"110101001",
  22881=>"001010001",
  22882=>"101100101",
  22883=>"110000000",
  22884=>"101111110",
  22885=>"011010100",
  22886=>"010010110",
  22887=>"101111110",
  22888=>"101011111",
  22889=>"111101110",
  22890=>"010100000",
  22891=>"011110101",
  22892=>"000101100",
  22893=>"010101011",
  22894=>"011111010",
  22895=>"000100001",
  22896=>"110111010",
  22897=>"111000000",
  22898=>"111010010",
  22899=>"011110010",
  22900=>"100001111",
  22901=>"010010010",
  22902=>"001101100",
  22903=>"001000101",
  22904=>"000001110",
  22905=>"100110111",
  22906=>"000100011",
  22907=>"110111101",
  22908=>"011100001",
  22909=>"101011100",
  22910=>"000101110",
  22911=>"000010010",
  22912=>"010001010",
  22913=>"101011001",
  22914=>"001000011",
  22915=>"100110000",
  22916=>"100001100",
  22917=>"111011000",
  22918=>"011000111",
  22919=>"101111111",
  22920=>"110000011",
  22921=>"010010010",
  22922=>"010110101",
  22923=>"001010011",
  22924=>"000001111",
  22925=>"111010010",
  22926=>"101101000",
  22927=>"110000011",
  22928=>"010101111",
  22929=>"000010001",
  22930=>"100000011",
  22931=>"010000101",
  22932=>"110010111",
  22933=>"101100101",
  22934=>"010111000",
  22935=>"010110110",
  22936=>"000101111",
  22937=>"011110100",
  22938=>"110010000",
  22939=>"000100100",
  22940=>"100001011",
  22941=>"010011000",
  22942=>"100010011",
  22943=>"011011100",
  22944=>"000001010",
  22945=>"000110111",
  22946=>"000111101",
  22947=>"111100100",
  22948=>"100010000",
  22949=>"001100001",
  22950=>"001111111",
  22951=>"001101100",
  22952=>"000011011",
  22953=>"010000101",
  22954=>"111001001",
  22955=>"100110010",
  22956=>"101111011",
  22957=>"111101111",
  22958=>"110111111",
  22959=>"010111110",
  22960=>"001011001",
  22961=>"010110011",
  22962=>"000100010",
  22963=>"100100101",
  22964=>"011111011",
  22965=>"000101011",
  22966=>"111110001",
  22967=>"001001000",
  22968=>"000010010",
  22969=>"010001001",
  22970=>"101100111",
  22971=>"001110111",
  22972=>"100001000",
  22973=>"000110111",
  22974=>"001100011",
  22975=>"010010001",
  22976=>"101100100",
  22977=>"001000111",
  22978=>"001110110",
  22979=>"011111100",
  22980=>"100011111",
  22981=>"011010101",
  22982=>"001101000",
  22983=>"011110111",
  22984=>"011001001",
  22985=>"000011110",
  22986=>"111100010",
  22987=>"111110001",
  22988=>"000001010",
  22989=>"010000000",
  22990=>"010001011",
  22991=>"101010011",
  22992=>"110000000",
  22993=>"010000010",
  22994=>"010101110",
  22995=>"111001111",
  22996=>"110001100",
  22997=>"110000010",
  22998=>"110111101",
  22999=>"110010110",
  23000=>"111101011",
  23001=>"011111010",
  23002=>"001110100",
  23003=>"010101111",
  23004=>"110000010",
  23005=>"001101110",
  23006=>"110111111",
  23007=>"000010100",
  23008=>"010000000",
  23009=>"111111000",
  23010=>"110110010",
  23011=>"101101011",
  23012=>"001111110",
  23013=>"010011010",
  23014=>"100010111",
  23015=>"011011011",
  23016=>"100101011",
  23017=>"100000110",
  23018=>"101110000",
  23019=>"001011110",
  23020=>"111010101",
  23021=>"010011101",
  23022=>"011011001",
  23023=>"010001011",
  23024=>"111110111",
  23025=>"110001111",
  23026=>"100010001",
  23027=>"010100111",
  23028=>"011001010",
  23029=>"001010100",
  23030=>"101100001",
  23031=>"111011011",
  23032=>"000001001",
  23033=>"001100010",
  23034=>"101010100",
  23035=>"001001110",
  23036=>"010000000",
  23037=>"010101000",
  23038=>"000011010",
  23039=>"011101100",
  23040=>"111011001",
  23041=>"010111100",
  23042=>"011010001",
  23043=>"000111011",
  23044=>"000000110",
  23045=>"111010100",
  23046=>"110010001",
  23047=>"001111100",
  23048=>"010111011",
  23049=>"110100100",
  23050=>"011011101",
  23051=>"110001010",
  23052=>"001011101",
  23053=>"101000111",
  23054=>"110110110",
  23055=>"100010001",
  23056=>"110010011",
  23057=>"010010010",
  23058=>"101100100",
  23059=>"000011001",
  23060=>"000110111",
  23061=>"100111101",
  23062=>"000000000",
  23063=>"010110010",
  23064=>"001010101",
  23065=>"110111100",
  23066=>"111100100",
  23067=>"001011001",
  23068=>"111000100",
  23069=>"010000101",
  23070=>"101000111",
  23071=>"100010011",
  23072=>"111010101",
  23073=>"011110011",
  23074=>"011001010",
  23075=>"011110111",
  23076=>"110111111",
  23077=>"111100010",
  23078=>"011001100",
  23079=>"110111100",
  23080=>"111101001",
  23081=>"100110111",
  23082=>"111011011",
  23083=>"101001110",
  23084=>"000101011",
  23085=>"011101100",
  23086=>"111011011",
  23087=>"111111111",
  23088=>"011010010",
  23089=>"111001011",
  23090=>"000011111",
  23091=>"110001001",
  23092=>"101000101",
  23093=>"101011100",
  23094=>"100011100",
  23095=>"011001100",
  23096=>"001001111",
  23097=>"000100111",
  23098=>"100111011",
  23099=>"010100000",
  23100=>"010100011",
  23101=>"000101101",
  23102=>"000010000",
  23103=>"101101101",
  23104=>"000101000",
  23105=>"010111000",
  23106=>"011111001",
  23107=>"111111010",
  23108=>"101100000",
  23109=>"000000111",
  23110=>"111111110",
  23111=>"011110010",
  23112=>"110100011",
  23113=>"011100010",
  23114=>"110000011",
  23115=>"000110010",
  23116=>"110111110",
  23117=>"101001101",
  23118=>"001010110",
  23119=>"010011010",
  23120=>"000001001",
  23121=>"100111010",
  23122=>"010011001",
  23123=>"011111010",
  23124=>"101011110",
  23125=>"111000010",
  23126=>"000101000",
  23127=>"000000010",
  23128=>"011100001",
  23129=>"101101000",
  23130=>"101101110",
  23131=>"001100110",
  23132=>"100111000",
  23133=>"011011000",
  23134=>"000001111",
  23135=>"111001101",
  23136=>"000001010",
  23137=>"100000001",
  23138=>"001100001",
  23139=>"011101110",
  23140=>"110111011",
  23141=>"001011100",
  23142=>"010111010",
  23143=>"111101010",
  23144=>"100110110",
  23145=>"010010110",
  23146=>"101110101",
  23147=>"011011010",
  23148=>"000011001",
  23149=>"011001000",
  23150=>"111101011",
  23151=>"101000000",
  23152=>"110000010",
  23153=>"101001011",
  23154=>"010011001",
  23155=>"110101100",
  23156=>"111010110",
  23157=>"111000110",
  23158=>"011010010",
  23159=>"111101100",
  23160=>"110101010",
  23161=>"000011110",
  23162=>"110000101",
  23163=>"100111111",
  23164=>"100101100",
  23165=>"101000011",
  23166=>"101001111",
  23167=>"110001101",
  23168=>"000000100",
  23169=>"011100110",
  23170=>"111000110",
  23171=>"000101111",
  23172=>"111010000",
  23173=>"001010001",
  23174=>"010011100",
  23175=>"000010010",
  23176=>"010001101",
  23177=>"000100000",
  23178=>"010101100",
  23179=>"000011111",
  23180=>"010011111",
  23181=>"011001001",
  23182=>"111100101",
  23183=>"101110011",
  23184=>"000100110",
  23185=>"101011011",
  23186=>"010010101",
  23187=>"101111010",
  23188=>"000100110",
  23189=>"011000001",
  23190=>"000001110",
  23191=>"110011110",
  23192=>"101011100",
  23193=>"000011001",
  23194=>"100010100",
  23195=>"000011011",
  23196=>"111110011",
  23197=>"100100110",
  23198=>"100001110",
  23199=>"110011101",
  23200=>"111101011",
  23201=>"010110111",
  23202=>"111000011",
  23203=>"000101100",
  23204=>"010011100",
  23205=>"000111010",
  23206=>"111000011",
  23207=>"001000000",
  23208=>"101001000",
  23209=>"011101001",
  23210=>"011001101",
  23211=>"000100010",
  23212=>"101000001",
  23213=>"110110010",
  23214=>"010100111",
  23215=>"000001000",
  23216=>"100001011",
  23217=>"101100101",
  23218=>"000001011",
  23219=>"111110010",
  23220=>"101111010",
  23221=>"000110011",
  23222=>"010110110",
  23223=>"110010100",
  23224=>"101011111",
  23225=>"010100101",
  23226=>"111010111",
  23227=>"110011110",
  23228=>"111011000",
  23229=>"101100010",
  23230=>"010001001",
  23231=>"100111000",
  23232=>"111000000",
  23233=>"100111011",
  23234=>"010010100",
  23235=>"111100111",
  23236=>"111101000",
  23237=>"111000100",
  23238=>"011000101",
  23239=>"011111000",
  23240=>"000011000",
  23241=>"100000111",
  23242=>"010110111",
  23243=>"001100010",
  23244=>"001001101",
  23245=>"001000000",
  23246=>"110000010",
  23247=>"011010001",
  23248=>"100110010",
  23249=>"000010010",
  23250=>"110100110",
  23251=>"011101100",
  23252=>"010000100",
  23253=>"011111101",
  23254=>"101000101",
  23255=>"000100010",
  23256=>"011111111",
  23257=>"000100001",
  23258=>"111001010",
  23259=>"110001110",
  23260=>"100001101",
  23261=>"111101011",
  23262=>"010000010",
  23263=>"010011001",
  23264=>"100101000",
  23265=>"100100010",
  23266=>"000111011",
  23267=>"101110010",
  23268=>"111111010",
  23269=>"110001111",
  23270=>"000110111",
  23271=>"110010101",
  23272=>"101110010",
  23273=>"100100100",
  23274=>"111010110",
  23275=>"000100010",
  23276=>"100111100",
  23277=>"110010101",
  23278=>"001001001",
  23279=>"111000111",
  23280=>"011011110",
  23281=>"111111001",
  23282=>"000001001",
  23283=>"011111100",
  23284=>"010011101",
  23285=>"110110101",
  23286=>"001110110",
  23287=>"000011110",
  23288=>"111000110",
  23289=>"001111111",
  23290=>"000100100",
  23291=>"111011001",
  23292=>"101101101",
  23293=>"000101010",
  23294=>"010000011",
  23295=>"000110111",
  23296=>"001011000",
  23297=>"100111000",
  23298=>"010010010",
  23299=>"001111100",
  23300=>"000001110",
  23301=>"111001101",
  23302=>"101101101",
  23303=>"011110100",
  23304=>"100111111",
  23305=>"000010011",
  23306=>"101011011",
  23307=>"011110111",
  23308=>"011001001",
  23309=>"110001000",
  23310=>"011110110",
  23311=>"000011111",
  23312=>"001100001",
  23313=>"100101011",
  23314=>"100110101",
  23315=>"010001111",
  23316=>"110001001",
  23317=>"100101111",
  23318=>"101011011",
  23319=>"111111010",
  23320=>"110011100",
  23321=>"101000110",
  23322=>"010010111",
  23323=>"100100001",
  23324=>"010011000",
  23325=>"100111111",
  23326=>"010101001",
  23327=>"001111011",
  23328=>"011000001",
  23329=>"000100001",
  23330=>"100001000",
  23331=>"000100010",
  23332=>"011001111",
  23333=>"001011000",
  23334=>"000111100",
  23335=>"111001111",
  23336=>"000010010",
  23337=>"001011101",
  23338=>"010001110",
  23339=>"010101111",
  23340=>"010011101",
  23341=>"111111110",
  23342=>"110101000",
  23343=>"100010000",
  23344=>"101010000",
  23345=>"100011001",
  23346=>"001001111",
  23347=>"010010100",
  23348=>"001000101",
  23349=>"110110111",
  23350=>"011111111",
  23351=>"000110100",
  23352=>"101110101",
  23353=>"011011101",
  23354=>"001101001",
  23355=>"011111101",
  23356=>"100100110",
  23357=>"111010001",
  23358=>"110111001",
  23359=>"000000110",
  23360=>"001000101",
  23361=>"000011001",
  23362=>"011101001",
  23363=>"101001011",
  23364=>"000010101",
  23365=>"101000001",
  23366=>"101111110",
  23367=>"111001111",
  23368=>"110001111",
  23369=>"010111101",
  23370=>"010101010",
  23371=>"101000101",
  23372=>"000011000",
  23373=>"010101110",
  23374=>"101100101",
  23375=>"011010101",
  23376=>"111000001",
  23377=>"011001001",
  23378=>"101101111",
  23379=>"011110011",
  23380=>"110111000",
  23381=>"101011011",
  23382=>"111111000",
  23383=>"111010001",
  23384=>"000110100",
  23385=>"101110001",
  23386=>"110100111",
  23387=>"101100111",
  23388=>"000110111",
  23389=>"010111001",
  23390=>"000010111",
  23391=>"101100110",
  23392=>"011111111",
  23393=>"010100100",
  23394=>"101001001",
  23395=>"101111100",
  23396=>"010110000",
  23397=>"000001000",
  23398=>"110110000",
  23399=>"010100101",
  23400=>"100000111",
  23401=>"000010111",
  23402=>"010011010",
  23403=>"000000101",
  23404=>"111101010",
  23405=>"000101001",
  23406=>"000011001",
  23407=>"111001111",
  23408=>"010101100",
  23409=>"100000101",
  23410=>"010111111",
  23411=>"111011011",
  23412=>"010000001",
  23413=>"000001100",
  23414=>"000001001",
  23415=>"111110000",
  23416=>"001001010",
  23417=>"000000111",
  23418=>"100100011",
  23419=>"001110010",
  23420=>"011010100",
  23421=>"111001101",
  23422=>"101111100",
  23423=>"001111011",
  23424=>"111000101",
  23425=>"001010111",
  23426=>"001100111",
  23427=>"101010110",
  23428=>"011011001",
  23429=>"010100100",
  23430=>"001111111",
  23431=>"110011111",
  23432=>"101001000",
  23433=>"101101100",
  23434=>"010111001",
  23435=>"101111001",
  23436=>"010100001",
  23437=>"100011111",
  23438=>"011110101",
  23439=>"000000000",
  23440=>"101101100",
  23441=>"101111001",
  23442=>"111000000",
  23443=>"100011111",
  23444=>"000010001",
  23445=>"110000000",
  23446=>"011111011",
  23447=>"100111001",
  23448=>"100111000",
  23449=>"101001110",
  23450=>"101110010",
  23451=>"100110101",
  23452=>"111100100",
  23453=>"110110000",
  23454=>"010000001",
  23455=>"011011011",
  23456=>"001101110",
  23457=>"010101100",
  23458=>"000110111",
  23459=>"010000111",
  23460=>"000110101",
  23461=>"101100001",
  23462=>"001001001",
  23463=>"111111011",
  23464=>"110000101",
  23465=>"100110111",
  23466=>"001001101",
  23467=>"100010000",
  23468=>"110111110",
  23469=>"000011111",
  23470=>"101000110",
  23471=>"101000110",
  23472=>"011111011",
  23473=>"111110111",
  23474=>"110000000",
  23475=>"111101000",
  23476=>"000010000",
  23477=>"110011011",
  23478=>"000010010",
  23479=>"101001000",
  23480=>"011000000",
  23481=>"010000000",
  23482=>"111011100",
  23483=>"011101000",
  23484=>"101101001",
  23485=>"010000001",
  23486=>"111000100",
  23487=>"000101100",
  23488=>"010010001",
  23489=>"001001001",
  23490=>"100110011",
  23491=>"111011111",
  23492=>"111010000",
  23493=>"101111011",
  23494=>"110010110",
  23495=>"001010100",
  23496=>"000110011",
  23497=>"110100101",
  23498=>"110100100",
  23499=>"010011000",
  23500=>"101100000",
  23501=>"011101011",
  23502=>"000100110",
  23503=>"001010001",
  23504=>"110111010",
  23505=>"110001110",
  23506=>"001110101",
  23507=>"110110001",
  23508=>"101100111",
  23509=>"001100100",
  23510=>"110111111",
  23511=>"011001100",
  23512=>"100001100",
  23513=>"010000011",
  23514=>"000110111",
  23515=>"000000001",
  23516=>"101100000",
  23517=>"010001011",
  23518=>"100111001",
  23519=>"000000010",
  23520=>"101101001",
  23521=>"101011111",
  23522=>"001010000",
  23523=>"100110111",
  23524=>"010110010",
  23525=>"011110110",
  23526=>"000011111",
  23527=>"100110101",
  23528=>"011101101",
  23529=>"010101010",
  23530=>"001100011",
  23531=>"110100010",
  23532=>"000110010",
  23533=>"101001000",
  23534=>"011011011",
  23535=>"001110100",
  23536=>"101101100",
  23537=>"101100110",
  23538=>"001000010",
  23539=>"111101101",
  23540=>"110110101",
  23541=>"100100100",
  23542=>"111111011",
  23543=>"101111100",
  23544=>"001001100",
  23545=>"011010001",
  23546=>"000001001",
  23547=>"100001001",
  23548=>"111110010",
  23549=>"101111010",
  23550=>"100100101",
  23551=>"000001101",
  23552=>"011111000",
  23553=>"000101111",
  23554=>"011100100",
  23555=>"101110111",
  23556=>"111000111",
  23557=>"110010111",
  23558=>"100000010",
  23559=>"111001001",
  23560=>"111010100",
  23561=>"011110100",
  23562=>"000011000",
  23563=>"010110101",
  23564=>"010100011",
  23565=>"011000110",
  23566=>"100100000",
  23567=>"010010100",
  23568=>"101011011",
  23569=>"000000101",
  23570=>"000010100",
  23571=>"011111101",
  23572=>"100000111",
  23573=>"010111001",
  23574=>"001011111",
  23575=>"101101110",
  23576=>"010110110",
  23577=>"111011000",
  23578=>"101001110",
  23579=>"100000100",
  23580=>"111110000",
  23581=>"111001010",
  23582=>"101110010",
  23583=>"101101111",
  23584=>"011010011",
  23585=>"010010110",
  23586=>"010111111",
  23587=>"001101000",
  23588=>"110110101",
  23589=>"000100111",
  23590=>"100100000",
  23591=>"010010001",
  23592=>"100010010",
  23593=>"110010001",
  23594=>"101001100",
  23595=>"001011110",
  23596=>"100100000",
  23597=>"011010011",
  23598=>"101111101",
  23599=>"010001100",
  23600=>"000000100",
  23601=>"010101000",
  23602=>"010110001",
  23603=>"010011111",
  23604=>"010111110",
  23605=>"010101001",
  23606=>"000000011",
  23607=>"001110010",
  23608=>"000100101",
  23609=>"101000100",
  23610=>"110011111",
  23611=>"011010101",
  23612=>"111101010",
  23613=>"111101100",
  23614=>"100101010",
  23615=>"001001001",
  23616=>"111000100",
  23617=>"000111000",
  23618=>"111111110",
  23619=>"011111011",
  23620=>"011001100",
  23621=>"000100001",
  23622=>"011100100",
  23623=>"001101110",
  23624=>"000111011",
  23625=>"001000101",
  23626=>"001000001",
  23627=>"010001000",
  23628=>"000100101",
  23629=>"000000011",
  23630=>"101001100",
  23631=>"010111110",
  23632=>"000001010",
  23633=>"101010000",
  23634=>"011100010",
  23635=>"011000001",
  23636=>"011011001",
  23637=>"011011101",
  23638=>"011001101",
  23639=>"000100001",
  23640=>"100101111",
  23641=>"000001100",
  23642=>"111010110",
  23643=>"100100000",
  23644=>"100101000",
  23645=>"101000010",
  23646=>"000000010",
  23647=>"110000100",
  23648=>"001010010",
  23649=>"001111110",
  23650=>"001111101",
  23651=>"001010000",
  23652=>"001010000",
  23653=>"010010000",
  23654=>"100000010",
  23655=>"111001011",
  23656=>"001100110",
  23657=>"001100000",
  23658=>"001101100",
  23659=>"110110101",
  23660=>"001001001",
  23661=>"000111010",
  23662=>"000111100",
  23663=>"111111001",
  23664=>"000000010",
  23665=>"011110111",
  23666=>"010101000",
  23667=>"110011011",
  23668=>"101010100",
  23669=>"100111001",
  23670=>"111011011",
  23671=>"100101100",
  23672=>"001101111",
  23673=>"110111100",
  23674=>"111000100",
  23675=>"010000010",
  23676=>"110101111",
  23677=>"011111000",
  23678=>"010100010",
  23679=>"110101110",
  23680=>"100000011",
  23681=>"101111011",
  23682=>"000101010",
  23683=>"100001010",
  23684=>"010000000",
  23685=>"001111001",
  23686=>"110001000",
  23687=>"111100110",
  23688=>"010011010",
  23689=>"111010001",
  23690=>"000010000",
  23691=>"101101011",
  23692=>"110110100",
  23693=>"000110010",
  23694=>"000101111",
  23695=>"000110011",
  23696=>"000101100",
  23697=>"000011101",
  23698=>"010101010",
  23699=>"011000011",
  23700=>"101100001",
  23701=>"101001111",
  23702=>"001111011",
  23703=>"110001100",
  23704=>"101101000",
  23705=>"011110011",
  23706=>"101111111",
  23707=>"001110000",
  23708=>"001010001",
  23709=>"011110111",
  23710=>"001110111",
  23711=>"000111100",
  23712=>"100110110",
  23713=>"111110111",
  23714=>"001010011",
  23715=>"111010100",
  23716=>"010011001",
  23717=>"000001100",
  23718=>"111101111",
  23719=>"001101110",
  23720=>"111000001",
  23721=>"100000011",
  23722=>"010110100",
  23723=>"100010011",
  23724=>"001110100",
  23725=>"000001001",
  23726=>"110011010",
  23727=>"100001010",
  23728=>"011101000",
  23729=>"100010101",
  23730=>"000100011",
  23731=>"011100101",
  23732=>"101110111",
  23733=>"110111110",
  23734=>"101101001",
  23735=>"111001001",
  23736=>"111110010",
  23737=>"101110100",
  23738=>"010011000",
  23739=>"000010111",
  23740=>"110110000",
  23741=>"001001100",
  23742=>"000011111",
  23743=>"100100011",
  23744=>"100110101",
  23745=>"110001111",
  23746=>"000101011",
  23747=>"010011100",
  23748=>"100111110",
  23749=>"000010011",
  23750=>"111001100",
  23751=>"010111000",
  23752=>"100011110",
  23753=>"001111000",
  23754=>"001011100",
  23755=>"001000101",
  23756=>"101001000",
  23757=>"011011010",
  23758=>"001100110",
  23759=>"111011100",
  23760=>"000001100",
  23761=>"011101110",
  23762=>"100010100",
  23763=>"100111011",
  23764=>"001000000",
  23765=>"010001101",
  23766=>"111100001",
  23767=>"101100110",
  23768=>"010110001",
  23769=>"110001001",
  23770=>"001000001",
  23771=>"010010110",
  23772=>"011110101",
  23773=>"011000100",
  23774=>"000010001",
  23775=>"100000010",
  23776=>"110100000",
  23777=>"011100000",
  23778=>"011010111",
  23779=>"001000000",
  23780=>"010000000",
  23781=>"001111100",
  23782=>"100011101",
  23783=>"100111010",
  23784=>"011000000",
  23785=>"100110101",
  23786=>"010111110",
  23787=>"011011100",
  23788=>"101101011",
  23789=>"111001110",
  23790=>"001000001",
  23791=>"110010110",
  23792=>"100000000",
  23793=>"010001000",
  23794=>"000000000",
  23795=>"100000111",
  23796=>"100001011",
  23797=>"110000100",
  23798=>"111100000",
  23799=>"011010001",
  23800=>"001001001",
  23801=>"001010111",
  23802=>"011101011",
  23803=>"101100100",
  23804=>"100000001",
  23805=>"101000011",
  23806=>"101111000",
  23807=>"111100110",
  23808=>"010110011",
  23809=>"111011111",
  23810=>"001100010",
  23811=>"111111010",
  23812=>"000010101",
  23813=>"101111101",
  23814=>"111000010",
  23815=>"111000010",
  23816=>"000000101",
  23817=>"110101001",
  23818=>"001100111",
  23819=>"110110011",
  23820=>"010011101",
  23821=>"010011011",
  23822=>"000011011",
  23823=>"111101100",
  23824=>"101000111",
  23825=>"011000110",
  23826=>"010011111",
  23827=>"100010101",
  23828=>"111001000",
  23829=>"101011010",
  23830=>"101100001",
  23831=>"110001000",
  23832=>"101011110",
  23833=>"111110101",
  23834=>"100100100",
  23835=>"110111011",
  23836=>"100100111",
  23837=>"011100100",
  23838=>"101010011",
  23839=>"111011011",
  23840=>"000100001",
  23841=>"000101011",
  23842=>"010000111",
  23843=>"101110111",
  23844=>"010010001",
  23845=>"100000001",
  23846=>"100001011",
  23847=>"010011011",
  23848=>"111001111",
  23849=>"100011101",
  23850=>"101010011",
  23851=>"010000011",
  23852=>"100110000",
  23853=>"010011000",
  23854=>"111011101",
  23855=>"001001001",
  23856=>"100110010",
  23857=>"110101100",
  23858=>"011001101",
  23859=>"011010010",
  23860=>"111111000",
  23861=>"000110010",
  23862=>"001110110",
  23863=>"111111110",
  23864=>"001110001",
  23865=>"010111011",
  23866=>"100000101",
  23867=>"010111001",
  23868=>"110000001",
  23869=>"011111111",
  23870=>"010000011",
  23871=>"000010010",
  23872=>"101100010",
  23873=>"011001001",
  23874=>"010100000",
  23875=>"011101101",
  23876=>"101000100",
  23877=>"001100001",
  23878=>"000111010",
  23879=>"000001101",
  23880=>"000100001",
  23881=>"100011000",
  23882=>"010110011",
  23883=>"101111100",
  23884=>"010000110",
  23885=>"100111100",
  23886=>"010101000",
  23887=>"111100011",
  23888=>"101011111",
  23889=>"001100111",
  23890=>"101111110",
  23891=>"100101101",
  23892=>"010011010",
  23893=>"010000110",
  23894=>"000000100",
  23895=>"010000011",
  23896=>"001010010",
  23897=>"001110111",
  23898=>"101011111",
  23899=>"100100000",
  23900=>"010001011",
  23901=>"000101111",
  23902=>"000011001",
  23903=>"101011011",
  23904=>"111001001",
  23905=>"100000010",
  23906=>"101011001",
  23907=>"100010000",
  23908=>"100100101",
  23909=>"011001111",
  23910=>"000111010",
  23911=>"010111000",
  23912=>"111100001",
  23913=>"110000101",
  23914=>"100001100",
  23915=>"100110111",
  23916=>"111001111",
  23917=>"011100010",
  23918=>"110001110",
  23919=>"111010001",
  23920=>"101111010",
  23921=>"010101010",
  23922=>"101111100",
  23923=>"101101110",
  23924=>"011000011",
  23925=>"010000010",
  23926=>"000100000",
  23927=>"000010000",
  23928=>"110110001",
  23929=>"100100001",
  23930=>"001010000",
  23931=>"111100100",
  23932=>"001110000",
  23933=>"110001010",
  23934=>"110000101",
  23935=>"010001010",
  23936=>"010100111",
  23937=>"110011110",
  23938=>"100010110",
  23939=>"111111011",
  23940=>"001111100",
  23941=>"110110100",
  23942=>"101110101",
  23943=>"011100110",
  23944=>"110010111",
  23945=>"100101101",
  23946=>"010101111",
  23947=>"011001100",
  23948=>"011000100",
  23949=>"101001001",
  23950=>"111100000",
  23951=>"001101111",
  23952=>"100010111",
  23953=>"011011101",
  23954=>"110000000",
  23955=>"111101101",
  23956=>"000011010",
  23957=>"111101011",
  23958=>"000100011",
  23959=>"110000100",
  23960=>"101100101",
  23961=>"100001000",
  23962=>"010101100",
  23963=>"000011000",
  23964=>"000010111",
  23965=>"111110110",
  23966=>"111111000",
  23967=>"000000010",
  23968=>"101011101",
  23969=>"000110010",
  23970=>"000101101",
  23971=>"000110101",
  23972=>"110101111",
  23973=>"100100000",
  23974=>"101110100",
  23975=>"110110000",
  23976=>"110001000",
  23977=>"100001010",
  23978=>"001101110",
  23979=>"000011010",
  23980=>"111000010",
  23981=>"101000010",
  23982=>"110111110",
  23983=>"110001010",
  23984=>"010010011",
  23985=>"011101010",
  23986=>"011110111",
  23987=>"100101001",
  23988=>"011110111",
  23989=>"110000110",
  23990=>"010110000",
  23991=>"101110010",
  23992=>"101011001",
  23993=>"001001000",
  23994=>"000101110",
  23995=>"000000010",
  23996=>"010000111",
  23997=>"001110010",
  23998=>"010110101",
  23999=>"110111010",
  24000=>"010100000",
  24001=>"011000010",
  24002=>"100001000",
  24003=>"001111111",
  24004=>"011000011",
  24005=>"000000001",
  24006=>"011001011",
  24007=>"101000000",
  24008=>"111001010",
  24009=>"101001011",
  24010=>"011010001",
  24011=>"110000011",
  24012=>"000010001",
  24013=>"100000011",
  24014=>"001101010",
  24015=>"111010001",
  24016=>"100010111",
  24017=>"111000001",
  24018=>"100100110",
  24019=>"100100111",
  24020=>"010001010",
  24021=>"110011000",
  24022=>"101110110",
  24023=>"000010010",
  24024=>"010001100",
  24025=>"111111100",
  24026=>"100100010",
  24027=>"100001110",
  24028=>"001101001",
  24029=>"000111110",
  24030=>"101110101",
  24031=>"111100101",
  24032=>"111011001",
  24033=>"100111011",
  24034=>"011101001",
  24035=>"011010110",
  24036=>"110111001",
  24037=>"110011010",
  24038=>"100100011",
  24039=>"100000011",
  24040=>"000010101",
  24041=>"001011100",
  24042=>"001010000",
  24043=>"110111100",
  24044=>"111101011",
  24045=>"110101101",
  24046=>"111100000",
  24047=>"010111110",
  24048=>"111001001",
  24049=>"101001110",
  24050=>"100110011",
  24051=>"100111100",
  24052=>"110001001",
  24053=>"011011001",
  24054=>"000000100",
  24055=>"101010001",
  24056=>"111011110",
  24057=>"101010100",
  24058=>"011111010",
  24059=>"101010011",
  24060=>"111011101",
  24061=>"111011100",
  24062=>"100000100",
  24063=>"001111000",
  24064=>"000111111",
  24065=>"011100011",
  24066=>"100101001",
  24067=>"010010110",
  24068=>"110111010",
  24069=>"111000111",
  24070=>"001001110",
  24071=>"100111001",
  24072=>"001001001",
  24073=>"011110111",
  24074=>"000100100",
  24075=>"100101000",
  24076=>"011010110",
  24077=>"010111101",
  24078=>"000010100",
  24079=>"100101001",
  24080=>"111001111",
  24081=>"001111111",
  24082=>"100000000",
  24083=>"001000011",
  24084=>"000001110",
  24085=>"111110101",
  24086=>"011100101",
  24087=>"110001101",
  24088=>"000010010",
  24089=>"110010010",
  24090=>"100101001",
  24091=>"001010010",
  24092=>"100010000",
  24093=>"000110100",
  24094=>"110010010",
  24095=>"111101001",
  24096=>"111011111",
  24097=>"101010000",
  24098=>"100111111",
  24099=>"110000101",
  24100=>"110000110",
  24101=>"000011010",
  24102=>"011001010",
  24103=>"111101100",
  24104=>"001001101",
  24105=>"011111110",
  24106=>"001110010",
  24107=>"011001000",
  24108=>"110011111",
  24109=>"111001111",
  24110=>"100010110",
  24111=>"001111001",
  24112=>"000000100",
  24113=>"000011110",
  24114=>"110100000",
  24115=>"010101100",
  24116=>"110100000",
  24117=>"100001000",
  24118=>"111010100",
  24119=>"010000100",
  24120=>"110011010",
  24121=>"010111111",
  24122=>"101011100",
  24123=>"011010111",
  24124=>"100101010",
  24125=>"000110000",
  24126=>"110110001",
  24127=>"101011010",
  24128=>"000100010",
  24129=>"101011111",
  24130=>"101110110",
  24131=>"011100010",
  24132=>"110010110",
  24133=>"011100101",
  24134=>"101111111",
  24135=>"111001000",
  24136=>"000011011",
  24137=>"010011101",
  24138=>"100111000",
  24139=>"101100000",
  24140=>"100100111",
  24141=>"001101011",
  24142=>"001111110",
  24143=>"110111111",
  24144=>"100010111",
  24145=>"111111100",
  24146=>"010110010",
  24147=>"001011001",
  24148=>"000111011",
  24149=>"000111000",
  24150=>"100100010",
  24151=>"001101101",
  24152=>"110011000",
  24153=>"000111000",
  24154=>"110111101",
  24155=>"001010001",
  24156=>"010001100",
  24157=>"101010011",
  24158=>"101001011",
  24159=>"100001110",
  24160=>"000000100",
  24161=>"001100111",
  24162=>"110110111",
  24163=>"100100111",
  24164=>"011010011",
  24165=>"011000110",
  24166=>"011100111",
  24167=>"000100011",
  24168=>"111110000",
  24169=>"111110100",
  24170=>"011100011",
  24171=>"000001011",
  24172=>"001101100",
  24173=>"011011011",
  24174=>"010000010",
  24175=>"111011011",
  24176=>"111011101",
  24177=>"000100100",
  24178=>"010101101",
  24179=>"110111010",
  24180=>"000111101",
  24181=>"010011011",
  24182=>"010111010",
  24183=>"000111000",
  24184=>"001010010",
  24185=>"111111011",
  24186=>"001101010",
  24187=>"101000000",
  24188=>"010111101",
  24189=>"100000101",
  24190=>"000111101",
  24191=>"101000110",
  24192=>"111001100",
  24193=>"010100101",
  24194=>"011000111",
  24195=>"111100000",
  24196=>"001101100",
  24197=>"110100101",
  24198=>"111011111",
  24199=>"000110011",
  24200=>"011111011",
  24201=>"000001101",
  24202=>"101111001",
  24203=>"001011011",
  24204=>"110101111",
  24205=>"100011010",
  24206=>"111101111",
  24207=>"010010000",
  24208=>"101111111",
  24209=>"000000001",
  24210=>"100011100",
  24211=>"001001001",
  24212=>"000111100",
  24213=>"110101001",
  24214=>"111100010",
  24215=>"010110010",
  24216=>"010010100",
  24217=>"000000111",
  24218=>"010010110",
  24219=>"010011110",
  24220=>"000011011",
  24221=>"111000100",
  24222=>"100101110",
  24223=>"001110010",
  24224=>"100110100",
  24225=>"001111010",
  24226=>"000101110",
  24227=>"011011011",
  24228=>"000001111",
  24229=>"010111011",
  24230=>"100000001",
  24231=>"000100011",
  24232=>"111010001",
  24233=>"010011111",
  24234=>"110111010",
  24235=>"100001101",
  24236=>"000011010",
  24237=>"100111110",
  24238=>"110100010",
  24239=>"111011111",
  24240=>"100000010",
  24241=>"111000011",
  24242=>"101110111",
  24243=>"101011011",
  24244=>"011110010",
  24245=>"101111011",
  24246=>"001000101",
  24247=>"101101010",
  24248=>"100010110",
  24249=>"010100000",
  24250=>"001010011",
  24251=>"110010010",
  24252=>"011011101",
  24253=>"000111100",
  24254=>"010110010",
  24255=>"100101111",
  24256=>"000000001",
  24257=>"110101110",
  24258=>"100010000",
  24259=>"110001000",
  24260=>"000110100",
  24261=>"110100111",
  24262=>"010110010",
  24263=>"001000101",
  24264=>"101111010",
  24265=>"001010010",
  24266=>"010100001",
  24267=>"010100100",
  24268=>"011100111",
  24269=>"101010100",
  24270=>"111110110",
  24271=>"011001111",
  24272=>"100100010",
  24273=>"100100110",
  24274=>"001000010",
  24275=>"000001001",
  24276=>"100110010",
  24277=>"000001011",
  24278=>"110011111",
  24279=>"001111011",
  24280=>"111111100",
  24281=>"110011011",
  24282=>"100110000",
  24283=>"010010001",
  24284=>"100011001",
  24285=>"010001000",
  24286=>"111011000",
  24287=>"001001101",
  24288=>"111111011",
  24289=>"000100100",
  24290=>"000111100",
  24291=>"011100101",
  24292=>"000011010",
  24293=>"111011111",
  24294=>"101000101",
  24295=>"101011111",
  24296=>"000101101",
  24297=>"110101000",
  24298=>"110110011",
  24299=>"100010111",
  24300=>"000010011",
  24301=>"100110001",
  24302=>"110010100",
  24303=>"001110100",
  24304=>"111000101",
  24305=>"000010011",
  24306=>"111110001",
  24307=>"000111100",
  24308=>"010100101",
  24309=>"101100111",
  24310=>"110111101",
  24311=>"111100110",
  24312=>"010011001",
  24313=>"001110010",
  24314=>"101001100",
  24315=>"000101010",
  24316=>"111110011",
  24317=>"110010100",
  24318=>"100110101",
  24319=>"000010011",
  24320=>"000010110",
  24321=>"110110001",
  24322=>"101111111",
  24323=>"100101000",
  24324=>"100110011",
  24325=>"111001001",
  24326=>"110100001",
  24327=>"100010110",
  24328=>"001011100",
  24329=>"100000010",
  24330=>"001100000",
  24331=>"111101001",
  24332=>"101011011",
  24333=>"101000000",
  24334=>"001010001",
  24335=>"010001110",
  24336=>"100010011",
  24337=>"010100010",
  24338=>"101000101",
  24339=>"000010111",
  24340=>"001011001",
  24341=>"100010101",
  24342=>"110010101",
  24343=>"111111001",
  24344=>"001101111",
  24345=>"101100111",
  24346=>"001000001",
  24347=>"010111010",
  24348=>"001100010",
  24349=>"010011000",
  24350=>"100000110",
  24351=>"101001010",
  24352=>"001110010",
  24353=>"111101000",
  24354=>"000000000",
  24355=>"000010100",
  24356=>"100100010",
  24357=>"001010000",
  24358=>"101111110",
  24359=>"011001110",
  24360=>"000100111",
  24361=>"100110001",
  24362=>"111001001",
  24363=>"110000011",
  24364=>"000000110",
  24365=>"101100001",
  24366=>"001101001",
  24367=>"111110100",
  24368=>"010110000",
  24369=>"101000011",
  24370=>"100010011",
  24371=>"010001011",
  24372=>"110011100",
  24373=>"011101101",
  24374=>"000100100",
  24375=>"111111111",
  24376=>"011100001",
  24377=>"011001100",
  24378=>"001011000",
  24379=>"001110001",
  24380=>"110001011",
  24381=>"010110001",
  24382=>"100110110",
  24383=>"001010001",
  24384=>"010000010",
  24385=>"010010011",
  24386=>"101011010",
  24387=>"101111011",
  24388=>"111100000",
  24389=>"011010111",
  24390=>"001011010",
  24391=>"011001101",
  24392=>"001001000",
  24393=>"010100110",
  24394=>"101101100",
  24395=>"010011000",
  24396=>"100000000",
  24397=>"000110010",
  24398=>"101110000",
  24399=>"100101010",
  24400=>"100001110",
  24401=>"011110001",
  24402=>"000001011",
  24403=>"100111011",
  24404=>"100010101",
  24405=>"110101011",
  24406=>"011001101",
  24407=>"111111110",
  24408=>"001001101",
  24409=>"001011000",
  24410=>"001101010",
  24411=>"101110100",
  24412=>"010001010",
  24413=>"101001111",
  24414=>"111111011",
  24415=>"111011010",
  24416=>"011011110",
  24417=>"110101011",
  24418=>"110100100",
  24419=>"100100001",
  24420=>"011100101",
  24421=>"010011000",
  24422=>"101011000",
  24423=>"111001010",
  24424=>"000110011",
  24425=>"001000000",
  24426=>"001011101",
  24427=>"100100000",
  24428=>"010110000",
  24429=>"111111010",
  24430=>"111011010",
  24431=>"111011010",
  24432=>"110101010",
  24433=>"011100000",
  24434=>"011110000",
  24435=>"010011110",
  24436=>"101100111",
  24437=>"000000011",
  24438=>"100000000",
  24439=>"100100101",
  24440=>"010101100",
  24441=>"101101101",
  24442=>"011101100",
  24443=>"110010110",
  24444=>"111111100",
  24445=>"000001110",
  24446=>"111100010",
  24447=>"011100001",
  24448=>"010000000",
  24449=>"000010001",
  24450=>"101111111",
  24451=>"011011011",
  24452=>"000001110",
  24453=>"011110101",
  24454=>"111011111",
  24455=>"000000111",
  24456=>"110110111",
  24457=>"000011000",
  24458=>"110100110",
  24459=>"010101010",
  24460=>"000111001",
  24461=>"101001110",
  24462=>"110111111",
  24463=>"011111011",
  24464=>"101100110",
  24465=>"010100111",
  24466=>"011010100",
  24467=>"100000001",
  24468=>"100010000",
  24469=>"000011101",
  24470=>"100111010",
  24471=>"111010110",
  24472=>"000011110",
  24473=>"010101111",
  24474=>"100110001",
  24475=>"101101110",
  24476=>"001111011",
  24477=>"111111101",
  24478=>"101000110",
  24479=>"011000011",
  24480=>"001110100",
  24481=>"100011000",
  24482=>"011010001",
  24483=>"010000110",
  24484=>"001111100",
  24485=>"111011101",
  24486=>"011000001",
  24487=>"100011001",
  24488=>"100001001",
  24489=>"101101111",
  24490=>"110111001",
  24491=>"101111111",
  24492=>"010100101",
  24493=>"010000001",
  24494=>"001100110",
  24495=>"000010001",
  24496=>"101000001",
  24497=>"111110110",
  24498=>"100111010",
  24499=>"001101011",
  24500=>"100110100",
  24501=>"111001001",
  24502=>"100111001",
  24503=>"011011000",
  24504=>"001001000",
  24505=>"000100010",
  24506=>"001010110",
  24507=>"000111101",
  24508=>"110010011",
  24509=>"110101000",
  24510=>"111100001",
  24511=>"101110110",
  24512=>"000000100",
  24513=>"110110111",
  24514=>"010101110",
  24515=>"011111100",
  24516=>"000010111",
  24517=>"010111010",
  24518=>"010101010",
  24519=>"010011101",
  24520=>"111001010",
  24521=>"000000010",
  24522=>"110001101",
  24523=>"011000110",
  24524=>"010010000",
  24525=>"111100100",
  24526=>"111100001",
  24527=>"001110010",
  24528=>"011011000",
  24529=>"110101111",
  24530=>"100110011",
  24531=>"111000101",
  24532=>"000001010",
  24533=>"001000111",
  24534=>"010001110",
  24535=>"100101000",
  24536=>"011001011",
  24537=>"111010101",
  24538=>"010111110",
  24539=>"000000011",
  24540=>"100010110",
  24541=>"000100011",
  24542=>"000000111",
  24543=>"111011100",
  24544=>"110100011",
  24545=>"010011011",
  24546=>"101000100",
  24547=>"010110110",
  24548=>"010110000",
  24549=>"000100001",
  24550=>"000010000",
  24551=>"111110111",
  24552=>"001101111",
  24553=>"111101000",
  24554=>"010000000",
  24555=>"000000011",
  24556=>"111101001",
  24557=>"100001110",
  24558=>"110000011",
  24559=>"011000001",
  24560=>"000100001",
  24561=>"100000111",
  24562=>"011000110",
  24563=>"010011011",
  24564=>"011110001",
  24565=>"111111000",
  24566=>"111111011",
  24567=>"111001000",
  24568=>"100100000",
  24569=>"010011001",
  24570=>"011001101",
  24571=>"000101000",
  24572=>"001111110",
  24573=>"101101000",
  24574=>"000001000",
  24575=>"000011011",
  24576=>"101001110",
  24577=>"100110011",
  24578=>"000101111",
  24579=>"100001001",
  24580=>"101110010",
  24581=>"011001000",
  24582=>"100100110",
  24583=>"011001001",
  24584=>"111110001",
  24585=>"010000101",
  24586=>"011110101",
  24587=>"100011101",
  24588=>"101101111",
  24589=>"011100010",
  24590=>"100011100",
  24591=>"010110101",
  24592=>"011111001",
  24593=>"011000101",
  24594=>"010011101",
  24595=>"111100011",
  24596=>"010010001",
  24597=>"001000010",
  24598=>"001111111",
  24599=>"100111011",
  24600=>"010000001",
  24601=>"100000100",
  24602=>"111000001",
  24603=>"101011111",
  24604=>"101011110",
  24605=>"011011010",
  24606=>"011111100",
  24607=>"010101010",
  24608=>"011110010",
  24609=>"000101101",
  24610=>"111010111",
  24611=>"111000111",
  24612=>"010101111",
  24613=>"100011001",
  24614=>"000000101",
  24615=>"100010000",
  24616=>"111100010",
  24617=>"000111000",
  24618=>"111010101",
  24619=>"110010010",
  24620=>"011010010",
  24621=>"111110110",
  24622=>"001000110",
  24623=>"111010110",
  24624=>"001110010",
  24625=>"001110011",
  24626=>"110001101",
  24627=>"001011101",
  24628=>"010101010",
  24629=>"110111110",
  24630=>"111110011",
  24631=>"110000111",
  24632=>"000001010",
  24633=>"011110001",
  24634=>"001111101",
  24635=>"010001000",
  24636=>"111111100",
  24637=>"100100100",
  24638=>"001010110",
  24639=>"101011010",
  24640=>"100100100",
  24641=>"010101001",
  24642=>"000100101",
  24643=>"001110010",
  24644=>"010100010",
  24645=>"011101101",
  24646=>"110101000",
  24647=>"000111000",
  24648=>"011010011",
  24649=>"101100010",
  24650=>"011101110",
  24651=>"101100110",
  24652=>"111010110",
  24653=>"010100011",
  24654=>"111011101",
  24655=>"101111101",
  24656=>"000110000",
  24657=>"101100101",
  24658=>"110110110",
  24659=>"011101011",
  24660=>"101110000",
  24661=>"010010001",
  24662=>"111100010",
  24663=>"001101001",
  24664=>"010010110",
  24665=>"000010100",
  24666=>"010010101",
  24667=>"001000011",
  24668=>"001011010",
  24669=>"001101110",
  24670=>"100011110",
  24671=>"001010111",
  24672=>"101001010",
  24673=>"100111000",
  24674=>"100101100",
  24675=>"000000101",
  24676=>"111001011",
  24677=>"101111110",
  24678=>"010101101",
  24679=>"100101000",
  24680=>"000010110",
  24681=>"110111000",
  24682=>"000001011",
  24683=>"100100100",
  24684=>"101001011",
  24685=>"001011110",
  24686=>"001010000",
  24687=>"011111111",
  24688=>"011000001",
  24689=>"000011000",
  24690=>"111100101",
  24691=>"111010100",
  24692=>"100100010",
  24693=>"000111010",
  24694=>"000001101",
  24695=>"000101101",
  24696=>"001000110",
  24697=>"011001100",
  24698=>"001000100",
  24699=>"000011001",
  24700=>"011000011",
  24701=>"100010011",
  24702=>"001000111",
  24703=>"111001001",
  24704=>"001000010",
  24705=>"010011001",
  24706=>"111100111",
  24707=>"011000111",
  24708=>"000000011",
  24709=>"000110010",
  24710=>"100000010",
  24711=>"000100011",
  24712=>"101001000",
  24713=>"110010111",
  24714=>"010101000",
  24715=>"000110011",
  24716=>"101101100",
  24717=>"010000100",
  24718=>"100001000",
  24719=>"110000100",
  24720=>"011101101",
  24721=>"110111110",
  24722=>"110001010",
  24723=>"111110111",
  24724=>"011010110",
  24725=>"011011110",
  24726=>"101000000",
  24727=>"010010110",
  24728=>"001011001",
  24729=>"101111110",
  24730=>"001010110",
  24731=>"010001100",
  24732=>"111000100",
  24733=>"000100101",
  24734=>"110000000",
  24735=>"001110101",
  24736=>"000110110",
  24737=>"001001101",
  24738=>"111010010",
  24739=>"000110100",
  24740=>"011010010",
  24741=>"000000010",
  24742=>"011000101",
  24743=>"000001000",
  24744=>"010001110",
  24745=>"001010000",
  24746=>"110000101",
  24747=>"001100011",
  24748=>"011111110",
  24749=>"111101001",
  24750=>"111100100",
  24751=>"100101011",
  24752=>"110000000",
  24753=>"101101011",
  24754=>"111010011",
  24755=>"110011100",
  24756=>"100001110",
  24757=>"000001000",
  24758=>"100101011",
  24759=>"101101000",
  24760=>"011001011",
  24761=>"001011010",
  24762=>"001010110",
  24763=>"101100111",
  24764=>"011111001",
  24765=>"011111011",
  24766=>"000100001",
  24767=>"110101011",
  24768=>"100010011",
  24769=>"100111101",
  24770=>"011011001",
  24771=>"010001110",
  24772=>"110110101",
  24773=>"000010001",
  24774=>"010000100",
  24775=>"011110100",
  24776=>"000100011",
  24777=>"010000001",
  24778=>"110100111",
  24779=>"010010010",
  24780=>"111100001",
  24781=>"101011110",
  24782=>"101001000",
  24783=>"111001011",
  24784=>"100010101",
  24785=>"110100101",
  24786=>"100100101",
  24787=>"000010010",
  24788=>"110111101",
  24789=>"001011101",
  24790=>"100010010",
  24791=>"000010111",
  24792=>"100110101",
  24793=>"010010010",
  24794=>"000100110",
  24795=>"001100111",
  24796=>"010100101",
  24797=>"101010000",
  24798=>"100101000",
  24799=>"111101111",
  24800=>"111011001",
  24801=>"011110000",
  24802=>"100110100",
  24803=>"010110101",
  24804=>"101011010",
  24805=>"011001110",
  24806=>"001001100",
  24807=>"100011001",
  24808=>"000001000",
  24809=>"011111000",
  24810=>"111001111",
  24811=>"011001101",
  24812=>"111100010",
  24813=>"000101111",
  24814=>"000110110",
  24815=>"011101111",
  24816=>"101110111",
  24817=>"000000101",
  24818=>"011000001",
  24819=>"000001111",
  24820=>"011101110",
  24821=>"001000110",
  24822=>"000011111",
  24823=>"000111110",
  24824=>"100101000",
  24825=>"110111100",
  24826=>"111010011",
  24827=>"000011110",
  24828=>"101010000",
  24829=>"100111111",
  24830=>"110101100",
  24831=>"111001110",
  24832=>"010110011",
  24833=>"100110110",
  24834=>"000101101",
  24835=>"000110101",
  24836=>"001111011",
  24837=>"100111000",
  24838=>"000000101",
  24839=>"110100000",
  24840=>"001010111",
  24841=>"011110011",
  24842=>"001001101",
  24843=>"100110100",
  24844=>"010001000",
  24845=>"001110101",
  24846=>"010001001",
  24847=>"110000010",
  24848=>"010111110",
  24849=>"000001100",
  24850=>"111110111",
  24851=>"100010100",
  24852=>"001000111",
  24853=>"101001110",
  24854=>"010111110",
  24855=>"111100110",
  24856=>"001101001",
  24857=>"011010011",
  24858=>"101100010",
  24859=>"010010001",
  24860=>"011010110",
  24861=>"010001001",
  24862=>"111010001",
  24863=>"000101111",
  24864=>"000110011",
  24865=>"011000100",
  24866=>"011001000",
  24867=>"011010110",
  24868=>"111001000",
  24869=>"111101001",
  24870=>"001000000",
  24871=>"100100100",
  24872=>"010001111",
  24873=>"101100111",
  24874=>"000011010",
  24875=>"010100010",
  24876=>"110010001",
  24877=>"101100111",
  24878=>"011001001",
  24879=>"000101010",
  24880=>"101101100",
  24881=>"011001010",
  24882=>"010011010",
  24883=>"000101011",
  24884=>"000000000",
  24885=>"011001101",
  24886=>"110000111",
  24887=>"010011000",
  24888=>"001100101",
  24889=>"000100100",
  24890=>"101011001",
  24891=>"111101101",
  24892=>"111000110",
  24893=>"111100001",
  24894=>"101001000",
  24895=>"000110110",
  24896=>"001100101",
  24897=>"110001011",
  24898=>"111111010",
  24899=>"001010011",
  24900=>"011100100",
  24901=>"011001101",
  24902=>"100011000",
  24903=>"010111111",
  24904=>"100011011",
  24905=>"111000110",
  24906=>"000101100",
  24907=>"111111010",
  24908=>"111011011",
  24909=>"110110011",
  24910=>"110000001",
  24911=>"010100111",
  24912=>"011100000",
  24913=>"000101110",
  24914=>"110001110",
  24915=>"000110101",
  24916=>"000111000",
  24917=>"011011101",
  24918=>"111100011",
  24919=>"110101110",
  24920=>"001000100",
  24921=>"100110100",
  24922=>"110101111",
  24923=>"001101001",
  24924=>"100000001",
  24925=>"100111110",
  24926=>"101111001",
  24927=>"010011111",
  24928=>"100110010",
  24929=>"001000111",
  24930=>"110110001",
  24931=>"011110010",
  24932=>"111000101",
  24933=>"101110010",
  24934=>"010010000",
  24935=>"001110101",
  24936=>"011110011",
  24937=>"000110101",
  24938=>"001010111",
  24939=>"000111101",
  24940=>"111110000",
  24941=>"101001111",
  24942=>"100111101",
  24943=>"100000111",
  24944=>"000010111",
  24945=>"110000001",
  24946=>"101111001",
  24947=>"001011010",
  24948=>"110001110",
  24949=>"110110000",
  24950=>"010001100",
  24951=>"000111100",
  24952=>"001101101",
  24953=>"000010100",
  24954=>"011101001",
  24955=>"001000001",
  24956=>"001101011",
  24957=>"011101100",
  24958=>"100000111",
  24959=>"010000111",
  24960=>"100111001",
  24961=>"011100100",
  24962=>"001011011",
  24963=>"011110101",
  24964=>"111111101",
  24965=>"010101100",
  24966=>"000010001",
  24967=>"000000110",
  24968=>"000110100",
  24969=>"000111101",
  24970=>"100111110",
  24971=>"101111010",
  24972=>"011101011",
  24973=>"011000010",
  24974=>"010111111",
  24975=>"001111111",
  24976=>"011000100",
  24977=>"111100010",
  24978=>"111100011",
  24979=>"000010110",
  24980=>"111000100",
  24981=>"001001011",
  24982=>"111101011",
  24983=>"000001110",
  24984=>"010111000",
  24985=>"001110001",
  24986=>"010111001",
  24987=>"101000110",
  24988=>"101100101",
  24989=>"011010110",
  24990=>"110110111",
  24991=>"010101000",
  24992=>"011100100",
  24993=>"101001011",
  24994=>"011110001",
  24995=>"001011111",
  24996=>"100100100",
  24997=>"110001011",
  24998=>"000001111",
  24999=>"010000010",
  25000=>"101011101",
  25001=>"001111011",
  25002=>"100010001",
  25003=>"000100100",
  25004=>"000001000",
  25005=>"001000000",
  25006=>"010011000",
  25007=>"000101101",
  25008=>"101100110",
  25009=>"110000101",
  25010=>"110100011",
  25011=>"111000011",
  25012=>"110100011",
  25013=>"110101000",
  25014=>"101111101",
  25015=>"111100011",
  25016=>"001000001",
  25017=>"001000010",
  25018=>"000000100",
  25019=>"000111011",
  25020=>"010101110",
  25021=>"100001111",
  25022=>"101101011",
  25023=>"010100111",
  25024=>"100100101",
  25025=>"100010110",
  25026=>"110001100",
  25027=>"111010101",
  25028=>"000011001",
  25029=>"010001010",
  25030=>"001000011",
  25031=>"110000000",
  25032=>"101000011",
  25033=>"011100010",
  25034=>"101110010",
  25035=>"010000111",
  25036=>"101110000",
  25037=>"010110010",
  25038=>"001100000",
  25039=>"111001000",
  25040=>"101001000",
  25041=>"111100111",
  25042=>"001010001",
  25043=>"000100101",
  25044=>"010001000",
  25045=>"000100111",
  25046=>"111110100",
  25047=>"010010000",
  25048=>"011110110",
  25049=>"101001000",
  25050=>"111101001",
  25051=>"010101111",
  25052=>"101000010",
  25053=>"110000010",
  25054=>"001000000",
  25055=>"000100110",
  25056=>"011101010",
  25057=>"100100101",
  25058=>"110111101",
  25059=>"011101101",
  25060=>"001111110",
  25061=>"111101110",
  25062=>"001000111",
  25063=>"101100000",
  25064=>"111111111",
  25065=>"111111010",
  25066=>"000000101",
  25067=>"111110100",
  25068=>"001011110",
  25069=>"001010010",
  25070=>"010100100",
  25071=>"000010010",
  25072=>"111001011",
  25073=>"011110011",
  25074=>"100111000",
  25075=>"000101000",
  25076=>"001111000",
  25077=>"111000011",
  25078=>"101000100",
  25079=>"101111110",
  25080=>"011001001",
  25081=>"011011010",
  25082=>"001011001",
  25083=>"110011000",
  25084=>"001010011",
  25085=>"010111001",
  25086=>"010100111",
  25087=>"000110010",
  25088=>"101011101",
  25089=>"100101100",
  25090=>"111101100",
  25091=>"001000001",
  25092=>"100101111",
  25093=>"111101001",
  25094=>"111101111",
  25095=>"011110110",
  25096=>"001010000",
  25097=>"110110111",
  25098=>"000110000",
  25099=>"000011001",
  25100=>"001100001",
  25101=>"100001110",
  25102=>"100101000",
  25103=>"011001100",
  25104=>"011001011",
  25105=>"011000100",
  25106=>"010110000",
  25107=>"001000001",
  25108=>"100101100",
  25109=>"010101010",
  25110=>"001101010",
  25111=>"011111001",
  25112=>"000010011",
  25113=>"100010001",
  25114=>"100111111",
  25115=>"000001000",
  25116=>"101000100",
  25117=>"001001001",
  25118=>"111001011",
  25119=>"011010000",
  25120=>"111010101",
  25121=>"111011111",
  25122=>"000000011",
  25123=>"101111110",
  25124=>"101011000",
  25125=>"100110101",
  25126=>"001011011",
  25127=>"100000101",
  25128=>"010000101",
  25129=>"001100110",
  25130=>"001110101",
  25131=>"100110101",
  25132=>"111010011",
  25133=>"100000000",
  25134=>"001011000",
  25135=>"010110101",
  25136=>"111111010",
  25137=>"111001101",
  25138=>"101111011",
  25139=>"010011101",
  25140=>"000010000",
  25141=>"011110101",
  25142=>"001110110",
  25143=>"000011100",
  25144=>"011010001",
  25145=>"010000100",
  25146=>"000001110",
  25147=>"011111110",
  25148=>"011101001",
  25149=>"100101111",
  25150=>"000101100",
  25151=>"111111111",
  25152=>"110100111",
  25153=>"010110111",
  25154=>"010001001",
  25155=>"010111001",
  25156=>"011001011",
  25157=>"100011010",
  25158=>"010010111",
  25159=>"001000000",
  25160=>"110001010",
  25161=>"001111101",
  25162=>"101011000",
  25163=>"101000001",
  25164=>"101010000",
  25165=>"110110010",
  25166=>"000011010",
  25167=>"001001000",
  25168=>"101100111",
  25169=>"001001100",
  25170=>"101111101",
  25171=>"010101011",
  25172=>"011001011",
  25173=>"010111000",
  25174=>"111111111",
  25175=>"010000110",
  25176=>"111110101",
  25177=>"000001110",
  25178=>"000000100",
  25179=>"101001111",
  25180=>"001010010",
  25181=>"011101111",
  25182=>"101110010",
  25183=>"111000100",
  25184=>"010011100",
  25185=>"010101110",
  25186=>"100111100",
  25187=>"000100101",
  25188=>"100101000",
  25189=>"001001111",
  25190=>"000000001",
  25191=>"101010011",
  25192=>"001010110",
  25193=>"100110101",
  25194=>"101111001",
  25195=>"111001110",
  25196=>"111100100",
  25197=>"010011101",
  25198=>"111100001",
  25199=>"011110111",
  25200=>"101111011",
  25201=>"110111110",
  25202=>"111111000",
  25203=>"000001011",
  25204=>"111010000",
  25205=>"001000100",
  25206=>"110101101",
  25207=>"101001100",
  25208=>"011010100",
  25209=>"001011101",
  25210=>"010010000",
  25211=>"101001011",
  25212=>"001000011",
  25213=>"101111101",
  25214=>"101101011",
  25215=>"101001001",
  25216=>"001101111",
  25217=>"011010100",
  25218=>"001011100",
  25219=>"100001100",
  25220=>"100011010",
  25221=>"011111001",
  25222=>"011111000",
  25223=>"000011000",
  25224=>"000010110",
  25225=>"110000100",
  25226=>"110110110",
  25227=>"010011101",
  25228=>"100010101",
  25229=>"111110011",
  25230=>"100000111",
  25231=>"000000000",
  25232=>"110011110",
  25233=>"111101101",
  25234=>"100110101",
  25235=>"011001100",
  25236=>"001000110",
  25237=>"011000001",
  25238=>"100001010",
  25239=>"110011011",
  25240=>"111010001",
  25241=>"110000111",
  25242=>"001000101",
  25243=>"111001101",
  25244=>"011011101",
  25245=>"110010000",
  25246=>"101110010",
  25247=>"110000101",
  25248=>"111011101",
  25249=>"000001110",
  25250=>"011111011",
  25251=>"011011010",
  25252=>"110010110",
  25253=>"000001010",
  25254=>"110001000",
  25255=>"000110011",
  25256=>"000011010",
  25257=>"110001010",
  25258=>"111111101",
  25259=>"000101010",
  25260=>"110010011",
  25261=>"001001101",
  25262=>"010010111",
  25263=>"110010011",
  25264=>"111101000",
  25265=>"110110100",
  25266=>"011111010",
  25267=>"000110010",
  25268=>"010010111",
  25269=>"110010001",
  25270=>"100010000",
  25271=>"100100011",
  25272=>"101000011",
  25273=>"110011101",
  25274=>"011111110",
  25275=>"111100011",
  25276=>"100100111",
  25277=>"001001110",
  25278=>"101100111",
  25279=>"000110011",
  25280=>"011011000",
  25281=>"111101001",
  25282=>"100101101",
  25283=>"100111111",
  25284=>"011011010",
  25285=>"100001011",
  25286=>"000100100",
  25287=>"010110101",
  25288=>"010001111",
  25289=>"100101100",
  25290=>"000011110",
  25291=>"101010100",
  25292=>"000110001",
  25293=>"011000011",
  25294=>"100000110",
  25295=>"110010110",
  25296=>"000100111",
  25297=>"110000011",
  25298=>"111110010",
  25299=>"101110000",
  25300=>"101000101",
  25301=>"000010001",
  25302=>"011101000",
  25303=>"010111001",
  25304=>"010001010",
  25305=>"111000111",
  25306=>"010001110",
  25307=>"101110011",
  25308=>"101001101",
  25309=>"110000111",
  25310=>"001000101",
  25311=>"000000100",
  25312=>"011110000",
  25313=>"101010011",
  25314=>"000111111",
  25315=>"000101101",
  25316=>"100010101",
  25317=>"001110001",
  25318=>"111110101",
  25319=>"101000000",
  25320=>"111110011",
  25321=>"000011000",
  25322=>"001011011",
  25323=>"001001000",
  25324=>"011101110",
  25325=>"110001100",
  25326=>"000011100",
  25327=>"001110011",
  25328=>"110100101",
  25329=>"011100000",
  25330=>"000110111",
  25331=>"100001101",
  25332=>"001101100",
  25333=>"111000001",
  25334=>"010010101",
  25335=>"011101100",
  25336=>"111011110",
  25337=>"110111101",
  25338=>"110000001",
  25339=>"001011001",
  25340=>"111110001",
  25341=>"000110000",
  25342=>"010010110",
  25343=>"000000110",
  25344=>"100101010",
  25345=>"001010111",
  25346=>"111001001",
  25347=>"001011111",
  25348=>"111011100",
  25349=>"000110010",
  25350=>"101110001",
  25351=>"010111110",
  25352=>"110010000",
  25353=>"110111100",
  25354=>"111010110",
  25355=>"000001101",
  25356=>"100110011",
  25357=>"111000000",
  25358=>"111110101",
  25359=>"001001111",
  25360=>"000001000",
  25361=>"010101011",
  25362=>"100010001",
  25363=>"001111001",
  25364=>"000110110",
  25365=>"100100100",
  25366=>"000001101",
  25367=>"001011101",
  25368=>"000000001",
  25369=>"100001100",
  25370=>"001110010",
  25371=>"011110000",
  25372=>"111011001",
  25373=>"010010110",
  25374=>"000001001",
  25375=>"011111001",
  25376=>"111110100",
  25377=>"111101111",
  25378=>"010011011",
  25379=>"111101010",
  25380=>"110100010",
  25381=>"111111001",
  25382=>"000000110",
  25383=>"010001110",
  25384=>"010111101",
  25385=>"011100100",
  25386=>"101100111",
  25387=>"111000000",
  25388=>"011000000",
  25389=>"101011101",
  25390=>"101101101",
  25391=>"101111000",
  25392=>"110010100",
  25393=>"111110000",
  25394=>"101111001",
  25395=>"100010000",
  25396=>"110111001",
  25397=>"001100111",
  25398=>"111010110",
  25399=>"001010111",
  25400=>"101011001",
  25401=>"000101100",
  25402=>"000000010",
  25403=>"011101100",
  25404=>"000101001",
  25405=>"110111110",
  25406=>"101001001",
  25407=>"000111010",
  25408=>"110101011",
  25409=>"110110111",
  25410=>"000100101",
  25411=>"100001010",
  25412=>"001110001",
  25413=>"000000001",
  25414=>"011001010",
  25415=>"100110011",
  25416=>"000110101",
  25417=>"101111010",
  25418=>"010001011",
  25419=>"000001101",
  25420=>"011110100",
  25421=>"011111001",
  25422=>"011000100",
  25423=>"001001000",
  25424=>"110100000",
  25425=>"011010100",
  25426=>"111001110",
  25427=>"001111011",
  25428=>"110111111",
  25429=>"111011101",
  25430=>"111001110",
  25431=>"110100100",
  25432=>"110101101",
  25433=>"001001101",
  25434=>"010110000",
  25435=>"101101100",
  25436=>"111001000",
  25437=>"110100011",
  25438=>"111111111",
  25439=>"001101001",
  25440=>"000001000",
  25441=>"111011000",
  25442=>"010101111",
  25443=>"010011011",
  25444=>"000001000",
  25445=>"010001100",
  25446=>"111000001",
  25447=>"111110100",
  25448=>"011111011",
  25449=>"111001101",
  25450=>"111111101",
  25451=>"010001000",
  25452=>"001000000",
  25453=>"111011011",
  25454=>"001101100",
  25455=>"110110011",
  25456=>"111100110",
  25457=>"100000010",
  25458=>"100111010",
  25459=>"001110010",
  25460=>"111001010",
  25461=>"101110010",
  25462=>"000010010",
  25463=>"110110101",
  25464=>"100101000",
  25465=>"100000010",
  25466=>"010010110",
  25467=>"100010100",
  25468=>"011111000",
  25469=>"110101011",
  25470=>"111111111",
  25471=>"011100010",
  25472=>"010111100",
  25473=>"100011100",
  25474=>"010100110",
  25475=>"101101010",
  25476=>"001011001",
  25477=>"110110000",
  25478=>"001011010",
  25479=>"011010000",
  25480=>"011101100",
  25481=>"101101111",
  25482=>"100101100",
  25483=>"011111001",
  25484=>"101110011",
  25485=>"010100001",
  25486=>"110101110",
  25487=>"111101111",
  25488=>"000011000",
  25489=>"100000001",
  25490=>"000011100",
  25491=>"111000101",
  25492=>"110111000",
  25493=>"101000111",
  25494=>"011000000",
  25495=>"101110011",
  25496=>"100010100",
  25497=>"011101110",
  25498=>"001110010",
  25499=>"111111111",
  25500=>"010010001",
  25501=>"001001001",
  25502=>"010101000",
  25503=>"001110101",
  25504=>"111111110",
  25505=>"110001100",
  25506=>"011010111",
  25507=>"001110010",
  25508=>"101001111",
  25509=>"010100100",
  25510=>"111001011",
  25511=>"110010010",
  25512=>"001011100",
  25513=>"010000110",
  25514=>"000011001",
  25515=>"111101110",
  25516=>"000000001",
  25517=>"100011011",
  25518=>"010111000",
  25519=>"011001101",
  25520=>"010100010",
  25521=>"111011111",
  25522=>"100101100",
  25523=>"000010101",
  25524=>"011110110",
  25525=>"010000000",
  25526=>"011000001",
  25527=>"111101010",
  25528=>"000101000",
  25529=>"000101111",
  25530=>"001111101",
  25531=>"001111110",
  25532=>"110000101",
  25533=>"011001010",
  25534=>"101111111",
  25535=>"000001111",
  25536=>"011111011",
  25537=>"011011111",
  25538=>"010100101",
  25539=>"100011011",
  25540=>"010000101",
  25541=>"100111101",
  25542=>"000111000",
  25543=>"111011001",
  25544=>"100000001",
  25545=>"100000100",
  25546=>"001010110",
  25547=>"100000011",
  25548=>"110010001",
  25549=>"001010011",
  25550=>"011000100",
  25551=>"001111010",
  25552=>"101010011",
  25553=>"000110000",
  25554=>"110000001",
  25555=>"001100011",
  25556=>"010111011",
  25557=>"101101101",
  25558=>"101111100",
  25559=>"110111100",
  25560=>"000110101",
  25561=>"000101101",
  25562=>"100010001",
  25563=>"100101101",
  25564=>"010001001",
  25565=>"010000010",
  25566=>"000011100",
  25567=>"111100001",
  25568=>"111100101",
  25569=>"000010101",
  25570=>"001101010",
  25571=>"110000000",
  25572=>"011001101",
  25573=>"100000000",
  25574=>"011011100",
  25575=>"100000110",
  25576=>"110111111",
  25577=>"100111100",
  25578=>"110111000",
  25579=>"010011100",
  25580=>"010000100",
  25581=>"100100010",
  25582=>"000000011",
  25583=>"110111100",
  25584=>"011101100",
  25585=>"101110010",
  25586=>"100011011",
  25587=>"011000110",
  25588=>"101100101",
  25589=>"101011000",
  25590=>"000101010",
  25591=>"000101110",
  25592=>"000001011",
  25593=>"101001010",
  25594=>"000001000",
  25595=>"101010100",
  25596=>"100011111",
  25597=>"100010010",
  25598=>"111011100",
  25599=>"010101101",
  25600=>"101001000",
  25601=>"000001111",
  25602=>"001101000",
  25603=>"000111011",
  25604=>"110011000",
  25605=>"011101100",
  25606=>"000111001",
  25607=>"011010010",
  25608=>"000000000",
  25609=>"101110111",
  25610=>"011000000",
  25611=>"110110011",
  25612=>"011110001",
  25613=>"000010001",
  25614=>"101010000",
  25615=>"001011000",
  25616=>"000100101",
  25617=>"110010011",
  25618=>"100111110",
  25619=>"010101000",
  25620=>"000000000",
  25621=>"101101111",
  25622=>"111011111",
  25623=>"001010101",
  25624=>"011001011",
  25625=>"011100011",
  25626=>"001110100",
  25627=>"101100100",
  25628=>"001110011",
  25629=>"010010110",
  25630=>"000000111",
  25631=>"001000000",
  25632=>"101001100",
  25633=>"100000110",
  25634=>"110111010",
  25635=>"110010111",
  25636=>"010110100",
  25637=>"010111111",
  25638=>"100100101",
  25639=>"011101111",
  25640=>"011110111",
  25641=>"111000111",
  25642=>"111011011",
  25643=>"100111011",
  25644=>"001000001",
  25645=>"001100000",
  25646=>"111010101",
  25647=>"110001011",
  25648=>"100001000",
  25649=>"010111011",
  25650=>"000011100",
  25651=>"000000111",
  25652=>"111110000",
  25653=>"100010010",
  25654=>"111100010",
  25655=>"110001001",
  25656=>"100010000",
  25657=>"000011010",
  25658=>"010100110",
  25659=>"110010110",
  25660=>"001001010",
  25661=>"011001000",
  25662=>"001011100",
  25663=>"010010001",
  25664=>"110000000",
  25665=>"101101101",
  25666=>"010011001",
  25667=>"100100000",
  25668=>"111001101",
  25669=>"111000000",
  25670=>"010010101",
  25671=>"111101001",
  25672=>"010100010",
  25673=>"100110000",
  25674=>"111000000",
  25675=>"110110011",
  25676=>"001000100",
  25677=>"000001000",
  25678=>"000101010",
  25679=>"100000010",
  25680=>"011011101",
  25681=>"011001110",
  25682=>"110001011",
  25683=>"111000111",
  25684=>"100001011",
  25685=>"111010111",
  25686=>"000000110",
  25687=>"001101100",
  25688=>"110000111",
  25689=>"101000110",
  25690=>"100001001",
  25691=>"100010000",
  25692=>"011001000",
  25693=>"011000101",
  25694=>"010110110",
  25695=>"100010001",
  25696=>"001001010",
  25697=>"001000001",
  25698=>"101101001",
  25699=>"111110111",
  25700=>"001000101",
  25701=>"001011101",
  25702=>"000011100",
  25703=>"000100010",
  25704=>"011101001",
  25705=>"111000111",
  25706=>"000000101",
  25707=>"101000101",
  25708=>"111001111",
  25709=>"000000010",
  25710=>"100100001",
  25711=>"110111000",
  25712=>"111100010",
  25713=>"110101101",
  25714=>"011000010",
  25715=>"000001000",
  25716=>"000101101",
  25717=>"000111111",
  25718=>"111110100",
  25719=>"101000111",
  25720=>"011010001",
  25721=>"100111110",
  25722=>"110110011",
  25723=>"101011110",
  25724=>"100010000",
  25725=>"000100101",
  25726=>"011000001",
  25727=>"101101000",
  25728=>"111100010",
  25729=>"111101001",
  25730=>"111011101",
  25731=>"010100100",
  25732=>"100101101",
  25733=>"000100100",
  25734=>"100111110",
  25735=>"101111011",
  25736=>"011010110",
  25737=>"101111000",
  25738=>"000011111",
  25739=>"100000101",
  25740=>"110001001",
  25741=>"010011000",
  25742=>"010111011",
  25743=>"001001100",
  25744=>"111001011",
  25745=>"001101010",
  25746=>"111010010",
  25747=>"111000110",
  25748=>"111000100",
  25749=>"111111100",
  25750=>"000111010",
  25751=>"010110011",
  25752=>"001010010",
  25753=>"100011101",
  25754=>"111111101",
  25755=>"001111101",
  25756=>"110000111",
  25757=>"000111100",
  25758=>"100101001",
  25759=>"000011110",
  25760=>"001000001",
  25761=>"011111010",
  25762=>"001111011",
  25763=>"000111111",
  25764=>"001000000",
  25765=>"000000001",
  25766=>"101000110",
  25767=>"000010001",
  25768=>"101111101",
  25769=>"001110101",
  25770=>"010001011",
  25771=>"110011000",
  25772=>"100100000",
  25773=>"101011100",
  25774=>"100001111",
  25775=>"010101110",
  25776=>"011100011",
  25777=>"111100110",
  25778=>"101010001",
  25779=>"010100110",
  25780=>"100011011",
  25781=>"110111110",
  25782=>"101000001",
  25783=>"010100100",
  25784=>"110000101",
  25785=>"010011001",
  25786=>"111111000",
  25787=>"000101010",
  25788=>"000010000",
  25789=>"101010011",
  25790=>"100001000",
  25791=>"011010111",
  25792=>"010001100",
  25793=>"010011110",
  25794=>"100101111",
  25795=>"111110110",
  25796=>"001101010",
  25797=>"110100101",
  25798=>"101010100",
  25799=>"011100011",
  25800=>"000111100",
  25801=>"001101100",
  25802=>"101001101",
  25803=>"011101011",
  25804=>"010111011",
  25805=>"001101101",
  25806=>"001000011",
  25807=>"110100110",
  25808=>"011100011",
  25809=>"001011010",
  25810=>"100111011",
  25811=>"011011001",
  25812=>"111101001",
  25813=>"111011001",
  25814=>"100111101",
  25815=>"011110010",
  25816=>"000000100",
  25817=>"111111001",
  25818=>"011010110",
  25819=>"110001101",
  25820=>"000011010",
  25821=>"000010110",
  25822=>"001001000",
  25823=>"111001100",
  25824=>"000100001",
  25825=>"001000000",
  25826=>"001001111",
  25827=>"000010010",
  25828=>"111110111",
  25829=>"110100011",
  25830=>"011010000",
  25831=>"011110100",
  25832=>"011111101",
  25833=>"010111110",
  25834=>"100111001",
  25835=>"000101110",
  25836=>"011010000",
  25837=>"011010101",
  25838=>"101010000",
  25839=>"001110011",
  25840=>"100100111",
  25841=>"100011010",
  25842=>"011101110",
  25843=>"100110000",
  25844=>"101011101",
  25845=>"000110000",
  25846=>"100000111",
  25847=>"110100000",
  25848=>"000101010",
  25849=>"000100110",
  25850=>"100101010",
  25851=>"100100001",
  25852=>"000101011",
  25853=>"111101010",
  25854=>"011011000",
  25855=>"110000101",
  25856=>"111110110",
  25857=>"000001110",
  25858=>"101111101",
  25859=>"001100110",
  25860=>"101110111",
  25861=>"111000010",
  25862=>"110011100",
  25863=>"100011010",
  25864=>"001001111",
  25865=>"111100011",
  25866=>"110010000",
  25867=>"100011010",
  25868=>"111001100",
  25869=>"010101011",
  25870=>"111010010",
  25871=>"001011000",
  25872=>"000001000",
  25873=>"111011110",
  25874=>"001001010",
  25875=>"111011000",
  25876=>"001110111",
  25877=>"010101000",
  25878=>"110000100",
  25879=>"110001001",
  25880=>"111001111",
  25881=>"001000001",
  25882=>"100101100",
  25883=>"110001100",
  25884=>"000000110",
  25885=>"011111001",
  25886=>"101011110",
  25887=>"010001000",
  25888=>"101001100",
  25889=>"000001000",
  25890=>"110100010",
  25891=>"011001010",
  25892=>"111011100",
  25893=>"100100110",
  25894=>"101011111",
  25895=>"100011111",
  25896=>"111110000",
  25897=>"100101110",
  25898=>"000000010",
  25899=>"010011001",
  25900=>"011100010",
  25901=>"111000000",
  25902=>"110110010",
  25903=>"101000001",
  25904=>"100111010",
  25905=>"000110111",
  25906=>"111011000",
  25907=>"111101011",
  25908=>"000010100",
  25909=>"100101101",
  25910=>"111010011",
  25911=>"111101111",
  25912=>"000000001",
  25913=>"010010011",
  25914=>"100001011",
  25915=>"000000011",
  25916=>"000000001",
  25917=>"101011011",
  25918=>"100111000",
  25919=>"110111111",
  25920=>"101110010",
  25921=>"100010011",
  25922=>"111110100",
  25923=>"000110101",
  25924=>"011001011",
  25925=>"111000001",
  25926=>"101000000",
  25927=>"000001001",
  25928=>"000100001",
  25929=>"111101000",
  25930=>"001001111",
  25931=>"000001111",
  25932=>"001110010",
  25933=>"010101000",
  25934=>"100101010",
  25935=>"111111011",
  25936=>"001010100",
  25937=>"011101100",
  25938=>"000110111",
  25939=>"011000101",
  25940=>"110001100",
  25941=>"100011001",
  25942=>"110101001",
  25943=>"000110101",
  25944=>"001010110",
  25945=>"001111101",
  25946=>"000000010",
  25947=>"111011001",
  25948=>"011101111",
  25949=>"001011001",
  25950=>"101001110",
  25951=>"010110010",
  25952=>"010111000",
  25953=>"011100100",
  25954=>"111101010",
  25955=>"110101111",
  25956=>"101100001",
  25957=>"010010000",
  25958=>"101011010",
  25959=>"011001011",
  25960=>"111001000",
  25961=>"111110110",
  25962=>"101101111",
  25963=>"010010011",
  25964=>"000101000",
  25965=>"011011010",
  25966=>"101011110",
  25967=>"000001011",
  25968=>"101011111",
  25969=>"110011100",
  25970=>"110010011",
  25971=>"010010110",
  25972=>"100000100",
  25973=>"101001100",
  25974=>"111010111",
  25975=>"010001110",
  25976=>"010001011",
  25977=>"100111000",
  25978=>"000001010",
  25979=>"110110111",
  25980=>"100010010",
  25981=>"000111111",
  25982=>"011110101",
  25983=>"001101110",
  25984=>"011011100",
  25985=>"010001001",
  25986=>"110110111",
  25987=>"001010111",
  25988=>"111111111",
  25989=>"100011101",
  25990=>"100100011",
  25991=>"111000001",
  25992=>"011110101",
  25993=>"110110011",
  25994=>"011101011",
  25995=>"111111010",
  25996=>"010000110",
  25997=>"110100011",
  25998=>"100011100",
  25999=>"010011101",
  26000=>"001001101",
  26001=>"001100010",
  26002=>"111010000",
  26003=>"111101100",
  26004=>"010010011",
  26005=>"010011110",
  26006=>"010111000",
  26007=>"101000110",
  26008=>"100010010",
  26009=>"110010101",
  26010=>"000100011",
  26011=>"111001110",
  26012=>"110011001",
  26013=>"000001000",
  26014=>"101001011",
  26015=>"101000000",
  26016=>"110000000",
  26017=>"010110000",
  26018=>"001100001",
  26019=>"011000001",
  26020=>"100110100",
  26021=>"110111011",
  26022=>"000010011",
  26023=>"110110110",
  26024=>"010010111",
  26025=>"011000110",
  26026=>"110000101",
  26027=>"100100011",
  26028=>"111010101",
  26029=>"000100101",
  26030=>"110111111",
  26031=>"101000010",
  26032=>"000011101",
  26033=>"010110000",
  26034=>"000010011",
  26035=>"000101000",
  26036=>"010010111",
  26037=>"110000001",
  26038=>"001101111",
  26039=>"101110010",
  26040=>"100010011",
  26041=>"001010000",
  26042=>"000100000",
  26043=>"111110110",
  26044=>"101010000",
  26045=>"001101111",
  26046=>"000000000",
  26047=>"010100110",
  26048=>"110110010",
  26049=>"010010001",
  26050=>"100101110",
  26051=>"001000011",
  26052=>"101000001",
  26053=>"000010001",
  26054=>"001111111",
  26055=>"000110101",
  26056=>"110001100",
  26057=>"001000011",
  26058=>"010111111",
  26059=>"001101001",
  26060=>"111101100",
  26061=>"101011111",
  26062=>"001001101",
  26063=>"000110100",
  26064=>"001111110",
  26065=>"010110010",
  26066=>"011001001",
  26067=>"011101011",
  26068=>"000110110",
  26069=>"000101011",
  26070=>"110101100",
  26071=>"111010101",
  26072=>"100100111",
  26073=>"010010100",
  26074=>"001010010",
  26075=>"101100010",
  26076=>"110100111",
  26077=>"100010001",
  26078=>"111101111",
  26079=>"111110000",
  26080=>"100001110",
  26081=>"111100000",
  26082=>"011101100",
  26083=>"111111100",
  26084=>"111010101",
  26085=>"101010000",
  26086=>"100001001",
  26087=>"010011100",
  26088=>"011110011",
  26089=>"111110000",
  26090=>"001110110",
  26091=>"110111000",
  26092=>"000010010",
  26093=>"110110101",
  26094=>"000001111",
  26095=>"011001001",
  26096=>"110100100",
  26097=>"101000101",
  26098=>"001100000",
  26099=>"011111001",
  26100=>"110100011",
  26101=>"110010101",
  26102=>"011111111",
  26103=>"100110111",
  26104=>"001110010",
  26105=>"001010110",
  26106=>"010110010",
  26107=>"101000000",
  26108=>"000011011",
  26109=>"011111111",
  26110=>"111010001",
  26111=>"010001111",
  26112=>"011100111",
  26113=>"000100101",
  26114=>"001010111",
  26115=>"000110100",
  26116=>"100111101",
  26117=>"000101100",
  26118=>"110100001",
  26119=>"010111100",
  26120=>"001001100",
  26121=>"101111111",
  26122=>"011010100",
  26123=>"111111000",
  26124=>"110001100",
  26125=>"101000101",
  26126=>"001000100",
  26127=>"101100000",
  26128=>"110010111",
  26129=>"111101011",
  26130=>"111010100",
  26131=>"011010101",
  26132=>"001101100",
  26133=>"010010011",
  26134=>"011110001",
  26135=>"110101110",
  26136=>"110101110",
  26137=>"111011010",
  26138=>"110010100",
  26139=>"001001011",
  26140=>"101100100",
  26141=>"001010100",
  26142=>"111101100",
  26143=>"001100010",
  26144=>"011011101",
  26145=>"001101011",
  26146=>"010001011",
  26147=>"000101001",
  26148=>"001110110",
  26149=>"111101100",
  26150=>"100010100",
  26151=>"001100101",
  26152=>"100000010",
  26153=>"101101010",
  26154=>"000110000",
  26155=>"001000100",
  26156=>"101000110",
  26157=>"011001011",
  26158=>"011000101",
  26159=>"001010000",
  26160=>"111101100",
  26161=>"101001001",
  26162=>"111011100",
  26163=>"101111111",
  26164=>"110110110",
  26165=>"100011110",
  26166=>"110011010",
  26167=>"111010111",
  26168=>"000101110",
  26169=>"100101110",
  26170=>"011101010",
  26171=>"011011100",
  26172=>"001110100",
  26173=>"001100101",
  26174=>"011010101",
  26175=>"110111101",
  26176=>"100100001",
  26177=>"100101011",
  26178=>"011000100",
  26179=>"001011010",
  26180=>"100000001",
  26181=>"100000001",
  26182=>"001001001",
  26183=>"010101110",
  26184=>"010111001",
  26185=>"110010101",
  26186=>"110110011",
  26187=>"010000100",
  26188=>"001111001",
  26189=>"000010100",
  26190=>"010110000",
  26191=>"100010100",
  26192=>"111010100",
  26193=>"010001111",
  26194=>"101000011",
  26195=>"000101001",
  26196=>"010100100",
  26197=>"100000101",
  26198=>"000111001",
  26199=>"111011101",
  26200=>"101011011",
  26201=>"010011011",
  26202=>"010010010",
  26203=>"010011111",
  26204=>"000000000",
  26205=>"010101001",
  26206=>"000001100",
  26207=>"011100000",
  26208=>"000100100",
  26209=>"000011011",
  26210=>"010011111",
  26211=>"111000001",
  26212=>"100111000",
  26213=>"111100110",
  26214=>"001010110",
  26215=>"010001000",
  26216=>"001110101",
  26217=>"100011111",
  26218=>"010110011",
  26219=>"101011100",
  26220=>"101010001",
  26221=>"110100000",
  26222=>"000010110",
  26223=>"111001011",
  26224=>"001001011",
  26225=>"100100101",
  26226=>"001111000",
  26227=>"100000000",
  26228=>"101101110",
  26229=>"110100100",
  26230=>"111111101",
  26231=>"100101011",
  26232=>"111111011",
  26233=>"110100001",
  26234=>"011111100",
  26235=>"000001001",
  26236=>"111000111",
  26237=>"101101000",
  26238=>"011000010",
  26239=>"011000111",
  26240=>"111000001",
  26241=>"111011101",
  26242=>"111000001",
  26243=>"101101111",
  26244=>"111110010",
  26245=>"100101110",
  26246=>"101100110",
  26247=>"010000110",
  26248=>"000011110",
  26249=>"000100100",
  26250=>"110001101",
  26251=>"001001011",
  26252=>"000011001",
  26253=>"110010010",
  26254=>"000011111",
  26255=>"010100000",
  26256=>"100110101",
  26257=>"111111010",
  26258=>"101111011",
  26259=>"101110110",
  26260=>"110101000",
  26261=>"110101111",
  26262=>"100010100",
  26263=>"010110101",
  26264=>"111000101",
  26265=>"011101100",
  26266=>"000100110",
  26267=>"011100111",
  26268=>"000110100",
  26269=>"000011100",
  26270=>"010011000",
  26271=>"000000111",
  26272=>"100000111",
  26273=>"000100111",
  26274=>"110001011",
  26275=>"111110101",
  26276=>"110011101",
  26277=>"000000001",
  26278=>"011010100",
  26279=>"100000101",
  26280=>"110011111",
  26281=>"101000100",
  26282=>"001100010",
  26283=>"111110111",
  26284=>"001101100",
  26285=>"100110101",
  26286=>"101011001",
  26287=>"001010110",
  26288=>"101010010",
  26289=>"100001011",
  26290=>"111101110",
  26291=>"111110111",
  26292=>"101100011",
  26293=>"001001111",
  26294=>"100110111",
  26295=>"100101101",
  26296=>"110101011",
  26297=>"100111011",
  26298=>"100101000",
  26299=>"110010101",
  26300=>"110011101",
  26301=>"111000001",
  26302=>"101110000",
  26303=>"100110001",
  26304=>"010000000",
  26305=>"100001101",
  26306=>"000000101",
  26307=>"100101110",
  26308=>"001011101",
  26309=>"000000011",
  26310=>"110111100",
  26311=>"101001011",
  26312=>"110000000",
  26313=>"111000011",
  26314=>"110001111",
  26315=>"111111100",
  26316=>"100001111",
  26317=>"011110011",
  26318=>"011001000",
  26319=>"011111101",
  26320=>"110110010",
  26321=>"010101110",
  26322=>"010000101",
  26323=>"010011001",
  26324=>"001111101",
  26325=>"111000111",
  26326=>"000000000",
  26327=>"000001100",
  26328=>"000000000",
  26329=>"100001111",
  26330=>"010111001",
  26331=>"110100000",
  26332=>"110001100",
  26333=>"010001001",
  26334=>"101111111",
  26335=>"001100010",
  26336=>"000110111",
  26337=>"001001001",
  26338=>"100001011",
  26339=>"010111000",
  26340=>"110001000",
  26341=>"001111000",
  26342=>"011010110",
  26343=>"010100100",
  26344=>"110010110",
  26345=>"111110010",
  26346=>"101110000",
  26347=>"000000101",
  26348=>"010100110",
  26349=>"100011110",
  26350=>"111001111",
  26351=>"000000000",
  26352=>"110111110",
  26353=>"101101000",
  26354=>"001000001",
  26355=>"010001000",
  26356=>"101010010",
  26357=>"101110101",
  26358=>"001001000",
  26359=>"011111111",
  26360=>"100000010",
  26361=>"100101101",
  26362=>"111110011",
  26363=>"100001010",
  26364=>"111100101",
  26365=>"101011001",
  26366=>"110101101",
  26367=>"101101111",
  26368=>"110000010",
  26369=>"110011010",
  26370=>"010101001",
  26371=>"111000001",
  26372=>"111111110",
  26373=>"000001111",
  26374=>"100011100",
  26375=>"110011110",
  26376=>"001001011",
  26377=>"011111001",
  26378=>"011100100",
  26379=>"100001000",
  26380=>"010011111",
  26381=>"111111010",
  26382=>"101001001",
  26383=>"110110101",
  26384=>"101000001",
  26385=>"001010101",
  26386=>"001000000",
  26387=>"100111101",
  26388=>"010010010",
  26389=>"111000100",
  26390=>"010111100",
  26391=>"011110001",
  26392=>"101001001",
  26393=>"001011100",
  26394=>"000000011",
  26395=>"011101110",
  26396=>"110001011",
  26397=>"100000010",
  26398=>"010010010",
  26399=>"100001010",
  26400=>"111011110",
  26401=>"000010100",
  26402=>"001100100",
  26403=>"101100100",
  26404=>"111110010",
  26405=>"010011000",
  26406=>"001010111",
  26407=>"001000000",
  26408=>"110111101",
  26409=>"100110010",
  26410=>"011100111",
  26411=>"001010000",
  26412=>"100011000",
  26413=>"000110111",
  26414=>"000101110",
  26415=>"001010010",
  26416=>"110001001",
  26417=>"010101000",
  26418=>"100100110",
  26419=>"001001000",
  26420=>"000111011",
  26421=>"101001010",
  26422=>"111001111",
  26423=>"110011110",
  26424=>"010111101",
  26425=>"000000001",
  26426=>"111100100",
  26427=>"110010111",
  26428=>"000111000",
  26429=>"001000100",
  26430=>"111000010",
  26431=>"001010100",
  26432=>"011100000",
  26433=>"001110111",
  26434=>"101010110",
  26435=>"000010000",
  26436=>"100111000",
  26437=>"010110101",
  26438=>"111010100",
  26439=>"100011110",
  26440=>"010000100",
  26441=>"101101100",
  26442=>"010011101",
  26443=>"010110100",
  26444=>"011011111",
  26445=>"011011111",
  26446=>"001010000",
  26447=>"011111001",
  26448=>"110001001",
  26449=>"000010111",
  26450=>"101101111",
  26451=>"001111001",
  26452=>"010101001",
  26453=>"000011011",
  26454=>"101111111",
  26455=>"100010100",
  26456=>"111011011",
  26457=>"111111010",
  26458=>"000110111",
  26459=>"011010101",
  26460=>"101011010",
  26461=>"011110101",
  26462=>"001001010",
  26463=>"000100010",
  26464=>"100001111",
  26465=>"001010011",
  26466=>"100000001",
  26467=>"010111111",
  26468=>"110011011",
  26469=>"011010111",
  26470=>"101001000",
  26471=>"100001111",
  26472=>"110100000",
  26473=>"000000001",
  26474=>"111010010",
  26475=>"010110000",
  26476=>"000001101",
  26477=>"100100001",
  26478=>"011010111",
  26479=>"011000111",
  26480=>"100001111",
  26481=>"110000011",
  26482=>"111110011",
  26483=>"110001001",
  26484=>"000001010",
  26485=>"011000100",
  26486=>"110001111",
  26487=>"001101101",
  26488=>"111101110",
  26489=>"000000111",
  26490=>"000001111",
  26491=>"100111000",
  26492=>"100001011",
  26493=>"100010100",
  26494=>"000000010",
  26495=>"011011110",
  26496=>"001000000",
  26497=>"101011011",
  26498=>"011101111",
  26499=>"000000101",
  26500=>"011000000",
  26501=>"010000010",
  26502=>"101101010",
  26503=>"101001010",
  26504=>"000110100",
  26505=>"000110011",
  26506=>"010111101",
  26507=>"000000000",
  26508=>"000111100",
  26509=>"000001111",
  26510=>"001000001",
  26511=>"100010100",
  26512=>"010010000",
  26513=>"111001100",
  26514=>"100101100",
  26515=>"000101111",
  26516=>"001111011",
  26517=>"100011100",
  26518=>"010000011",
  26519=>"100010001",
  26520=>"000001010",
  26521=>"000010110",
  26522=>"100011100",
  26523=>"000100001",
  26524=>"010111101",
  26525=>"011111101",
  26526=>"000001101",
  26527=>"001000100",
  26528=>"000000110",
  26529=>"100010101",
  26530=>"001000011",
  26531=>"010100101",
  26532=>"001000010",
  26533=>"000000010",
  26534=>"110000110",
  26535=>"011010100",
  26536=>"010011000",
  26537=>"110100111",
  26538=>"101010000",
  26539=>"101101000",
  26540=>"111011000",
  26541=>"101000101",
  26542=>"110110110",
  26543=>"011111110",
  26544=>"001011001",
  26545=>"000111111",
  26546=>"110100101",
  26547=>"011100001",
  26548=>"110111110",
  26549=>"011101001",
  26550=>"011000011",
  26551=>"001001010",
  26552=>"110001011",
  26553=>"010100000",
  26554=>"010111111",
  26555=>"011110100",
  26556=>"110110100",
  26557=>"000000011",
  26558=>"100010111",
  26559=>"000000011",
  26560=>"110111001",
  26561=>"011001111",
  26562=>"000001011",
  26563=>"000000110",
  26564=>"011111100",
  26565=>"101010111",
  26566=>"011110000",
  26567=>"110001101",
  26568=>"000000000",
  26569=>"001010110",
  26570=>"100010111",
  26571=>"011101101",
  26572=>"001010111",
  26573=>"010010111",
  26574=>"001110011",
  26575=>"111101101",
  26576=>"001100001",
  26577=>"001000110",
  26578=>"000110000",
  26579=>"011101000",
  26580=>"111111011",
  26581=>"111010110",
  26582=>"111001001",
  26583=>"010001110",
  26584=>"100011001",
  26585=>"010001010",
  26586=>"011110010",
  26587=>"010101101",
  26588=>"111110101",
  26589=>"001000101",
  26590=>"001101011",
  26591=>"111011101",
  26592=>"011100011",
  26593=>"100111101",
  26594=>"011101100",
  26595=>"101000000",
  26596=>"010000000",
  26597=>"011000100",
  26598=>"101110110",
  26599=>"011100100",
  26600=>"000010010",
  26601=>"111001010",
  26602=>"000110110",
  26603=>"001011000",
  26604=>"110000110",
  26605=>"001110100",
  26606=>"111000001",
  26607=>"110011110",
  26608=>"000010111",
  26609=>"000000000",
  26610=>"010000010",
  26611=>"001100111",
  26612=>"011110101",
  26613=>"001010111",
  26614=>"100011101",
  26615=>"010000010",
  26616=>"111010001",
  26617=>"011110111",
  26618=>"011011101",
  26619=>"001011001",
  26620=>"001001100",
  26621=>"000111010",
  26622=>"110111101",
  26623=>"001001011",
  26624=>"111010001",
  26625=>"100000100",
  26626=>"110101100",
  26627=>"000000101",
  26628=>"111101010",
  26629=>"000000001",
  26630=>"010101001",
  26631=>"000111000",
  26632=>"111110111",
  26633=>"101100111",
  26634=>"000001111",
  26635=>"000111001",
  26636=>"110010011",
  26637=>"001010111",
  26638=>"110100111",
  26639=>"010010010",
  26640=>"111100000",
  26641=>"001000010",
  26642=>"110100101",
  26643=>"000100000",
  26644=>"000010110",
  26645=>"100011101",
  26646=>"100111001",
  26647=>"110110010",
  26648=>"010000111",
  26649=>"000000001",
  26650=>"111110101",
  26651=>"011010101",
  26652=>"110100100",
  26653=>"011110100",
  26654=>"101100110",
  26655=>"101000110",
  26656=>"001010111",
  26657=>"101100111",
  26658=>"001011100",
  26659=>"111010110",
  26660=>"001000000",
  26661=>"011110010",
  26662=>"000011011",
  26663=>"111100100",
  26664=>"101111101",
  26665=>"100111010",
  26666=>"100010010",
  26667=>"001110111",
  26668=>"001100011",
  26669=>"011011111",
  26670=>"000011111",
  26671=>"000101101",
  26672=>"111111001",
  26673=>"010001111",
  26674=>"000000001",
  26675=>"011011010",
  26676=>"000000000",
  26677=>"101000100",
  26678=>"010100000",
  26679=>"010110011",
  26680=>"110100111",
  26681=>"000000100",
  26682=>"001100000",
  26683=>"000010110",
  26684=>"101101110",
  26685=>"001110111",
  26686=>"110001100",
  26687=>"000011000",
  26688=>"001001111",
  26689=>"001110000",
  26690=>"100100010",
  26691=>"101000111",
  26692=>"111111111",
  26693=>"010010101",
  26694=>"110011011",
  26695=>"110110000",
  26696=>"111000111",
  26697=>"100101110",
  26698=>"001110000",
  26699=>"000010010",
  26700=>"101100111",
  26701=>"000110110",
  26702=>"010001011",
  26703=>"110000011",
  26704=>"000111001",
  26705=>"010010110",
  26706=>"001010001",
  26707=>"101011101",
  26708=>"111011101",
  26709=>"111101100",
  26710=>"010101010",
  26711=>"001001101",
  26712=>"101011110",
  26713=>"001100101",
  26714=>"001101110",
  26715=>"000100110",
  26716=>"111010110",
  26717=>"000001100",
  26718=>"110110010",
  26719=>"101110000",
  26720=>"001100010",
  26721=>"011000101",
  26722=>"001010100",
  26723=>"010001001",
  26724=>"000000000",
  26725=>"101001100",
  26726=>"111111111",
  26727=>"110101100",
  26728=>"110000101",
  26729=>"101100111",
  26730=>"000100111",
  26731=>"001111101",
  26732=>"111000000",
  26733=>"000110000",
  26734=>"110001011",
  26735=>"100100111",
  26736=>"110000000",
  26737=>"000000010",
  26738=>"000101110",
  26739=>"100100010",
  26740=>"000010110",
  26741=>"010111001",
  26742=>"011010010",
  26743=>"111101011",
  26744=>"011110001",
  26745=>"011111100",
  26746=>"111010110",
  26747=>"111000100",
  26748=>"011111110",
  26749=>"000011110",
  26750=>"010110011",
  26751=>"110100110",
  26752=>"000000010",
  26753=>"000110001",
  26754=>"001001011",
  26755=>"110010000",
  26756=>"001111000",
  26757=>"001000110",
  26758=>"010010011",
  26759=>"011000001",
  26760=>"100010010",
  26761=>"010000001",
  26762=>"000001010",
  26763=>"110111001",
  26764=>"111100101",
  26765=>"110100111",
  26766=>"110100010",
  26767=>"001100010",
  26768=>"101100011",
  26769=>"110011100",
  26770=>"111011101",
  26771=>"111000011",
  26772=>"101011111",
  26773=>"010111011",
  26774=>"000001001",
  26775=>"011000100",
  26776=>"010000011",
  26777=>"011101101",
  26778=>"110111001",
  26779=>"100110010",
  26780=>"101101000",
  26781=>"101101011",
  26782=>"100110011",
  26783=>"011111100",
  26784=>"001100010",
  26785=>"011011001",
  26786=>"111111110",
  26787=>"000111001",
  26788=>"010000001",
  26789=>"010101111",
  26790=>"000101000",
  26791=>"110011100",
  26792=>"000101100",
  26793=>"100110011",
  26794=>"110111101",
  26795=>"001100101",
  26796=>"100110110",
  26797=>"010010011",
  26798=>"100110011",
  26799=>"101101111",
  26800=>"010100101",
  26801=>"110100100",
  26802=>"011001111",
  26803=>"101011101",
  26804=>"000001001",
  26805=>"111101100",
  26806=>"001010011",
  26807=>"000111010",
  26808=>"010011010",
  26809=>"101111101",
  26810=>"000000101",
  26811=>"111110101",
  26812=>"101101000",
  26813=>"011000011",
  26814=>"011000110",
  26815=>"110110110",
  26816=>"001010110",
  26817=>"100001000",
  26818=>"111110100",
  26819=>"010000001",
  26820=>"000010101",
  26821=>"111100110",
  26822=>"011000000",
  26823=>"001001101",
  26824=>"000101100",
  26825=>"011100000",
  26826=>"111011010",
  26827=>"010111011",
  26828=>"011010101",
  26829=>"111101100",
  26830=>"100100001",
  26831=>"011010010",
  26832=>"101010000",
  26833=>"101011101",
  26834=>"100101000",
  26835=>"111100100",
  26836=>"001101011",
  26837=>"101100111",
  26838=>"100011010",
  26839=>"010101001",
  26840=>"000111111",
  26841=>"011111111",
  26842=>"110100011",
  26843=>"001100000",
  26844=>"101001110",
  26845=>"110100101",
  26846=>"000100101",
  26847=>"110010100",
  26848=>"100010001",
  26849=>"101111111",
  26850=>"001010010",
  26851=>"000110000",
  26852=>"011000011",
  26853=>"010111110",
  26854=>"001000100",
  26855=>"011010010",
  26856=>"000111010",
  26857=>"100010011",
  26858=>"000101010",
  26859=>"000011000",
  26860=>"111111101",
  26861=>"010011010",
  26862=>"000001101",
  26863=>"011010000",
  26864=>"111010000",
  26865=>"001100111",
  26866=>"111110010",
  26867=>"110000000",
  26868=>"010000011",
  26869=>"011111100",
  26870=>"010011100",
  26871=>"000010010",
  26872=>"000000101",
  26873=>"100001111",
  26874=>"111110111",
  26875=>"010110110",
  26876=>"110000001",
  26877=>"010001110",
  26878=>"111111000",
  26879=>"100101111",
  26880=>"001111011",
  26881=>"001101010",
  26882=>"011001111",
  26883=>"010001110",
  26884=>"010000111",
  26885=>"011100111",
  26886=>"001010100",
  26887=>"100110110",
  26888=>"011101111",
  26889=>"100011001",
  26890=>"110010001",
  26891=>"011101101",
  26892=>"010011101",
  26893=>"001011010",
  26894=>"100110100",
  26895=>"011110111",
  26896=>"101010000",
  26897=>"110000011",
  26898=>"110010111",
  26899=>"100111110",
  26900=>"110110011",
  26901=>"011000001",
  26902=>"011111001",
  26903=>"000000100",
  26904=>"100101001",
  26905=>"010000001",
  26906=>"000011101",
  26907=>"111011100",
  26908=>"000110110",
  26909=>"110100000",
  26910=>"110111110",
  26911=>"001010101",
  26912=>"001000111",
  26913=>"001001010",
  26914=>"100000111",
  26915=>"111111001",
  26916=>"111011010",
  26917=>"001100101",
  26918=>"001000111",
  26919=>"111011011",
  26920=>"000001011",
  26921=>"010110010",
  26922=>"011011000",
  26923=>"100010001",
  26924=>"110011111",
  26925=>"101011110",
  26926=>"000000111",
  26927=>"010011111",
  26928=>"110001011",
  26929=>"100000111",
  26930=>"011010111",
  26931=>"000010101",
  26932=>"001110010",
  26933=>"100010100",
  26934=>"000111001",
  26935=>"101011100",
  26936=>"010000100",
  26937=>"001100011",
  26938=>"100110111",
  26939=>"010100111",
  26940=>"110000111",
  26941=>"111111101",
  26942=>"010100010",
  26943=>"000101100",
  26944=>"010110001",
  26945=>"001101001",
  26946=>"111011101",
  26947=>"101101001",
  26948=>"001010001",
  26949=>"111101001",
  26950=>"110001011",
  26951=>"010000110",
  26952=>"110011111",
  26953=>"101100000",
  26954=>"111101110",
  26955=>"000010000",
  26956=>"110111111",
  26957=>"110000000",
  26958=>"000100110",
  26959=>"110000001",
  26960=>"010010101",
  26961=>"001111110",
  26962=>"001100000",
  26963=>"110100101",
  26964=>"110010001",
  26965=>"111000010",
  26966=>"111001111",
  26967=>"110111101",
  26968=>"000001101",
  26969=>"000001000",
  26970=>"111111100",
  26971=>"000000011",
  26972=>"010011001",
  26973=>"001100010",
  26974=>"011010001",
  26975=>"001110001",
  26976=>"011000010",
  26977=>"100001110",
  26978=>"001000111",
  26979=>"001101001",
  26980=>"101001010",
  26981=>"001011111",
  26982=>"011001101",
  26983=>"111000000",
  26984=>"000001000",
  26985=>"000000000",
  26986=>"100001010",
  26987=>"000101111",
  26988=>"001010010",
  26989=>"000100010",
  26990=>"000000110",
  26991=>"011001000",
  26992=>"000101111",
  26993=>"000100010",
  26994=>"010101100",
  26995=>"010111011",
  26996=>"000110110",
  26997=>"101000000",
  26998=>"010001010",
  26999=>"000011111",
  27000=>"011011010",
  27001=>"000000000",
  27002=>"110011000",
  27003=>"001001010",
  27004=>"010000100",
  27005=>"011100010",
  27006=>"100010101",
  27007=>"100000000",
  27008=>"000111100",
  27009=>"011000111",
  27010=>"110001101",
  27011=>"100011111",
  27012=>"001000011",
  27013=>"100001011",
  27014=>"100101100",
  27015=>"100100101",
  27016=>"101001000",
  27017=>"011010000",
  27018=>"100010111",
  27019=>"001001111",
  27020=>"100100101",
  27021=>"010010001",
  27022=>"111101101",
  27023=>"010100001",
  27024=>"000000011",
  27025=>"000000010",
  27026=>"001010111",
  27027=>"010000100",
  27028=>"101011001",
  27029=>"101110100",
  27030=>"101111111",
  27031=>"101110001",
  27032=>"010011111",
  27033=>"001011100",
  27034=>"111001001",
  27035=>"010000101",
  27036=>"000101101",
  27037=>"100011000",
  27038=>"100111111",
  27039=>"111010000",
  27040=>"110100110",
  27041=>"001000100",
  27042=>"010010010",
  27043=>"001000001",
  27044=>"110111100",
  27045=>"110000000",
  27046=>"010001011",
  27047=>"111010110",
  27048=>"101010110",
  27049=>"000110100",
  27050=>"101001101",
  27051=>"101010101",
  27052=>"011110101",
  27053=>"101010111",
  27054=>"001100010",
  27055=>"100001011",
  27056=>"010110101",
  27057=>"111001110",
  27058=>"001010101",
  27059=>"111011001",
  27060=>"001001011",
  27061=>"001000000",
  27062=>"001100111",
  27063=>"010001101",
  27064=>"001011000",
  27065=>"000000110",
  27066=>"001101001",
  27067=>"101110000",
  27068=>"010111100",
  27069=>"111010011",
  27070=>"010110110",
  27071=>"010010000",
  27072=>"000000000",
  27073=>"011111111",
  27074=>"000000010",
  27075=>"111001111",
  27076=>"110101010",
  27077=>"010101010",
  27078=>"001011001",
  27079=>"111110100",
  27080=>"101111101",
  27081=>"100100110",
  27082=>"010110000",
  27083=>"100110001",
  27084=>"101010011",
  27085=>"110110011",
  27086=>"101001010",
  27087=>"011111010",
  27088=>"111011001",
  27089=>"010001100",
  27090=>"001111000",
  27091=>"011111111",
  27092=>"011001100",
  27093=>"001111101",
  27094=>"011111000",
  27095=>"011101101",
  27096=>"010000011",
  27097=>"000111001",
  27098=>"001111101",
  27099=>"111100010",
  27100=>"110110101",
  27101=>"111100111",
  27102=>"010111011",
  27103=>"111010100",
  27104=>"110100001",
  27105=>"110110110",
  27106=>"101111111",
  27107=>"011011100",
  27108=>"010110110",
  27109=>"101011001",
  27110=>"100111011",
  27111=>"100110001",
  27112=>"011011100",
  27113=>"111111101",
  27114=>"100011010",
  27115=>"111111010",
  27116=>"111111000",
  27117=>"110100010",
  27118=>"001010000",
  27119=>"000000011",
  27120=>"111011001",
  27121=>"100111110",
  27122=>"101000010",
  27123=>"000000100",
  27124=>"010001010",
  27125=>"000000101",
  27126=>"101011010",
  27127=>"110000111",
  27128=>"110101111",
  27129=>"001000000",
  27130=>"101110001",
  27131=>"001111111",
  27132=>"110101101",
  27133=>"111101011",
  27134=>"001100110",
  27135=>"111001101",
  27136=>"011000001",
  27137=>"001011110",
  27138=>"010001101",
  27139=>"101011010",
  27140=>"111010111",
  27141=>"111110010",
  27142=>"111100111",
  27143=>"111010111",
  27144=>"111000000",
  27145=>"110100001",
  27146=>"001001100",
  27147=>"000010100",
  27148=>"010111000",
  27149=>"100111001",
  27150=>"101000100",
  27151=>"101011010",
  27152=>"010001100",
  27153=>"101011100",
  27154=>"001000001",
  27155=>"001000011",
  27156=>"000101010",
  27157=>"011000010",
  27158=>"111000101",
  27159=>"010011001",
  27160=>"100010101",
  27161=>"100010011",
  27162=>"000001000",
  27163=>"011000101",
  27164=>"100001100",
  27165=>"011101100",
  27166=>"111010110",
  27167=>"111110001",
  27168=>"100101000",
  27169=>"001000100",
  27170=>"110001011",
  27171=>"011110101",
  27172=>"111011101",
  27173=>"011111101",
  27174=>"000110010",
  27175=>"111010010",
  27176=>"010100101",
  27177=>"100001000",
  27178=>"011001100",
  27179=>"000001001",
  27180=>"000000001",
  27181=>"101001000",
  27182=>"100000011",
  27183=>"000100010",
  27184=>"101110101",
  27185=>"010100101",
  27186=>"100100101",
  27187=>"000100010",
  27188=>"001111111",
  27189=>"000000100",
  27190=>"101110100",
  27191=>"010101010",
  27192=>"010011010",
  27193=>"000001111",
  27194=>"110000100",
  27195=>"000010111",
  27196=>"000101010",
  27197=>"110100000",
  27198=>"010111100",
  27199=>"100110011",
  27200=>"000101111",
  27201=>"000100000",
  27202=>"110011001",
  27203=>"110100110",
  27204=>"110101111",
  27205=>"011011100",
  27206=>"110000000",
  27207=>"100010100",
  27208=>"001101100",
  27209=>"101000000",
  27210=>"101111000",
  27211=>"010011011",
  27212=>"110010111",
  27213=>"111001101",
  27214=>"101101011",
  27215=>"100101000",
  27216=>"110001010",
  27217=>"000000100",
  27218=>"101101111",
  27219=>"010101010",
  27220=>"111101010",
  27221=>"000100010",
  27222=>"100100111",
  27223=>"110110011",
  27224=>"111001011",
  27225=>"111000000",
  27226=>"000111001",
  27227=>"001000000",
  27228=>"111000000",
  27229=>"000000100",
  27230=>"010100010",
  27231=>"011110101",
  27232=>"001000010",
  27233=>"010010100",
  27234=>"110001010",
  27235=>"001010000",
  27236=>"010110111",
  27237=>"101100101",
  27238=>"110000001",
  27239=>"100011111",
  27240=>"100001110",
  27241=>"101011101",
  27242=>"101110111",
  27243=>"100100101",
  27244=>"100111011",
  27245=>"101001001",
  27246=>"010110000",
  27247=>"001010111",
  27248=>"010011100",
  27249=>"101000000",
  27250=>"110010000",
  27251=>"011001111",
  27252=>"101111100",
  27253=>"010011001",
  27254=>"000011110",
  27255=>"001111100",
  27256=>"101000111",
  27257=>"110010000",
  27258=>"010111110",
  27259=>"111001010",
  27260=>"101010000",
  27261=>"000010000",
  27262=>"111101100",
  27263=>"111110110",
  27264=>"101000110",
  27265=>"101100100",
  27266=>"000001011",
  27267=>"100010000",
  27268=>"011110100",
  27269=>"011001000",
  27270=>"101100100",
  27271=>"001010000",
  27272=>"100010110",
  27273=>"101110110",
  27274=>"010111111",
  27275=>"000011011",
  27276=>"010111101",
  27277=>"100100011",
  27278=>"111100010",
  27279=>"100001101",
  27280=>"110100101",
  27281=>"100101110",
  27282=>"110110001",
  27283=>"011101110",
  27284=>"100010100",
  27285=>"100011010",
  27286=>"100000011",
  27287=>"101001001",
  27288=>"011111101",
  27289=>"000101011",
  27290=>"110111010",
  27291=>"010000110",
  27292=>"100011111",
  27293=>"101101010",
  27294=>"001111110",
  27295=>"011000011",
  27296=>"001111111",
  27297=>"101110101",
  27298=>"101100111",
  27299=>"100101001",
  27300=>"001101110",
  27301=>"110100101",
  27302=>"100100010",
  27303=>"111011101",
  27304=>"001101010",
  27305=>"100001011",
  27306=>"101011110",
  27307=>"011011001",
  27308=>"010111011",
  27309=>"101100001",
  27310=>"111101011",
  27311=>"011001100",
  27312=>"000000010",
  27313=>"001111101",
  27314=>"010111000",
  27315=>"000010101",
  27316=>"000000010",
  27317=>"100001101",
  27318=>"001011000",
  27319=>"111111111",
  27320=>"010001100",
  27321=>"010001010",
  27322=>"101001011",
  27323=>"100011001",
  27324=>"110100101",
  27325=>"001000110",
  27326=>"100100110",
  27327=>"010010101",
  27328=>"010100001",
  27329=>"001101000",
  27330=>"001001110",
  27331=>"001110100",
  27332=>"001000110",
  27333=>"101111100",
  27334=>"100100011",
  27335=>"110111111",
  27336=>"111111101",
  27337=>"011101111",
  27338=>"011110100",
  27339=>"001010101",
  27340=>"011100111",
  27341=>"011011110",
  27342=>"010000000",
  27343=>"111010001",
  27344=>"110001000",
  27345=>"101100100",
  27346=>"001011100",
  27347=>"001111001",
  27348=>"010100111",
  27349=>"000000110",
  27350=>"011101001",
  27351=>"101000111",
  27352=>"100100101",
  27353=>"011000011",
  27354=>"001110100",
  27355=>"010101011",
  27356=>"000100000",
  27357=>"000101000",
  27358=>"110111000",
  27359=>"100101100",
  27360=>"010111011",
  27361=>"101000100",
  27362=>"111101010",
  27363=>"100100001",
  27364=>"100110111",
  27365=>"000011100",
  27366=>"110001101",
  27367=>"100110011",
  27368=>"000010100",
  27369=>"110100010",
  27370=>"110110100",
  27371=>"010000010",
  27372=>"000001101",
  27373=>"100100010",
  27374=>"011110101",
  27375=>"010010001",
  27376=>"010101101",
  27377=>"001011110",
  27378=>"000010000",
  27379=>"110100010",
  27380=>"011000100",
  27381=>"001111001",
  27382=>"101110001",
  27383=>"111000000",
  27384=>"101110001",
  27385=>"011000000",
  27386=>"010000000",
  27387=>"111001010",
  27388=>"001000100",
  27389=>"001000111",
  27390=>"100011001",
  27391=>"100010011",
  27392=>"011001100",
  27393=>"011011011",
  27394=>"110101111",
  27395=>"011000010",
  27396=>"101011110",
  27397=>"000000010",
  27398=>"000101000",
  27399=>"000001001",
  27400=>"100011001",
  27401=>"011010010",
  27402=>"011100010",
  27403=>"111111110",
  27404=>"101110110",
  27405=>"110001010",
  27406=>"011010000",
  27407=>"000011100",
  27408=>"001011001",
  27409=>"001110000",
  27410=>"100111000",
  27411=>"111001111",
  27412=>"110000010",
  27413=>"110100010",
  27414=>"000000000",
  27415=>"000001110",
  27416=>"101110111",
  27417=>"111101001",
  27418=>"001111100",
  27419=>"010110000",
  27420=>"110110000",
  27421=>"010000101",
  27422=>"110100010",
  27423=>"101101110",
  27424=>"100000101",
  27425=>"101011101",
  27426=>"111110100",
  27427=>"110110101",
  27428=>"100011010",
  27429=>"000000010",
  27430=>"101001010",
  27431=>"001001111",
  27432=>"110000111",
  27433=>"101100000",
  27434=>"100101111",
  27435=>"110111100",
  27436=>"010010101",
  27437=>"100001010",
  27438=>"101100110",
  27439=>"111100100",
  27440=>"011110010",
  27441=>"000010000",
  27442=>"111000000",
  27443=>"010010111",
  27444=>"101111101",
  27445=>"111011110",
  27446=>"000000110",
  27447=>"101101010",
  27448=>"011000111",
  27449=>"111000111",
  27450=>"010111110",
  27451=>"011100001",
  27452=>"000001001",
  27453=>"111001010",
  27454=>"001000001",
  27455=>"100111001",
  27456=>"001111111",
  27457=>"101010101",
  27458=>"111110000",
  27459=>"111110101",
  27460=>"001111101",
  27461=>"101010001",
  27462=>"101000001",
  27463=>"101001101",
  27464=>"111010000",
  27465=>"010001000",
  27466=>"001011000",
  27467=>"100110001",
  27468=>"101111010",
  27469=>"001011010",
  27470=>"010010000",
  27471=>"011010011",
  27472=>"111111001",
  27473=>"000001110",
  27474=>"101011110",
  27475=>"011101101",
  27476=>"011000100",
  27477=>"100110111",
  27478=>"011011110",
  27479=>"000011101",
  27480=>"001110010",
  27481=>"000011011",
  27482=>"110001011",
  27483=>"010110110",
  27484=>"011001001",
  27485=>"011111010",
  27486=>"110111111",
  27487=>"000000011",
  27488=>"010001000",
  27489=>"111101110",
  27490=>"001000001",
  27491=>"111011010",
  27492=>"101010100",
  27493=>"011110000",
  27494=>"101111010",
  27495=>"110010111",
  27496=>"010011000",
  27497=>"001111110",
  27498=>"010010011",
  27499=>"111010101",
  27500=>"111101001",
  27501=>"110110011",
  27502=>"110100010",
  27503=>"100101100",
  27504=>"011010000",
  27505=>"001011100",
  27506=>"011000000",
  27507=>"111100111",
  27508=>"100110100",
  27509=>"110101110",
  27510=>"110100011",
  27511=>"110000000",
  27512=>"110110010",
  27513=>"010011011",
  27514=>"111101000",
  27515=>"000100111",
  27516=>"010011101",
  27517=>"010100000",
  27518=>"100110110",
  27519=>"110011111",
  27520=>"111011101",
  27521=>"101011100",
  27522=>"111000001",
  27523=>"000110101",
  27524=>"000110101",
  27525=>"000100011",
  27526=>"001101001",
  27527=>"000110010",
  27528=>"111111101",
  27529=>"110111011",
  27530=>"010001001",
  27531=>"000000010",
  27532=>"011010000",
  27533=>"011111110",
  27534=>"000101101",
  27535=>"101000100",
  27536=>"010011001",
  27537=>"001001100",
  27538=>"001000100",
  27539=>"001000110",
  27540=>"101000111",
  27541=>"101111010",
  27542=>"111001000",
  27543=>"111001000",
  27544=>"000110010",
  27545=>"111101001",
  27546=>"110110001",
  27547=>"001110110",
  27548=>"011011011",
  27549=>"111000100",
  27550=>"110001010",
  27551=>"001100000",
  27552=>"111001111",
  27553=>"111110100",
  27554=>"100010111",
  27555=>"000101010",
  27556=>"000011101",
  27557=>"101001001",
  27558=>"100111110",
  27559=>"111010001",
  27560=>"010100111",
  27561=>"000001000",
  27562=>"001011011",
  27563=>"001010011",
  27564=>"101011010",
  27565=>"100011000",
  27566=>"000101110",
  27567=>"111101010",
  27568=>"011011111",
  27569=>"111011010",
  27570=>"001001010",
  27571=>"101001011",
  27572=>"010100001",
  27573=>"011011001",
  27574=>"001101111",
  27575=>"110011100",
  27576=>"110100011",
  27577=>"011111001",
  27578=>"100110001",
  27579=>"000000110",
  27580=>"000000000",
  27581=>"111101101",
  27582=>"101101011",
  27583=>"101100100",
  27584=>"111110101",
  27585=>"011111000",
  27586=>"000010011",
  27587=>"010111010",
  27588=>"000000000",
  27589=>"010101111",
  27590=>"010111100",
  27591=>"110100001",
  27592=>"100110000",
  27593=>"000101001",
  27594=>"100011001",
  27595=>"110110110",
  27596=>"011101101",
  27597=>"101100100",
  27598=>"100001111",
  27599=>"110101001",
  27600=>"001110110",
  27601=>"001100100",
  27602=>"100000000",
  27603=>"011011010",
  27604=>"010111010",
  27605=>"010001111",
  27606=>"101100010",
  27607=>"101001010",
  27608=>"111010101",
  27609=>"011100101",
  27610=>"011001101",
  27611=>"011010000",
  27612=>"101101010",
  27613=>"000101001",
  27614=>"000110001",
  27615=>"100010001",
  27616=>"110111111",
  27617=>"000000100",
  27618=>"111011011",
  27619=>"110111001",
  27620=>"101110010",
  27621=>"011010111",
  27622=>"111110000",
  27623=>"010101100",
  27624=>"101011000",
  27625=>"110111000",
  27626=>"100001100",
  27627=>"010000111",
  27628=>"000000010",
  27629=>"010001001",
  27630=>"010000011",
  27631=>"011110000",
  27632=>"010110011",
  27633=>"001111110",
  27634=>"111010000",
  27635=>"001101000",
  27636=>"110011000",
  27637=>"111100100",
  27638=>"001011000",
  27639=>"010001001",
  27640=>"011001100",
  27641=>"110011010",
  27642=>"100000100",
  27643=>"111111011",
  27644=>"011011001",
  27645=>"110111010",
  27646=>"000001011",
  27647=>"110011000",
  27648=>"011101000",
  27649=>"111100010",
  27650=>"011101011",
  27651=>"011100101",
  27652=>"000001100",
  27653=>"000000000",
  27654=>"011011001",
  27655=>"111110110",
  27656=>"010111001",
  27657=>"000011110",
  27658=>"011100000",
  27659=>"101100010",
  27660=>"110101100",
  27661=>"011000101",
  27662=>"010000001",
  27663=>"111101111",
  27664=>"001001001",
  27665=>"100001000",
  27666=>"111001111",
  27667=>"001010110",
  27668=>"001001010",
  27669=>"101110001",
  27670=>"000011110",
  27671=>"100000011",
  27672=>"001011001",
  27673=>"111011101",
  27674=>"010110001",
  27675=>"110001110",
  27676=>"111000010",
  27677=>"000111111",
  27678=>"011000011",
  27679=>"110101010",
  27680=>"011100110",
  27681=>"011001000",
  27682=>"001110010",
  27683=>"001011001",
  27684=>"111100100",
  27685=>"101101001",
  27686=>"101101110",
  27687=>"000010100",
  27688=>"000000101",
  27689=>"100011110",
  27690=>"011101000",
  27691=>"001001010",
  27692=>"111101101",
  27693=>"001110100",
  27694=>"001000000",
  27695=>"010110001",
  27696=>"001011111",
  27697=>"001011000",
  27698=>"101110101",
  27699=>"100100110",
  27700=>"001101110",
  27701=>"001101000",
  27702=>"110101111",
  27703=>"100110111",
  27704=>"011101000",
  27705=>"000000111",
  27706=>"001100001",
  27707=>"011011111",
  27708=>"100100010",
  27709=>"100000100",
  27710=>"101110110",
  27711=>"000010011",
  27712=>"110001001",
  27713=>"101011010",
  27714=>"000111111",
  27715=>"100011000",
  27716=>"111011011",
  27717=>"010001110",
  27718=>"000100000",
  27719=>"010010001",
  27720=>"000110001",
  27721=>"010100100",
  27722=>"001011110",
  27723=>"101000111",
  27724=>"001010100",
  27725=>"101001110",
  27726=>"000110001",
  27727=>"001111110",
  27728=>"101000101",
  27729=>"101001110",
  27730=>"100001100",
  27731=>"011110101",
  27732=>"101111110",
  27733=>"010010111",
  27734=>"011101110",
  27735=>"101101000",
  27736=>"010110101",
  27737=>"001110110",
  27738=>"101100111",
  27739=>"000011001",
  27740=>"000000000",
  27741=>"101110101",
  27742=>"000001011",
  27743=>"011100101",
  27744=>"001000111",
  27745=>"010110110",
  27746=>"001001110",
  27747=>"011110111",
  27748=>"110011100",
  27749=>"100010010",
  27750=>"010100011",
  27751=>"010011100",
  27752=>"011010100",
  27753=>"101111001",
  27754=>"011000100",
  27755=>"101010110",
  27756=>"000001010",
  27757=>"111101011",
  27758=>"100010111",
  27759=>"011001100",
  27760=>"100100010",
  27761=>"001000001",
  27762=>"111111001",
  27763=>"000011011",
  27764=>"101110110",
  27765=>"100110100",
  27766=>"111011101",
  27767=>"011011000",
  27768=>"000100000",
  27769=>"111100111",
  27770=>"000000100",
  27771=>"111110010",
  27772=>"010000101",
  27773=>"110100100",
  27774=>"101010000",
  27775=>"000110001",
  27776=>"101011111",
  27777=>"100000011",
  27778=>"000111111",
  27779=>"111001011",
  27780=>"011010001",
  27781=>"000001101",
  27782=>"010010001",
  27783=>"011111010",
  27784=>"001010101",
  27785=>"010001100",
  27786=>"011001100",
  27787=>"010001000",
  27788=>"111001011",
  27789=>"000001010",
  27790=>"111001111",
  27791=>"011100100",
  27792=>"001000111",
  27793=>"101000111",
  27794=>"000101000",
  27795=>"100011010",
  27796=>"000000101",
  27797=>"100100000",
  27798=>"010001111",
  27799=>"101110010",
  27800=>"001001000",
  27801=>"000100000",
  27802=>"011110010",
  27803=>"111000100",
  27804=>"100110101",
  27805=>"100000000",
  27806=>"010001001",
  27807=>"000100010",
  27808=>"111000111",
  27809=>"011111100",
  27810=>"111011110",
  27811=>"110001010",
  27812=>"101010000",
  27813=>"100110010",
  27814=>"000000000",
  27815=>"111000100",
  27816=>"010010110",
  27817=>"001001101",
  27818=>"100101110",
  27819=>"011111010",
  27820=>"010110110",
  27821=>"111100100",
  27822=>"111100101",
  27823=>"101010001",
  27824=>"011110000",
  27825=>"000000000",
  27826=>"100010101",
  27827=>"100110001",
  27828=>"001100111",
  27829=>"100110010",
  27830=>"100000101",
  27831=>"000110101",
  27832=>"000100100",
  27833=>"001010001",
  27834=>"101100100",
  27835=>"010111011",
  27836=>"111110101",
  27837=>"000100110",
  27838=>"011000110",
  27839=>"101010010",
  27840=>"000001101",
  27841=>"101100000",
  27842=>"001011001",
  27843=>"110101000",
  27844=>"110111100",
  27845=>"011111101",
  27846=>"011101011",
  27847=>"111101001",
  27848=>"011010010",
  27849=>"000101100",
  27850=>"001001010",
  27851=>"100000010",
  27852=>"100011111",
  27853=>"110101101",
  27854=>"000111000",
  27855=>"111010011",
  27856=>"100111101",
  27857=>"001100100",
  27858=>"000100101",
  27859=>"110111101",
  27860=>"101011001",
  27861=>"000111111",
  27862=>"010001111",
  27863=>"110001110",
  27864=>"000010000",
  27865=>"001100100",
  27866=>"100110101",
  27867=>"001110111",
  27868=>"010000111",
  27869=>"110011101",
  27870=>"001100000",
  27871=>"101001111",
  27872=>"100100011",
  27873=>"111010101",
  27874=>"111101010",
  27875=>"111011100",
  27876=>"001000001",
  27877=>"001011101",
  27878=>"100011111",
  27879=>"000011001",
  27880=>"010100101",
  27881=>"001100001",
  27882=>"110101111",
  27883=>"010001010",
  27884=>"110110111",
  27885=>"111011101",
  27886=>"100110100",
  27887=>"000100010",
  27888=>"101111001",
  27889=>"100110010",
  27890=>"100101101",
  27891=>"000000000",
  27892=>"001001101",
  27893=>"000011110",
  27894=>"100111110",
  27895=>"000101011",
  27896=>"010010100",
  27897=>"100101010",
  27898=>"111001011",
  27899=>"100100110",
  27900=>"010001100",
  27901=>"100001101",
  27902=>"111110011",
  27903=>"101110111",
  27904=>"011001001",
  27905=>"010011110",
  27906=>"100011000",
  27907=>"010100000",
  27908=>"010010011",
  27909=>"111111010",
  27910=>"001100001",
  27911=>"000100001",
  27912=>"011100011",
  27913=>"111001110",
  27914=>"110001111",
  27915=>"110101010",
  27916=>"010110000",
  27917=>"000000110",
  27918=>"000011101",
  27919=>"000000000",
  27920=>"101011001",
  27921=>"011101101",
  27922=>"011101010",
  27923=>"100011110",
  27924=>"000010101",
  27925=>"100011000",
  27926=>"010000100",
  27927=>"101111000",
  27928=>"101011001",
  27929=>"001000111",
  27930=>"010000011",
  27931=>"100010010",
  27932=>"110001010",
  27933=>"001011111",
  27934=>"110111110",
  27935=>"100000110",
  27936=>"111100100",
  27937=>"011110001",
  27938=>"101100100",
  27939=>"011100011",
  27940=>"101101101",
  27941=>"001000010",
  27942=>"010010000",
  27943=>"010011011",
  27944=>"101110010",
  27945=>"010001100",
  27946=>"111001001",
  27947=>"100001010",
  27948=>"101111011",
  27949=>"110001000",
  27950=>"010101111",
  27951=>"000011011",
  27952=>"111010001",
  27953=>"000011101",
  27954=>"001011111",
  27955=>"100010110",
  27956=>"000110111",
  27957=>"110111000",
  27958=>"010000001",
  27959=>"101110101",
  27960=>"000000110",
  27961=>"110010011",
  27962=>"011111110",
  27963=>"100011011",
  27964=>"000001001",
  27965=>"100000101",
  27966=>"010011100",
  27967=>"100110000",
  27968=>"011101000",
  27969=>"000010110",
  27970=>"010111111",
  27971=>"010111010",
  27972=>"000001111",
  27973=>"001010101",
  27974=>"000100010",
  27975=>"000000111",
  27976=>"101000100",
  27977=>"011001110",
  27978=>"111010000",
  27979=>"001111100",
  27980=>"110010001",
  27981=>"110110111",
  27982=>"110000011",
  27983=>"011001011",
  27984=>"111001000",
  27985=>"101101100",
  27986=>"101110011",
  27987=>"110001011",
  27988=>"101111101",
  27989=>"110011000",
  27990=>"110101001",
  27991=>"100010110",
  27992=>"100010011",
  27993=>"000000110",
  27994=>"011111011",
  27995=>"010001111",
  27996=>"101111101",
  27997=>"010010101",
  27998=>"111111000",
  27999=>"000010110",
  28000=>"010011101",
  28001=>"100111111",
  28002=>"110000000",
  28003=>"101100010",
  28004=>"101111111",
  28005=>"010001000",
  28006=>"010100101",
  28007=>"010111010",
  28008=>"110010001",
  28009=>"001000111",
  28010=>"000001100",
  28011=>"000101011",
  28012=>"011010010",
  28013=>"101110101",
  28014=>"100001001",
  28015=>"100001110",
  28016=>"100111100",
  28017=>"001111010",
  28018=>"101111001",
  28019=>"101011111",
  28020=>"011011101",
  28021=>"011101101",
  28022=>"000000011",
  28023=>"111010011",
  28024=>"110101001",
  28025=>"101100111",
  28026=>"011010001",
  28027=>"101010101",
  28028=>"111011111",
  28029=>"000101011",
  28030=>"110111101",
  28031=>"110101110",
  28032=>"001110110",
  28033=>"101001010",
  28034=>"100100011",
  28035=>"110101111",
  28036=>"110010011",
  28037=>"011111010",
  28038=>"010111011",
  28039=>"000110111",
  28040=>"010011111",
  28041=>"110111011",
  28042=>"000101000",
  28043=>"101111011",
  28044=>"100011101",
  28045=>"011001001",
  28046=>"011101000",
  28047=>"000100011",
  28048=>"001010111",
  28049=>"000010100",
  28050=>"010110011",
  28051=>"001001100",
  28052=>"000111111",
  28053=>"111101101",
  28054=>"101111110",
  28055=>"101011100",
  28056=>"100011000",
  28057=>"110011100",
  28058=>"011010001",
  28059=>"100110000",
  28060=>"111001110",
  28061=>"000010000",
  28062=>"000011011",
  28063=>"111110100",
  28064=>"011110100",
  28065=>"110111001",
  28066=>"100010010",
  28067=>"000000111",
  28068=>"010011101",
  28069=>"011010000",
  28070=>"111000100",
  28071=>"100101110",
  28072=>"110111101",
  28073=>"001010010",
  28074=>"000101110",
  28075=>"101000010",
  28076=>"010110101",
  28077=>"010001010",
  28078=>"111111101",
  28079=>"001111011",
  28080=>"000101010",
  28081=>"011011110",
  28082=>"010011111",
  28083=>"111101100",
  28084=>"101101101",
  28085=>"000111101",
  28086=>"010010001",
  28087=>"000001011",
  28088=>"010101010",
  28089=>"000110010",
  28090=>"001001001",
  28091=>"001000000",
  28092=>"010110110",
  28093=>"011000000",
  28094=>"111100001",
  28095=>"110001000",
  28096=>"111111101",
  28097=>"100000111",
  28098=>"001111001",
  28099=>"110101110",
  28100=>"011001101",
  28101=>"111111001",
  28102=>"101110111",
  28103=>"100010110",
  28104=>"101100011",
  28105=>"011111011",
  28106=>"010000001",
  28107=>"001110101",
  28108=>"011110010",
  28109=>"000111000",
  28110=>"011001001",
  28111=>"000000110",
  28112=>"111011011",
  28113=>"111000100",
  28114=>"100111011",
  28115=>"000100010",
  28116=>"011011100",
  28117=>"011001001",
  28118=>"001110001",
  28119=>"110010100",
  28120=>"110110011",
  28121=>"011000001",
  28122=>"001000100",
  28123=>"000000000",
  28124=>"011011001",
  28125=>"001110011",
  28126=>"110010001",
  28127=>"101111111",
  28128=>"010000011",
  28129=>"111000001",
  28130=>"010100000",
  28131=>"011001011",
  28132=>"111100101",
  28133=>"110111111",
  28134=>"001010001",
  28135=>"111100100",
  28136=>"011101001",
  28137=>"000101000",
  28138=>"111011010",
  28139=>"100010001",
  28140=>"000100011",
  28141=>"111000000",
  28142=>"000111010",
  28143=>"011101000",
  28144=>"000100001",
  28145=>"111100001",
  28146=>"011000000",
  28147=>"000001101",
  28148=>"100110111",
  28149=>"110110011",
  28150=>"000001111",
  28151=>"110110100",
  28152=>"001100010",
  28153=>"010001010",
  28154=>"110000010",
  28155=>"011011011",
  28156=>"011111001",
  28157=>"100000000",
  28158=>"010110010",
  28159=>"011101111",
  28160=>"000010000",
  28161=>"111010001",
  28162=>"100100101",
  28163=>"101111001",
  28164=>"101010110",
  28165=>"000111010",
  28166=>"001000101",
  28167=>"010100101",
  28168=>"000111000",
  28169=>"100111011",
  28170=>"100011011",
  28171=>"000011100",
  28172=>"001101011",
  28173=>"100111100",
  28174=>"111000101",
  28175=>"100010111",
  28176=>"000111010",
  28177=>"100111111",
  28178=>"100011001",
  28179=>"101001111",
  28180=>"000111011",
  28181=>"100110000",
  28182=>"000100110",
  28183=>"000010000",
  28184=>"001001101",
  28185=>"001110010",
  28186=>"001100110",
  28187=>"000010001",
  28188=>"101000000",
  28189=>"001111111",
  28190=>"110011100",
  28191=>"101001010",
  28192=>"110001111",
  28193=>"100001101",
  28194=>"111011001",
  28195=>"100000100",
  28196=>"000011101",
  28197=>"000100011",
  28198=>"010100011",
  28199=>"001110111",
  28200=>"000010001",
  28201=>"101101100",
  28202=>"010101111",
  28203=>"110110110",
  28204=>"001011011",
  28205=>"001100110",
  28206=>"110101101",
  28207=>"010001111",
  28208=>"000000011",
  28209=>"111000011",
  28210=>"011101011",
  28211=>"111110110",
  28212=>"100011110",
  28213=>"001101110",
  28214=>"011010100",
  28215=>"110000001",
  28216=>"100000000",
  28217=>"110010111",
  28218=>"011011011",
  28219=>"011101010",
  28220=>"110011111",
  28221=>"101100111",
  28222=>"110001000",
  28223=>"011101111",
  28224=>"100101010",
  28225=>"000001110",
  28226=>"000000000",
  28227=>"000011110",
  28228=>"000110100",
  28229=>"110100011",
  28230=>"100001001",
  28231=>"010000000",
  28232=>"110010010",
  28233=>"010010101",
  28234=>"010010100",
  28235=>"111001100",
  28236=>"111001000",
  28237=>"111001001",
  28238=>"011110000",
  28239=>"011010110",
  28240=>"101111011",
  28241=>"000110111",
  28242=>"101001010",
  28243=>"110000111",
  28244=>"001010000",
  28245=>"111100111",
  28246=>"000110110",
  28247=>"010000011",
  28248=>"000000010",
  28249=>"110000010",
  28250=>"011010011",
  28251=>"010001111",
  28252=>"101010110",
  28253=>"101110111",
  28254=>"001011100",
  28255=>"000000100",
  28256=>"101101101",
  28257=>"010001111",
  28258=>"100011001",
  28259=>"010010000",
  28260=>"000100011",
  28261=>"110010110",
  28262=>"011110000",
  28263=>"000111110",
  28264=>"011110111",
  28265=>"011111000",
  28266=>"001110001",
  28267=>"000000001",
  28268=>"011001110",
  28269=>"001110011",
  28270=>"110100111",
  28271=>"011001101",
  28272=>"100011011",
  28273=>"000010001",
  28274=>"010001000",
  28275=>"101101001",
  28276=>"010011110",
  28277=>"010100100",
  28278=>"011110000",
  28279=>"010110001",
  28280=>"111110001",
  28281=>"010001000",
  28282=>"001011011",
  28283=>"011110010",
  28284=>"100100101",
  28285=>"101000011",
  28286=>"111010010",
  28287=>"101100011",
  28288=>"001000010",
  28289=>"010010000",
  28290=>"000110000",
  28291=>"000101100",
  28292=>"111001111",
  28293=>"101011011",
  28294=>"111110110",
  28295=>"100100100",
  28296=>"111011011",
  28297=>"110011001",
  28298=>"000111011",
  28299=>"010001010",
  28300=>"010010101",
  28301=>"101010101",
  28302=>"001000000",
  28303=>"010100010",
  28304=>"001111101",
  28305=>"111101000",
  28306=>"111010101",
  28307=>"111111011",
  28308=>"001000010",
  28309=>"000100001",
  28310=>"100100001",
  28311=>"100001001",
  28312=>"101110000",
  28313=>"101111110",
  28314=>"110111010",
  28315=>"100110110",
  28316=>"100111111",
  28317=>"110111100",
  28318=>"111100111",
  28319=>"000000001",
  28320=>"111011100",
  28321=>"001010001",
  28322=>"111011101",
  28323=>"000001010",
  28324=>"110110000",
  28325=>"011110000",
  28326=>"000001000",
  28327=>"001100110",
  28328=>"101111000",
  28329=>"010101001",
  28330=>"100011010",
  28331=>"110000111",
  28332=>"010001110",
  28333=>"000001101",
  28334=>"111100001",
  28335=>"010000011",
  28336=>"001010001",
  28337=>"110001101",
  28338=>"001111011",
  28339=>"000110110",
  28340=>"100101100",
  28341=>"000001100",
  28342=>"100110111",
  28343=>"001000110",
  28344=>"110110111",
  28345=>"010100100",
  28346=>"101111001",
  28347=>"011100111",
  28348=>"001000001",
  28349=>"100100111",
  28350=>"011000111",
  28351=>"111100010",
  28352=>"101110110",
  28353=>"101011011",
  28354=>"100000110",
  28355=>"101001111",
  28356=>"101000111",
  28357=>"110100000",
  28358=>"001111101",
  28359=>"010011000",
  28360=>"001111001",
  28361=>"000110010",
  28362=>"100100010",
  28363=>"100111110",
  28364=>"000101001",
  28365=>"000100011",
  28366=>"010110010",
  28367=>"001101000",
  28368=>"000110000",
  28369=>"000000111",
  28370=>"010011001",
  28371=>"000000001",
  28372=>"110011001",
  28373=>"010000111",
  28374=>"011010101",
  28375=>"100001001",
  28376=>"010100010",
  28377=>"010011011",
  28378=>"011010000",
  28379=>"110110010",
  28380=>"011000011",
  28381=>"011101101",
  28382=>"110010100",
  28383=>"110000000",
  28384=>"000110111",
  28385=>"001101011",
  28386=>"101100001",
  28387=>"001110111",
  28388=>"100011111",
  28389=>"000111111",
  28390=>"011010001",
  28391=>"100101011",
  28392=>"100100000",
  28393=>"110111001",
  28394=>"010010101",
  28395=>"010110011",
  28396=>"000111111",
  28397=>"000000010",
  28398=>"101010110",
  28399=>"111000010",
  28400=>"001011110",
  28401=>"101000111",
  28402=>"000011011",
  28403=>"111101011",
  28404=>"000111001",
  28405=>"110010101",
  28406=>"110100010",
  28407=>"011101011",
  28408=>"101000010",
  28409=>"101000111",
  28410=>"010101010",
  28411=>"011001011",
  28412=>"110001111",
  28413=>"011011001",
  28414=>"010001000",
  28415=>"000010010",
  28416=>"110101001",
  28417=>"101000001",
  28418=>"000010000",
  28419=>"110001101",
  28420=>"001110101",
  28421=>"000000011",
  28422=>"010111110",
  28423=>"000011011",
  28424=>"001110110",
  28425=>"100110101",
  28426=>"011000111",
  28427=>"111000101",
  28428=>"101011011",
  28429=>"010110101",
  28430=>"100110010",
  28431=>"010000011",
  28432=>"010101101",
  28433=>"110100001",
  28434=>"011110100",
  28435=>"001011001",
  28436=>"001101100",
  28437=>"000010110",
  28438=>"100011010",
  28439=>"110111110",
  28440=>"111100000",
  28441=>"011011011",
  28442=>"010110010",
  28443=>"000111001",
  28444=>"000011110",
  28445=>"100010100",
  28446=>"011011001",
  28447=>"000111100",
  28448=>"110010000",
  28449=>"101101000",
  28450=>"010111010",
  28451=>"110110110",
  28452=>"000101011",
  28453=>"101110110",
  28454=>"111111010",
  28455=>"000110101",
  28456=>"011001100",
  28457=>"101110110",
  28458=>"111101110",
  28459=>"111001010",
  28460=>"000000001",
  28461=>"010100100",
  28462=>"100111000",
  28463=>"001000011",
  28464=>"111000100",
  28465=>"110000010",
  28466=>"101001100",
  28467=>"010100000",
  28468=>"001010101",
  28469=>"100000100",
  28470=>"101100110",
  28471=>"011111001",
  28472=>"100000001",
  28473=>"111101100",
  28474=>"110010111",
  28475=>"101100111",
  28476=>"011111000",
  28477=>"001010010",
  28478=>"110011001",
  28479=>"000000111",
  28480=>"100000110",
  28481=>"010101010",
  28482=>"001001010",
  28483=>"101000101",
  28484=>"000110111",
  28485=>"110000101",
  28486=>"111101110",
  28487=>"110010100",
  28488=>"100011110",
  28489=>"111110011",
  28490=>"001000100",
  28491=>"101010111",
  28492=>"001001101",
  28493=>"010001010",
  28494=>"111010010",
  28495=>"001010001",
  28496=>"001100010",
  28497=>"010100111",
  28498=>"110111101",
  28499=>"001001000",
  28500=>"111101010",
  28501=>"001100010",
  28502=>"010111001",
  28503=>"011011011",
  28504=>"010010111",
  28505=>"011010000",
  28506=>"110011001",
  28507=>"110110110",
  28508=>"110011111",
  28509=>"100001011",
  28510=>"000100001",
  28511=>"111010000",
  28512=>"110110111",
  28513=>"000011111",
  28514=>"100111111",
  28515=>"011110100",
  28516=>"000011101",
  28517=>"001111010",
  28518=>"010110110",
  28519=>"001011011",
  28520=>"101000100",
  28521=>"011110011",
  28522=>"000100110",
  28523=>"011000010",
  28524=>"010011101",
  28525=>"101001100",
  28526=>"011001111",
  28527=>"001100111",
  28528=>"101001111",
  28529=>"101001110",
  28530=>"111111100",
  28531=>"111100010",
  28532=>"000101111",
  28533=>"110111011",
  28534=>"101000111",
  28535=>"000001100",
  28536=>"101110000",
  28537=>"111110010",
  28538=>"111010101",
  28539=>"110111101",
  28540=>"101100111",
  28541=>"110100111",
  28542=>"000111010",
  28543=>"010100101",
  28544=>"110111000",
  28545=>"001000000",
  28546=>"110001010",
  28547=>"110000011",
  28548=>"100100001",
  28549=>"110101011",
  28550=>"011010001",
  28551=>"111111100",
  28552=>"111110110",
  28553=>"010010001",
  28554=>"111010001",
  28555=>"110011100",
  28556=>"100001011",
  28557=>"011010000",
  28558=>"100001001",
  28559=>"110011011",
  28560=>"000110011",
  28561=>"000000011",
  28562=>"000100101",
  28563=>"010011010",
  28564=>"101100100",
  28565=>"011011000",
  28566=>"000110011",
  28567=>"000011011",
  28568=>"100111110",
  28569=>"010001000",
  28570=>"011011100",
  28571=>"010001010",
  28572=>"010000000",
  28573=>"111010111",
  28574=>"111000000",
  28575=>"111000100",
  28576=>"100001110",
  28577=>"111100100",
  28578=>"111111111",
  28579=>"100011110",
  28580=>"010111110",
  28581=>"101000011",
  28582=>"011100011",
  28583=>"001000000",
  28584=>"011011101",
  28585=>"100101000",
  28586=>"111110001",
  28587=>"101010100",
  28588=>"111111100",
  28589=>"111001010",
  28590=>"001110111",
  28591=>"011101011",
  28592=>"011111001",
  28593=>"001111001",
  28594=>"010100111",
  28595=>"011100110",
  28596=>"000010111",
  28597=>"110000100",
  28598=>"111101000",
  28599=>"111100101",
  28600=>"001001101",
  28601=>"011110101",
  28602=>"010010010",
  28603=>"001110000",
  28604=>"000100010",
  28605=>"011010001",
  28606=>"001110101",
  28607=>"001110010",
  28608=>"000101000",
  28609=>"111100011",
  28610=>"000100100",
  28611=>"000010110",
  28612=>"101010000",
  28613=>"010110110",
  28614=>"000101111",
  28615=>"010111001",
  28616=>"000111111",
  28617=>"011100011",
  28618=>"000000111",
  28619=>"101010001",
  28620=>"111101111",
  28621=>"111000111",
  28622=>"101101100",
  28623=>"101000000",
  28624=>"111011111",
  28625=>"001100000",
  28626=>"011111001",
  28627=>"100011010",
  28628=>"110111111",
  28629=>"111100010",
  28630=>"100110110",
  28631=>"100111000",
  28632=>"001011111",
  28633=>"011011111",
  28634=>"001001100",
  28635=>"001110010",
  28636=>"011111100",
  28637=>"111110101",
  28638=>"011000111",
  28639=>"001000001",
  28640=>"001000001",
  28641=>"111001001",
  28642=>"101001010",
  28643=>"001001010",
  28644=>"111001011",
  28645=>"111010001",
  28646=>"101000100",
  28647=>"101101110",
  28648=>"010011001",
  28649=>"101101001",
  28650=>"001110110",
  28651=>"001101110",
  28652=>"011111001",
  28653=>"010100110",
  28654=>"100010010",
  28655=>"101000010",
  28656=>"000100100",
  28657=>"000001101",
  28658=>"111100100",
  28659=>"010010011",
  28660=>"011111111",
  28661=>"000111110",
  28662=>"111110100",
  28663=>"001000001",
  28664=>"011001111",
  28665=>"111110100",
  28666=>"010001000",
  28667=>"100010000",
  28668=>"000000011",
  28669=>"011111001",
  28670=>"111000100",
  28671=>"111010100",
  28672=>"101111100",
  28673=>"000001101",
  28674=>"010010100",
  28675=>"110010111",
  28676=>"000000101",
  28677=>"101101011",
  28678=>"001001001",
  28679=>"100000111",
  28680=>"010100101",
  28681=>"000001100",
  28682=>"001011111",
  28683=>"100111111",
  28684=>"100110011",
  28685=>"110011110",
  28686=>"111010001",
  28687=>"000111000",
  28688=>"100100001",
  28689=>"001110101",
  28690=>"111011110",
  28691=>"010100000",
  28692=>"001110100",
  28693=>"110000000",
  28694=>"111001111",
  28695=>"010100111",
  28696=>"101100011",
  28697=>"100100100",
  28698=>"110100100",
  28699=>"000011111",
  28700=>"110001001",
  28701=>"101000011",
  28702=>"000110110",
  28703=>"011101000",
  28704=>"010101000",
  28705=>"011100111",
  28706=>"001000100",
  28707=>"101100100",
  28708=>"011011010",
  28709=>"100110011",
  28710=>"001100100",
  28711=>"010010100",
  28712=>"011110100",
  28713=>"001011011",
  28714=>"110111000",
  28715=>"101101000",
  28716=>"010101100",
  28717=>"000111101",
  28718=>"011101110",
  28719=>"110000000",
  28720=>"111111111",
  28721=>"110001001",
  28722=>"001000001",
  28723=>"111011111",
  28724=>"001000010",
  28725=>"000101011",
  28726=>"101101000",
  28727=>"010000101",
  28728=>"100000100",
  28729=>"010110101",
  28730=>"111001001",
  28731=>"110011000",
  28732=>"000000000",
  28733=>"100010110",
  28734=>"001011100",
  28735=>"011100000",
  28736=>"011100010",
  28737=>"110100000",
  28738=>"001000010",
  28739=>"011101000",
  28740=>"001010110",
  28741=>"001100010",
  28742=>"100100101",
  28743=>"011100000",
  28744=>"101111100",
  28745=>"110000101",
  28746=>"000111101",
  28747=>"010001100",
  28748=>"101101101",
  28749=>"000110110",
  28750=>"111111000",
  28751=>"001010010",
  28752=>"011110011",
  28753=>"100001100",
  28754=>"111111101",
  28755=>"110110111",
  28756=>"111111111",
  28757=>"101100000",
  28758=>"011010000",
  28759=>"001011101",
  28760=>"100101011",
  28761=>"011100000",
  28762=>"110100000",
  28763=>"001100101",
  28764=>"001010100",
  28765=>"100011111",
  28766=>"110100111",
  28767=>"010100000",
  28768=>"001001011",
  28769=>"110100100",
  28770=>"111110111",
  28771=>"010010001",
  28772=>"011101111",
  28773=>"111111110",
  28774=>"001111000",
  28775=>"011110100",
  28776=>"011110100",
  28777=>"001110000",
  28778=>"010111010",
  28779=>"100010101",
  28780=>"011001010",
  28781=>"001010100",
  28782=>"011000101",
  28783=>"100000110",
  28784=>"011000001",
  28785=>"000001010",
  28786=>"011001000",
  28787=>"101101011",
  28788=>"010000111",
  28789=>"010010100",
  28790=>"101001000",
  28791=>"110101110",
  28792=>"001110010",
  28793=>"010110011",
  28794=>"000111000",
  28795=>"000100010",
  28796=>"010001111",
  28797=>"101111101",
  28798=>"110100110",
  28799=>"010100010",
  28800=>"000100011",
  28801=>"011100101",
  28802=>"000101111",
  28803=>"000001001",
  28804=>"111101110",
  28805=>"011111101",
  28806=>"100101011",
  28807=>"100100010",
  28808=>"110111001",
  28809=>"101111111",
  28810=>"001000010",
  28811=>"010011110",
  28812=>"001110001",
  28813=>"100111011",
  28814=>"000110100",
  28815=>"101010001",
  28816=>"000010000",
  28817=>"101110000",
  28818=>"100111100",
  28819=>"100101111",
  28820=>"110001000",
  28821=>"111100101",
  28822=>"001000101",
  28823=>"010011101",
  28824=>"110101010",
  28825=>"101011001",
  28826=>"000000111",
  28827=>"110001011",
  28828=>"000001110",
  28829=>"100110100",
  28830=>"110101100",
  28831=>"001100001",
  28832=>"101111001",
  28833=>"101011011",
  28834=>"111110110",
  28835=>"111010100",
  28836=>"111101101",
  28837=>"000111001",
  28838=>"100110100",
  28839=>"011010100",
  28840=>"011010011",
  28841=>"001011011",
  28842=>"000000111",
  28843=>"110100100",
  28844=>"111100001",
  28845=>"111101110",
  28846=>"010011011",
  28847=>"101101110",
  28848=>"011001001",
  28849=>"101000010",
  28850=>"111011011",
  28851=>"000000101",
  28852=>"000010110",
  28853=>"111100110",
  28854=>"001101110",
  28855=>"100111111",
  28856=>"110000101",
  28857=>"101101001",
  28858=>"010001010",
  28859=>"101010001",
  28860=>"011001100",
  28861=>"011010000",
  28862=>"100010000",
  28863=>"110000001",
  28864=>"001100000",
  28865=>"000000010",
  28866=>"111100000",
  28867=>"011111111",
  28868=>"010011000",
  28869=>"001100101",
  28870=>"001011011",
  28871=>"100101010",
  28872=>"110111101",
  28873=>"111000011",
  28874=>"111000001",
  28875=>"111000001",
  28876=>"010010011",
  28877=>"010111111",
  28878=>"010011011",
  28879=>"101101100",
  28880=>"100000001",
  28881=>"010100000",
  28882=>"100110101",
  28883=>"011000011",
  28884=>"001010111",
  28885=>"010100110",
  28886=>"100001010",
  28887=>"000011100",
  28888=>"110111100",
  28889=>"000011100",
  28890=>"100011010",
  28891=>"110000000",
  28892=>"011001111",
  28893=>"001100100",
  28894=>"000001100",
  28895=>"011110011",
  28896=>"110101001",
  28897=>"101100110",
  28898=>"111011101",
  28899=>"001101111",
  28900=>"101101101",
  28901=>"111010000",
  28902=>"110110001",
  28903=>"000001111",
  28904=>"001001010",
  28905=>"011111100",
  28906=>"011001111",
  28907=>"011001111",
  28908=>"111001000",
  28909=>"101011110",
  28910=>"001010110",
  28911=>"010101110",
  28912=>"011001010",
  28913=>"101010111",
  28914=>"101000010",
  28915=>"011101000",
  28916=>"101100100",
  28917=>"110111011",
  28918=>"001000010",
  28919=>"010111001",
  28920=>"100101001",
  28921=>"110110001",
  28922=>"100010100",
  28923=>"101100100",
  28924=>"101000110",
  28925=>"010101011",
  28926=>"111101010",
  28927=>"100010100",
  28928=>"010010111",
  28929=>"011110000",
  28930=>"001000110",
  28931=>"100001011",
  28932=>"110011111",
  28933=>"101100110",
  28934=>"001000011",
  28935=>"101110010",
  28936=>"110000000",
  28937=>"010111101",
  28938=>"110111110",
  28939=>"010000001",
  28940=>"010010011",
  28941=>"100111011",
  28942=>"100000011",
  28943=>"000100110",
  28944=>"110110111",
  28945=>"110011010",
  28946=>"100111110",
  28947=>"101000010",
  28948=>"010100011",
  28949=>"111001010",
  28950=>"000000010",
  28951=>"100011000",
  28952=>"000000000",
  28953=>"110001011",
  28954=>"101011001",
  28955=>"001000110",
  28956=>"011110101",
  28957=>"111100011",
  28958=>"011111100",
  28959=>"110001010",
  28960=>"111110111",
  28961=>"011000110",
  28962=>"111000001",
  28963=>"000110001",
  28964=>"100110110",
  28965=>"010001110",
  28966=>"010100100",
  28967=>"111101001",
  28968=>"000001000",
  28969=>"001001000",
  28970=>"010111111",
  28971=>"010101010",
  28972=>"010010001",
  28973=>"011111111",
  28974=>"000000000",
  28975=>"101011111",
  28976=>"111100110",
  28977=>"001111010",
  28978=>"000010001",
  28979=>"111011101",
  28980=>"111100011",
  28981=>"001001100",
  28982=>"001101000",
  28983=>"111010110",
  28984=>"000101110",
  28985=>"010011111",
  28986=>"100101101",
  28987=>"111011011",
  28988=>"101011110",
  28989=>"111101001",
  28990=>"110100100",
  28991=>"010001011",
  28992=>"111111110",
  28993=>"000010101",
  28994=>"010101010",
  28995=>"011101001",
  28996=>"110111011",
  28997=>"000011011",
  28998=>"101011000",
  28999=>"000100000",
  29000=>"110001100",
  29001=>"000000001",
  29002=>"101010101",
  29003=>"100000010",
  29004=>"010101101",
  29005=>"000101110",
  29006=>"000000111",
  29007=>"101010000",
  29008=>"011110110",
  29009=>"011010101",
  29010=>"011010111",
  29011=>"101001110",
  29012=>"100101101",
  29013=>"111011111",
  29014=>"001100000",
  29015=>"110000000",
  29016=>"011100111",
  29017=>"011111101",
  29018=>"110101010",
  29019=>"001000001",
  29020=>"010101011",
  29021=>"000111010",
  29022=>"111000110",
  29023=>"111000110",
  29024=>"101001001",
  29025=>"110010010",
  29026=>"010100010",
  29027=>"111110101",
  29028=>"110111111",
  29029=>"011110111",
  29030=>"000001001",
  29031=>"110111101",
  29032=>"000000110",
  29033=>"011101101",
  29034=>"110001011",
  29035=>"001110001",
  29036=>"100000110",
  29037=>"011010011",
  29038=>"010111110",
  29039=>"101011111",
  29040=>"111010101",
  29041=>"001100101",
  29042=>"101001000",
  29043=>"010011101",
  29044=>"100100011",
  29045=>"110110000",
  29046=>"100011010",
  29047=>"000001111",
  29048=>"101111101",
  29049=>"011001100",
  29050=>"010101010",
  29051=>"001100110",
  29052=>"101100111",
  29053=>"011000101",
  29054=>"110111111",
  29055=>"100001100",
  29056=>"010011010",
  29057=>"000100011",
  29058=>"110111011",
  29059=>"110110101",
  29060=>"101110010",
  29061=>"100011100",
  29062=>"101000010",
  29063=>"000001111",
  29064=>"001011000",
  29065=>"011101101",
  29066=>"010101001",
  29067=>"000101001",
  29068=>"000100000",
  29069=>"111011011",
  29070=>"100111001",
  29071=>"101011100",
  29072=>"011100000",
  29073=>"011010100",
  29074=>"001001110",
  29075=>"111110110",
  29076=>"101001110",
  29077=>"011000010",
  29078=>"110101101",
  29079=>"001001011",
  29080=>"101101010",
  29081=>"111011001",
  29082=>"001000111",
  29083=>"010100110",
  29084=>"101111011",
  29085=>"101101000",
  29086=>"111110110",
  29087=>"010000010",
  29088=>"111111101",
  29089=>"010001001",
  29090=>"011110100",
  29091=>"000100011",
  29092=>"110000000",
  29093=>"011000110",
  29094=>"111001110",
  29095=>"101111101",
  29096=>"010101010",
  29097=>"101001111",
  29098=>"101101000",
  29099=>"101111100",
  29100=>"110110101",
  29101=>"010110001",
  29102=>"110101101",
  29103=>"011011101",
  29104=>"101001100",
  29105=>"111000100",
  29106=>"000100100",
  29107=>"001001010",
  29108=>"011101101",
  29109=>"011100001",
  29110=>"110010101",
  29111=>"011101101",
  29112=>"111000001",
  29113=>"011011110",
  29114=>"101000010",
  29115=>"100000001",
  29116=>"100001000",
  29117=>"111111100",
  29118=>"100101010",
  29119=>"110110101",
  29120=>"001010111",
  29121=>"100101011",
  29122=>"011100010",
  29123=>"010111100",
  29124=>"011001001",
  29125=>"111110000",
  29126=>"000100010",
  29127=>"010100100",
  29128=>"111100010",
  29129=>"100011010",
  29130=>"010010000",
  29131=>"101000111",
  29132=>"011101011",
  29133=>"101011000",
  29134=>"010101001",
  29135=>"100110000",
  29136=>"111001000",
  29137=>"010111111",
  29138=>"000110011",
  29139=>"000100101",
  29140=>"010111111",
  29141=>"000011010",
  29142=>"111010110",
  29143=>"001110100",
  29144=>"111101001",
  29145=>"110001111",
  29146=>"000001110",
  29147=>"011000110",
  29148=>"101110111",
  29149=>"010000100",
  29150=>"101110010",
  29151=>"010110100",
  29152=>"011111111",
  29153=>"110110000",
  29154=>"101110010",
  29155=>"101000001",
  29156=>"001100100",
  29157=>"000000110",
  29158=>"101011110",
  29159=>"000100101",
  29160=>"011011011",
  29161=>"110101110",
  29162=>"100101000",
  29163=>"110001011",
  29164=>"010010001",
  29165=>"100010010",
  29166=>"111011011",
  29167=>"010001000",
  29168=>"110111000",
  29169=>"111001000",
  29170=>"111011000",
  29171=>"011010100",
  29172=>"000010000",
  29173=>"101000100",
  29174=>"111100011",
  29175=>"110010100",
  29176=>"000101101",
  29177=>"001100010",
  29178=>"110000100",
  29179=>"001110011",
  29180=>"000011111",
  29181=>"000100011",
  29182=>"110110100",
  29183=>"111110110",
  29184=>"111010100",
  29185=>"011110011",
  29186=>"100110110",
  29187=>"100101101",
  29188=>"101001000",
  29189=>"000001011",
  29190=>"110101001",
  29191=>"000000100",
  29192=>"000010111",
  29193=>"000110011",
  29194=>"101101110",
  29195=>"110111011",
  29196=>"100011101",
  29197=>"100000000",
  29198=>"001011000",
  29199=>"010101010",
  29200=>"001010100",
  29201=>"001100101",
  29202=>"010110011",
  29203=>"101000111",
  29204=>"011011001",
  29205=>"000001001",
  29206=>"100111001",
  29207=>"101101111",
  29208=>"100000111",
  29209=>"001111111",
  29210=>"011000100",
  29211=>"110000011",
  29212=>"100000000",
  29213=>"011110111",
  29214=>"011000001",
  29215=>"110111101",
  29216=>"000010001",
  29217=>"111011001",
  29218=>"010000011",
  29219=>"101100110",
  29220=>"001010101",
  29221=>"111001101",
  29222=>"100101010",
  29223=>"110010110",
  29224=>"111100100",
  29225=>"001100011",
  29226=>"100000000",
  29227=>"001011010",
  29228=>"001000100",
  29229=>"001100010",
  29230=>"000010000",
  29231=>"000001001",
  29232=>"000011001",
  29233=>"010111001",
  29234=>"110111100",
  29235=>"101101110",
  29236=>"011011001",
  29237=>"011011101",
  29238=>"000011100",
  29239=>"111010110",
  29240=>"001100111",
  29241=>"001111000",
  29242=>"001000001",
  29243=>"001111010",
  29244=>"010011111",
  29245=>"110001100",
  29246=>"001011111",
  29247=>"110001100",
  29248=>"001011001",
  29249=>"110000000",
  29250=>"001100101",
  29251=>"001110110",
  29252=>"000011000",
  29253=>"011100110",
  29254=>"010100111",
  29255=>"101111011",
  29256=>"010000000",
  29257=>"101101001",
  29258=>"000001000",
  29259=>"000111000",
  29260=>"001011011",
  29261=>"000110000",
  29262=>"001000101",
  29263=>"111000111",
  29264=>"001000100",
  29265=>"100011000",
  29266=>"000110110",
  29267=>"110110101",
  29268=>"111110001",
  29269=>"110010100",
  29270=>"111000000",
  29271=>"001101101",
  29272=>"101100111",
  29273=>"010010001",
  29274=>"001110000",
  29275=>"100001000",
  29276=>"000000000",
  29277=>"110110110",
  29278=>"010111000",
  29279=>"001001110",
  29280=>"101000010",
  29281=>"101011100",
  29282=>"000001110",
  29283=>"000100001",
  29284=>"010010000",
  29285=>"111010110",
  29286=>"000111111",
  29287=>"010100010",
  29288=>"110000011",
  29289=>"000010110",
  29290=>"011010010",
  29291=>"101100101",
  29292=>"100000010",
  29293=>"111111111",
  29294=>"100011011",
  29295=>"101111000",
  29296=>"011001000",
  29297=>"101011001",
  29298=>"110100010",
  29299=>"010011000",
  29300=>"101001101",
  29301=>"111110000",
  29302=>"111111000",
  29303=>"011110010",
  29304=>"110111100",
  29305=>"011000001",
  29306=>"101000010",
  29307=>"001011011",
  29308=>"000001010",
  29309=>"001000011",
  29310=>"101001111",
  29311=>"010101010",
  29312=>"111001100",
  29313=>"001110001",
  29314=>"010110010",
  29315=>"111101111",
  29316=>"011110000",
  29317=>"010101000",
  29318=>"001101110",
  29319=>"010101010",
  29320=>"110000110",
  29321=>"100000000",
  29322=>"110111110",
  29323=>"101011001",
  29324=>"101111111",
  29325=>"111100010",
  29326=>"011001010",
  29327=>"101101101",
  29328=>"111000100",
  29329=>"100010110",
  29330=>"110110101",
  29331=>"111101001",
  29332=>"000100100",
  29333=>"111001000",
  29334=>"001011101",
  29335=>"111011000",
  29336=>"101111101",
  29337=>"111001100",
  29338=>"001010100",
  29339=>"011101000",
  29340=>"010101100",
  29341=>"100111100",
  29342=>"011010100",
  29343=>"111101010",
  29344=>"011000101",
  29345=>"111101001",
  29346=>"000111001",
  29347=>"011010001",
  29348=>"101011001",
  29349=>"100110110",
  29350=>"100110001",
  29351=>"000000001",
  29352=>"100100110",
  29353=>"000010100",
  29354=>"000101101",
  29355=>"001100100",
  29356=>"001000011",
  29357=>"011111110",
  29358=>"010011110",
  29359=>"010001010",
  29360=>"000110111",
  29361=>"111001000",
  29362=>"111010100",
  29363=>"011001011",
  29364=>"111000001",
  29365=>"001000001",
  29366=>"010111100",
  29367=>"000101001",
  29368=>"110110111",
  29369=>"101110100",
  29370=>"110101111",
  29371=>"100110101",
  29372=>"101101001",
  29373=>"001111101",
  29374=>"101010101",
  29375=>"100101011",
  29376=>"010100111",
  29377=>"010111111",
  29378=>"001011011",
  29379=>"011110111",
  29380=>"101010101",
  29381=>"000111100",
  29382=>"100100001",
  29383=>"010111000",
  29384=>"000000100",
  29385=>"011001010",
  29386=>"010000101",
  29387=>"001001100",
  29388=>"001010011",
  29389=>"000000111",
  29390=>"111110011",
  29391=>"100010100",
  29392=>"101111111",
  29393=>"000111111",
  29394=>"110000110",
  29395=>"000001011",
  29396=>"011111111",
  29397=>"101111111",
  29398=>"010000001",
  29399=>"111010010",
  29400=>"000100000",
  29401=>"000100010",
  29402=>"111000110",
  29403=>"001001000",
  29404=>"011011010",
  29405=>"101001100",
  29406=>"000010100",
  29407=>"100111001",
  29408=>"011111100",
  29409=>"011111101",
  29410=>"110000101",
  29411=>"011001010",
  29412=>"001000100",
  29413=>"110001010",
  29414=>"000100100",
  29415=>"011110101",
  29416=>"001011100",
  29417=>"001101000",
  29418=>"001001010",
  29419=>"010001100",
  29420=>"001000001",
  29421=>"010100010",
  29422=>"100000010",
  29423=>"110101110",
  29424=>"111001011",
  29425=>"111101100",
  29426=>"101100100",
  29427=>"011001011",
  29428=>"001110111",
  29429=>"000000101",
  29430=>"010010101",
  29431=>"111101000",
  29432=>"111010100",
  29433=>"000000000",
  29434=>"001011001",
  29435=>"001000010",
  29436=>"001111011",
  29437=>"100110111",
  29438=>"000100111",
  29439=>"001100001",
  29440=>"101111101",
  29441=>"010001001",
  29442=>"011001110",
  29443=>"110111111",
  29444=>"000111010",
  29445=>"110100101",
  29446=>"010110001",
  29447=>"110101001",
  29448=>"100100010",
  29449=>"000110001",
  29450=>"000001111",
  29451=>"000100011",
  29452=>"011000001",
  29453=>"010011010",
  29454=>"100101101",
  29455=>"001100001",
  29456=>"110001100",
  29457=>"000100110",
  29458=>"010011110",
  29459=>"001111101",
  29460=>"010110101",
  29461=>"000000110",
  29462=>"000100000",
  29463=>"010000010",
  29464=>"001011000",
  29465=>"111001000",
  29466=>"000110010",
  29467=>"110101111",
  29468=>"001011000",
  29469=>"000001100",
  29470=>"101001110",
  29471=>"011111101",
  29472=>"101110110",
  29473=>"000101010",
  29474=>"011010110",
  29475=>"000100010",
  29476=>"110100011",
  29477=>"000001011",
  29478=>"010001110",
  29479=>"011001001",
  29480=>"011111011",
  29481=>"000100000",
  29482=>"111101110",
  29483=>"001001101",
  29484=>"101001100",
  29485=>"001101101",
  29486=>"100001011",
  29487=>"110101111",
  29488=>"001100110",
  29489=>"000100000",
  29490=>"011101001",
  29491=>"110010010",
  29492=>"001010111",
  29493=>"011111011",
  29494=>"000101100",
  29495=>"100001011",
  29496=>"010100111",
  29497=>"101101100",
  29498=>"001000111",
  29499=>"001110001",
  29500=>"001010101",
  29501=>"100000110",
  29502=>"001010111",
  29503=>"111001101",
  29504=>"010110010",
  29505=>"100000100",
  29506=>"000000110",
  29507=>"100010010",
  29508=>"001100100",
  29509=>"011111101",
  29510=>"110101001",
  29511=>"001101100",
  29512=>"101000010",
  29513=>"000000101",
  29514=>"111101110",
  29515=>"000000011",
  29516=>"011110001",
  29517=>"110011101",
  29518=>"001011100",
  29519=>"001010000",
  29520=>"100111110",
  29521=>"000011101",
  29522=>"100101000",
  29523=>"010101111",
  29524=>"000011110",
  29525=>"010100001",
  29526=>"001101000",
  29527=>"111110101",
  29528=>"111110010",
  29529=>"101101010",
  29530=>"000001001",
  29531=>"101011111",
  29532=>"110010000",
  29533=>"110011011",
  29534=>"011001011",
  29535=>"100011000",
  29536=>"000011111",
  29537=>"001001000",
  29538=>"011100100",
  29539=>"000100001",
  29540=>"001010010",
  29541=>"001100011",
  29542=>"100111110",
  29543=>"100101110",
  29544=>"010100111",
  29545=>"100011011",
  29546=>"111001011",
  29547=>"110010110",
  29548=>"111001110",
  29549=>"001000101",
  29550=>"100000110",
  29551=>"111001111",
  29552=>"111101100",
  29553=>"110001110",
  29554=>"000111011",
  29555=>"111110100",
  29556=>"001100100",
  29557=>"111000010",
  29558=>"100110011",
  29559=>"100111101",
  29560=>"001111011",
  29561=>"100011101",
  29562=>"110000000",
  29563=>"000100110",
  29564=>"000000111",
  29565=>"001010101",
  29566=>"111100100",
  29567=>"010101111",
  29568=>"100100000",
  29569=>"110000100",
  29570=>"100000101",
  29571=>"101001100",
  29572=>"000010110",
  29573=>"111010011",
  29574=>"101000011",
  29575=>"010100111",
  29576=>"100000001",
  29577=>"011010000",
  29578=>"000010111",
  29579=>"101000101",
  29580=>"011001110",
  29581=>"110001000",
  29582=>"001011000",
  29583=>"101000101",
  29584=>"111110000",
  29585=>"111110111",
  29586=>"001111100",
  29587=>"110000111",
  29588=>"100011001",
  29589=>"101110101",
  29590=>"000001111",
  29591=>"011101100",
  29592=>"101010000",
  29593=>"100101000",
  29594=>"010111011",
  29595=>"010111100",
  29596=>"011100001",
  29597=>"101111101",
  29598=>"111000011",
  29599=>"010011000",
  29600=>"000101000",
  29601=>"011111100",
  29602=>"001010010",
  29603=>"110011001",
  29604=>"011111100",
  29605=>"111110110",
  29606=>"000010110",
  29607=>"001010010",
  29608=>"011110001",
  29609=>"101101011",
  29610=>"100101011",
  29611=>"101111100",
  29612=>"001000110",
  29613=>"100011111",
  29614=>"111011010",
  29615=>"101111100",
  29616=>"110010110",
  29617=>"000001111",
  29618=>"011011101",
  29619=>"100001001",
  29620=>"000110010",
  29621=>"001111100",
  29622=>"101110100",
  29623=>"001111001",
  29624=>"000101001",
  29625=>"101110000",
  29626=>"000110001",
  29627=>"010001110",
  29628=>"001011011",
  29629=>"001001010",
  29630=>"101100100",
  29631=>"000110101",
  29632=>"101110001",
  29633=>"001011011",
  29634=>"100111111",
  29635=>"011001111",
  29636=>"100001001",
  29637=>"110001111",
  29638=>"101110111",
  29639=>"000111111",
  29640=>"000011100",
  29641=>"011000101",
  29642=>"010101111",
  29643=>"001011101",
  29644=>"011001100",
  29645=>"010100000",
  29646=>"000011010",
  29647=>"001101001",
  29648=>"001101110",
  29649=>"001010000",
  29650=>"101000000",
  29651=>"110111101",
  29652=>"101100110",
  29653=>"000011101",
  29654=>"000001111",
  29655=>"110001100",
  29656=>"111110010",
  29657=>"110111110",
  29658=>"010001000",
  29659=>"100001001",
  29660=>"000001001",
  29661=>"111101001",
  29662=>"000010001",
  29663=>"000100100",
  29664=>"100100011",
  29665=>"101011111",
  29666=>"101001001",
  29667=>"001110010",
  29668=>"010001110",
  29669=>"000101111",
  29670=>"110100110",
  29671=>"101000011",
  29672=>"001101110",
  29673=>"010000101",
  29674=>"110110001",
  29675=>"011000100",
  29676=>"100001010",
  29677=>"000110100",
  29678=>"000010100",
  29679=>"111010011",
  29680=>"000001100",
  29681=>"010101101",
  29682=>"011001111",
  29683=>"100100111",
  29684=>"101101011",
  29685=>"010011000",
  29686=>"100011000",
  29687=>"100101011",
  29688=>"001011010",
  29689=>"010111111",
  29690=>"101000010",
  29691=>"100000010",
  29692=>"001101100",
  29693=>"011111111",
  29694=>"111000011",
  29695=>"111111000",
  29696=>"010000011",
  29697=>"000010111",
  29698=>"101110011",
  29699=>"100000110",
  29700=>"101101000",
  29701=>"110110010",
  29702=>"011011010",
  29703=>"001011010",
  29704=>"110000010",
  29705=>"110000001",
  29706=>"111101100",
  29707=>"100001010",
  29708=>"001111000",
  29709=>"111000110",
  29710=>"011110110",
  29711=>"000110000",
  29712=>"000101000",
  29713=>"000000010",
  29714=>"011100111",
  29715=>"100111001",
  29716=>"111011000",
  29717=>"110110110",
  29718=>"101100001",
  29719=>"100101101",
  29720=>"110011111",
  29721=>"100100110",
  29722=>"111111000",
  29723=>"011111110",
  29724=>"101011111",
  29725=>"011101101",
  29726=>"101001001",
  29727=>"111111111",
  29728=>"001000000",
  29729=>"111101011",
  29730=>"101111011",
  29731=>"001101110",
  29732=>"010110000",
  29733=>"100110101",
  29734=>"111011111",
  29735=>"001110100",
  29736=>"110011000",
  29737=>"110101000",
  29738=>"111101010",
  29739=>"111111010",
  29740=>"010101101",
  29741=>"000110110",
  29742=>"010111110",
  29743=>"010011010",
  29744=>"100110110",
  29745=>"101001101",
  29746=>"000010110",
  29747=>"001100111",
  29748=>"010010011",
  29749=>"011110011",
  29750=>"011100111",
  29751=>"100001111",
  29752=>"010100100",
  29753=>"100010010",
  29754=>"001001110",
  29755=>"111011011",
  29756=>"000111000",
  29757=>"010010001",
  29758=>"001110000",
  29759=>"101101111",
  29760=>"001101110",
  29761=>"011111000",
  29762=>"101100000",
  29763=>"000110101",
  29764=>"000100001",
  29765=>"110010011",
  29766=>"001001100",
  29767=>"001001100",
  29768=>"101101111",
  29769=>"000101110",
  29770=>"010111000",
  29771=>"011101001",
  29772=>"101111010",
  29773=>"100101001",
  29774=>"000110001",
  29775=>"110100001",
  29776=>"000001000",
  29777=>"110101110",
  29778=>"011111100",
  29779=>"010000101",
  29780=>"111111001",
  29781=>"010110111",
  29782=>"011100111",
  29783=>"100010011",
  29784=>"100111101",
  29785=>"001101001",
  29786=>"100011101",
  29787=>"000101010",
  29788=>"010011100",
  29789=>"111001111",
  29790=>"111010010",
  29791=>"110010110",
  29792=>"010100011",
  29793=>"111000011",
  29794=>"001011111",
  29795=>"010010101",
  29796=>"100100101",
  29797=>"001011101",
  29798=>"000100011",
  29799=>"111101011",
  29800=>"010011111",
  29801=>"011101000",
  29802=>"001010110",
  29803=>"100011110",
  29804=>"100111000",
  29805=>"010001011",
  29806=>"111001010",
  29807=>"100100100",
  29808=>"111111011",
  29809=>"111110011",
  29810=>"010111001",
  29811=>"101111111",
  29812=>"011011101",
  29813=>"010010010",
  29814=>"011001001",
  29815=>"110000001",
  29816=>"000110010",
  29817=>"101111010",
  29818=>"100011111",
  29819=>"000000110",
  29820=>"100001100",
  29821=>"001001001",
  29822=>"011001011",
  29823=>"111011110",
  29824=>"010001011",
  29825=>"010101000",
  29826=>"000100101",
  29827=>"101000101",
  29828=>"000011011",
  29829=>"011111111",
  29830=>"011001111",
  29831=>"000110010",
  29832=>"000001011",
  29833=>"111100010",
  29834=>"110011110",
  29835=>"100010010",
  29836=>"001111110",
  29837=>"011111001",
  29838=>"000100101",
  29839=>"011000001",
  29840=>"100110110",
  29841=>"010111100",
  29842=>"001001111",
  29843=>"111110010",
  29844=>"100010001",
  29845=>"100100111",
  29846=>"000000001",
  29847=>"110011111",
  29848=>"011000110",
  29849=>"100011111",
  29850=>"100111101",
  29851=>"110110111",
  29852=>"100101111",
  29853=>"010011010",
  29854=>"001100000",
  29855=>"101010101",
  29856=>"001100001",
  29857=>"110111010",
  29858=>"100110100",
  29859=>"111101000",
  29860=>"111110110",
  29861=>"111100101",
  29862=>"010011001",
  29863=>"010000001",
  29864=>"101111100",
  29865=>"110100111",
  29866=>"110100000",
  29867=>"010110101",
  29868=>"010110100",
  29869=>"001001011",
  29870=>"001101001",
  29871=>"000001000",
  29872=>"001000000",
  29873=>"011100100",
  29874=>"011001000",
  29875=>"010100010",
  29876=>"101000010",
  29877=>"011001000",
  29878=>"110110100",
  29879=>"010110010",
  29880=>"010001001",
  29881=>"010001111",
  29882=>"001001100",
  29883=>"000111101",
  29884=>"110111101",
  29885=>"101000111",
  29886=>"111101100",
  29887=>"110110101",
  29888=>"110100001",
  29889=>"000010110",
  29890=>"110000101",
  29891=>"100100010",
  29892=>"001101000",
  29893=>"010011101",
  29894=>"110111010",
  29895=>"011000010",
  29896=>"001000110",
  29897=>"000000000",
  29898=>"000011001",
  29899=>"011111010",
  29900=>"101110011",
  29901=>"011100111",
  29902=>"110101001",
  29903=>"000001100",
  29904=>"100000010",
  29905=>"010001011",
  29906=>"010100001",
  29907=>"010111101",
  29908=>"100001010",
  29909=>"001011001",
  29910=>"111001101",
  29911=>"111011001",
  29912=>"000011011",
  29913=>"110110100",
  29914=>"010000100",
  29915=>"110001110",
  29916=>"111011001",
  29917=>"011101000",
  29918=>"000010001",
  29919=>"000000010",
  29920=>"000110000",
  29921=>"000011100",
  29922=>"011110010",
  29923=>"100001000",
  29924=>"101100000",
  29925=>"110001010",
  29926=>"000000101",
  29927=>"000000110",
  29928=>"001010001",
  29929=>"000101001",
  29930=>"100001001",
  29931=>"011111101",
  29932=>"011001010",
  29933=>"000011001",
  29934=>"111101001",
  29935=>"011100001",
  29936=>"111111001",
  29937=>"111110101",
  29938=>"110001010",
  29939=>"100011101",
  29940=>"101000101",
  29941=>"100011000",
  29942=>"110101111",
  29943=>"010101101",
  29944=>"100111000",
  29945=>"111100111",
  29946=>"100001001",
  29947=>"110010000",
  29948=>"110001101",
  29949=>"001111110",
  29950=>"010011001",
  29951=>"000010101",
  29952=>"111001110",
  29953=>"110100111",
  29954=>"110100110",
  29955=>"101010000",
  29956=>"100011111",
  29957=>"101000111",
  29958=>"011011111",
  29959=>"011110100",
  29960=>"011000111",
  29961=>"001000111",
  29962=>"010010000",
  29963=>"010101111",
  29964=>"001011110",
  29965=>"001010110",
  29966=>"010001011",
  29967=>"000010010",
  29968=>"010100100",
  29969=>"010011000",
  29970=>"100000110",
  29971=>"001010111",
  29972=>"001011011",
  29973=>"001000010",
  29974=>"001010100",
  29975=>"001100111",
  29976=>"101001010",
  29977=>"101100111",
  29978=>"101011110",
  29979=>"000011101",
  29980=>"100100101",
  29981=>"110111010",
  29982=>"110000100",
  29983=>"001000110",
  29984=>"000100010",
  29985=>"000100110",
  29986=>"100101001",
  29987=>"111010111",
  29988=>"100000001",
  29989=>"101110000",
  29990=>"010010110",
  29991=>"101000000",
  29992=>"110000001",
  29993=>"101110001",
  29994=>"011011011",
  29995=>"000101010",
  29996=>"100111100",
  29997=>"000010100",
  29998=>"001000000",
  29999=>"010000111",
  30000=>"110000110",
  30001=>"000010000",
  30002=>"001111001",
  30003=>"101001111",
  30004=>"011011010",
  30005=>"110100101",
  30006=>"011101110",
  30007=>"000000111",
  30008=>"001111110",
  30009=>"110011010",
  30010=>"001110111",
  30011=>"110101110",
  30012=>"011010101",
  30013=>"011111100",
  30014=>"010110010",
  30015=>"000001011",
  30016=>"111110011",
  30017=>"100000101",
  30018=>"000111111",
  30019=>"100111111",
  30020=>"011101010",
  30021=>"000001100",
  30022=>"100010110",
  30023=>"101000101",
  30024=>"111010000",
  30025=>"100011000",
  30026=>"100010111",
  30027=>"110010011",
  30028=>"001011000",
  30029=>"100000011",
  30030=>"101100110",
  30031=>"011011101",
  30032=>"000001110",
  30033=>"100000010",
  30034=>"000101001",
  30035=>"111011100",
  30036=>"001101001",
  30037=>"111110111",
  30038=>"101111011",
  30039=>"100100100",
  30040=>"000001000",
  30041=>"000100111",
  30042=>"001010010",
  30043=>"100110101",
  30044=>"100000111",
  30045=>"101111010",
  30046=>"001100101",
  30047=>"011011000",
  30048=>"010100010",
  30049=>"000111101",
  30050=>"111100101",
  30051=>"011010011",
  30052=>"100001010",
  30053=>"100000000",
  30054=>"111101111",
  30055=>"011111100",
  30056=>"000100111",
  30057=>"110010110",
  30058=>"101001101",
  30059=>"111100110",
  30060=>"001101100",
  30061=>"001011010",
  30062=>"100000000",
  30063=>"001000000",
  30064=>"101101100",
  30065=>"110100000",
  30066=>"011011000",
  30067=>"100010110",
  30068=>"111001100",
  30069=>"100001111",
  30070=>"101110100",
  30071=>"100111110",
  30072=>"100110011",
  30073=>"110011001",
  30074=>"101111101",
  30075=>"110111101",
  30076=>"011110010",
  30077=>"100010110",
  30078=>"111001000",
  30079=>"011110010",
  30080=>"010000110",
  30081=>"011101110",
  30082=>"010011101",
  30083=>"100010111",
  30084=>"100010000",
  30085=>"111100100",
  30086=>"101110001",
  30087=>"111011111",
  30088=>"111001101",
  30089=>"001011011",
  30090=>"010010011",
  30091=>"001000101",
  30092=>"111101111",
  30093=>"011101100",
  30094=>"101100101",
  30095=>"100010000",
  30096=>"001011111",
  30097=>"001000110",
  30098=>"001111001",
  30099=>"011110100",
  30100=>"111110000",
  30101=>"100000010",
  30102=>"111010010",
  30103=>"111100110",
  30104=>"010110101",
  30105=>"000000011",
  30106=>"100111101",
  30107=>"000000000",
  30108=>"010111100",
  30109=>"101011101",
  30110=>"000100001",
  30111=>"111011111",
  30112=>"000101011",
  30113=>"001110001",
  30114=>"010000010",
  30115=>"111101011",
  30116=>"110011010",
  30117=>"001001110",
  30118=>"111111111",
  30119=>"010000110",
  30120=>"100010001",
  30121=>"100111111",
  30122=>"000011100",
  30123=>"100010001",
  30124=>"100010010",
  30125=>"000110000",
  30126=>"010011101",
  30127=>"101110111",
  30128=>"111001001",
  30129=>"001011011",
  30130=>"101110101",
  30131=>"001111001",
  30132=>"001011100",
  30133=>"100101100",
  30134=>"010110010",
  30135=>"100011111",
  30136=>"100101001",
  30137=>"111001011",
  30138=>"110011111",
  30139=>"010111000",
  30140=>"100101100",
  30141=>"010010111",
  30142=>"000001010",
  30143=>"100110111",
  30144=>"100101111",
  30145=>"000011110",
  30146=>"100010110",
  30147=>"101101110",
  30148=>"111011111",
  30149=>"001101110",
  30150=>"001000110",
  30151=>"110110010",
  30152=>"111110001",
  30153=>"100000101",
  30154=>"001011000",
  30155=>"000111000",
  30156=>"101111101",
  30157=>"000100000",
  30158=>"010001110",
  30159=>"010101101",
  30160=>"001001101",
  30161=>"010011101",
  30162=>"111100011",
  30163=>"101011000",
  30164=>"101100111",
  30165=>"100110010",
  30166=>"001010101",
  30167=>"000000110",
  30168=>"110101111",
  30169=>"100010010",
  30170=>"000010000",
  30171=>"000001010",
  30172=>"110010001",
  30173=>"101110111",
  30174=>"000110010",
  30175=>"101011000",
  30176=>"111001110",
  30177=>"110100111",
  30178=>"111111110",
  30179=>"011100000",
  30180=>"100011111",
  30181=>"101101010",
  30182=>"110000110",
  30183=>"011011101",
  30184=>"111110110",
  30185=>"010111011",
  30186=>"111010000",
  30187=>"001111010",
  30188=>"101111010",
  30189=>"010011111",
  30190=>"010100111",
  30191=>"110000001",
  30192=>"001101100",
  30193=>"100010100",
  30194=>"110011010",
  30195=>"110101001",
  30196=>"100010001",
  30197=>"000101101",
  30198=>"110100001",
  30199=>"110110010",
  30200=>"001011001",
  30201=>"000100010",
  30202=>"100111100",
  30203=>"000110100",
  30204=>"000011001",
  30205=>"101011001",
  30206=>"010011000",
  30207=>"111110001",
  30208=>"010101110",
  30209=>"100001011",
  30210=>"100011010",
  30211=>"000000101",
  30212=>"010000010",
  30213=>"101011001",
  30214=>"100111011",
  30215=>"010100101",
  30216=>"000001001",
  30217=>"101000001",
  30218=>"100111100",
  30219=>"100001111",
  30220=>"011110100",
  30221=>"100111010",
  30222=>"000001111",
  30223=>"000100111",
  30224=>"010011101",
  30225=>"000100010",
  30226=>"000001101",
  30227=>"101101010",
  30228=>"101010001",
  30229=>"100001010",
  30230=>"001101000",
  30231=>"001000101",
  30232=>"110100101",
  30233=>"110110010",
  30234=>"001100110",
  30235=>"011011001",
  30236=>"110010100",
  30237=>"011110001",
  30238=>"000001100",
  30239=>"010000111",
  30240=>"110010101",
  30241=>"001111100",
  30242=>"111001110",
  30243=>"101100100",
  30244=>"000101111",
  30245=>"011101101",
  30246=>"110011000",
  30247=>"100100011",
  30248=>"100011000",
  30249=>"100100001",
  30250=>"001010000",
  30251=>"010110111",
  30252=>"110010110",
  30253=>"110001011",
  30254=>"101101110",
  30255=>"010101001",
  30256=>"010011100",
  30257=>"111101111",
  30258=>"111010011",
  30259=>"010100111",
  30260=>"100101011",
  30261=>"000000100",
  30262=>"001001001",
  30263=>"110111110",
  30264=>"001110011",
  30265=>"111000101",
  30266=>"111001110",
  30267=>"101100001",
  30268=>"111001001",
  30269=>"000001110",
  30270=>"101110110",
  30271=>"010111110",
  30272=>"101010010",
  30273=>"011110000",
  30274=>"001101010",
  30275=>"000100011",
  30276=>"001011000",
  30277=>"000011110",
  30278=>"001010000",
  30279=>"100110000",
  30280=>"000001100",
  30281=>"101110100",
  30282=>"101010010",
  30283=>"100110110",
  30284=>"011100011",
  30285=>"100000000",
  30286=>"011100000",
  30287=>"110101111",
  30288=>"111100010",
  30289=>"011101111",
  30290=>"100000010",
  30291=>"011001110",
  30292=>"110000101",
  30293=>"011001101",
  30294=>"101010111",
  30295=>"011111111",
  30296=>"011000011",
  30297=>"101110111",
  30298=>"011110111",
  30299=>"111110101",
  30300=>"000101101",
  30301=>"110101001",
  30302=>"110011100",
  30303=>"100000010",
  30304=>"000000101",
  30305=>"111001000",
  30306=>"001100110",
  30307=>"000001110",
  30308=>"010100111",
  30309=>"110111111",
  30310=>"100000011",
  30311=>"111010111",
  30312=>"100011011",
  30313=>"110110111",
  30314=>"011010011",
  30315=>"000001000",
  30316=>"110110100",
  30317=>"100000011",
  30318=>"011111011",
  30319=>"100000110",
  30320=>"110001110",
  30321=>"111111100",
  30322=>"011100010",
  30323=>"110101011",
  30324=>"010111101",
  30325=>"010111110",
  30326=>"111000000",
  30327=>"100101000",
  30328=>"100010101",
  30329=>"011010111",
  30330=>"001011111",
  30331=>"011110001",
  30332=>"000011100",
  30333=>"000001111",
  30334=>"100011000",
  30335=>"000110011",
  30336=>"000100000",
  30337=>"101001111",
  30338=>"001100001",
  30339=>"110111111",
  30340=>"010110010",
  30341=>"000111100",
  30342=>"011000000",
  30343=>"001110001",
  30344=>"111001010",
  30345=>"111110111",
  30346=>"101001101",
  30347=>"110011001",
  30348=>"101011100",
  30349=>"110011110",
  30350=>"111000010",
  30351=>"000000101",
  30352=>"100010011",
  30353=>"111111110",
  30354=>"110100100",
  30355=>"001111000",
  30356=>"000000110",
  30357=>"000110100",
  30358=>"101001101",
  30359=>"001110010",
  30360=>"000110110",
  30361=>"101001100",
  30362=>"010000001",
  30363=>"001111101",
  30364=>"000101001",
  30365=>"011001010",
  30366=>"110100010",
  30367=>"011001111",
  30368=>"000100111",
  30369=>"100100111",
  30370=>"000110010",
  30371=>"001001001",
  30372=>"001011001",
  30373=>"111001110",
  30374=>"100110111",
  30375=>"000000110",
  30376=>"001100111",
  30377=>"000000101",
  30378=>"101101110",
  30379=>"000001001",
  30380=>"000101111",
  30381=>"000010111",
  30382=>"100011010",
  30383=>"001100000",
  30384=>"001010011",
  30385=>"110001110",
  30386=>"001001100",
  30387=>"011100001",
  30388=>"111101010",
  30389=>"001110000",
  30390=>"100000010",
  30391=>"111001000",
  30392=>"111010101",
  30393=>"011101110",
  30394=>"000011001",
  30395=>"000001001",
  30396=>"001100111",
  30397=>"101111011",
  30398=>"101110100",
  30399=>"001001001",
  30400=>"011101100",
  30401=>"000100111",
  30402=>"101011000",
  30403=>"000001000",
  30404=>"101011011",
  30405=>"000001000",
  30406=>"101011000",
  30407=>"001000001",
  30408=>"110101011",
  30409=>"110010011",
  30410=>"000000010",
  30411=>"110010101",
  30412=>"000000001",
  30413=>"111111101",
  30414=>"101010101",
  30415=>"011100011",
  30416=>"011011100",
  30417=>"100111001",
  30418=>"010010000",
  30419=>"011111010",
  30420=>"101001101",
  30421=>"101100110",
  30422=>"111000010",
  30423=>"100000101",
  30424=>"101101100",
  30425=>"000011101",
  30426=>"001011010",
  30427=>"111011000",
  30428=>"011110100",
  30429=>"110110000",
  30430=>"000001111",
  30431=>"011011101",
  30432=>"010000110",
  30433=>"001000010",
  30434=>"001111111",
  30435=>"010110001",
  30436=>"010100101",
  30437=>"000100101",
  30438=>"111101110",
  30439=>"101010110",
  30440=>"001110111",
  30441=>"010011100",
  30442=>"011100011",
  30443=>"100000000",
  30444=>"000100111",
  30445=>"101101110",
  30446=>"101110101",
  30447=>"001110100",
  30448=>"100001010",
  30449=>"111100111",
  30450=>"010101110",
  30451=>"110011111",
  30452=>"101100101",
  30453=>"111010110",
  30454=>"001000100",
  30455=>"110000100",
  30456=>"011101011",
  30457=>"100110101",
  30458=>"001111110",
  30459=>"110101011",
  30460=>"100011110",
  30461=>"010100010",
  30462=>"000000110",
  30463=>"010011000",
  30464=>"110011010",
  30465=>"001000010",
  30466=>"111101100",
  30467=>"100010010",
  30468=>"001001100",
  30469=>"110000010",
  30470=>"100011100",
  30471=>"001001010",
  30472=>"000000100",
  30473=>"111110010",
  30474=>"110001101",
  30475=>"111111011",
  30476=>"011000000",
  30477=>"110111111",
  30478=>"000011110",
  30479=>"010101111",
  30480=>"000011000",
  30481=>"011000001",
  30482=>"011100100",
  30483=>"111011000",
  30484=>"001001011",
  30485=>"010001010",
  30486=>"101000010",
  30487=>"100101110",
  30488=>"001101111",
  30489=>"101000101",
  30490=>"111001111",
  30491=>"000101100",
  30492=>"101000000",
  30493=>"010100001",
  30494=>"100010111",
  30495=>"011101111",
  30496=>"110100010",
  30497=>"000010001",
  30498=>"101010001",
  30499=>"110111111",
  30500=>"111001111",
  30501=>"001110001",
  30502=>"000000011",
  30503=>"011010011",
  30504=>"110110000",
  30505=>"010011010",
  30506=>"111101001",
  30507=>"101000100",
  30508=>"011111010",
  30509=>"101101111",
  30510=>"110001100",
  30511=>"101111110",
  30512=>"010010010",
  30513=>"000100000",
  30514=>"100001111",
  30515=>"001001100",
  30516=>"000101011",
  30517=>"010111100",
  30518=>"111101001",
  30519=>"100001111",
  30520=>"011011001",
  30521=>"011011101",
  30522=>"111111000",
  30523=>"111110011",
  30524=>"000100011",
  30525=>"010000101",
  30526=>"110011101",
  30527=>"011110101",
  30528=>"110100001",
  30529=>"000011010",
  30530=>"100001000",
  30531=>"001101001",
  30532=>"000000001",
  30533=>"101000011",
  30534=>"000111010",
  30535=>"110011001",
  30536=>"110111010",
  30537=>"010011100",
  30538=>"001101000",
  30539=>"010100111",
  30540=>"101110100",
  30541=>"111110101",
  30542=>"001001100",
  30543=>"011001000",
  30544=>"001110001",
  30545=>"111011011",
  30546=>"111111110",
  30547=>"000001100",
  30548=>"001100100",
  30549=>"100001011",
  30550=>"101100001",
  30551=>"001100000",
  30552=>"100111101",
  30553=>"101010110",
  30554=>"101101010",
  30555=>"000000100",
  30556=>"011001011",
  30557=>"010011001",
  30558=>"011010101",
  30559=>"011101000",
  30560=>"010111011",
  30561=>"100101000",
  30562=>"100000001",
  30563=>"110011001",
  30564=>"011111110",
  30565=>"100011000",
  30566=>"111000111",
  30567=>"110010011",
  30568=>"111001000",
  30569=>"111110001",
  30570=>"011100010",
  30571=>"010010111",
  30572=>"001101011",
  30573=>"101000001",
  30574=>"111011010",
  30575=>"010110110",
  30576=>"010110101",
  30577=>"000101100",
  30578=>"000110100",
  30579=>"111001000",
  30580=>"101000100",
  30581=>"010101010",
  30582=>"001000011",
  30583=>"100010100",
  30584=>"011000110",
  30585=>"110111100",
  30586=>"011100011",
  30587=>"000111011",
  30588=>"010101000",
  30589=>"101100100",
  30590=>"111000011",
  30591=>"111011111",
  30592=>"010110100",
  30593=>"101010001",
  30594=>"111001001",
  30595=>"011001100",
  30596=>"110010010",
  30597=>"101010110",
  30598=>"000011110",
  30599=>"101111001",
  30600=>"100111010",
  30601=>"000010011",
  30602=>"111100010",
  30603=>"110000000",
  30604=>"101100101",
  30605=>"101100111",
  30606=>"100100101",
  30607=>"010011001",
  30608=>"101001111",
  30609=>"111000100",
  30610=>"110111100",
  30611=>"000111001",
  30612=>"111110000",
  30613=>"010010100",
  30614=>"010010111",
  30615=>"011110100",
  30616=>"000011101",
  30617=>"111110000",
  30618=>"100000001",
  30619=>"110101000",
  30620=>"001100010",
  30621=>"100011001",
  30622=>"000011000",
  30623=>"111011111",
  30624=>"111111111",
  30625=>"101111010",
  30626=>"110011110",
  30627=>"101001000",
  30628=>"011110001",
  30629=>"100000011",
  30630=>"101011000",
  30631=>"010111010",
  30632=>"000001110",
  30633=>"111110111",
  30634=>"011010111",
  30635=>"000100011",
  30636=>"000011000",
  30637=>"110001110",
  30638=>"100110001",
  30639=>"110110100",
  30640=>"101010101",
  30641=>"000110111",
  30642=>"010011001",
  30643=>"100111001",
  30644=>"111011001",
  30645=>"111101101",
  30646=>"111101101",
  30647=>"101000000",
  30648=>"000001110",
  30649=>"000100010",
  30650=>"010101111",
  30651=>"100111011",
  30652=>"011000110",
  30653=>"100101000",
  30654=>"010101010",
  30655=>"101110000",
  30656=>"010101101",
  30657=>"101000101",
  30658=>"111010010",
  30659=>"110001001",
  30660=>"111110101",
  30661=>"011011100",
  30662=>"101111101",
  30663=>"001001001",
  30664=>"011001001",
  30665=>"111110001",
  30666=>"100011000",
  30667=>"010100000",
  30668=>"101101010",
  30669=>"001001000",
  30670=>"111110000",
  30671=>"010011100",
  30672=>"100000100",
  30673=>"111001001",
  30674=>"001001000",
  30675=>"001011010",
  30676=>"000000011",
  30677=>"110011001",
  30678=>"111010111",
  30679=>"111100101",
  30680=>"010101011",
  30681=>"100110101",
  30682=>"101111110",
  30683=>"101000001",
  30684=>"000101001",
  30685=>"001111011",
  30686=>"000011111",
  30687=>"000101000",
  30688=>"000000000",
  30689=>"001101001",
  30690=>"000001101",
  30691=>"010000101",
  30692=>"000111101",
  30693=>"011001010",
  30694=>"000001010",
  30695=>"110001110",
  30696=>"001010110",
  30697=>"100100011",
  30698=>"111100010",
  30699=>"000010100",
  30700=>"101010011",
  30701=>"000010010",
  30702=>"101000011",
  30703=>"111111101",
  30704=>"100101001",
  30705=>"010000000",
  30706=>"100010101",
  30707=>"001000101",
  30708=>"001000000",
  30709=>"110001011",
  30710=>"010101100",
  30711=>"010000100",
  30712=>"111000101",
  30713=>"111010110",
  30714=>"110100111",
  30715=>"001111001",
  30716=>"000011001",
  30717=>"101100011",
  30718=>"110110110",
  30719=>"000100010",
  30720=>"000101001",
  30721=>"001010010",
  30722=>"001101101",
  30723=>"001111000",
  30724=>"011000101",
  30725=>"111001010",
  30726=>"110101010",
  30727=>"101010110",
  30728=>"111100000",
  30729=>"000011101",
  30730=>"001100010",
  30731=>"010001001",
  30732=>"001111111",
  30733=>"101110111",
  30734=>"000000010",
  30735=>"010000111",
  30736=>"110001011",
  30737=>"000000101",
  30738=>"110010100",
  30739=>"111000101",
  30740=>"000111010",
  30741=>"110000111",
  30742=>"101101110",
  30743=>"011111111",
  30744=>"000011101",
  30745=>"111100101",
  30746=>"101101101",
  30747=>"111000111",
  30748=>"001101100",
  30749=>"110110111",
  30750=>"111100101",
  30751=>"110101110",
  30752=>"110010111",
  30753=>"011110011",
  30754=>"101000110",
  30755=>"011001110",
  30756=>"000001010",
  30757=>"001100100",
  30758=>"000001101",
  30759=>"100111101",
  30760=>"101000010",
  30761=>"001111110",
  30762=>"111011011",
  30763=>"111100001",
  30764=>"000001110",
  30765=>"101001110",
  30766=>"010000101",
  30767=>"110110010",
  30768=>"111100100",
  30769=>"100011000",
  30770=>"111110010",
  30771=>"011000001",
  30772=>"110101000",
  30773=>"000000110",
  30774=>"001100111",
  30775=>"110101001",
  30776=>"101100011",
  30777=>"111111001",
  30778=>"111111111",
  30779=>"110000001",
  30780=>"111000110",
  30781=>"001010100",
  30782=>"101011011",
  30783=>"111100100",
  30784=>"000011011",
  30785=>"010100110",
  30786=>"101011000",
  30787=>"101000101",
  30788=>"100010011",
  30789=>"100100100",
  30790=>"111010111",
  30791=>"111111100",
  30792=>"000101100",
  30793=>"000101100",
  30794=>"100001010",
  30795=>"100010100",
  30796=>"001001001",
  30797=>"100010000",
  30798=>"101000110",
  30799=>"100011111",
  30800=>"110110110",
  30801=>"110101000",
  30802=>"110001110",
  30803=>"000000011",
  30804=>"001001110",
  30805=>"111110011",
  30806=>"100111011",
  30807=>"001001111",
  30808=>"101100100",
  30809=>"001111010",
  30810=>"110101001",
  30811=>"000101100",
  30812=>"110111111",
  30813=>"110101000",
  30814=>"110110101",
  30815=>"111011011",
  30816=>"110011010",
  30817=>"000010101",
  30818=>"011101101",
  30819=>"000001011",
  30820=>"001111001",
  30821=>"001100101",
  30822=>"101011100",
  30823=>"000010100",
  30824=>"111001011",
  30825=>"111001000",
  30826=>"011100000",
  30827=>"100100000",
  30828=>"110101111",
  30829=>"110001100",
  30830=>"001011110",
  30831=>"101010000",
  30832=>"000011010",
  30833=>"011010100",
  30834=>"111111111",
  30835=>"101001001",
  30836=>"111110110",
  30837=>"110010011",
  30838=>"011111110",
  30839=>"101000011",
  30840=>"111011110",
  30841=>"110111010",
  30842=>"000111001",
  30843=>"001001100",
  30844=>"011111100",
  30845=>"010101111",
  30846=>"000010010",
  30847=>"110101111",
  30848=>"001001000",
  30849=>"101010001",
  30850=>"001010010",
  30851=>"001101100",
  30852=>"111111101",
  30853=>"100001101",
  30854=>"000011100",
  30855=>"101010101",
  30856=>"011000110",
  30857=>"000111000",
  30858=>"111001100",
  30859=>"110101110",
  30860=>"001110110",
  30861=>"111010111",
  30862=>"101111001",
  30863=>"000011100",
  30864=>"000111011",
  30865=>"110110101",
  30866=>"010111110",
  30867=>"011010101",
  30868=>"101011111",
  30869=>"110101101",
  30870=>"000111000",
  30871=>"001000011",
  30872=>"100100010",
  30873=>"110010111",
  30874=>"100011111",
  30875=>"000111011",
  30876=>"011101111",
  30877=>"100010111",
  30878=>"111001110",
  30879=>"000011000",
  30880=>"001010100",
  30881=>"100101101",
  30882=>"001111011",
  30883=>"111100100",
  30884=>"110111101",
  30885=>"110100101",
  30886=>"101001110",
  30887=>"000000100",
  30888=>"111001101",
  30889=>"000011111",
  30890=>"000001000",
  30891=>"100010001",
  30892=>"100110011",
  30893=>"011100001",
  30894=>"101111001",
  30895=>"000000000",
  30896=>"101111010",
  30897=>"000001100",
  30898=>"100101111",
  30899=>"001100111",
  30900=>"000000001",
  30901=>"111110101",
  30902=>"101101101",
  30903=>"010001110",
  30904=>"111100100",
  30905=>"111001110",
  30906=>"000010100",
  30907=>"011010100",
  30908=>"110010110",
  30909=>"110111110",
  30910=>"100010000",
  30911=>"110010000",
  30912=>"001111101",
  30913=>"000011000",
  30914=>"111111101",
  30915=>"111110010",
  30916=>"100010100",
  30917=>"000010101",
  30918=>"100111111",
  30919=>"101100000",
  30920=>"010101001",
  30921=>"000111010",
  30922=>"110011111",
  30923=>"011011111",
  30924=>"100010110",
  30925=>"111101100",
  30926=>"101110100",
  30927=>"011010100",
  30928=>"000111000",
  30929=>"101110111",
  30930=>"101011011",
  30931=>"110011000",
  30932=>"001100001",
  30933=>"010011111",
  30934=>"101110101",
  30935=>"011110010",
  30936=>"110100101",
  30937=>"111001000",
  30938=>"001100100",
  30939=>"101010101",
  30940=>"111011100",
  30941=>"100000100",
  30942=>"000000100",
  30943=>"011100000",
  30944=>"111101000",
  30945=>"000001010",
  30946=>"101010111",
  30947=>"010010111",
  30948=>"100101000",
  30949=>"111000010",
  30950=>"100101010",
  30951=>"110000011",
  30952=>"010111111",
  30953=>"001010110",
  30954=>"010111110",
  30955=>"000011001",
  30956=>"011111101",
  30957=>"100000001",
  30958=>"101010111",
  30959=>"110100111",
  30960=>"001101001",
  30961=>"011000011",
  30962=>"000000000",
  30963=>"111011010",
  30964=>"111000011",
  30965=>"010011010",
  30966=>"100110111",
  30967=>"111111101",
  30968=>"100010011",
  30969=>"011000101",
  30970=>"110110000",
  30971=>"001010111",
  30972=>"101111011",
  30973=>"111011101",
  30974=>"010100100",
  30975=>"000111111",
  30976=>"001001010",
  30977=>"101001111",
  30978=>"011010011",
  30979=>"111111110",
  30980=>"001010001",
  30981=>"101000010",
  30982=>"111001111",
  30983=>"110110000",
  30984=>"101001001",
  30985=>"000101011",
  30986=>"001010110",
  30987=>"001110111",
  30988=>"011110111",
  30989=>"101101111",
  30990=>"110000010",
  30991=>"001100000",
  30992=>"101011101",
  30993=>"110010110",
  30994=>"110100001",
  30995=>"111100000",
  30996=>"101010100",
  30997=>"010000000",
  30998=>"000001001",
  30999=>"000011100",
  31000=>"001000111",
  31001=>"011101010",
  31002=>"110100010",
  31003=>"111011100",
  31004=>"111101111",
  31005=>"001011111",
  31006=>"100010100",
  31007=>"111110011",
  31008=>"101111001",
  31009=>"111101010",
  31010=>"001110000",
  31011=>"111000101",
  31012=>"011001100",
  31013=>"111110110",
  31014=>"110010011",
  31015=>"010001000",
  31016=>"100101101",
  31017=>"010010111",
  31018=>"111111111",
  31019=>"111101100",
  31020=>"111000000",
  31021=>"100001000",
  31022=>"101010001",
  31023=>"001001001",
  31024=>"010100111",
  31025=>"000110000",
  31026=>"011111110",
  31027=>"100110111",
  31028=>"001011011",
  31029=>"000000101",
  31030=>"111101000",
  31031=>"010101101",
  31032=>"000011101",
  31033=>"100101100",
  31034=>"100000000",
  31035=>"001110000",
  31036=>"010011010",
  31037=>"110001111",
  31038=>"100000000",
  31039=>"110110111",
  31040=>"000000101",
  31041=>"010110101",
  31042=>"010001001",
  31043=>"101011001",
  31044=>"010100000",
  31045=>"100101100",
  31046=>"100011000",
  31047=>"100100101",
  31048=>"010010101",
  31049=>"110110111",
  31050=>"010110011",
  31051=>"100000011",
  31052=>"100011001",
  31053=>"010000010",
  31054=>"111110001",
  31055=>"011001010",
  31056=>"011100000",
  31057=>"010110100",
  31058=>"100110011",
  31059=>"011111000",
  31060=>"111010001",
  31061=>"111101010",
  31062=>"110011000",
  31063=>"011000101",
  31064=>"100011010",
  31065=>"010001011",
  31066=>"100001000",
  31067=>"101001111",
  31068=>"110100011",
  31069=>"110111011",
  31070=>"010000011",
  31071=>"100000100",
  31072=>"101100111",
  31073=>"101100011",
  31074=>"101001110",
  31075=>"000010001",
  31076=>"100111001",
  31077=>"110001011",
  31078=>"011010011",
  31079=>"111011101",
  31080=>"000111111",
  31081=>"111010101",
  31082=>"110110111",
  31083=>"111001111",
  31084=>"111000000",
  31085=>"000001101",
  31086=>"101001011",
  31087=>"001010100",
  31088=>"001110101",
  31089=>"010100101",
  31090=>"110011101",
  31091=>"000001100",
  31092=>"100111111",
  31093=>"001110000",
  31094=>"100101100",
  31095=>"111111101",
  31096=>"110010010",
  31097=>"010000101",
  31098=>"101110000",
  31099=>"011101111",
  31100=>"010011110",
  31101=>"111100011",
  31102=>"001110001",
  31103=>"111111001",
  31104=>"111011000",
  31105=>"010001110",
  31106=>"111000100",
  31107=>"000000111",
  31108=>"010111010",
  31109=>"001101110",
  31110=>"000011110",
  31111=>"101010010",
  31112=>"011111001",
  31113=>"000001110",
  31114=>"101011100",
  31115=>"111111000",
  31116=>"111010001",
  31117=>"001001001",
  31118=>"101001011",
  31119=>"001010100",
  31120=>"111001111",
  31121=>"100000001",
  31122=>"101001111",
  31123=>"000010101",
  31124=>"101111101",
  31125=>"001010101",
  31126=>"111010101",
  31127=>"100100111",
  31128=>"111000000",
  31129=>"000111000",
  31130=>"111110000",
  31131=>"101011001",
  31132=>"010010001",
  31133=>"010000011",
  31134=>"010100111",
  31135=>"111001110",
  31136=>"111111100",
  31137=>"000111011",
  31138=>"110010011",
  31139=>"101110000",
  31140=>"100000001",
  31141=>"100010100",
  31142=>"001110111",
  31143=>"000100010",
  31144=>"010111000",
  31145=>"011011011",
  31146=>"001000111",
  31147=>"010000111",
  31148=>"011110000",
  31149=>"110101111",
  31150=>"000100011",
  31151=>"000011101",
  31152=>"001101011",
  31153=>"110111110",
  31154=>"010110011",
  31155=>"111000011",
  31156=>"001010101",
  31157=>"110111111",
  31158=>"001110111",
  31159=>"010110000",
  31160=>"010001101",
  31161=>"111001001",
  31162=>"110011101",
  31163=>"110101110",
  31164=>"100010000",
  31165=>"100010011",
  31166=>"100000000",
  31167=>"011011011",
  31168=>"011111001",
  31169=>"010001110",
  31170=>"100100101",
  31171=>"111000000",
  31172=>"011111111",
  31173=>"000010011",
  31174=>"110111010",
  31175=>"110000001",
  31176=>"100011100",
  31177=>"000110000",
  31178=>"110110010",
  31179=>"101011101",
  31180=>"001101011",
  31181=>"000101001",
  31182=>"000110000",
  31183=>"011101101",
  31184=>"110011010",
  31185=>"011100100",
  31186=>"100000100",
  31187=>"111001101",
  31188=>"110110100",
  31189=>"111010011",
  31190=>"011111101",
  31191=>"110001100",
  31192=>"111010110",
  31193=>"100100001",
  31194=>"111100111",
  31195=>"101001100",
  31196=>"000101110",
  31197=>"000100101",
  31198=>"000111011",
  31199=>"010011101",
  31200=>"101100100",
  31201=>"100000110",
  31202=>"101001010",
  31203=>"010001010",
  31204=>"011111111",
  31205=>"010010000",
  31206=>"110011001",
  31207=>"101100001",
  31208=>"100000100",
  31209=>"110010101",
  31210=>"000000110",
  31211=>"001110010",
  31212=>"010011001",
  31213=>"110100100",
  31214=>"100101101",
  31215=>"101101011",
  31216=>"000010000",
  31217=>"111001000",
  31218=>"000111110",
  31219=>"101000010",
  31220=>"011110011",
  31221=>"000000110",
  31222=>"011011100",
  31223=>"011011111",
  31224=>"110110001",
  31225=>"011010001",
  31226=>"000001000",
  31227=>"011100000",
  31228=>"000010100",
  31229=>"010110110",
  31230=>"110111000",
  31231=>"000101101",
  31232=>"100101100",
  31233=>"000010101",
  31234=>"001110100",
  31235=>"111000000",
  31236=>"111000001",
  31237=>"111011001",
  31238=>"111101101",
  31239=>"010110110",
  31240=>"100100111",
  31241=>"000110111",
  31242=>"000011011",
  31243=>"001001001",
  31244=>"010000111",
  31245=>"111111011",
  31246=>"010111001",
  31247=>"110100001",
  31248=>"010011000",
  31249=>"100101001",
  31250=>"101100100",
  31251=>"100010001",
  31252=>"001101111",
  31253=>"111100100",
  31254=>"111010101",
  31255=>"111011011",
  31256=>"010010101",
  31257=>"111011010",
  31258=>"111000000",
  31259=>"010001101",
  31260=>"001111101",
  31261=>"111010100",
  31262=>"011010000",
  31263=>"011111111",
  31264=>"010001001",
  31265=>"101001011",
  31266=>"001110100",
  31267=>"110111100",
  31268=>"101001000",
  31269=>"000110011",
  31270=>"110000111",
  31271=>"010000110",
  31272=>"101001010",
  31273=>"100111111",
  31274=>"101010011",
  31275=>"111011110",
  31276=>"110110001",
  31277=>"111000001",
  31278=>"101101100",
  31279=>"011001000",
  31280=>"100100011",
  31281=>"101000001",
  31282=>"101111100",
  31283=>"100100000",
  31284=>"000010011",
  31285=>"101010111",
  31286=>"100001101",
  31287=>"101111000",
  31288=>"000010110",
  31289=>"011100110",
  31290=>"101110010",
  31291=>"010001110",
  31292=>"010010011",
  31293=>"110101011",
  31294=>"101100011",
  31295=>"101000101",
  31296=>"100011111",
  31297=>"011101000",
  31298=>"001001010",
  31299=>"101010000",
  31300=>"010011100",
  31301=>"100110001",
  31302=>"000111011",
  31303=>"010111110",
  31304=>"011001101",
  31305=>"011110111",
  31306=>"000111101",
  31307=>"101010100",
  31308=>"111000101",
  31309=>"101000111",
  31310=>"010000101",
  31311=>"000111110",
  31312=>"001011101",
  31313=>"011100100",
  31314=>"001111101",
  31315=>"100000110",
  31316=>"010010001",
  31317=>"000000000",
  31318=>"000100001",
  31319=>"000110101",
  31320=>"111111111",
  31321=>"101010000",
  31322=>"010011010",
  31323=>"101001001",
  31324=>"011110101",
  31325=>"110110110",
  31326=>"011101011",
  31327=>"000000000",
  31328=>"010000100",
  31329=>"011000111",
  31330=>"111101011",
  31331=>"111001100",
  31332=>"100100100",
  31333=>"001100000",
  31334=>"011101101",
  31335=>"010011101",
  31336=>"000101000",
  31337=>"000011001",
  31338=>"000000111",
  31339=>"001000000",
  31340=>"011011001",
  31341=>"010000100",
  31342=>"111010001",
  31343=>"000111011",
  31344=>"000110100",
  31345=>"111100000",
  31346=>"111101111",
  31347=>"111100011",
  31348=>"001101010",
  31349=>"100110001",
  31350=>"000100110",
  31351=>"010101100",
  31352=>"000010110",
  31353=>"000101000",
  31354=>"011111110",
  31355=>"100101101",
  31356=>"010001111",
  31357=>"110100111",
  31358=>"111100000",
  31359=>"111011001",
  31360=>"101100000",
  31361=>"111110100",
  31362=>"100000100",
  31363=>"100000110",
  31364=>"000110001",
  31365=>"010110011",
  31366=>"000101000",
  31367=>"001110001",
  31368=>"010010011",
  31369=>"111000110",
  31370=>"111100100",
  31371=>"101100000",
  31372=>"011000110",
  31373=>"010101000",
  31374=>"101100010",
  31375=>"000100001",
  31376=>"100010000",
  31377=>"011100000",
  31378=>"000000111",
  31379=>"000101000",
  31380=>"111000011",
  31381=>"000101111",
  31382=>"011110000",
  31383=>"111000101",
  31384=>"010111101",
  31385=>"000000000",
  31386=>"001111010",
  31387=>"111010101",
  31388=>"000110010",
  31389=>"100101110",
  31390=>"000110001",
  31391=>"010011010",
  31392=>"000110010",
  31393=>"110000110",
  31394=>"101110110",
  31395=>"100100000",
  31396=>"100001101",
  31397=>"011010100",
  31398=>"001111110",
  31399=>"001111000",
  31400=>"000100010",
  31401=>"111101111",
  31402=>"010110000",
  31403=>"010110111",
  31404=>"111011011",
  31405=>"001110110",
  31406=>"011000100",
  31407=>"111111011",
  31408=>"101100010",
  31409=>"111111000",
  31410=>"011111000",
  31411=>"110111111",
  31412=>"101111101",
  31413=>"001010001",
  31414=>"000001110",
  31415=>"000000001",
  31416=>"100000110",
  31417=>"000000110",
  31418=>"001110011",
  31419=>"010000000",
  31420=>"110010010",
  31421=>"000110011",
  31422=>"100110101",
  31423=>"010101111",
  31424=>"001100011",
  31425=>"001001101",
  31426=>"001100100",
  31427=>"110000101",
  31428=>"101100111",
  31429=>"001000100",
  31430=>"100000110",
  31431=>"101101100",
  31432=>"110101001",
  31433=>"010111000",
  31434=>"111110000",
  31435=>"110100010",
  31436=>"101001100",
  31437=>"111010101",
  31438=>"001111111",
  31439=>"011010001",
  31440=>"100001000",
  31441=>"000001111",
  31442=>"010010000",
  31443=>"001011010",
  31444=>"010001101",
  31445=>"000111000",
  31446=>"101011001",
  31447=>"001000010",
  31448=>"110100000",
  31449=>"100000110",
  31450=>"110111000",
  31451=>"100101001",
  31452=>"101010010",
  31453=>"000101011",
  31454=>"001010111",
  31455=>"011001010",
  31456=>"111110000",
  31457=>"110100101",
  31458=>"000111110",
  31459=>"001001001",
  31460=>"100000010",
  31461=>"101100001",
  31462=>"011101011",
  31463=>"110110110",
  31464=>"100111110",
  31465=>"110111000",
  31466=>"011011011",
  31467=>"010000010",
  31468=>"001101111",
  31469=>"100001101",
  31470=>"101011011",
  31471=>"100111100",
  31472=>"100000001",
  31473=>"101010001",
  31474=>"100010111",
  31475=>"001110110",
  31476=>"001111101",
  31477=>"100111001",
  31478=>"000111110",
  31479=>"100001101",
  31480=>"111111100",
  31481=>"001111111",
  31482=>"001001100",
  31483=>"001000111",
  31484=>"000110100",
  31485=>"010001111",
  31486=>"100011001",
  31487=>"111100111",
  31488=>"011001100",
  31489=>"101010000",
  31490=>"011010110",
  31491=>"000101100",
  31492=>"101111111",
  31493=>"101000110",
  31494=>"011011101",
  31495=>"101111010",
  31496=>"001110101",
  31497=>"001001100",
  31498=>"101010111",
  31499=>"100110101",
  31500=>"000001111",
  31501=>"010001011",
  31502=>"010101010",
  31503=>"110100111",
  31504=>"000001011",
  31505=>"010100000",
  31506=>"101111010",
  31507=>"111001000",
  31508=>"010000010",
  31509=>"100101110",
  31510=>"000011010",
  31511=>"111010010",
  31512=>"101001001",
  31513=>"001111100",
  31514=>"100101011",
  31515=>"100110010",
  31516=>"101000100",
  31517=>"111011000",
  31518=>"011100110",
  31519=>"100000111",
  31520=>"010000101",
  31521=>"010110101",
  31522=>"111111110",
  31523=>"010010000",
  31524=>"110111000",
  31525=>"011110000",
  31526=>"010011000",
  31527=>"011000000",
  31528=>"111100011",
  31529=>"100011001",
  31530=>"011101011",
  31531=>"101001101",
  31532=>"011001110",
  31533=>"111010000",
  31534=>"000010001",
  31535=>"001110110",
  31536=>"110111101",
  31537=>"111101101",
  31538=>"001111100",
  31539=>"100010111",
  31540=>"111101011",
  31541=>"110011011",
  31542=>"001010101",
  31543=>"111000111",
  31544=>"001001011",
  31545=>"111011000",
  31546=>"110101010",
  31547=>"100000000",
  31548=>"001001111",
  31549=>"101111000",
  31550=>"111110101",
  31551=>"111110000",
  31552=>"001110010",
  31553=>"111000110",
  31554=>"110001001",
  31555=>"111101110",
  31556=>"100000100",
  31557=>"001101100",
  31558=>"111000110",
  31559=>"100001011",
  31560=>"010000010",
  31561=>"011100010",
  31562=>"111011110",
  31563=>"011001011",
  31564=>"101110101",
  31565=>"011100011",
  31566=>"010001000",
  31567=>"110101000",
  31568=>"110000010",
  31569=>"100000010",
  31570=>"011110000",
  31571=>"100110010",
  31572=>"010000101",
  31573=>"111010000",
  31574=>"100001001",
  31575=>"101110011",
  31576=>"001010100",
  31577=>"010000100",
  31578=>"011000001",
  31579=>"100000000",
  31580=>"111011111",
  31581=>"000010101",
  31582=>"110101000",
  31583=>"111110001",
  31584=>"111001101",
  31585=>"000101111",
  31586=>"010000010",
  31587=>"100001010",
  31588=>"010100010",
  31589=>"100100110",
  31590=>"110011101",
  31591=>"101100000",
  31592=>"010111000",
  31593=>"010111100",
  31594=>"011100001",
  31595=>"100111011",
  31596=>"000010000",
  31597=>"111000111",
  31598=>"000100110",
  31599=>"010010111",
  31600=>"000000100",
  31601=>"101001100",
  31602=>"011010100",
  31603=>"100101111",
  31604=>"000011010",
  31605=>"110010001",
  31606=>"110000001",
  31607=>"001001010",
  31608=>"010010111",
  31609=>"000001001",
  31610=>"100110000",
  31611=>"101000111",
  31612=>"100101111",
  31613=>"110000110",
  31614=>"100111110",
  31615=>"101100011",
  31616=>"010101110",
  31617=>"100110110",
  31618=>"011101011",
  31619=>"101000001",
  31620=>"001111111",
  31621=>"011111000",
  31622=>"011000100",
  31623=>"000001000",
  31624=>"111111000",
  31625=>"111010010",
  31626=>"111101010",
  31627=>"010110100",
  31628=>"010010000",
  31629=>"000110000",
  31630=>"100010111",
  31631=>"110110101",
  31632=>"101110011",
  31633=>"000000110",
  31634=>"101100001",
  31635=>"010011100",
  31636=>"110111100",
  31637=>"001110010",
  31638=>"101000001",
  31639=>"001001011",
  31640=>"011011001",
  31641=>"011101010",
  31642=>"101001100",
  31643=>"101001111",
  31644=>"111101011",
  31645=>"010011001",
  31646=>"100100101",
  31647=>"000010101",
  31648=>"000000011",
  31649=>"011111111",
  31650=>"010001100",
  31651=>"010100101",
  31652=>"111110110",
  31653=>"001010111",
  31654=>"000100001",
  31655=>"001001000",
  31656=>"101111101",
  31657=>"000000001",
  31658=>"000011000",
  31659=>"110000000",
  31660=>"000000110",
  31661=>"110111110",
  31662=>"111111110",
  31663=>"000001101",
  31664=>"011110101",
  31665=>"001000000",
  31666=>"011000100",
  31667=>"001001100",
  31668=>"001011101",
  31669=>"011111111",
  31670=>"010011001",
  31671=>"010101000",
  31672=>"001100000",
  31673=>"010011001",
  31674=>"010101011",
  31675=>"000011000",
  31676=>"101110100",
  31677=>"110010110",
  31678=>"110000110",
  31679=>"101111100",
  31680=>"000110000",
  31681=>"100111010",
  31682=>"011100011",
  31683=>"000010110",
  31684=>"111111100",
  31685=>"101111011",
  31686=>"111001000",
  31687=>"101101010",
  31688=>"110100101",
  31689=>"011000000",
  31690=>"001101110",
  31691=>"100111111",
  31692=>"000010110",
  31693=>"000111100",
  31694=>"010100100",
  31695=>"111111010",
  31696=>"011000110",
  31697=>"101110100",
  31698=>"000010011",
  31699=>"000000010",
  31700=>"010101000",
  31701=>"100000101",
  31702=>"111001100",
  31703=>"111001000",
  31704=>"010100001",
  31705=>"000001110",
  31706=>"111100110",
  31707=>"101100111",
  31708=>"000100010",
  31709=>"010100001",
  31710=>"110000111",
  31711=>"111011010",
  31712=>"111011100",
  31713=>"110100000",
  31714=>"100011001",
  31715=>"101011111",
  31716=>"010111100",
  31717=>"101011001",
  31718=>"111000001",
  31719=>"001010100",
  31720=>"101101001",
  31721=>"100111001",
  31722=>"000000000",
  31723=>"110110001",
  31724=>"000011000",
  31725=>"100111100",
  31726=>"000100101",
  31727=>"000110010",
  31728=>"100111001",
  31729=>"100000011",
  31730=>"000010100",
  31731=>"000110010",
  31732=>"011111110",
  31733=>"000011100",
  31734=>"000000000",
  31735=>"001101100",
  31736=>"101101100",
  31737=>"001001010",
  31738=>"010001011",
  31739=>"111101100",
  31740=>"111000111",
  31741=>"111101001",
  31742=>"100100011",
  31743=>"001010010",
  31744=>"111101001",
  31745=>"110101111",
  31746=>"100001111",
  31747=>"001100111",
  31748=>"001000011",
  31749=>"001101011",
  31750=>"001011101",
  31751=>"001100110",
  31752=>"000101001",
  31753=>"000110000",
  31754=>"001001000",
  31755=>"001001010",
  31756=>"000111111",
  31757=>"101011010",
  31758=>"010001001",
  31759=>"011110110",
  31760=>"011100001",
  31761=>"000110010",
  31762=>"100010000",
  31763=>"011010000",
  31764=>"011100011",
  31765=>"011100111",
  31766=>"001011000",
  31767=>"001111110",
  31768=>"011001110",
  31769=>"010010001",
  31770=>"101000100",
  31771=>"011110101",
  31772=>"110100101",
  31773=>"010101101",
  31774=>"000000110",
  31775=>"010000100",
  31776=>"011110111",
  31777=>"011010100",
  31778=>"110111110",
  31779=>"000100010",
  31780=>"110001101",
  31781=>"001011110",
  31782=>"010110000",
  31783=>"000011111",
  31784=>"110010000",
  31785=>"010001000",
  31786=>"100000000",
  31787=>"010111011",
  31788=>"100001010",
  31789=>"100001100",
  31790=>"010011110",
  31791=>"001011000",
  31792=>"000101001",
  31793=>"100101110",
  31794=>"010110001",
  31795=>"010000110",
  31796=>"111101100",
  31797=>"010100011",
  31798=>"001000010",
  31799=>"100001110",
  31800=>"100000000",
  31801=>"100010111",
  31802=>"010000111",
  31803=>"000101001",
  31804=>"110100001",
  31805=>"010110101",
  31806=>"010100011",
  31807=>"101100101",
  31808=>"001100100",
  31809=>"001000101",
  31810=>"101011111",
  31811=>"010111000",
  31812=>"101011010",
  31813=>"100011111",
  31814=>"010010111",
  31815=>"000110110",
  31816=>"001100011",
  31817=>"101111100",
  31818=>"110100100",
  31819=>"001010010",
  31820=>"001010110",
  31821=>"110000011",
  31822=>"111110000",
  31823=>"100100110",
  31824=>"101111010",
  31825=>"000011111",
  31826=>"001000110",
  31827=>"101101111",
  31828=>"110101111",
  31829=>"110011000",
  31830=>"011110000",
  31831=>"111011111",
  31832=>"011100111",
  31833=>"010101111",
  31834=>"101011100",
  31835=>"010011000",
  31836=>"001101010",
  31837=>"110100000",
  31838=>"000010000",
  31839=>"011011010",
  31840=>"010010001",
  31841=>"100110011",
  31842=>"001010101",
  31843=>"111110101",
  31844=>"011100101",
  31845=>"001000011",
  31846=>"110101010",
  31847=>"111011111",
  31848=>"110110001",
  31849=>"111110111",
  31850=>"010100100",
  31851=>"001000010",
  31852=>"001010010",
  31853=>"100010010",
  31854=>"100110110",
  31855=>"010000000",
  31856=>"111110011",
  31857=>"001001010",
  31858=>"110011000",
  31859=>"011100000",
  31860=>"101000010",
  31861=>"100001001",
  31862=>"001011101",
  31863=>"011000011",
  31864=>"010011111",
  31865=>"001000111",
  31866=>"100011010",
  31867=>"011001111",
  31868=>"011011010",
  31869=>"010101010",
  31870=>"101111111",
  31871=>"110011110",
  31872=>"010100001",
  31873=>"001011011",
  31874=>"010101000",
  31875=>"101000010",
  31876=>"100100000",
  31877=>"000001100",
  31878=>"101010110",
  31879=>"001101111",
  31880=>"000110100",
  31881=>"010010011",
  31882=>"011011001",
  31883=>"001010100",
  31884=>"000100001",
  31885=>"000010101",
  31886=>"100110110",
  31887=>"111101111",
  31888=>"111000101",
  31889=>"101100101",
  31890=>"011001110",
  31891=>"001101110",
  31892=>"101100111",
  31893=>"111100000",
  31894=>"101100100",
  31895=>"111010110",
  31896=>"101110000",
  31897=>"001001100",
  31898=>"000110001",
  31899=>"011111100",
  31900=>"001000010",
  31901=>"000001011",
  31902=>"011000110",
  31903=>"000101011",
  31904=>"100101001",
  31905=>"100010110",
  31906=>"001010011",
  31907=>"001011001",
  31908=>"101100001",
  31909=>"000111011",
  31910=>"000100000",
  31911=>"110000000",
  31912=>"111010101",
  31913=>"110010101",
  31914=>"110110001",
  31915=>"010101011",
  31916=>"100011000",
  31917=>"101110001",
  31918=>"110010100",
  31919=>"001010111",
  31920=>"000000110",
  31921=>"000010000",
  31922=>"010100110",
  31923=>"101100110",
  31924=>"001010010",
  31925=>"000100000",
  31926=>"111011000",
  31927=>"001010000",
  31928=>"001001100",
  31929=>"111010111",
  31930=>"111011010",
  31931=>"100100011",
  31932=>"001110010",
  31933=>"111111100",
  31934=>"000010001",
  31935=>"100110000",
  31936=>"111100110",
  31937=>"000011110",
  31938=>"100001101",
  31939=>"010101001",
  31940=>"011110001",
  31941=>"111110001",
  31942=>"101110101",
  31943=>"001010110",
  31944=>"000110110",
  31945=>"011111100",
  31946=>"010100001",
  31947=>"100100000",
  31948=>"011001110",
  31949=>"001011001",
  31950=>"010111011",
  31951=>"010000010",
  31952=>"110101110",
  31953=>"001001100",
  31954=>"001011000",
  31955=>"001000110",
  31956=>"001000000",
  31957=>"101001010",
  31958=>"110101110",
  31959=>"001100110",
  31960=>"101000110",
  31961=>"011111011",
  31962=>"001101100",
  31963=>"110011011",
  31964=>"000110111",
  31965=>"000010101",
  31966=>"100011000",
  31967=>"101110000",
  31968=>"010100100",
  31969=>"001011010",
  31970=>"101101110",
  31971=>"000000011",
  31972=>"110100000",
  31973=>"010101101",
  31974=>"011011101",
  31975=>"001000100",
  31976=>"111011010",
  31977=>"100010111",
  31978=>"111000110",
  31979=>"110010000",
  31980=>"010101110",
  31981=>"111101101",
  31982=>"110010100",
  31983=>"010000111",
  31984=>"011010001",
  31985=>"100111000",
  31986=>"000110000",
  31987=>"100100011",
  31988=>"000110110",
  31989=>"101110101",
  31990=>"001100110",
  31991=>"000110000",
  31992=>"101111111",
  31993=>"100001011",
  31994=>"001110111",
  31995=>"100110110",
  31996=>"000010000",
  31997=>"100110101",
  31998=>"101101000",
  31999=>"011110110",
  32000=>"100111011",
  32001=>"000100101",
  32002=>"001110111",
  32003=>"111101000",
  32004=>"100001100",
  32005=>"010101000",
  32006=>"110100000",
  32007=>"111101110",
  32008=>"011111001",
  32009=>"011101101",
  32010=>"000101010",
  32011=>"000001011",
  32012=>"100001000",
  32013=>"000101011",
  32014=>"000001001",
  32015=>"000111100",
  32016=>"110010011",
  32017=>"100101100",
  32018=>"010110110",
  32019=>"010100100",
  32020=>"011111101",
  32021=>"100101001",
  32022=>"100101010",
  32023=>"111110000",
  32024=>"001011010",
  32025=>"101111111",
  32026=>"101111000",
  32027=>"110101111",
  32028=>"010010100",
  32029=>"000000011",
  32030=>"100110011",
  32031=>"101000001",
  32032=>"100011011",
  32033=>"001011011",
  32034=>"000001101",
  32035=>"010011010",
  32036=>"100101111",
  32037=>"000111010",
  32038=>"010010100",
  32039=>"001101001",
  32040=>"110010111",
  32041=>"101100010",
  32042=>"100001000",
  32043=>"000101101",
  32044=>"000001110",
  32045=>"001111000",
  32046=>"100111011",
  32047=>"110111011",
  32048=>"111010111",
  32049=>"011100100",
  32050=>"010111101",
  32051=>"000001001",
  32052=>"001010101",
  32053=>"000111101",
  32054=>"001110000",
  32055=>"001010111",
  32056=>"110101111",
  32057=>"111001000",
  32058=>"000101111",
  32059=>"000010001",
  32060=>"001100010",
  32061=>"001110011",
  32062=>"001100001",
  32063=>"011110111",
  32064=>"110100111",
  32065=>"110111011",
  32066=>"111000011",
  32067=>"000110110",
  32068=>"011101011",
  32069=>"110100010",
  32070=>"010000010",
  32071=>"011110110",
  32072=>"100001110",
  32073=>"101100100",
  32074=>"000010010",
  32075=>"010100000",
  32076=>"001111110",
  32077=>"011100000",
  32078=>"111110000",
  32079=>"001001111",
  32080=>"001111001",
  32081=>"110111100",
  32082=>"100011111",
  32083=>"111110001",
  32084=>"010110100",
  32085=>"011010011",
  32086=>"011011101",
  32087=>"101101110",
  32088=>"111010000",
  32089=>"010100010",
  32090=>"011011001",
  32091=>"101000100",
  32092=>"010110111",
  32093=>"001010101",
  32094=>"000100000",
  32095=>"000011101",
  32096=>"001100111",
  32097=>"101110100",
  32098=>"111000111",
  32099=>"110110011",
  32100=>"000001010",
  32101=>"001101011",
  32102=>"111000010",
  32103=>"110101001",
  32104=>"100011111",
  32105=>"101111000",
  32106=>"111010001",
  32107=>"010001001",
  32108=>"000100010",
  32109=>"010000011",
  32110=>"010011000",
  32111=>"010110011",
  32112=>"101111010",
  32113=>"000011001",
  32114=>"111011011",
  32115=>"110100101",
  32116=>"011001100",
  32117=>"111111011",
  32118=>"000100111",
  32119=>"010010101",
  32120=>"110011110",
  32121=>"101100010",
  32122=>"010011010",
  32123=>"111001100",
  32124=>"111110110",
  32125=>"101100010",
  32126=>"101000100",
  32127=>"110101111",
  32128=>"111001100",
  32129=>"100001101",
  32130=>"101011011",
  32131=>"101000101",
  32132=>"001111100",
  32133=>"010001000",
  32134=>"110001010",
  32135=>"000111000",
  32136=>"011010100",
  32137=>"001010101",
  32138=>"001011101",
  32139=>"001101010",
  32140=>"001100011",
  32141=>"100111000",
  32142=>"100001000",
  32143=>"110111011",
  32144=>"101100100",
  32145=>"111011001",
  32146=>"000101001",
  32147=>"110100110",
  32148=>"110100010",
  32149=>"000110011",
  32150=>"101010111",
  32151=>"100011111",
  32152=>"100000100",
  32153=>"100000000",
  32154=>"111111011",
  32155=>"110001010",
  32156=>"001100100",
  32157=>"001010101",
  32158=>"101100011",
  32159=>"000010001",
  32160=>"011001110",
  32161=>"001000111",
  32162=>"010011100",
  32163=>"100010101",
  32164=>"001100010",
  32165=>"111011101",
  32166=>"011110000",
  32167=>"101001000",
  32168=>"111100100",
  32169=>"100010010",
  32170=>"010011111",
  32171=>"110101100",
  32172=>"001000101",
  32173=>"110100001",
  32174=>"110111101",
  32175=>"111000110",
  32176=>"100111110",
  32177=>"110100010",
  32178=>"111000000",
  32179=>"011000110",
  32180=>"111111110",
  32181=>"111010111",
  32182=>"000101111",
  32183=>"011101100",
  32184=>"101111010",
  32185=>"101010100",
  32186=>"000011011",
  32187=>"111001111",
  32188=>"000011000",
  32189=>"001111111",
  32190=>"101011010",
  32191=>"011000111",
  32192=>"000011011",
  32193=>"001000010",
  32194=>"000001010",
  32195=>"001001110",
  32196=>"101001110",
  32197=>"100000001",
  32198=>"000111010",
  32199=>"001010010",
  32200=>"001001000",
  32201=>"110011000",
  32202=>"101000010",
  32203=>"001010010",
  32204=>"101100000",
  32205=>"010011010",
  32206=>"111110011",
  32207=>"101100000",
  32208=>"100000010",
  32209=>"001010010",
  32210=>"000010100",
  32211=>"010111110",
  32212=>"001010010",
  32213=>"001111111",
  32214=>"010011101",
  32215=>"000001010",
  32216=>"011001001",
  32217=>"010101111",
  32218=>"110000101",
  32219=>"001001010",
  32220=>"010110010",
  32221=>"110000110",
  32222=>"001111000",
  32223=>"111101101",
  32224=>"000000111",
  32225=>"100011101",
  32226=>"111111001",
  32227=>"001000110",
  32228=>"101110001",
  32229=>"110101110",
  32230=>"011110111",
  32231=>"110110100",
  32232=>"100101110",
  32233=>"100011101",
  32234=>"110011110",
  32235=>"101111001",
  32236=>"001111010",
  32237=>"011111110",
  32238=>"111010101",
  32239=>"100110011",
  32240=>"001000111",
  32241=>"010000110",
  32242=>"111110001",
  32243=>"001000111",
  32244=>"011111001",
  32245=>"011110011",
  32246=>"110000000",
  32247=>"000101111",
  32248=>"011101111",
  32249=>"010100000",
  32250=>"010111111",
  32251=>"111011111",
  32252=>"000000000",
  32253=>"000000010",
  32254=>"110111110",
  32255=>"110010111",
  32256=>"001000100",
  32257=>"100001001",
  32258=>"011100110",
  32259=>"011101111",
  32260=>"101000101",
  32261=>"011010101",
  32262=>"001000111",
  32263=>"001100110",
  32264=>"100010110",
  32265=>"001101111",
  32266=>"101010011",
  32267=>"001001101",
  32268=>"010011111",
  32269=>"001111110",
  32270=>"101100010",
  32271=>"011011010",
  32272=>"001011111",
  32273=>"011011000",
  32274=>"111000100",
  32275=>"110010011",
  32276=>"010111110",
  32277=>"001110111",
  32278=>"101001011",
  32279=>"110011110",
  32280=>"000110010",
  32281=>"101100101",
  32282=>"000110110",
  32283=>"001110100",
  32284=>"001000010",
  32285=>"010010010",
  32286=>"010011000",
  32287=>"100001000",
  32288=>"000011100",
  32289=>"111000010",
  32290=>"101001011",
  32291=>"010001000",
  32292=>"101010011",
  32293=>"101000001",
  32294=>"111111101",
  32295=>"000000110",
  32296=>"010001111",
  32297=>"010011101",
  32298=>"001010010",
  32299=>"111010100",
  32300=>"001001000",
  32301=>"001101100",
  32302=>"011100110",
  32303=>"000010011",
  32304=>"110000101",
  32305=>"110110111",
  32306=>"000110111",
  32307=>"100010101",
  32308=>"101111010",
  32309=>"001111100",
  32310=>"000010110",
  32311=>"100000010",
  32312=>"011110010",
  32313=>"000000011",
  32314=>"001101011",
  32315=>"111111100",
  32316=>"010011001",
  32317=>"110111101",
  32318=>"101101000",
  32319=>"111000000",
  32320=>"110011110",
  32321=>"101010100",
  32322=>"000100000",
  32323=>"011100000",
  32324=>"101110100",
  32325=>"101110001",
  32326=>"001011100",
  32327=>"100101100",
  32328=>"010001100",
  32329=>"010111101",
  32330=>"001001101",
  32331=>"000001100",
  32332=>"001001111",
  32333=>"001111000",
  32334=>"010001011",
  32335=>"010010101",
  32336=>"110011101",
  32337=>"111101001",
  32338=>"110111101",
  32339=>"011101010",
  32340=>"010100100",
  32341=>"011110000",
  32342=>"000101110",
  32343=>"100001100",
  32344=>"111010110",
  32345=>"111001000",
  32346=>"010010110",
  32347=>"000100001",
  32348=>"000110011",
  32349=>"001000010",
  32350=>"011101011",
  32351=>"001011111",
  32352=>"011101100",
  32353=>"001011001",
  32354=>"111011001",
  32355=>"010000110",
  32356=>"110111100",
  32357=>"011000110",
  32358=>"110000100",
  32359=>"100111011",
  32360=>"000001010",
  32361=>"100100010",
  32362=>"000100100",
  32363=>"000110101",
  32364=>"111000000",
  32365=>"010010101",
  32366=>"111000001",
  32367=>"100010011",
  32368=>"001100110",
  32369=>"001101111",
  32370=>"111101011",
  32371=>"101111100",
  32372=>"101000101",
  32373=>"000111111",
  32374=>"011001110",
  32375=>"101011101",
  32376=>"011111110",
  32377=>"000011010",
  32378=>"011101111",
  32379=>"000101101",
  32380=>"110001010",
  32381=>"111100111",
  32382=>"100101100",
  32383=>"100010110",
  32384=>"110110110",
  32385=>"000110011",
  32386=>"101010001",
  32387=>"101110000",
  32388=>"011011011",
  32389=>"100100000",
  32390=>"011101100",
  32391=>"001000011",
  32392=>"011111001",
  32393=>"000101001",
  32394=>"011100001",
  32395=>"010101001",
  32396=>"001101000",
  32397=>"101101011",
  32398=>"101001001",
  32399=>"011110111",
  32400=>"111100111",
  32401=>"000010010",
  32402=>"110111110",
  32403=>"101110010",
  32404=>"000110011",
  32405=>"001001000",
  32406=>"110010101",
  32407=>"100010000",
  32408=>"110000000",
  32409=>"100000001",
  32410=>"000101000",
  32411=>"111101111",
  32412=>"111010111",
  32413=>"010000000",
  32414=>"100110100",
  32415=>"000000011",
  32416=>"111011011",
  32417=>"001001111",
  32418=>"011100100",
  32419=>"001010111",
  32420=>"001110000",
  32421=>"100001111",
  32422=>"010110010",
  32423=>"110010001",
  32424=>"000000010",
  32425=>"000111001",
  32426=>"101111000",
  32427=>"101100111",
  32428=>"110110111",
  32429=>"111100000",
  32430=>"100110001",
  32431=>"100010111",
  32432=>"110110101",
  32433=>"000000010",
  32434=>"101010101",
  32435=>"111010101",
  32436=>"001000000",
  32437=>"111000110",
  32438=>"000111110",
  32439=>"111101000",
  32440=>"111101101",
  32441=>"111001000",
  32442=>"011111001",
  32443=>"011000011",
  32444=>"001000111",
  32445=>"010000011",
  32446=>"110111001",
  32447=>"111010001",
  32448=>"010000000",
  32449=>"010010011",
  32450=>"000010110",
  32451=>"011101101",
  32452=>"110001001",
  32453=>"000010110",
  32454=>"011011111",
  32455=>"000111001",
  32456=>"110101000",
  32457=>"100101111",
  32458=>"000011001",
  32459=>"011110001",
  32460=>"100010011",
  32461=>"001111011",
  32462=>"100101000",
  32463=>"101101101",
  32464=>"000011110",
  32465=>"110000010",
  32466=>"001101110",
  32467=>"110011110",
  32468=>"001110101",
  32469=>"110011100",
  32470=>"101100000",
  32471=>"100000001",
  32472=>"010000110",
  32473=>"111111101",
  32474=>"000000011",
  32475=>"101001100",
  32476=>"001010111",
  32477=>"000001001",
  32478=>"110111111",
  32479=>"011001001",
  32480=>"100110111",
  32481=>"001101000",
  32482=>"110011100",
  32483=>"001011000",
  32484=>"000000101",
  32485=>"001100010",
  32486=>"100111110",
  32487=>"101111110",
  32488=>"010001101",
  32489=>"010001110",
  32490=>"001001111",
  32491=>"110100000",
  32492=>"110100011",
  32493=>"000101000",
  32494=>"111001101",
  32495=>"101101011",
  32496=>"110110101",
  32497=>"110101101",
  32498=>"101110010",
  32499=>"000100111",
  32500=>"011001000",
  32501=>"011101101",
  32502=>"100111001",
  32503=>"001100111",
  32504=>"001001000",
  32505=>"110001100",
  32506=>"110110011",
  32507=>"000010001",
  32508=>"000001000",
  32509=>"000000101",
  32510=>"111011101",
  32511=>"000011111",
  32512=>"101000111",
  32513=>"111110011",
  32514=>"000111000",
  32515=>"111100101",
  32516=>"101011100",
  32517=>"111110010",
  32518=>"110111111",
  32519=>"010100110",
  32520=>"010010111",
  32521=>"110001000",
  32522=>"101100101",
  32523=>"111100001",
  32524=>"110110011",
  32525=>"101110000",
  32526=>"100101100",
  32527=>"111101110",
  32528=>"100010011",
  32529=>"000100100",
  32530=>"110110010",
  32531=>"100010000",
  32532=>"000011000",
  32533=>"110010100",
  32534=>"001001111",
  32535=>"011110011",
  32536=>"101111110",
  32537=>"111110100",
  32538=>"101010100",
  32539=>"110111110",
  32540=>"111101101",
  32541=>"110000000",
  32542=>"111011011",
  32543=>"000000011",
  32544=>"111000010",
  32545=>"110110110",
  32546=>"101100100",
  32547=>"000111000",
  32548=>"111111010",
  32549=>"001010110",
  32550=>"000001011",
  32551=>"001010110",
  32552=>"111111101",
  32553=>"100101110",
  32554=>"010010111",
  32555=>"010011110",
  32556=>"100100010",
  32557=>"001010011",
  32558=>"000010010",
  32559=>"111001011",
  32560=>"101000110",
  32561=>"001111110",
  32562=>"101111101",
  32563=>"011000001",
  32564=>"000000001",
  32565=>"111100000",
  32566=>"011101100",
  32567=>"111001011",
  32568=>"110101101",
  32569=>"111011110",
  32570=>"001001101",
  32571=>"110000001",
  32572=>"111101100",
  32573=>"100010100",
  32574=>"000010001",
  32575=>"110110101",
  32576=>"001100100",
  32577=>"000111111",
  32578=>"101101110",
  32579=>"101111100",
  32580=>"100101010",
  32581=>"110011000",
  32582=>"000101010",
  32583=>"000000101",
  32584=>"000100010",
  32585=>"000011100",
  32586=>"100010101",
  32587=>"010001100",
  32588=>"011000101",
  32589=>"111110111",
  32590=>"000101010",
  32591=>"101000100",
  32592=>"000111010",
  32593=>"110100110",
  32594=>"101101101",
  32595=>"000000010",
  32596=>"101011001",
  32597=>"100110010",
  32598=>"000011010",
  32599=>"100011100",
  32600=>"111110011",
  32601=>"101000101",
  32602=>"011111011",
  32603=>"000101100",
  32604=>"000100101",
  32605=>"111011011",
  32606=>"111000000",
  32607=>"000100101",
  32608=>"110001001",
  32609=>"100010111",
  32610=>"001001100",
  32611=>"110000011",
  32612=>"011010100",
  32613=>"100001011",
  32614=>"011101110",
  32615=>"001101110",
  32616=>"100010000",
  32617=>"110101110",
  32618=>"011111100",
  32619=>"000001100",
  32620=>"111011100",
  32621=>"111110000",
  32622=>"111011000",
  32623=>"110010001",
  32624=>"011001010",
  32625=>"110110110",
  32626=>"100100010",
  32627=>"011100100",
  32628=>"100000010",
  32629=>"110101011",
  32630=>"001101001",
  32631=>"000110011",
  32632=>"001100111",
  32633=>"011001110",
  32634=>"110001000",
  32635=>"010111001",
  32636=>"000110100",
  32637=>"101111000",
  32638=>"111111011",
  32639=>"101001101",
  32640=>"110000110",
  32641=>"101010111",
  32642=>"010001111",
  32643=>"110001110",
  32644=>"010100111",
  32645=>"000001110",
  32646=>"010001010",
  32647=>"011011011",
  32648=>"010000010",
  32649=>"111111110",
  32650=>"111100110",
  32651=>"010100001",
  32652=>"001000000",
  32653=>"010000011",
  32654=>"000110011",
  32655=>"100110101",
  32656=>"111011101",
  32657=>"100101010",
  32658=>"001110101",
  32659=>"010111111",
  32660=>"101001000",
  32661=>"100100011",
  32662=>"010000001",
  32663=>"101110011",
  32664=>"000010101",
  32665=>"111101101",
  32666=>"111111010",
  32667=>"010110100",
  32668=>"011111000",
  32669=>"101101010",
  32670=>"001101011",
  32671=>"111001011",
  32672=>"000000011",
  32673=>"100110111",
  32674=>"101001001",
  32675=>"101110100",
  32676=>"100011110",
  32677=>"000110100",
  32678=>"001000110",
  32679=>"100000110",
  32680=>"101110110",
  32681=>"000000000",
  32682=>"101100100",
  32683=>"111001100",
  32684=>"010100111",
  32685=>"010100110",
  32686=>"101101110",
  32687=>"010110010",
  32688=>"111111001",
  32689=>"100010011",
  32690=>"000011011",
  32691=>"010111011",
  32692=>"000110100",
  32693=>"100000100",
  32694=>"111001111",
  32695=>"000011010",
  32696=>"001111100",
  32697=>"000100110",
  32698=>"100011110",
  32699=>"001110010",
  32700=>"011011110",
  32701=>"100000110",
  32702=>"111111111",
  32703=>"101000000",
  32704=>"010000001",
  32705=>"111000100",
  32706=>"001001001",
  32707=>"110101111",
  32708=>"001001100",
  32709=>"011001111",
  32710=>"111101101",
  32711=>"100010100",
  32712=>"001001001",
  32713=>"100000011",
  32714=>"011001001",
  32715=>"101001110",
  32716=>"111011101",
  32717=>"101101011",
  32718=>"000111111",
  32719=>"010100011",
  32720=>"110101110",
  32721=>"000100001",
  32722=>"100000011",
  32723=>"110011100",
  32724=>"001100000",
  32725=>"010001010",
  32726=>"101011100",
  32727=>"010010001",
  32728=>"111111011",
  32729=>"011001110",
  32730=>"101000010",
  32731=>"111000011",
  32732=>"101001100",
  32733=>"101111000",
  32734=>"000111011",
  32735=>"111011010",
  32736=>"110101100",
  32737=>"001101110",
  32738=>"110100011",
  32739=>"001010110",
  32740=>"010111000",
  32741=>"000000111",
  32742=>"001111010",
  32743=>"000010100",
  32744=>"011010000",
  32745=>"100000010",
  32746=>"101000010",
  32747=>"000110010",
  32748=>"000100000",
  32749=>"010100011",
  32750=>"100101010",
  32751=>"101110000",
  32752=>"001110001",
  32753=>"010110101",
  32754=>"010101100",
  32755=>"101011001",
  32756=>"110001110",
  32757=>"111000001",
  32758=>"110110001",
  32759=>"001010011",
  32760=>"100000010",
  32761=>"111000000",
  32762=>"100110010",
  32763=>"101101111",
  32764=>"010000111",
  32765=>"010001100",
  32766=>"001011011",
  32767=>"000111010",
  32768=>"001000001",
  32769=>"011110000",
  32770=>"100100101",
  32771=>"111010001",
  32772=>"101100000",
  32773=>"000101111",
  32774=>"000100110",
  32775=>"100001100",
  32776=>"110100110",
  32777=>"010110011",
  32778=>"001110000",
  32779=>"101111010",
  32780=>"010111111",
  32781=>"010000000",
  32782=>"010110011",
  32783=>"010010111",
  32784=>"010110011",
  32785=>"010101000",
  32786=>"110111101",
  32787=>"010000101",
  32788=>"001110011",
  32789=>"000111101",
  32790=>"000001110",
  32791=>"011100110",
  32792=>"001001010",
  32793=>"100011000",
  32794=>"000101001",
  32795=>"011110010",
  32796=>"001110000",
  32797=>"011001011",
  32798=>"100011001",
  32799=>"010001010",
  32800=>"101110010",
  32801=>"001010011",
  32802=>"101011011",
  32803=>"101011100",
  32804=>"111101100",
  32805=>"100110111",
  32806=>"000001100",
  32807=>"110011001",
  32808=>"010010000",
  32809=>"111110110",
  32810=>"101010000",
  32811=>"011010111",
  32812=>"101011000",
  32813=>"100001101",
  32814=>"010011100",
  32815=>"110001110",
  32816=>"101111010",
  32817=>"010011011",
  32818=>"010001101",
  32819=>"000010110",
  32820=>"111100000",
  32821=>"011100001",
  32822=>"110010110",
  32823=>"101101100",
  32824=>"001000001",
  32825=>"101111101",
  32826=>"111010000",
  32827=>"100101011",
  32828=>"000001010",
  32829=>"001000000",
  32830=>"101000101",
  32831=>"011000110",
  32832=>"110010100",
  32833=>"001100111",
  32834=>"100101110",
  32835=>"101001011",
  32836=>"001110011",
  32837=>"100001101",
  32838=>"101111101",
  32839=>"100010011",
  32840=>"001000111",
  32841=>"100110010",
  32842=>"110100010",
  32843=>"011110010",
  32844=>"101000010",
  32845=>"111111010",
  32846=>"101111000",
  32847=>"110101111",
  32848=>"100111110",
  32849=>"010100110",
  32850=>"010101100",
  32851=>"011111000",
  32852=>"101101101",
  32853=>"001010101",
  32854=>"101100011",
  32855=>"100000001",
  32856=>"100101111",
  32857=>"110000110",
  32858=>"000100001",
  32859=>"000001111",
  32860=>"011000010",
  32861=>"000110010",
  32862=>"011000010",
  32863=>"000011111",
  32864=>"001110110",
  32865=>"001111000",
  32866=>"011100100",
  32867=>"000000000",
  32868=>"010001010",
  32869=>"101100100",
  32870=>"011100100",
  32871=>"011111101",
  32872=>"100000011",
  32873=>"111111101",
  32874=>"110000110",
  32875=>"001100110",
  32876=>"010111110",
  32877=>"010100100",
  32878=>"100011101",
  32879=>"100011000",
  32880=>"111001100",
  32881=>"111010011",
  32882=>"111000000",
  32883=>"011111011",
  32884=>"001011110",
  32885=>"100111000",
  32886=>"111010101",
  32887=>"111001000",
  32888=>"000100111",
  32889=>"010001101",
  32890=>"010110110",
  32891=>"101111100",
  32892=>"010001011",
  32893=>"111100101",
  32894=>"100110000",
  32895=>"010110001",
  32896=>"100100010",
  32897=>"011100000",
  32898=>"011001101",
  32899=>"001110010",
  32900=>"010010011",
  32901=>"000101010",
  32902=>"000100100",
  32903=>"101111101",
  32904=>"000011000",
  32905=>"011010001",
  32906=>"010010000",
  32907=>"000110000",
  32908=>"111111110",
  32909=>"101111100",
  32910=>"010001000",
  32911=>"111000101",
  32912=>"010001000",
  32913=>"110101001",
  32914=>"011110111",
  32915=>"111000110",
  32916=>"111111111",
  32917=>"101101000",
  32918=>"010100010",
  32919=>"010100011",
  32920=>"110000011",
  32921=>"011101100",
  32922=>"011110101",
  32923=>"110010101",
  32924=>"010100111",
  32925=>"001000110",
  32926=>"010100110",
  32927=>"110110110",
  32928=>"011001010",
  32929=>"100100010",
  32930=>"111111001",
  32931=>"000100110",
  32932=>"111100011",
  32933=>"001110010",
  32934=>"010100001",
  32935=>"011010011",
  32936=>"111001111",
  32937=>"000000010",
  32938=>"010010000",
  32939=>"011001100",
  32940=>"100000100",
  32941=>"110101111",
  32942=>"110001000",
  32943=>"000001011",
  32944=>"000101101",
  32945=>"111111001",
  32946=>"000000010",
  32947=>"001100101",
  32948=>"100001000",
  32949=>"111010010",
  32950=>"100100111",
  32951=>"110000011",
  32952=>"010000111",
  32953=>"000100100",
  32954=>"101010101",
  32955=>"000110101",
  32956=>"101101010",
  32957=>"001000111",
  32958=>"001101001",
  32959=>"101111001",
  32960=>"001011011",
  32961=>"010010011",
  32962=>"101010010",
  32963=>"001001111",
  32964=>"111110110",
  32965=>"000000010",
  32966=>"011111110",
  32967=>"001111001",
  32968=>"101101001",
  32969=>"010011011",
  32970=>"001011011",
  32971=>"100011010",
  32972=>"101110110",
  32973=>"110010100",
  32974=>"001111101",
  32975=>"001101010",
  32976=>"110101010",
  32977=>"000010010",
  32978=>"001001110",
  32979=>"101111110",
  32980=>"011101011",
  32981=>"110001100",
  32982=>"100110010",
  32983=>"011001101",
  32984=>"100110111",
  32985=>"111101101",
  32986=>"101101111",
  32987=>"011111101",
  32988=>"101010001",
  32989=>"010100100",
  32990=>"011001100",
  32991=>"100100011",
  32992=>"101111110",
  32993=>"000010111",
  32994=>"010011100",
  32995=>"100110111",
  32996=>"000000111",
  32997=>"000111010",
  32998=>"000001001",
  32999=>"010100111",
  33000=>"011010111",
  33001=>"000100010",
  33002=>"010110011",
  33003=>"110101001",
  33004=>"111111111",
  33005=>"111010110",
  33006=>"011111011",
  33007=>"101001000",
  33008=>"100100010",
  33009=>"011010011",
  33010=>"111000000",
  33011=>"111010000",
  33012=>"110101001",
  33013=>"111110111",
  33014=>"100000100",
  33015=>"110001101",
  33016=>"110010101",
  33017=>"111101000",
  33018=>"000000100",
  33019=>"101010101",
  33020=>"110111100",
  33021=>"101111011",
  33022=>"010101111",
  33023=>"101101101",
  33024=>"011010001",
  33025=>"101110001",
  33026=>"011101110",
  33027=>"100011011",
  33028=>"100011010",
  33029=>"101101101",
  33030=>"111011110",
  33031=>"100010000",
  33032=>"010100000",
  33033=>"111000011",
  33034=>"111000100",
  33035=>"100001000",
  33036=>"110100010",
  33037=>"010011010",
  33038=>"000101111",
  33039=>"111100001",
  33040=>"000110000",
  33041=>"010001110",
  33042=>"111001100",
  33043=>"000111011",
  33044=>"110101110",
  33045=>"000111000",
  33046=>"100001010",
  33047=>"001101100",
  33048=>"101110000",
  33049=>"110010111",
  33050=>"001101110",
  33051=>"110100100",
  33052=>"100001000",
  33053=>"100010111",
  33054=>"100111110",
  33055=>"111001111",
  33056=>"100011100",
  33057=>"111000010",
  33058=>"111101010",
  33059=>"001101000",
  33060=>"001011001",
  33061=>"011101101",
  33062=>"110011111",
  33063=>"110010000",
  33064=>"110010001",
  33065=>"110111110",
  33066=>"010010010",
  33067=>"010000101",
  33068=>"011011001",
  33069=>"000101100",
  33070=>"000000000",
  33071=>"101100011",
  33072=>"011001010",
  33073=>"011111111",
  33074=>"101001010",
  33075=>"010110110",
  33076=>"010101101",
  33077=>"011110000",
  33078=>"011010010",
  33079=>"101111101",
  33080=>"101001011",
  33081=>"000001011",
  33082=>"000110110",
  33083=>"011001011",
  33084=>"111011000",
  33085=>"001110110",
  33086=>"011000111",
  33087=>"010000000",
  33088=>"010011001",
  33089=>"101100000",
  33090=>"101111001",
  33091=>"010011100",
  33092=>"111001010",
  33093=>"011111101",
  33094=>"001101111",
  33095=>"011000111",
  33096=>"110101010",
  33097=>"001101110",
  33098=>"010111110",
  33099=>"101000111",
  33100=>"110000110",
  33101=>"110000011",
  33102=>"111110110",
  33103=>"011111111",
  33104=>"000000100",
  33105=>"100101000",
  33106=>"000000011",
  33107=>"111010101",
  33108=>"010011000",
  33109=>"100011001",
  33110=>"101011111",
  33111=>"101110011",
  33112=>"000001101",
  33113=>"110101001",
  33114=>"010110001",
  33115=>"011011001",
  33116=>"011000011",
  33117=>"110001001",
  33118=>"100110001",
  33119=>"011111100",
  33120=>"000111000",
  33121=>"111110001",
  33122=>"010011000",
  33123=>"001100110",
  33124=>"000100011",
  33125=>"100011101",
  33126=>"111110100",
  33127=>"001110011",
  33128=>"000111100",
  33129=>"110000001",
  33130=>"010111100",
  33131=>"100111010",
  33132=>"111001110",
  33133=>"000000110",
  33134=>"001010111",
  33135=>"111101101",
  33136=>"101110000",
  33137=>"111101011",
  33138=>"110001000",
  33139=>"111111011",
  33140=>"111101000",
  33141=>"111111101",
  33142=>"111101011",
  33143=>"101111110",
  33144=>"010011000",
  33145=>"111000010",
  33146=>"110011000",
  33147=>"001010011",
  33148=>"100111000",
  33149=>"101001110",
  33150=>"010101101",
  33151=>"000011010",
  33152=>"010011111",
  33153=>"000110010",
  33154=>"010111001",
  33155=>"000010110",
  33156=>"110000100",
  33157=>"100101001",
  33158=>"101000001",
  33159=>"011001111",
  33160=>"001110110",
  33161=>"101101110",
  33162=>"010000111",
  33163=>"111011011",
  33164=>"001001001",
  33165=>"101001001",
  33166=>"101110000",
  33167=>"101111000",
  33168=>"101101100",
  33169=>"000101011",
  33170=>"111111111",
  33171=>"001000001",
  33172=>"011010101",
  33173=>"110000100",
  33174=>"111010001",
  33175=>"001100110",
  33176=>"010100011",
  33177=>"101010100",
  33178=>"100011010",
  33179=>"001101001",
  33180=>"101001001",
  33181=>"001110101",
  33182=>"000110101",
  33183=>"011000101",
  33184=>"010000011",
  33185=>"010100000",
  33186=>"001011011",
  33187=>"110001010",
  33188=>"001001001",
  33189=>"100000000",
  33190=>"101110100",
  33191=>"100110101",
  33192=>"011001011",
  33193=>"111001011",
  33194=>"111100011",
  33195=>"001000001",
  33196=>"101010001",
  33197=>"001100010",
  33198=>"110100010",
  33199=>"111110001",
  33200=>"100110011",
  33201=>"100110000",
  33202=>"000111101",
  33203=>"001100101",
  33204=>"000100001",
  33205=>"100001111",
  33206=>"000111101",
  33207=>"110110110",
  33208=>"010100011",
  33209=>"001010101",
  33210=>"001111101",
  33211=>"110010111",
  33212=>"011010100",
  33213=>"100101010",
  33214=>"101100100",
  33215=>"100100001",
  33216=>"000000010",
  33217=>"100001111",
  33218=>"010110100",
  33219=>"111001011",
  33220=>"011011101",
  33221=>"001100011",
  33222=>"011101110",
  33223=>"011011111",
  33224=>"101101001",
  33225=>"000000100",
  33226=>"001111010",
  33227=>"111001111",
  33228=>"100000111",
  33229=>"111010101",
  33230=>"000100111",
  33231=>"010011000",
  33232=>"111010011",
  33233=>"111111001",
  33234=>"010101000",
  33235=>"111100100",
  33236=>"111101010",
  33237=>"000010000",
  33238=>"011010010",
  33239=>"111101000",
  33240=>"010000111",
  33241=>"110000100",
  33242=>"101011100",
  33243=>"111110100",
  33244=>"111110111",
  33245=>"101110110",
  33246=>"010001001",
  33247=>"111110101",
  33248=>"001100111",
  33249=>"111011011",
  33250=>"011111101",
  33251=>"110110010",
  33252=>"100101001",
  33253=>"100000101",
  33254=>"011011011",
  33255=>"100011001",
  33256=>"010000001",
  33257=>"110110000",
  33258=>"011101110",
  33259=>"001001010",
  33260=>"100011100",
  33261=>"011010000",
  33262=>"000100011",
  33263=>"000010010",
  33264=>"111010111",
  33265=>"011111110",
  33266=>"101110111",
  33267=>"011111001",
  33268=>"000101111",
  33269=>"000101100",
  33270=>"111101100",
  33271=>"110011101",
  33272=>"000000101",
  33273=>"111111101",
  33274=>"000101001",
  33275=>"100010111",
  33276=>"011111111",
  33277=>"001011001",
  33278=>"010100011",
  33279=>"001000010",
  33280=>"001111010",
  33281=>"010100000",
  33282=>"101011010",
  33283=>"001101010",
  33284=>"101000101",
  33285=>"111101111",
  33286=>"010000001",
  33287=>"001000000",
  33288=>"101100000",
  33289=>"010010100",
  33290=>"011010010",
  33291=>"011001000",
  33292=>"100101111",
  33293=>"010101011",
  33294=>"000010101",
  33295=>"111010101",
  33296=>"000100011",
  33297=>"100110110",
  33298=>"100000011",
  33299=>"000001111",
  33300=>"101001110",
  33301=>"011010101",
  33302=>"100010001",
  33303=>"110111000",
  33304=>"111011000",
  33305=>"000011001",
  33306=>"001001101",
  33307=>"111111111",
  33308=>"000100110",
  33309=>"111111011",
  33310=>"011110100",
  33311=>"110000001",
  33312=>"100110001",
  33313=>"011011110",
  33314=>"011010101",
  33315=>"001011111",
  33316=>"110111011",
  33317=>"100101010",
  33318=>"001000111",
  33319=>"100101110",
  33320=>"010010000",
  33321=>"001111110",
  33322=>"110100101",
  33323=>"010100011",
  33324=>"110110010",
  33325=>"011000111",
  33326=>"010100011",
  33327=>"000101101",
  33328=>"011000010",
  33329=>"110111111",
  33330=>"111101101",
  33331=>"100110011",
  33332=>"000100011",
  33333=>"011111100",
  33334=>"100010101",
  33335=>"111001101",
  33336=>"101100001",
  33337=>"110010101",
  33338=>"010111100",
  33339=>"110010011",
  33340=>"001011101",
  33341=>"010101110",
  33342=>"111100010",
  33343=>"011110111",
  33344=>"000100010",
  33345=>"110011111",
  33346=>"011001010",
  33347=>"110111101",
  33348=>"111111111",
  33349=>"111010000",
  33350=>"000101111",
  33351=>"000001010",
  33352=>"010100010",
  33353=>"110000000",
  33354=>"000101001",
  33355=>"111011011",
  33356=>"101010111",
  33357=>"100010011",
  33358=>"011110111",
  33359=>"000001001",
  33360=>"100101100",
  33361=>"111010010",
  33362=>"011001110",
  33363=>"110000011",
  33364=>"001001001",
  33365=>"110110100",
  33366=>"100111010",
  33367=>"101010010",
  33368=>"001110010",
  33369=>"000101110",
  33370=>"100101110",
  33371=>"000000100",
  33372=>"000010101",
  33373=>"001101101",
  33374=>"011111101",
  33375=>"000000110",
  33376=>"011000111",
  33377=>"101110000",
  33378=>"000101111",
  33379=>"001110100",
  33380=>"110111011",
  33381=>"001000011",
  33382=>"111101011",
  33383=>"100000010",
  33384=>"000000010",
  33385=>"110010100",
  33386=>"010100111",
  33387=>"000101110",
  33388=>"111010000",
  33389=>"110101000",
  33390=>"010110111",
  33391=>"001001101",
  33392=>"011111111",
  33393=>"001110110",
  33394=>"001111010",
  33395=>"011101111",
  33396=>"000011101",
  33397=>"001000101",
  33398=>"111110110",
  33399=>"111110011",
  33400=>"010010111",
  33401=>"011010110",
  33402=>"011111000",
  33403=>"111110111",
  33404=>"111001000",
  33405=>"101000000",
  33406=>"111010011",
  33407=>"001000010",
  33408=>"001001000",
  33409=>"111100001",
  33410=>"011010000",
  33411=>"100000111",
  33412=>"111100001",
  33413=>"111101100",
  33414=>"100111110",
  33415=>"000100001",
  33416=>"100001011",
  33417=>"100111100",
  33418=>"110100101",
  33419=>"101111110",
  33420=>"011000000",
  33421=>"010101111",
  33422=>"111111100",
  33423=>"111101010",
  33424=>"111110100",
  33425=>"111010010",
  33426=>"100010001",
  33427=>"110100000",
  33428=>"000000110",
  33429=>"001110101",
  33430=>"000001001",
  33431=>"000001111",
  33432=>"001000011",
  33433=>"010001001",
  33434=>"110001000",
  33435=>"101100110",
  33436=>"100110110",
  33437=>"111000100",
  33438=>"110000001",
  33439=>"000110011",
  33440=>"011000010",
  33441=>"000011000",
  33442=>"011001111",
  33443=>"000111110",
  33444=>"011001110",
  33445=>"111101001",
  33446=>"111011011",
  33447=>"111000101",
  33448=>"110111100",
  33449=>"010101101",
  33450=>"000111011",
  33451=>"111010000",
  33452=>"010011011",
  33453=>"000011010",
  33454=>"100000101",
  33455=>"010101111",
  33456=>"011000011",
  33457=>"001011010",
  33458=>"011001001",
  33459=>"110110000",
  33460=>"010010100",
  33461=>"000111000",
  33462=>"001110001",
  33463=>"000111111",
  33464=>"011000011",
  33465=>"010000110",
  33466=>"010101011",
  33467=>"111010010",
  33468=>"001001111",
  33469=>"101001101",
  33470=>"001101010",
  33471=>"110100100",
  33472=>"011010010",
  33473=>"111100010",
  33474=>"101010000",
  33475=>"111100001",
  33476=>"110010100",
  33477=>"110010111",
  33478=>"000111010",
  33479=>"001011110",
  33480=>"110101100",
  33481=>"010100111",
  33482=>"100000110",
  33483=>"100111110",
  33484=>"110110010",
  33485=>"000000001",
  33486=>"100011000",
  33487=>"000011110",
  33488=>"011001100",
  33489=>"111001101",
  33490=>"010111000",
  33491=>"101000110",
  33492=>"001100011",
  33493=>"001011110",
  33494=>"010010001",
  33495=>"100011011",
  33496=>"000111000",
  33497=>"111011110",
  33498=>"011101011",
  33499=>"111111110",
  33500=>"100101010",
  33501=>"011010101",
  33502=>"100101011",
  33503=>"110000011",
  33504=>"001100011",
  33505=>"010100100",
  33506=>"100011110",
  33507=>"100111110",
  33508=>"101110101",
  33509=>"110010010",
  33510=>"010101110",
  33511=>"001000011",
  33512=>"100000011",
  33513=>"101000011",
  33514=>"000011000",
  33515=>"001010101",
  33516=>"000000010",
  33517=>"000000110",
  33518=>"110101000",
  33519=>"110010001",
  33520=>"001111100",
  33521=>"111100000",
  33522=>"111000000",
  33523=>"111001001",
  33524=>"111111011",
  33525=>"110010111",
  33526=>"000100010",
  33527=>"011100101",
  33528=>"011010010",
  33529=>"101010100",
  33530=>"110011100",
  33531=>"001011010",
  33532=>"110101111",
  33533=>"000101000",
  33534=>"001000001",
  33535=>"110000001",
  33536=>"000001011",
  33537=>"110010100",
  33538=>"101101000",
  33539=>"011000000",
  33540=>"111101101",
  33541=>"101001110",
  33542=>"010010000",
  33543=>"001110110",
  33544=>"101011001",
  33545=>"111001110",
  33546=>"110010100",
  33547=>"001011001",
  33548=>"001001100",
  33549=>"111100110",
  33550=>"110010100",
  33551=>"001011110",
  33552=>"100110001",
  33553=>"100010011",
  33554=>"010010011",
  33555=>"010011110",
  33556=>"101101001",
  33557=>"011010000",
  33558=>"000011110",
  33559=>"010010000",
  33560=>"101110000",
  33561=>"000011000",
  33562=>"010100111",
  33563=>"010111001",
  33564=>"101100010",
  33565=>"010100011",
  33566=>"010010011",
  33567=>"010101101",
  33568=>"100100001",
  33569=>"101010110",
  33570=>"001000101",
  33571=>"011110010",
  33572=>"110001100",
  33573=>"010000011",
  33574=>"110000001",
  33575=>"010010100",
  33576=>"111111101",
  33577=>"000111100",
  33578=>"100100100",
  33579=>"010100010",
  33580=>"101101101",
  33581=>"110111011",
  33582=>"000101010",
  33583=>"001000100",
  33584=>"001101100",
  33585=>"011000001",
  33586=>"001110100",
  33587=>"111000101",
  33588=>"011101101",
  33589=>"010101111",
  33590=>"101101111",
  33591=>"100100010",
  33592=>"111110111",
  33593=>"100001000",
  33594=>"110110100",
  33595=>"111000111",
  33596=>"111000110",
  33597=>"100110001",
  33598=>"100100001",
  33599=>"011011000",
  33600=>"011010111",
  33601=>"100101101",
  33602=>"011001111",
  33603=>"011011001",
  33604=>"011111001",
  33605=>"100000001",
  33606=>"001100000",
  33607=>"010110010",
  33608=>"000110101",
  33609=>"110110000",
  33610=>"111111011",
  33611=>"010010110",
  33612=>"000001001",
  33613=>"011111101",
  33614=>"000100010",
  33615=>"111110011",
  33616=>"011101010",
  33617=>"000100110",
  33618=>"011000000",
  33619=>"001001100",
  33620=>"000011101",
  33621=>"000000011",
  33622=>"111000000",
  33623=>"101011000",
  33624=>"101100111",
  33625=>"000000001",
  33626=>"000100000",
  33627=>"100110000",
  33628=>"000000100",
  33629=>"100111111",
  33630=>"011010000",
  33631=>"010100111",
  33632=>"101010111",
  33633=>"010110110",
  33634=>"110100011",
  33635=>"100000110",
  33636=>"110101010",
  33637=>"001000111",
  33638=>"010111100",
  33639=>"011010111",
  33640=>"111101001",
  33641=>"011111010",
  33642=>"100000100",
  33643=>"001110000",
  33644=>"010110010",
  33645=>"010011010",
  33646=>"111111000",
  33647=>"101001011",
  33648=>"110110000",
  33649=>"011000000",
  33650=>"110000010",
  33651=>"100011101",
  33652=>"101111100",
  33653=>"001111000",
  33654=>"001101100",
  33655=>"110011000",
  33656=>"100010010",
  33657=>"111110100",
  33658=>"100110001",
  33659=>"110110111",
  33660=>"110011000",
  33661=>"001010100",
  33662=>"010010000",
  33663=>"010011000",
  33664=>"001101001",
  33665=>"100010101",
  33666=>"100000111",
  33667=>"010100011",
  33668=>"000001000",
  33669=>"111001010",
  33670=>"100111101",
  33671=>"010101001",
  33672=>"110000001",
  33673=>"001001001",
  33674=>"111010011",
  33675=>"000101000",
  33676=>"000001110",
  33677=>"110000100",
  33678=>"001010010",
  33679=>"100111111",
  33680=>"011000100",
  33681=>"100000001",
  33682=>"000011110",
  33683=>"100000011",
  33684=>"001000001",
  33685=>"100111100",
  33686=>"010110100",
  33687=>"001100101",
  33688=>"101010100",
  33689=>"000111100",
  33690=>"100001001",
  33691=>"110010010",
  33692=>"001011111",
  33693=>"101101000",
  33694=>"010100111",
  33695=>"011100011",
  33696=>"000010011",
  33697=>"000100101",
  33698=>"010100110",
  33699=>"110110100",
  33700=>"010110000",
  33701=>"001001011",
  33702=>"111111011",
  33703=>"110101011",
  33704=>"000100000",
  33705=>"000110100",
  33706=>"110100100",
  33707=>"100110111",
  33708=>"000000010",
  33709=>"011111011",
  33710=>"001000011",
  33711=>"110101011",
  33712=>"111001100",
  33713=>"011011101",
  33714=>"011011101",
  33715=>"000000010",
  33716=>"001011011",
  33717=>"111100001",
  33718=>"101111100",
  33719=>"001010000",
  33720=>"010100100",
  33721=>"101101111",
  33722=>"011000010",
  33723=>"001010000",
  33724=>"111101100",
  33725=>"010110010",
  33726=>"011010111",
  33727=>"111001110",
  33728=>"100011011",
  33729=>"000001000",
  33730=>"000011001",
  33731=>"111110010",
  33732=>"001111111",
  33733=>"000110010",
  33734=>"110100001",
  33735=>"101100110",
  33736=>"110000101",
  33737=>"101100110",
  33738=>"000011110",
  33739=>"011111111",
  33740=>"001010110",
  33741=>"100000010",
  33742=>"110111100",
  33743=>"001000010",
  33744=>"011100110",
  33745=>"001011011",
  33746=>"011000000",
  33747=>"000001000",
  33748=>"100000110",
  33749=>"100001101",
  33750=>"110011100",
  33751=>"010111111",
  33752=>"000000011",
  33753=>"000010010",
  33754=>"001000100",
  33755=>"000001011",
  33756=>"100010011",
  33757=>"011110101",
  33758=>"000110111",
  33759=>"000101001",
  33760=>"010110111",
  33761=>"100010000",
  33762=>"101110010",
  33763=>"111110110",
  33764=>"010001010",
  33765=>"000011010",
  33766=>"110001101",
  33767=>"001110000",
  33768=>"101001111",
  33769=>"101001001",
  33770=>"001110010",
  33771=>"110111111",
  33772=>"111101001",
  33773=>"111110101",
  33774=>"111000001",
  33775=>"010010110",
  33776=>"010111100",
  33777=>"110111011",
  33778=>"001101000",
  33779=>"011101110",
  33780=>"110110001",
  33781=>"101111110",
  33782=>"011111111",
  33783=>"111100001",
  33784=>"100111010",
  33785=>"001111011",
  33786=>"101100011",
  33787=>"101111101",
  33788=>"000100011",
  33789=>"101110010",
  33790=>"011011101",
  33791=>"001100111",
  33792=>"000000110",
  33793=>"101111101",
  33794=>"010000100",
  33795=>"100000101",
  33796=>"000011011",
  33797=>"101011111",
  33798=>"011101110",
  33799=>"001111111",
  33800=>"010110001",
  33801=>"010111110",
  33802=>"001110011",
  33803=>"001101101",
  33804=>"111011101",
  33805=>"000000000",
  33806=>"111010001",
  33807=>"111000110",
  33808=>"001011100",
  33809=>"111100111",
  33810=>"101101010",
  33811=>"101000110",
  33812=>"101001100",
  33813=>"100100110",
  33814=>"000000001",
  33815=>"101001100",
  33816=>"110110110",
  33817=>"010110100",
  33818=>"110101111",
  33819=>"011101101",
  33820=>"000001011",
  33821=>"010111011",
  33822=>"101111101",
  33823=>"000010110",
  33824=>"000011101",
  33825=>"001100100",
  33826=>"011000011",
  33827=>"001110001",
  33828=>"011100100",
  33829=>"001010011",
  33830=>"000011110",
  33831=>"101111000",
  33832=>"001101010",
  33833=>"110011100",
  33834=>"000110001",
  33835=>"110001110",
  33836=>"101101001",
  33837=>"011111101",
  33838=>"000001010",
  33839=>"001000000",
  33840=>"101100000",
  33841=>"011100000",
  33842=>"000001011",
  33843=>"111100001",
  33844=>"101011111",
  33845=>"110010101",
  33846=>"000011010",
  33847=>"001010001",
  33848=>"111101010",
  33849=>"100010001",
  33850=>"001101011",
  33851=>"111111010",
  33852=>"110101010",
  33853=>"001011000",
  33854=>"110110001",
  33855=>"111110011",
  33856=>"101011100",
  33857=>"101100010",
  33858=>"000111011",
  33859=>"010001010",
  33860=>"100010110",
  33861=>"010100010",
  33862=>"100110001",
  33863=>"000101101",
  33864=>"001001001",
  33865=>"101111011",
  33866=>"001100011",
  33867=>"011101000",
  33868=>"010000000",
  33869=>"001000000",
  33870=>"000110000",
  33871=>"001001101",
  33872=>"001011010",
  33873=>"010000000",
  33874=>"110010011",
  33875=>"100000011",
  33876=>"010000111",
  33877=>"111010110",
  33878=>"111001000",
  33879=>"111010101",
  33880=>"011110001",
  33881=>"111111001",
  33882=>"011100011",
  33883=>"011111011",
  33884=>"111111010",
  33885=>"101110000",
  33886=>"000000000",
  33887=>"011110110",
  33888=>"001000111",
  33889=>"001111000",
  33890=>"000010010",
  33891=>"001001001",
  33892=>"001100101",
  33893=>"011000101",
  33894=>"000111111",
  33895=>"010000001",
  33896=>"000000000",
  33897=>"111000111",
  33898=>"001111111",
  33899=>"001011110",
  33900=>"100110001",
  33901=>"111001100",
  33902=>"000000110",
  33903=>"100000100",
  33904=>"000100010",
  33905=>"011011100",
  33906=>"011010000",
  33907=>"000010110",
  33908=>"011100000",
  33909=>"100000001",
  33910=>"010101011",
  33911=>"110110100",
  33912=>"101001100",
  33913=>"111100100",
  33914=>"000011010",
  33915=>"101101100",
  33916=>"111110001",
  33917=>"011100000",
  33918=>"101001110",
  33919=>"110000111",
  33920=>"001111010",
  33921=>"111110010",
  33922=>"010011111",
  33923=>"101010011",
  33924=>"110110011",
  33925=>"101100111",
  33926=>"001110101",
  33927=>"000010111",
  33928=>"000111100",
  33929=>"101111100",
  33930=>"111101101",
  33931=>"000101000",
  33932=>"111111011",
  33933=>"001100011",
  33934=>"010110001",
  33935=>"110000101",
  33936=>"111010001",
  33937=>"111110110",
  33938=>"001010111",
  33939=>"110101111",
  33940=>"101000110",
  33941=>"010100110",
  33942=>"000101010",
  33943=>"000101111",
  33944=>"000110111",
  33945=>"000001101",
  33946=>"000001011",
  33947=>"000011001",
  33948=>"111111101",
  33949=>"110110001",
  33950=>"001110011",
  33951=>"011001111",
  33952=>"011001010",
  33953=>"000001100",
  33954=>"110011000",
  33955=>"110011011",
  33956=>"111100000",
  33957=>"111010110",
  33958=>"110111111",
  33959=>"111111001",
  33960=>"010100111",
  33961=>"101111100",
  33962=>"100000111",
  33963=>"000011010",
  33964=>"001001100",
  33965=>"011111110",
  33966=>"011110000",
  33967=>"100011101",
  33968=>"011101000",
  33969=>"010101011",
  33970=>"101100001",
  33971=>"110001010",
  33972=>"100010000",
  33973=>"110110010",
  33974=>"010000010",
  33975=>"111011101",
  33976=>"000000101",
  33977=>"110011110",
  33978=>"001101101",
  33979=>"101111000",
  33980=>"010110101",
  33981=>"111101111",
  33982=>"110001000",
  33983=>"000001110",
  33984=>"111011000",
  33985=>"100111101",
  33986=>"000000010",
  33987=>"000000011",
  33988=>"000001000",
  33989=>"111110111",
  33990=>"000111011",
  33991=>"101100101",
  33992=>"111011001",
  33993=>"101000101",
  33994=>"100111001",
  33995=>"101110110",
  33996=>"010101110",
  33997=>"100000100",
  33998=>"000010011",
  33999=>"100110010",
  34000=>"101000011",
  34001=>"111100101",
  34002=>"001110111",
  34003=>"001000110",
  34004=>"010100000",
  34005=>"010010111",
  34006=>"100101010",
  34007=>"000110000",
  34008=>"010000000",
  34009=>"000101011",
  34010=>"001010100",
  34011=>"000010010",
  34012=>"010110011",
  34013=>"101111010",
  34014=>"011010101",
  34015=>"001111110",
  34016=>"010111000",
  34017=>"101011100",
  34018=>"101100001",
  34019=>"101000001",
  34020=>"011110010",
  34021=>"010101010",
  34022=>"000011110",
  34023=>"011010001",
  34024=>"011110001",
  34025=>"101011100",
  34026=>"110100000",
  34027=>"110100110",
  34028=>"111110010",
  34029=>"000111011",
  34030=>"000001101",
  34031=>"010100000",
  34032=>"010000110",
  34033=>"000011111",
  34034=>"111001111",
  34035=>"001110101",
  34036=>"110001010",
  34037=>"110111100",
  34038=>"001100011",
  34039=>"100001001",
  34040=>"010011110",
  34041=>"101111101",
  34042=>"101111110",
  34043=>"011011100",
  34044=>"010100000",
  34045=>"110111001",
  34046=>"011000001",
  34047=>"110000010",
  34048=>"111110001",
  34049=>"111001111",
  34050=>"111101111",
  34051=>"110000100",
  34052=>"011000000",
  34053=>"101001011",
  34054=>"011011111",
  34055=>"101110010",
  34056=>"111010110",
  34057=>"001000101",
  34058=>"000111110",
  34059=>"000110011",
  34060=>"111101110",
  34061=>"111011111",
  34062=>"011111101",
  34063=>"111111011",
  34064=>"101010101",
  34065=>"111101011",
  34066=>"010110101",
  34067=>"000010110",
  34068=>"110000110",
  34069=>"101101100",
  34070=>"110110010",
  34071=>"100100011",
  34072=>"001001001",
  34073=>"011011010",
  34074=>"110001111",
  34075=>"110011101",
  34076=>"010011001",
  34077=>"100001010",
  34078=>"001110010",
  34079=>"101110110",
  34080=>"111010111",
  34081=>"100111010",
  34082=>"110010011",
  34083=>"001101010",
  34084=>"100111010",
  34085=>"100011001",
  34086=>"110101001",
  34087=>"010111101",
  34088=>"101111111",
  34089=>"111000111",
  34090=>"011011100",
  34091=>"100110010",
  34092=>"110001111",
  34093=>"101010010",
  34094=>"111111100",
  34095=>"001000000",
  34096=>"111011110",
  34097=>"000001101",
  34098=>"111110100",
  34099=>"100010001",
  34100=>"101001010",
  34101=>"111101101",
  34102=>"111011111",
  34103=>"111110101",
  34104=>"000011111",
  34105=>"100001001",
  34106=>"111111101",
  34107=>"111100101",
  34108=>"100111101",
  34109=>"100001000",
  34110=>"101010100",
  34111=>"011100011",
  34112=>"111110100",
  34113=>"101110011",
  34114=>"010111110",
  34115=>"100101111",
  34116=>"100011100",
  34117=>"100110110",
  34118=>"110001011",
  34119=>"010001000",
  34120=>"101000110",
  34121=>"011000000",
  34122=>"110011100",
  34123=>"000000001",
  34124=>"000101110",
  34125=>"101010000",
  34126=>"011100110",
  34127=>"011000111",
  34128=>"000100110",
  34129=>"001111001",
  34130=>"000111100",
  34131=>"111000110",
  34132=>"011100011",
  34133=>"110000010",
  34134=>"011000100",
  34135=>"100111100",
  34136=>"111101110",
  34137=>"101011100",
  34138=>"110110011",
  34139=>"000010101",
  34140=>"110111110",
  34141=>"001000100",
  34142=>"101100101",
  34143=>"001011000",
  34144=>"001000010",
  34145=>"000001011",
  34146=>"010000100",
  34147=>"111110101",
  34148=>"001111101",
  34149=>"011011011",
  34150=>"011101000",
  34151=>"101111000",
  34152=>"111111001",
  34153=>"101110111",
  34154=>"011010111",
  34155=>"110010110",
  34156=>"100011101",
  34157=>"010110101",
  34158=>"101110011",
  34159=>"101111011",
  34160=>"111010100",
  34161=>"100101000",
  34162=>"000110110",
  34163=>"001111100",
  34164=>"011110000",
  34165=>"100011011",
  34166=>"100100100",
  34167=>"010100111",
  34168=>"000110001",
  34169=>"101011000",
  34170=>"100100001",
  34171=>"111011011",
  34172=>"111100000",
  34173=>"110101000",
  34174=>"100010101",
  34175=>"110011000",
  34176=>"110110000",
  34177=>"100000100",
  34178=>"100110001",
  34179=>"111110011",
  34180=>"011110010",
  34181=>"010001101",
  34182=>"101000000",
  34183=>"001100000",
  34184=>"000111000",
  34185=>"001110100",
  34186=>"111001001",
  34187=>"110111000",
  34188=>"010101011",
  34189=>"011011011",
  34190=>"110011110",
  34191=>"010010101",
  34192=>"000110101",
  34193=>"101010111",
  34194=>"000111001",
  34195=>"011000100",
  34196=>"100110011",
  34197=>"001010100",
  34198=>"010000110",
  34199=>"011000100",
  34200=>"101110101",
  34201=>"011000001",
  34202=>"011100101",
  34203=>"101110011",
  34204=>"110011101",
  34205=>"111011111",
  34206=>"000110100",
  34207=>"100100010",
  34208=>"110111010",
  34209=>"110011100",
  34210=>"001001100",
  34211=>"100101100",
  34212=>"100011010",
  34213=>"001110000",
  34214=>"011110100",
  34215=>"001101100",
  34216=>"000101110",
  34217=>"100000001",
  34218=>"010011111",
  34219=>"001110100",
  34220=>"000111000",
  34221=>"100001101",
  34222=>"101011011",
  34223=>"101111011",
  34224=>"111000010",
  34225=>"000110110",
  34226=>"111000100",
  34227=>"111001011",
  34228=>"111001011",
  34229=>"100100101",
  34230=>"100101110",
  34231=>"101111011",
  34232=>"010111000",
  34233=>"110110110",
  34234=>"000100111",
  34235=>"011100011",
  34236=>"000000110",
  34237=>"101011011",
  34238=>"000000100",
  34239=>"000010011",
  34240=>"110111011",
  34241=>"000111011",
  34242=>"111000000",
  34243=>"100011111",
  34244=>"001001000",
  34245=>"111111101",
  34246=>"011011111",
  34247=>"011011110",
  34248=>"100000110",
  34249=>"111011000",
  34250=>"100111000",
  34251=>"110001111",
  34252=>"101000100",
  34253=>"010000100",
  34254=>"010001010",
  34255=>"001110110",
  34256=>"111100000",
  34257=>"010000001",
  34258=>"010100110",
  34259=>"000001010",
  34260=>"100111000",
  34261=>"011001001",
  34262=>"101101101",
  34263=>"111000101",
  34264=>"110000000",
  34265=>"011101111",
  34266=>"110101010",
  34267=>"111101110",
  34268=>"011110010",
  34269=>"100100110",
  34270=>"100011010",
  34271=>"100010100",
  34272=>"101000110",
  34273=>"111111111",
  34274=>"110111010",
  34275=>"100101000",
  34276=>"110101111",
  34277=>"111000101",
  34278=>"101110010",
  34279=>"000010000",
  34280=>"100010001",
  34281=>"111100100",
  34282=>"011011100",
  34283=>"111010011",
  34284=>"101010100",
  34285=>"010000110",
  34286=>"111011010",
  34287=>"001101000",
  34288=>"011011111",
  34289=>"110100001",
  34290=>"011010100",
  34291=>"011100001",
  34292=>"101100101",
  34293=>"110111010",
  34294=>"100010111",
  34295=>"000001111",
  34296=>"011111101",
  34297=>"010001101",
  34298=>"001111111",
  34299=>"001010001",
  34300=>"110001110",
  34301=>"101101011",
  34302=>"110111000",
  34303=>"000010000",
  34304=>"101110000",
  34305=>"000101111",
  34306=>"101111101",
  34307=>"010100111",
  34308=>"100011011",
  34309=>"010100110",
  34310=>"110001111",
  34311=>"101100100",
  34312=>"011001000",
  34313=>"110100110",
  34314=>"110111001",
  34315=>"101110110",
  34316=>"100100111",
  34317=>"111110001",
  34318=>"101100110",
  34319=>"011100110",
  34320=>"111001100",
  34321=>"000101111",
  34322=>"011010101",
  34323=>"100110101",
  34324=>"100001101",
  34325=>"011000100",
  34326=>"000110010",
  34327=>"010001010",
  34328=>"000110010",
  34329=>"010000110",
  34330=>"110111011",
  34331=>"100101000",
  34332=>"000000110",
  34333=>"000010001",
  34334=>"001100001",
  34335=>"100010110",
  34336=>"100010001",
  34337=>"001010011",
  34338=>"010000000",
  34339=>"100011011",
  34340=>"001110101",
  34341=>"000011110",
  34342=>"001011101",
  34343=>"000001100",
  34344=>"100001111",
  34345=>"101111001",
  34346=>"011100011",
  34347=>"100110000",
  34348=>"000111100",
  34349=>"011011101",
  34350=>"010110111",
  34351=>"011011111",
  34352=>"001010110",
  34353=>"111011100",
  34354=>"001101011",
  34355=>"010111011",
  34356=>"111110100",
  34357=>"011001010",
  34358=>"100011011",
  34359=>"001010111",
  34360=>"110011100",
  34361=>"101010001",
  34362=>"110111011",
  34363=>"000000011",
  34364=>"010111011",
  34365=>"011010101",
  34366=>"001110011",
  34367=>"001010001",
  34368=>"101011110",
  34369=>"111110111",
  34370=>"001100111",
  34371=>"111010011",
  34372=>"100010111",
  34373=>"101101100",
  34374=>"111011010",
  34375=>"010111111",
  34376=>"010010001",
  34377=>"011000011",
  34378=>"001111110",
  34379=>"000111101",
  34380=>"001101110",
  34381=>"110100011",
  34382=>"100011110",
  34383=>"000111101",
  34384=>"011011011",
  34385=>"000001100",
  34386=>"001110001",
  34387=>"111111010",
  34388=>"000100010",
  34389=>"011100001",
  34390=>"000111101",
  34391=>"111111010",
  34392=>"000111110",
  34393=>"110101111",
  34394=>"101111011",
  34395=>"010000011",
  34396=>"100110100",
  34397=>"111101011",
  34398=>"100001111",
  34399=>"001101101",
  34400=>"000000101",
  34401=>"111101101",
  34402=>"100100011",
  34403=>"011111000",
  34404=>"010001101",
  34405=>"000010011",
  34406=>"110010011",
  34407=>"011101110",
  34408=>"100001101",
  34409=>"001101011",
  34410=>"010001011",
  34411=>"010000100",
  34412=>"001100101",
  34413=>"000110110",
  34414=>"101000100",
  34415=>"101010010",
  34416=>"001100111",
  34417=>"111010100",
  34418=>"011110100",
  34419=>"001011110",
  34420=>"110110111",
  34421=>"001111101",
  34422=>"011000000",
  34423=>"011110011",
  34424=>"100010011",
  34425=>"010011111",
  34426=>"000000111",
  34427=>"011011101",
  34428=>"011000001",
  34429=>"111101100",
  34430=>"001011110",
  34431=>"101010110",
  34432=>"100100011",
  34433=>"011110110",
  34434=>"100001000",
  34435=>"000011001",
  34436=>"000110110",
  34437=>"000001101",
  34438=>"100000110",
  34439=>"011111101",
  34440=>"110011000",
  34441=>"111011100",
  34442=>"011010001",
  34443=>"000110001",
  34444=>"000010111",
  34445=>"101100110",
  34446=>"110110110",
  34447=>"110110100",
  34448=>"111111101",
  34449=>"110111001",
  34450=>"000110010",
  34451=>"010100001",
  34452=>"010111101",
  34453=>"111100000",
  34454=>"001110000",
  34455=>"010001010",
  34456=>"010101000",
  34457=>"101101001",
  34458=>"100000000",
  34459=>"011110001",
  34460=>"011001100",
  34461=>"111111010",
  34462=>"110101010",
  34463=>"111001100",
  34464=>"100001100",
  34465=>"101000001",
  34466=>"011100111",
  34467=>"001000011",
  34468=>"111101000",
  34469=>"011110010",
  34470=>"101000001",
  34471=>"011101000",
  34472=>"110011101",
  34473=>"100000100",
  34474=>"101010000",
  34475=>"101110110",
  34476=>"110010010",
  34477=>"000101110",
  34478=>"111010010",
  34479=>"110100011",
  34480=>"010011110",
  34481=>"001001000",
  34482=>"001110000",
  34483=>"011110000",
  34484=>"000000111",
  34485=>"001110010",
  34486=>"111001001",
  34487=>"011111110",
  34488=>"010111110",
  34489=>"001011000",
  34490=>"001110101",
  34491=>"100101001",
  34492=>"100000010",
  34493=>"100001110",
  34494=>"111001100",
  34495=>"000010111",
  34496=>"111111000",
  34497=>"110111100",
  34498=>"000010100",
  34499=>"000110110",
  34500=>"110100001",
  34501=>"010010110",
  34502=>"111011001",
  34503=>"000111110",
  34504=>"111110100",
  34505=>"111100000",
  34506=>"011101110",
  34507=>"100101011",
  34508=>"100101100",
  34509=>"000000100",
  34510=>"011110110",
  34511=>"101110110",
  34512=>"110101110",
  34513=>"100010111",
  34514=>"100000110",
  34515=>"110101011",
  34516=>"100100000",
  34517=>"000000100",
  34518=>"100011010",
  34519=>"001010011",
  34520=>"100111011",
  34521=>"000100101",
  34522=>"000111000",
  34523=>"100011010",
  34524=>"010000111",
  34525=>"110001001",
  34526=>"000110010",
  34527=>"111011011",
  34528=>"101110101",
  34529=>"111010010",
  34530=>"100001101",
  34531=>"010000100",
  34532=>"011010010",
  34533=>"011110010",
  34534=>"010010000",
  34535=>"000000010",
  34536=>"010001010",
  34537=>"010011101",
  34538=>"111011100",
  34539=>"110100000",
  34540=>"000111111",
  34541=>"011101100",
  34542=>"100011010",
  34543=>"111101000",
  34544=>"001100100",
  34545=>"001010010",
  34546=>"000011111",
  34547=>"111101110",
  34548=>"010110110",
  34549=>"000010001",
  34550=>"000010110",
  34551=>"111110101",
  34552=>"101100110",
  34553=>"110100001",
  34554=>"101011101",
  34555=>"111100000",
  34556=>"111111011",
  34557=>"111000111",
  34558=>"111011000",
  34559=>"010110010",
  34560=>"111001001",
  34561=>"000100111",
  34562=>"001001011",
  34563=>"100010000",
  34564=>"001101000",
  34565=>"010010000",
  34566=>"110010110",
  34567=>"100000100",
  34568=>"000010010",
  34569=>"100111001",
  34570=>"000010111",
  34571=>"001010001",
  34572=>"101011111",
  34573=>"010000110",
  34574=>"000011111",
  34575=>"101100110",
  34576=>"111111101",
  34577=>"001110001",
  34578=>"100100001",
  34579=>"110111100",
  34580=>"001011000",
  34581=>"001100110",
  34582=>"000000010",
  34583=>"110101000",
  34584=>"000011101",
  34585=>"001000100",
  34586=>"010001000",
  34587=>"011010001",
  34588=>"001100101",
  34589=>"000101100",
  34590=>"110110011",
  34591=>"001001101",
  34592=>"100000110",
  34593=>"011111000",
  34594=>"010000001",
  34595=>"000000111",
  34596=>"100000100",
  34597=>"010111101",
  34598=>"010111001",
  34599=>"010100011",
  34600=>"111000010",
  34601=>"001101001",
  34602=>"001010011",
  34603=>"001111101",
  34604=>"000101100",
  34605=>"001101001",
  34606=>"101101001",
  34607=>"001100101",
  34608=>"111110000",
  34609=>"111011100",
  34610=>"111010010",
  34611=>"010101000",
  34612=>"101010100",
  34613=>"010100010",
  34614=>"010011000",
  34615=>"010011011",
  34616=>"111001101",
  34617=>"111010011",
  34618=>"110110001",
  34619=>"110111111",
  34620=>"011001010",
  34621=>"111111111",
  34622=>"110010101",
  34623=>"011000001",
  34624=>"110100110",
  34625=>"011001011",
  34626=>"010000010",
  34627=>"110011010",
  34628=>"100100101",
  34629=>"111000001",
  34630=>"010010001",
  34631=>"000111110",
  34632=>"101110010",
  34633=>"111001000",
  34634=>"010011100",
  34635=>"101100100",
  34636=>"101001001",
  34637=>"110101001",
  34638=>"000100101",
  34639=>"011010010",
  34640=>"001010010",
  34641=>"111001000",
  34642=>"111010000",
  34643=>"100100110",
  34644=>"111000101",
  34645=>"101001111",
  34646=>"101110001",
  34647=>"111110101",
  34648=>"001010100",
  34649=>"100010011",
  34650=>"001011111",
  34651=>"111110010",
  34652=>"110000000",
  34653=>"110000011",
  34654=>"000101110",
  34655=>"100100001",
  34656=>"110000000",
  34657=>"010011101",
  34658=>"010111111",
  34659=>"010110110",
  34660=>"011100101",
  34661=>"011111001",
  34662=>"001100011",
  34663=>"011101011",
  34664=>"011100000",
  34665=>"000101001",
  34666=>"111111001",
  34667=>"100110001",
  34668=>"101100100",
  34669=>"011000110",
  34670=>"000111000",
  34671=>"100110011",
  34672=>"001111011",
  34673=>"111101001",
  34674=>"011110100",
  34675=>"111110010",
  34676=>"000011110",
  34677=>"100001000",
  34678=>"111010100",
  34679=>"011011010",
  34680=>"010000010",
  34681=>"010100110",
  34682=>"110011110",
  34683=>"000101000",
  34684=>"001011010",
  34685=>"010111111",
  34686=>"000110101",
  34687=>"110111001",
  34688=>"011100111",
  34689=>"000110010",
  34690=>"111000111",
  34691=>"100101000",
  34692=>"011100011",
  34693=>"010011001",
  34694=>"011011000",
  34695=>"001010110",
  34696=>"010100001",
  34697=>"001111110",
  34698=>"011100001",
  34699=>"101101000",
  34700=>"000110110",
  34701=>"101011100",
  34702=>"011001100",
  34703=>"000111111",
  34704=>"000000111",
  34705=>"000110111",
  34706=>"111000110",
  34707=>"101010011",
  34708=>"010001100",
  34709=>"010101010",
  34710=>"111010111",
  34711=>"011001011",
  34712=>"010111010",
  34713=>"001010010",
  34714=>"010101100",
  34715=>"100010000",
  34716=>"011011001",
  34717=>"001101100",
  34718=>"011100011",
  34719=>"011010000",
  34720=>"000100111",
  34721=>"001010001",
  34722=>"011111000",
  34723=>"000001100",
  34724=>"011010000",
  34725=>"001000000",
  34726=>"000111010",
  34727=>"101101111",
  34728=>"111000000",
  34729=>"011100000",
  34730=>"111010111",
  34731=>"000101111",
  34732=>"110000001",
  34733=>"000101100",
  34734=>"110011011",
  34735=>"000010100",
  34736=>"001111010",
  34737=>"101000010",
  34738=>"011100100",
  34739=>"110011010",
  34740=>"011010111",
  34741=>"000000000",
  34742=>"000101101",
  34743=>"000110010",
  34744=>"111000100",
  34745=>"111001011",
  34746=>"010101010",
  34747=>"100110000",
  34748=>"100000011",
  34749=>"110000100",
  34750=>"001101011",
  34751=>"001000101",
  34752=>"000100110",
  34753=>"101010110",
  34754=>"111110000",
  34755=>"111100011",
  34756=>"010111110",
  34757=>"010101111",
  34758=>"101111111",
  34759=>"110011010",
  34760=>"111100010",
  34761=>"000110111",
  34762=>"110001001",
  34763=>"010000001",
  34764=>"000101001",
  34765=>"101011001",
  34766=>"010111001",
  34767=>"101010100",
  34768=>"111001011",
  34769=>"000001001",
  34770=>"011001100",
  34771=>"000101000",
  34772=>"001111000",
  34773=>"011110011",
  34774=>"110011101",
  34775=>"010101100",
  34776=>"100100111",
  34777=>"101000100",
  34778=>"011000001",
  34779=>"111000100",
  34780=>"010110001",
  34781=>"110101010",
  34782=>"011111101",
  34783=>"111111010",
  34784=>"100110111",
  34785=>"100000111",
  34786=>"101111011",
  34787=>"011011101",
  34788=>"110100100",
  34789=>"111111111",
  34790=>"111011100",
  34791=>"010010000",
  34792=>"110010010",
  34793=>"011101011",
  34794=>"111011111",
  34795=>"100111110",
  34796=>"010011110",
  34797=>"100001100",
  34798=>"111011101",
  34799=>"001100100",
  34800=>"000010100",
  34801=>"111110100",
  34802=>"110111001",
  34803=>"001000000",
  34804=>"110010011",
  34805=>"101110000",
  34806=>"111011000",
  34807=>"010100110",
  34808=>"011101001",
  34809=>"000011100",
  34810=>"011000111",
  34811=>"011010111",
  34812=>"100000000",
  34813=>"001100010",
  34814=>"110100011",
  34815=>"111110110",
  34816=>"100000101",
  34817=>"010000111",
  34818=>"111110001",
  34819=>"110011001",
  34820=>"011110001",
  34821=>"110111000",
  34822=>"011000000",
  34823=>"000100101",
  34824=>"110110001",
  34825=>"111101001",
  34826=>"011010111",
  34827=>"101101110",
  34828=>"011110100",
  34829=>"010001111",
  34830=>"010100010",
  34831=>"110010111",
  34832=>"100010110",
  34833=>"010011001",
  34834=>"111111010",
  34835=>"010000000",
  34836=>"101100101",
  34837=>"010001100",
  34838=>"110111111",
  34839=>"000010001",
  34840=>"100011100",
  34841=>"101110001",
  34842=>"101011101",
  34843=>"101110100",
  34844=>"110000101",
  34845=>"100110000",
  34846=>"110010000",
  34847=>"110101011",
  34848=>"001010011",
  34849=>"110101111",
  34850=>"000011011",
  34851=>"010101100",
  34852=>"001111011",
  34853=>"001101011",
  34854=>"100100000",
  34855=>"011111111",
  34856=>"011010110",
  34857=>"110110000",
  34858=>"011101011",
  34859=>"100010010",
  34860=>"110010001",
  34861=>"111000110",
  34862=>"100001111",
  34863=>"001111100",
  34864=>"111101011",
  34865=>"111001010",
  34866=>"001110000",
  34867=>"010001000",
  34868=>"110000001",
  34869=>"011111010",
  34870=>"000100110",
  34871=>"111011111",
  34872=>"101100011",
  34873=>"011000101",
  34874=>"111001000",
  34875=>"101000110",
  34876=>"011011110",
  34877=>"100000101",
  34878=>"000101101",
  34879=>"011101110",
  34880=>"101101011",
  34881=>"000111001",
  34882=>"001011110",
  34883=>"001100010",
  34884=>"011100000",
  34885=>"000011010",
  34886=>"111010000",
  34887=>"110100010",
  34888=>"100101101",
  34889=>"001100000",
  34890=>"111101001",
  34891=>"011110010",
  34892=>"000111001",
  34893=>"100100111",
  34894=>"110100111",
  34895=>"010111010",
  34896=>"110100000",
  34897=>"010000010",
  34898=>"000000110",
  34899=>"011011001",
  34900=>"110011100",
  34901=>"011101010",
  34902=>"000000001",
  34903=>"011111111",
  34904=>"101100111",
  34905=>"110100010",
  34906=>"011100101",
  34907=>"010000000",
  34908=>"010110110",
  34909=>"110011110",
  34910=>"011010111",
  34911=>"100000000",
  34912=>"000101101",
  34913=>"100000010",
  34914=>"100001101",
  34915=>"110000010",
  34916=>"001101111",
  34917=>"100101110",
  34918=>"000010001",
  34919=>"000111011",
  34920=>"110011011",
  34921=>"100111011",
  34922=>"111101101",
  34923=>"000100111",
  34924=>"000001100",
  34925=>"011111000",
  34926=>"010001001",
  34927=>"000101010",
  34928=>"111001010",
  34929=>"001011111",
  34930=>"100001100",
  34931=>"011100011",
  34932=>"011111001",
  34933=>"111001110",
  34934=>"100100000",
  34935=>"010011110",
  34936=>"111000010",
  34937=>"001000111",
  34938=>"101011100",
  34939=>"111111100",
  34940=>"001001101",
  34941=>"101100111",
  34942=>"001011000",
  34943=>"001001011",
  34944=>"110111001",
  34945=>"001001001",
  34946=>"000101000",
  34947=>"011010101",
  34948=>"111100011",
  34949=>"111000111",
  34950=>"011001110",
  34951=>"011110100",
  34952=>"111100101",
  34953=>"110101100",
  34954=>"001001000",
  34955=>"011110000",
  34956=>"111011010",
  34957=>"001000010",
  34958=>"110010101",
  34959=>"110011011",
  34960=>"101011100",
  34961=>"101001001",
  34962=>"110011000",
  34963=>"010001101",
  34964=>"100000100",
  34965=>"011011001",
  34966=>"001010000",
  34967=>"101001001",
  34968=>"000010011",
  34969=>"010001110",
  34970=>"011110000",
  34971=>"100100111",
  34972=>"011101001",
  34973=>"100000010",
  34974=>"011001100",
  34975=>"111111011",
  34976=>"110110110",
  34977=>"100011010",
  34978=>"110111101",
  34979=>"000100100",
  34980=>"010010101",
  34981=>"001110010",
  34982=>"101000100",
  34983=>"101001000",
  34984=>"000100000",
  34985=>"101000100",
  34986=>"111011111",
  34987=>"010000101",
  34988=>"011111101",
  34989=>"111011010",
  34990=>"010010000",
  34991=>"100111101",
  34992=>"001100010",
  34993=>"010110011",
  34994=>"001001111",
  34995=>"011110100",
  34996=>"000101101",
  34997=>"101101111",
  34998=>"000110011",
  34999=>"100000001",
  35000=>"011010010",
  35001=>"000001000",
  35002=>"110000111",
  35003=>"001111100",
  35004=>"110000001",
  35005=>"011011000",
  35006=>"100000000",
  35007=>"001111101",
  35008=>"000110101",
  35009=>"110100101",
  35010=>"110110100",
  35011=>"000101100",
  35012=>"000111100",
  35013=>"000110111",
  35014=>"010010011",
  35015=>"111111011",
  35016=>"000101000",
  35017=>"001101011",
  35018=>"000100101",
  35019=>"110011101",
  35020=>"000100001",
  35021=>"001110001",
  35022=>"001110001",
  35023=>"111111110",
  35024=>"011110111",
  35025=>"110110010",
  35026=>"110000010",
  35027=>"001001100",
  35028=>"011110100",
  35029=>"011000011",
  35030=>"010011000",
  35031=>"100001011",
  35032=>"111001010",
  35033=>"111010100",
  35034=>"000000100",
  35035=>"110101011",
  35036=>"010001111",
  35037=>"001010100",
  35038=>"000110000",
  35039=>"010001100",
  35040=>"111000001",
  35041=>"010100101",
  35042=>"101011001",
  35043=>"001001001",
  35044=>"000011100",
  35045=>"011101011",
  35046=>"011110101",
  35047=>"001010000",
  35048=>"010011100",
  35049=>"001010100",
  35050=>"011110100",
  35051=>"010010110",
  35052=>"011100001",
  35053=>"101001101",
  35054=>"001000100",
  35055=>"010101010",
  35056=>"100111000",
  35057=>"111111111",
  35058=>"100010000",
  35059=>"110100000",
  35060=>"001101010",
  35061=>"101100001",
  35062=>"101101010",
  35063=>"100000100",
  35064=>"000110111",
  35065=>"011000100",
  35066=>"100101100",
  35067=>"100000000",
  35068=>"111001100",
  35069=>"100010100",
  35070=>"011111100",
  35071=>"000011011",
  35072=>"101001001",
  35073=>"111101110",
  35074=>"001100011",
  35075=>"111110100",
  35076=>"101111011",
  35077=>"100111000",
  35078=>"100100001",
  35079=>"111010101",
  35080=>"000101010",
  35081=>"101000010",
  35082=>"011001000",
  35083=>"011000000",
  35084=>"000011010",
  35085=>"000101101",
  35086=>"000110010",
  35087=>"010100000",
  35088=>"111011011",
  35089=>"101000111",
  35090=>"100000000",
  35091=>"001100000",
  35092=>"001011000",
  35093=>"010010011",
  35094=>"001100110",
  35095=>"110110110",
  35096=>"101010011",
  35097=>"001011010",
  35098=>"001011110",
  35099=>"010001000",
  35100=>"001000111",
  35101=>"110100110",
  35102=>"110011100",
  35103=>"010001000",
  35104=>"111100111",
  35105=>"010101111",
  35106=>"010111101",
  35107=>"110101011",
  35108=>"111000111",
  35109=>"111011001",
  35110=>"001001000",
  35111=>"010000110",
  35112=>"011000100",
  35113=>"111000010",
  35114=>"100001001",
  35115=>"100110111",
  35116=>"100100100",
  35117=>"001101011",
  35118=>"101011101",
  35119=>"110101101",
  35120=>"110011000",
  35121=>"001011000",
  35122=>"001101010",
  35123=>"101101001",
  35124=>"110010100",
  35125=>"101101110",
  35126=>"011010111",
  35127=>"010011111",
  35128=>"111001010",
  35129=>"100000011",
  35130=>"100010101",
  35131=>"001100111",
  35132=>"001001110",
  35133=>"101110011",
  35134=>"101111011",
  35135=>"011000111",
  35136=>"111111001",
  35137=>"110111101",
  35138=>"101110011",
  35139=>"111100000",
  35140=>"110100011",
  35141=>"010010010",
  35142=>"100001010",
  35143=>"100101000",
  35144=>"011011001",
  35145=>"100011001",
  35146=>"001010100",
  35147=>"000011011",
  35148=>"001100000",
  35149=>"100101011",
  35150=>"111101010",
  35151=>"000101001",
  35152=>"100100011",
  35153=>"100000000",
  35154=>"111011101",
  35155=>"101110010",
  35156=>"110100000",
  35157=>"101001110",
  35158=>"111011101",
  35159=>"110011110",
  35160=>"000000010",
  35161=>"111000000",
  35162=>"000110000",
  35163=>"101000011",
  35164=>"101100100",
  35165=>"011111101",
  35166=>"000100111",
  35167=>"111111010",
  35168=>"101111111",
  35169=>"011000011",
  35170=>"101100111",
  35171=>"100101011",
  35172=>"001110000",
  35173=>"110000101",
  35174=>"101101011",
  35175=>"101100010",
  35176=>"001110001",
  35177=>"110010110",
  35178=>"100010010",
  35179=>"010100000",
  35180=>"000111101",
  35181=>"001110111",
  35182=>"010101110",
  35183=>"100000000",
  35184=>"000100101",
  35185=>"010010101",
  35186=>"101100100",
  35187=>"011000000",
  35188=>"010010000",
  35189=>"001011011",
  35190=>"010101100",
  35191=>"110001110",
  35192=>"001101011",
  35193=>"001110010",
  35194=>"111100011",
  35195=>"000101011",
  35196=>"001100011",
  35197=>"111000111",
  35198=>"100100011",
  35199=>"000000101",
  35200=>"111111011",
  35201=>"111110101",
  35202=>"000011010",
  35203=>"111111100",
  35204=>"110101111",
  35205=>"110001001",
  35206=>"010001001",
  35207=>"111001101",
  35208=>"111100100",
  35209=>"001100011",
  35210=>"001100111",
  35211=>"000101111",
  35212=>"111101000",
  35213=>"101000001",
  35214=>"110101100",
  35215=>"010110000",
  35216=>"010001000",
  35217=>"001110111",
  35218=>"100111001",
  35219=>"111110001",
  35220=>"001000000",
  35221=>"001000111",
  35222=>"000111001",
  35223=>"110100010",
  35224=>"110111111",
  35225=>"000001100",
  35226=>"011001011",
  35227=>"100010001",
  35228=>"111011100",
  35229=>"001010001",
  35230=>"000000100",
  35231=>"011101010",
  35232=>"000100110",
  35233=>"111000010",
  35234=>"110011101",
  35235=>"000010001",
  35236=>"110100011",
  35237=>"000011110",
  35238=>"110110110",
  35239=>"000101010",
  35240=>"101111101",
  35241=>"101110001",
  35242=>"001010011",
  35243=>"111101101",
  35244=>"001111010",
  35245=>"011000000",
  35246=>"110101110",
  35247=>"100000100",
  35248=>"101111111",
  35249=>"101011001",
  35250=>"011111110",
  35251=>"000111010",
  35252=>"010100010",
  35253=>"111000110",
  35254=>"111111001",
  35255=>"111111110",
  35256=>"011011110",
  35257=>"111000101",
  35258=>"100000000",
  35259=>"101001010",
  35260=>"100100100",
  35261=>"101010001",
  35262=>"000001001",
  35263=>"100000100",
  35264=>"111000011",
  35265=>"110100111",
  35266=>"011110111",
  35267=>"011110110",
  35268=>"110100010",
  35269=>"101000001",
  35270=>"011000101",
  35271=>"010010111",
  35272=>"010101000",
  35273=>"100011111",
  35274=>"000101101",
  35275=>"101010101",
  35276=>"111100101",
  35277=>"101100100",
  35278=>"111111001",
  35279=>"001110100",
  35280=>"101101010",
  35281=>"110101100",
  35282=>"101011010",
  35283=>"101001111",
  35284=>"101110111",
  35285=>"111000011",
  35286=>"110000100",
  35287=>"000011000",
  35288=>"100101110",
  35289=>"111001110",
  35290=>"000101010",
  35291=>"011001000",
  35292=>"101011111",
  35293=>"000001111",
  35294=>"010100011",
  35295=>"010110000",
  35296=>"010101011",
  35297=>"111000000",
  35298=>"111101111",
  35299=>"001011110",
  35300=>"000010101",
  35301=>"001110001",
  35302=>"000011111",
  35303=>"111111001",
  35304=>"010101110",
  35305=>"001110011",
  35306=>"011100000",
  35307=>"111110110",
  35308=>"010111000",
  35309=>"101000001",
  35310=>"100011001",
  35311=>"111010000",
  35312=>"110001111",
  35313=>"001000111",
  35314=>"010001010",
  35315=>"011110011",
  35316=>"011000100",
  35317=>"010000111",
  35318=>"000110000",
  35319=>"100000000",
  35320=>"010100111",
  35321=>"011111000",
  35322=>"011011100",
  35323=>"100111000",
  35324=>"101001100",
  35325=>"101011000",
  35326=>"111111001",
  35327=>"011000010",
  35328=>"101101100",
  35329=>"010100001",
  35330=>"001101111",
  35331=>"110011111",
  35332=>"100001000",
  35333=>"100110001",
  35334=>"110101000",
  35335=>"101100101",
  35336=>"111100110",
  35337=>"101100111",
  35338=>"011110101",
  35339=>"101110011",
  35340=>"000100010",
  35341=>"000100101",
  35342=>"010111100",
  35343=>"010100101",
  35344=>"000111110",
  35345=>"110110100",
  35346=>"001100111",
  35347=>"011110001",
  35348=>"101110001",
  35349=>"001100000",
  35350=>"100001111",
  35351=>"101111111",
  35352=>"100010010",
  35353=>"100110000",
  35354=>"111011010",
  35355=>"100101111",
  35356=>"011000101",
  35357=>"001111001",
  35358=>"100001110",
  35359=>"111001011",
  35360=>"001010100",
  35361=>"100011101",
  35362=>"001001011",
  35363=>"111101100",
  35364=>"111110010",
  35365=>"100111100",
  35366=>"011010100",
  35367=>"110000001",
  35368=>"001100000",
  35369=>"110101000",
  35370=>"101110011",
  35371=>"100001000",
  35372=>"000110111",
  35373=>"100010111",
  35374=>"011001010",
  35375=>"100011101",
  35376=>"100011000",
  35377=>"111101000",
  35378=>"000100100",
  35379=>"100010100",
  35380=>"010100110",
  35381=>"101100111",
  35382=>"010110110",
  35383=>"011000101",
  35384=>"001011010",
  35385=>"100111101",
  35386=>"010010101",
  35387=>"011111101",
  35388=>"110011001",
  35389=>"011101001",
  35390=>"001101101",
  35391=>"110010111",
  35392=>"000010000",
  35393=>"100110001",
  35394=>"001011100",
  35395=>"110100101",
  35396=>"101100011",
  35397=>"101011111",
  35398=>"101101011",
  35399=>"001001000",
  35400=>"011000100",
  35401=>"001000000",
  35402=>"100110011",
  35403=>"101100111",
  35404=>"000011010",
  35405=>"001110110",
  35406=>"011111111",
  35407=>"100011110",
  35408=>"110010110",
  35409=>"101100101",
  35410=>"100011100",
  35411=>"101010110",
  35412=>"111110011",
  35413=>"000011111",
  35414=>"000001001",
  35415=>"010111101",
  35416=>"100100010",
  35417=>"011101000",
  35418=>"010111010",
  35419=>"010000101",
  35420=>"010010010",
  35421=>"001000000",
  35422=>"000100011",
  35423=>"010101011",
  35424=>"011001000",
  35425=>"010000011",
  35426=>"011010100",
  35427=>"110000010",
  35428=>"111100111",
  35429=>"010101011",
  35430=>"100110000",
  35431=>"000010010",
  35432=>"011010000",
  35433=>"001110011",
  35434=>"011100000",
  35435=>"111110111",
  35436=>"000111110",
  35437=>"110001011",
  35438=>"000111001",
  35439=>"111110100",
  35440=>"110111110",
  35441=>"100000001",
  35442=>"111101001",
  35443=>"110000000",
  35444=>"010011110",
  35445=>"110001000",
  35446=>"100110111",
  35447=>"101001110",
  35448=>"001110111",
  35449=>"001110000",
  35450=>"010110101",
  35451=>"000100001",
  35452=>"011100000",
  35453=>"101101100",
  35454=>"011101110",
  35455=>"110100010",
  35456=>"001101010",
  35457=>"011101011",
  35458=>"101001001",
  35459=>"101101101",
  35460=>"011111001",
  35461=>"001000101",
  35462=>"011100000",
  35463=>"100111110",
  35464=>"111100000",
  35465=>"111011111",
  35466=>"001000000",
  35467=>"001110101",
  35468=>"111001001",
  35469=>"100001010",
  35470=>"101101000",
  35471=>"100110101",
  35472=>"001000101",
  35473=>"111101110",
  35474=>"001001101",
  35475=>"011111011",
  35476=>"000001001",
  35477=>"011110000",
  35478=>"100000011",
  35479=>"000001000",
  35480=>"010101111",
  35481=>"010110000",
  35482=>"101010101",
  35483=>"110101010",
  35484=>"001101001",
  35485=>"001110001",
  35486=>"110000100",
  35487=>"000011001",
  35488=>"101011011",
  35489=>"010111000",
  35490=>"000011000",
  35491=>"011100010",
  35492=>"011011011",
  35493=>"010101111",
  35494=>"101001010",
  35495=>"001000001",
  35496=>"111011001",
  35497=>"011110110",
  35498=>"001011010",
  35499=>"001010100",
  35500=>"000000001",
  35501=>"111111101",
  35502=>"000110010",
  35503=>"011011100",
  35504=>"000011001",
  35505=>"000101000",
  35506=>"000101000",
  35507=>"111000110",
  35508=>"001001000",
  35509=>"000111101",
  35510=>"111011111",
  35511=>"001011101",
  35512=>"011010111",
  35513=>"000001110",
  35514=>"010011110",
  35515=>"000010011",
  35516=>"010101000",
  35517=>"101011111",
  35518=>"000011010",
  35519=>"111101011",
  35520=>"010010000",
  35521=>"100111110",
  35522=>"000011011",
  35523=>"111111001",
  35524=>"100110111",
  35525=>"100100111",
  35526=>"111111111",
  35527=>"011010011",
  35528=>"010101010",
  35529=>"011011100",
  35530=>"011001110",
  35531=>"001100001",
  35532=>"011010011",
  35533=>"101011010",
  35534=>"111001010",
  35535=>"001000111",
  35536=>"001111000",
  35537=>"000100100",
  35538=>"110100111",
  35539=>"011011101",
  35540=>"010110000",
  35541=>"011000101",
  35542=>"111100011",
  35543=>"000010011",
  35544=>"000100100",
  35545=>"010010011",
  35546=>"000001011",
  35547=>"010101001",
  35548=>"011101110",
  35549=>"100110110",
  35550=>"111111101",
  35551=>"111101101",
  35552=>"000101110",
  35553=>"010111111",
  35554=>"000101111",
  35555=>"111011111",
  35556=>"000110100",
  35557=>"111010111",
  35558=>"001000001",
  35559=>"111000110",
  35560=>"000101001",
  35561=>"110001101",
  35562=>"000110010",
  35563=>"110111000",
  35564=>"010111000",
  35565=>"100101001",
  35566=>"110100000",
  35567=>"101001000",
  35568=>"000000100",
  35569=>"001110011",
  35570=>"011000110",
  35571=>"101101001",
  35572=>"101010111",
  35573=>"011101001",
  35574=>"101011110",
  35575=>"101011001",
  35576=>"000001001",
  35577=>"110100010",
  35578=>"010010100",
  35579=>"100010001",
  35580=>"100111100",
  35581=>"011010010",
  35582=>"111101001",
  35583=>"101101111",
  35584=>"111110000",
  35585=>"011000001",
  35586=>"010110111",
  35587=>"110000010",
  35588=>"100100001",
  35589=>"010010010",
  35590=>"101000110",
  35591=>"010011000",
  35592=>"111100000",
  35593=>"111100000",
  35594=>"101001111",
  35595=>"000101101",
  35596=>"100001101",
  35597=>"010110011",
  35598=>"010100111",
  35599=>"101000001",
  35600=>"001100111",
  35601=>"001101101",
  35602=>"000111101",
  35603=>"010110010",
  35604=>"100110101",
  35605=>"001101000",
  35606=>"101100110",
  35607=>"111000001",
  35608=>"000010111",
  35609=>"011011100",
  35610=>"010011011",
  35611=>"110000100",
  35612=>"101010110",
  35613=>"100110100",
  35614=>"000000111",
  35615=>"001000000",
  35616=>"100111110",
  35617=>"111011101",
  35618=>"101001010",
  35619=>"000110100",
  35620=>"000101111",
  35621=>"101111000",
  35622=>"000000001",
  35623=>"110000000",
  35624=>"101000010",
  35625=>"100000010",
  35626=>"000000000",
  35627=>"011100111",
  35628=>"111011010",
  35629=>"000100101",
  35630=>"000011010",
  35631=>"101011011",
  35632=>"110000001",
  35633=>"111000100",
  35634=>"111010001",
  35635=>"100111110",
  35636=>"001110111",
  35637=>"101001100",
  35638=>"000110100",
  35639=>"110110000",
  35640=>"001100000",
  35641=>"100100110",
  35642=>"010010000",
  35643=>"001100010",
  35644=>"000010011",
  35645=>"111111011",
  35646=>"111000110",
  35647=>"110000000",
  35648=>"110111011",
  35649=>"100010010",
  35650=>"010110011",
  35651=>"100001011",
  35652=>"000110000",
  35653=>"110101000",
  35654=>"000110010",
  35655=>"101101011",
  35656=>"011101101",
  35657=>"101000001",
  35658=>"001101010",
  35659=>"111001100",
  35660=>"000010000",
  35661=>"010010010",
  35662=>"011001110",
  35663=>"000100010",
  35664=>"011001000",
  35665=>"111101001",
  35666=>"011001011",
  35667=>"110010100",
  35668=>"001011001",
  35669=>"010101001",
  35670=>"010010010",
  35671=>"110011101",
  35672=>"010010010",
  35673=>"000100000",
  35674=>"100111010",
  35675=>"011100111",
  35676=>"011010111",
  35677=>"000001000",
  35678=>"000101001",
  35679=>"001000100",
  35680=>"000011100",
  35681=>"010010001",
  35682=>"101111101",
  35683=>"011001111",
  35684=>"101100101",
  35685=>"011101101",
  35686=>"111000011",
  35687=>"101010101",
  35688=>"001100001",
  35689=>"011111000",
  35690=>"001010100",
  35691=>"111111010",
  35692=>"100010101",
  35693=>"001101101",
  35694=>"100100010",
  35695=>"101111011",
  35696=>"010100100",
  35697=>"111001000",
  35698=>"101101000",
  35699=>"000111110",
  35700=>"100010000",
  35701=>"111011101",
  35702=>"100001010",
  35703=>"000010110",
  35704=>"111011010",
  35705=>"011000011",
  35706=>"111110101",
  35707=>"011111010",
  35708=>"010100000",
  35709=>"101000110",
  35710=>"010100100",
  35711=>"010010000",
  35712=>"011000010",
  35713=>"110111110",
  35714=>"101001010",
  35715=>"010101010",
  35716=>"011010010",
  35717=>"001101100",
  35718=>"100001010",
  35719=>"011100000",
  35720=>"001011100",
  35721=>"000110100",
  35722=>"110110110",
  35723=>"000010010",
  35724=>"011001000",
  35725=>"011110010",
  35726=>"011100001",
  35727=>"110110011",
  35728=>"011111000",
  35729=>"100111111",
  35730=>"000111000",
  35731=>"111011100",
  35732=>"110001001",
  35733=>"011010011",
  35734=>"000001011",
  35735=>"010001010",
  35736=>"110110110",
  35737=>"100000000",
  35738=>"111111101",
  35739=>"100101101",
  35740=>"011010101",
  35741=>"010110100",
  35742=>"100011011",
  35743=>"110010011",
  35744=>"000100011",
  35745=>"011011011",
  35746=>"100111110",
  35747=>"011000111",
  35748=>"100001001",
  35749=>"011110001",
  35750=>"101011001",
  35751=>"111001010",
  35752=>"101001001",
  35753=>"001001101",
  35754=>"001001100",
  35755=>"111111100",
  35756=>"000101111",
  35757=>"110101111",
  35758=>"001000010",
  35759=>"000010110",
  35760=>"111011101",
  35761=>"010111101",
  35762=>"001010111",
  35763=>"011000010",
  35764=>"111111011",
  35765=>"101100011",
  35766=>"000000011",
  35767=>"000001110",
  35768=>"110011000",
  35769=>"110000111",
  35770=>"010101010",
  35771=>"111011100",
  35772=>"011100111",
  35773=>"000100011",
  35774=>"111111110",
  35775=>"110100110",
  35776=>"011110000",
  35777=>"010010110",
  35778=>"001000000",
  35779=>"111010110",
  35780=>"101010111",
  35781=>"000000101",
  35782=>"010110110",
  35783=>"001101011",
  35784=>"110110100",
  35785=>"001001100",
  35786=>"101110111",
  35787=>"101000010",
  35788=>"111001100",
  35789=>"001111110",
  35790=>"110111111",
  35791=>"001000000",
  35792=>"111001001",
  35793=>"111110111",
  35794=>"101000110",
  35795=>"111010001",
  35796=>"000101010",
  35797=>"010000001",
  35798=>"001101001",
  35799=>"111110100",
  35800=>"100011001",
  35801=>"100010000",
  35802=>"111010001",
  35803=>"100011001",
  35804=>"101100011",
  35805=>"000010101",
  35806=>"110100001",
  35807=>"011100101",
  35808=>"001111011",
  35809=>"110111110",
  35810=>"011010011",
  35811=>"110110010",
  35812=>"100011000",
  35813=>"000000010",
  35814=>"000111110",
  35815=>"100010010",
  35816=>"100001110",
  35817=>"000111101",
  35818=>"111101011",
  35819=>"011101110",
  35820=>"100110001",
  35821=>"010001000",
  35822=>"101010111",
  35823=>"101111011",
  35824=>"011010001",
  35825=>"000001101",
  35826=>"000010110",
  35827=>"000100111",
  35828=>"100000110",
  35829=>"100011111",
  35830=>"001111110",
  35831=>"101100001",
  35832=>"010111110",
  35833=>"000001111",
  35834=>"000100101",
  35835=>"101011110",
  35836=>"001100100",
  35837=>"100011110",
  35838=>"000000110",
  35839=>"111110000",
  35840=>"111000100",
  35841=>"101010101",
  35842=>"101110110",
  35843=>"100111111",
  35844=>"100111101",
  35845=>"010011111",
  35846=>"010010110",
  35847=>"001111111",
  35848=>"000001111",
  35849=>"000111010",
  35850=>"000000110",
  35851=>"110001011",
  35852=>"100011000",
  35853=>"010110001",
  35854=>"101011001",
  35855=>"000100011",
  35856=>"100000001",
  35857=>"010000000",
  35858=>"110101100",
  35859=>"001001101",
  35860=>"110101110",
  35861=>"001111111",
  35862=>"101111000",
  35863=>"111010110",
  35864=>"110110000",
  35865=>"111000000",
  35866=>"000100110",
  35867=>"011100011",
  35868=>"100101111",
  35869=>"101000110",
  35870=>"111101111",
  35871=>"110101101",
  35872=>"110011010",
  35873=>"001001001",
  35874=>"101010011",
  35875=>"110101110",
  35876=>"010001000",
  35877=>"111101010",
  35878=>"011110111",
  35879=>"101001111",
  35880=>"010111010",
  35881=>"100110100",
  35882=>"010110111",
  35883=>"000010001",
  35884=>"000111100",
  35885=>"000000000",
  35886=>"110001100",
  35887=>"110110000",
  35888=>"000001001",
  35889=>"110001001",
  35890=>"010011011",
  35891=>"100000111",
  35892=>"001001001",
  35893=>"011011010",
  35894=>"000000001",
  35895=>"110011001",
  35896=>"111111010",
  35897=>"000111011",
  35898=>"011010110",
  35899=>"000111101",
  35900=>"001101001",
  35901=>"101111010",
  35902=>"101001001",
  35903=>"011111010",
  35904=>"100000010",
  35905=>"000110010",
  35906=>"100011100",
  35907=>"000110000",
  35908=>"100010000",
  35909=>"100111010",
  35910=>"100001001",
  35911=>"100000000",
  35912=>"111000011",
  35913=>"001010100",
  35914=>"100111101",
  35915=>"000011000",
  35916=>"000000010",
  35917=>"110100010",
  35918=>"111111001",
  35919=>"011000111",
  35920=>"110101111",
  35921=>"011111110",
  35922=>"000111111",
  35923=>"100000010",
  35924=>"011101111",
  35925=>"001001011",
  35926=>"101001100",
  35927=>"001011011",
  35928=>"111111001",
  35929=>"111100010",
  35930=>"000000010",
  35931=>"111001001",
  35932=>"001111110",
  35933=>"010100101",
  35934=>"011111000",
  35935=>"010100101",
  35936=>"000001010",
  35937=>"100010001",
  35938=>"010111110",
  35939=>"111111100",
  35940=>"111100010",
  35941=>"101011110",
  35942=>"100001001",
  35943=>"010011010",
  35944=>"111000111",
  35945=>"001101100",
  35946=>"110000010",
  35947=>"001001000",
  35948=>"001001010",
  35949=>"100101001",
  35950=>"101111111",
  35951=>"010110010",
  35952=>"110001111",
  35953=>"100100001",
  35954=>"111100110",
  35955=>"100010001",
  35956=>"010001010",
  35957=>"110110011",
  35958=>"100101100",
  35959=>"110001100",
  35960=>"100101111",
  35961=>"000110110",
  35962=>"111100100",
  35963=>"101010000",
  35964=>"010110110",
  35965=>"111000111",
  35966=>"010010111",
  35967=>"000000111",
  35968=>"111110100",
  35969=>"000010000",
  35970=>"010110100",
  35971=>"010111000",
  35972=>"111011111",
  35973=>"011111101",
  35974=>"000111100",
  35975=>"110001000",
  35976=>"001111100",
  35977=>"111000010",
  35978=>"010111111",
  35979=>"100100101",
  35980=>"010000000",
  35981=>"010101111",
  35982=>"111101111",
  35983=>"001001010",
  35984=>"001101111",
  35985=>"011110000",
  35986=>"001101110",
  35987=>"111100111",
  35988=>"000010111",
  35989=>"000000001",
  35990=>"000010010",
  35991=>"011101000",
  35992=>"001001001",
  35993=>"000100010",
  35994=>"001010100",
  35995=>"101110110",
  35996=>"011001110",
  35997=>"111110101",
  35998=>"011110111",
  35999=>"100010000",
  36000=>"010110010",
  36001=>"100010001",
  36002=>"000111010",
  36003=>"111011001",
  36004=>"111101001",
  36005=>"100000011",
  36006=>"111001010",
  36007=>"010101001",
  36008=>"000010001",
  36009=>"000000111",
  36010=>"100101111",
  36011=>"010001001",
  36012=>"100101001",
  36013=>"000010001",
  36014=>"010001111",
  36015=>"010010101",
  36016=>"101010111",
  36017=>"001001000",
  36018=>"101110101",
  36019=>"000100100",
  36020=>"110110101",
  36021=>"100101000",
  36022=>"000001011",
  36023=>"111000000",
  36024=>"110100110",
  36025=>"001001101",
  36026=>"111110011",
  36027=>"010001010",
  36028=>"110010101",
  36029=>"110110111",
  36030=>"111010111",
  36031=>"011110111",
  36032=>"010101000",
  36033=>"001010010",
  36034=>"001100000",
  36035=>"101110100",
  36036=>"001010001",
  36037=>"101111011",
  36038=>"100111111",
  36039=>"100001111",
  36040=>"100100000",
  36041=>"011111101",
  36042=>"111000110",
  36043=>"000000001",
  36044=>"000000100",
  36045=>"001001110",
  36046=>"001010101",
  36047=>"011111110",
  36048=>"111101111",
  36049=>"001101011",
  36050=>"011011111",
  36051=>"000101001",
  36052=>"110101010",
  36053=>"001011010",
  36054=>"101011010",
  36055=>"011011100",
  36056=>"011001000",
  36057=>"101100001",
  36058=>"111110001",
  36059=>"110101110",
  36060=>"110101101",
  36061=>"101011000",
  36062=>"111011000",
  36063=>"001111111",
  36064=>"101100111",
  36065=>"010001110",
  36066=>"100011100",
  36067=>"111110111",
  36068=>"000010011",
  36069=>"000001100",
  36070=>"001110101",
  36071=>"101010001",
  36072=>"110110000",
  36073=>"111001111",
  36074=>"101010111",
  36075=>"100101001",
  36076=>"001100000",
  36077=>"101101101",
  36078=>"101110100",
  36079=>"000101011",
  36080=>"110011011",
  36081=>"000100011",
  36082=>"011000101",
  36083=>"010000000",
  36084=>"011010110",
  36085=>"110111110",
  36086=>"100000111",
  36087=>"111011110",
  36088=>"101001000",
  36089=>"110001110",
  36090=>"101100000",
  36091=>"100001000",
  36092=>"001100100",
  36093=>"101110011",
  36094=>"101100101",
  36095=>"011110101",
  36096=>"000010000",
  36097=>"001001111",
  36098=>"010101101",
  36099=>"010010011",
  36100=>"011100001",
  36101=>"001000100",
  36102=>"111100000",
  36103=>"111000010",
  36104=>"000001011",
  36105=>"001110101",
  36106=>"110010100",
  36107=>"110000011",
  36108=>"110101100",
  36109=>"111110010",
  36110=>"000110111",
  36111=>"000100011",
  36112=>"101000010",
  36113=>"011000111",
  36114=>"110101001",
  36115=>"100001010",
  36116=>"000010000",
  36117=>"010010100",
  36118=>"100011101",
  36119=>"110011011",
  36120=>"001001011",
  36121=>"100111101",
  36122=>"101001101",
  36123=>"101000011",
  36124=>"101101011",
  36125=>"101011001",
  36126=>"011100010",
  36127=>"110101000",
  36128=>"011011110",
  36129=>"111111010",
  36130=>"110011010",
  36131=>"101000101",
  36132=>"001110101",
  36133=>"010100101",
  36134=>"110000001",
  36135=>"100110000",
  36136=>"010111100",
  36137=>"000110110",
  36138=>"101001110",
  36139=>"110111001",
  36140=>"010010110",
  36141=>"111110101",
  36142=>"110110010",
  36143=>"011100001",
  36144=>"000010011",
  36145=>"000101010",
  36146=>"111111101",
  36147=>"101000011",
  36148=>"110000100",
  36149=>"010000101",
  36150=>"001001110",
  36151=>"100011010",
  36152=>"011100111",
  36153=>"100101010",
  36154=>"000000110",
  36155=>"110110001",
  36156=>"010010101",
  36157=>"100110100",
  36158=>"011000100",
  36159=>"010111001",
  36160=>"101010100",
  36161=>"111111100",
  36162=>"101001001",
  36163=>"001111101",
  36164=>"101111111",
  36165=>"010010111",
  36166=>"110010010",
  36167=>"011101001",
  36168=>"010010001",
  36169=>"100100110",
  36170=>"001100001",
  36171=>"001100000",
  36172=>"011110011",
  36173=>"010000011",
  36174=>"101001000",
  36175=>"001011011",
  36176=>"111000100",
  36177=>"000100101",
  36178=>"111100100",
  36179=>"000001111",
  36180=>"100010011",
  36181=>"101110001",
  36182=>"000111000",
  36183=>"111110000",
  36184=>"011101010",
  36185=>"101110000",
  36186=>"010000100",
  36187=>"010010100",
  36188=>"100111100",
  36189=>"011010011",
  36190=>"110100000",
  36191=>"000111000",
  36192=>"101000100",
  36193=>"010000000",
  36194=>"111000111",
  36195=>"000101111",
  36196=>"111110111",
  36197=>"101110011",
  36198=>"110110101",
  36199=>"110001111",
  36200=>"010100100",
  36201=>"011100111",
  36202=>"000000000",
  36203=>"010101100",
  36204=>"010010100",
  36205=>"100111111",
  36206=>"010111101",
  36207=>"101111010",
  36208=>"011111010",
  36209=>"110101101",
  36210=>"100111010",
  36211=>"110001100",
  36212=>"101001000",
  36213=>"111011110",
  36214=>"001101111",
  36215=>"000001001",
  36216=>"111011110",
  36217=>"000111011",
  36218=>"110111101",
  36219=>"000001010",
  36220=>"000001110",
  36221=>"001110010",
  36222=>"110100100",
  36223=>"011111111",
  36224=>"011011000",
  36225=>"011000010",
  36226=>"111110011",
  36227=>"001000110",
  36228=>"101000111",
  36229=>"101011100",
  36230=>"000100101",
  36231=>"100000101",
  36232=>"000000101",
  36233=>"100101001",
  36234=>"010000110",
  36235=>"000010011",
  36236=>"011101101",
  36237=>"111011010",
  36238=>"001000010",
  36239=>"011010010",
  36240=>"100111111",
  36241=>"011000011",
  36242=>"110100100",
  36243=>"110010000",
  36244=>"100111100",
  36245=>"000000101",
  36246=>"110101111",
  36247=>"010000000",
  36248=>"000001000",
  36249=>"000011000",
  36250=>"101001011",
  36251=>"101110000",
  36252=>"010000100",
  36253=>"101100101",
  36254=>"110010001",
  36255=>"001101110",
  36256=>"000001001",
  36257=>"110110111",
  36258=>"100111101",
  36259=>"011010100",
  36260=>"111000011",
  36261=>"101001000",
  36262=>"111101111",
  36263=>"010000111",
  36264=>"001001110",
  36265=>"101000101",
  36266=>"001101001",
  36267=>"111110010",
  36268=>"010100001",
  36269=>"001111100",
  36270=>"011000111",
  36271=>"101111011",
  36272=>"011001010",
  36273=>"010010110",
  36274=>"010000111",
  36275=>"100011011",
  36276=>"011110010",
  36277=>"011010001",
  36278=>"000010011",
  36279=>"001010111",
  36280=>"001001001",
  36281=>"101011001",
  36282=>"011110100",
  36283=>"101000010",
  36284=>"010111110",
  36285=>"100001101",
  36286=>"111001100",
  36287=>"011011010",
  36288=>"111111100",
  36289=>"111111010",
  36290=>"000011011",
  36291=>"100011111",
  36292=>"100010000",
  36293=>"000001111",
  36294=>"110010110",
  36295=>"010110110",
  36296=>"100000011",
  36297=>"100000110",
  36298=>"110100110",
  36299=>"001000101",
  36300=>"000100011",
  36301=>"111110000",
  36302=>"000111001",
  36303=>"011110010",
  36304=>"110011110",
  36305=>"111000001",
  36306=>"011101001",
  36307=>"111100111",
  36308=>"000000000",
  36309=>"011010010",
  36310=>"101010111",
  36311=>"011101000",
  36312=>"000110010",
  36313=>"101010010",
  36314=>"010111111",
  36315=>"110111100",
  36316=>"011011010",
  36317=>"011001010",
  36318=>"001011100",
  36319=>"000000001",
  36320=>"000110000",
  36321=>"111011100",
  36322=>"101111011",
  36323=>"010100110",
  36324=>"100101101",
  36325=>"001010110",
  36326=>"111101110",
  36327=>"011110011",
  36328=>"000100101",
  36329=>"000010010",
  36330=>"000011000",
  36331=>"110110100",
  36332=>"001111101",
  36333=>"110111111",
  36334=>"111000001",
  36335=>"110000010",
  36336=>"000001100",
  36337=>"100111010",
  36338=>"000111010",
  36339=>"111111001",
  36340=>"101011001",
  36341=>"111111000",
  36342=>"011100110",
  36343=>"110010000",
  36344=>"011100011",
  36345=>"100111101",
  36346=>"111011110",
  36347=>"100000111",
  36348=>"100111010",
  36349=>"101110011",
  36350=>"111111011",
  36351=>"101110010",
  36352=>"101000011",
  36353=>"000000101",
  36354=>"011010001",
  36355=>"000001001",
  36356=>"001011100",
  36357=>"111110001",
  36358=>"001000010",
  36359=>"111100110",
  36360=>"000101111",
  36361=>"111100101",
  36362=>"100001100",
  36363=>"010001111",
  36364=>"101101110",
  36365=>"111001000",
  36366=>"001000000",
  36367=>"010010010",
  36368=>"100111000",
  36369=>"001010000",
  36370=>"011101111",
  36371=>"110000000",
  36372=>"100111101",
  36373=>"000010101",
  36374=>"111100110",
  36375=>"010111110",
  36376=>"101011111",
  36377=>"111010011",
  36378=>"111011110",
  36379=>"011101000",
  36380=>"001000000",
  36381=>"110110011",
  36382=>"000111000",
  36383=>"001100000",
  36384=>"001011100",
  36385=>"000110110",
  36386=>"100001010",
  36387=>"011001000",
  36388=>"101001001",
  36389=>"100000111",
  36390=>"110001111",
  36391=>"011111000",
  36392=>"010111111",
  36393=>"100110010",
  36394=>"001111111",
  36395=>"111101000",
  36396=>"101111100",
  36397=>"110000010",
  36398=>"100110001",
  36399=>"011000111",
  36400=>"010100111",
  36401=>"010011001",
  36402=>"110111100",
  36403=>"111110101",
  36404=>"010011000",
  36405=>"111111111",
  36406=>"001111010",
  36407=>"001100011",
  36408=>"110011001",
  36409=>"110001011",
  36410=>"000100001",
  36411=>"001011000",
  36412=>"001010100",
  36413=>"100010111",
  36414=>"101101011",
  36415=>"100000110",
  36416=>"000101000",
  36417=>"100011101",
  36418=>"110101110",
  36419=>"110011111",
  36420=>"100000100",
  36421=>"001000010",
  36422=>"010011011",
  36423=>"100001001",
  36424=>"100100000",
  36425=>"110111101",
  36426=>"100000010",
  36427=>"001011000",
  36428=>"111000000",
  36429=>"000111111",
  36430=>"001101001",
  36431=>"111110011",
  36432=>"101100001",
  36433=>"100101000",
  36434=>"010000000",
  36435=>"000000011",
  36436=>"010100001",
  36437=>"010111100",
  36438=>"101001100",
  36439=>"101001000",
  36440=>"011010110",
  36441=>"000111001",
  36442=>"010011000",
  36443=>"111011100",
  36444=>"010000010",
  36445=>"101000101",
  36446=>"000101111",
  36447=>"000101110",
  36448=>"000110000",
  36449=>"101011111",
  36450=>"100110111",
  36451=>"100111111",
  36452=>"110000000",
  36453=>"100011000",
  36454=>"101010100",
  36455=>"010000010",
  36456=>"110000010",
  36457=>"101101010",
  36458=>"010000010",
  36459=>"100110101",
  36460=>"000011011",
  36461=>"001010110",
  36462=>"001010010",
  36463=>"000001011",
  36464=>"010110001",
  36465=>"111101100",
  36466=>"111100001",
  36467=>"111010110",
  36468=>"101010111",
  36469=>"001001100",
  36470=>"101010001",
  36471=>"000000100",
  36472=>"100110101",
  36473=>"010111101",
  36474=>"101010110",
  36475=>"011011001",
  36476=>"011011100",
  36477=>"101011001",
  36478=>"001100011",
  36479=>"111001000",
  36480=>"001110101",
  36481=>"111000001",
  36482=>"010000010",
  36483=>"101001001",
  36484=>"010101111",
  36485=>"111011100",
  36486=>"000110111",
  36487=>"001001010",
  36488=>"011110100",
  36489=>"100100100",
  36490=>"010100101",
  36491=>"010010011",
  36492=>"000100011",
  36493=>"111010110",
  36494=>"011101011",
  36495=>"010000000",
  36496=>"100000111",
  36497=>"000100100",
  36498=>"111001111",
  36499=>"100111001",
  36500=>"011001100",
  36501=>"101010111",
  36502=>"010001000",
  36503=>"000010110",
  36504=>"011101010",
  36505=>"010111100",
  36506=>"001110101",
  36507=>"101110001",
  36508=>"101001111",
  36509=>"111111101",
  36510=>"100100111",
  36511=>"110110110",
  36512=>"101111011",
  36513=>"001011011",
  36514=>"001100111",
  36515=>"111001110",
  36516=>"011001001",
  36517=>"100100000",
  36518=>"100101001",
  36519=>"011001011",
  36520=>"111111100",
  36521=>"110000000",
  36522=>"110111011",
  36523=>"100011100",
  36524=>"101111101",
  36525=>"010111000",
  36526=>"111101000",
  36527=>"101011111",
  36528=>"000010001",
  36529=>"000111100",
  36530=>"001100010",
  36531=>"101100101",
  36532=>"110111000",
  36533=>"001100010",
  36534=>"111001110",
  36535=>"111110101",
  36536=>"011101000",
  36537=>"100010111",
  36538=>"111010101",
  36539=>"101011010",
  36540=>"000000001",
  36541=>"001011010",
  36542=>"111101010",
  36543=>"111010010",
  36544=>"100110010",
  36545=>"100011111",
  36546=>"010100111",
  36547=>"101111000",
  36548=>"011011011",
  36549=>"010011110",
  36550=>"100001110",
  36551=>"001111100",
  36552=>"100011111",
  36553=>"000011101",
  36554=>"011100100",
  36555=>"010101000",
  36556=>"011010100",
  36557=>"000010000",
  36558=>"001010110",
  36559=>"011010010",
  36560=>"101110111",
  36561=>"000100011",
  36562=>"000001011",
  36563=>"001111111",
  36564=>"100101111",
  36565=>"001101110",
  36566=>"111010101",
  36567=>"000001111",
  36568=>"000001000",
  36569=>"001011000",
  36570=>"011010111",
  36571=>"110110111",
  36572=>"110101010",
  36573=>"101101010",
  36574=>"100100001",
  36575=>"010001000",
  36576=>"010101110",
  36577=>"010101001",
  36578=>"000001010",
  36579=>"110001011",
  36580=>"101000010",
  36581=>"010001000",
  36582=>"111111111",
  36583=>"110000000",
  36584=>"001101001",
  36585=>"100101110",
  36586=>"110001111",
  36587=>"100110101",
  36588=>"011101100",
  36589=>"111001010",
  36590=>"001100101",
  36591=>"111011111",
  36592=>"111100111",
  36593=>"010010101",
  36594=>"110001001",
  36595=>"100101000",
  36596=>"001110100",
  36597=>"000110000",
  36598=>"100011111",
  36599=>"110110001",
  36600=>"100010111",
  36601=>"010100000",
  36602=>"110110111",
  36603=>"111110110",
  36604=>"101100001",
  36605=>"001101101",
  36606=>"111101110",
  36607=>"100101100",
  36608=>"001110111",
  36609=>"110010011",
  36610=>"010111010",
  36611=>"111100000",
  36612=>"000001011",
  36613=>"011110011",
  36614=>"011111011",
  36615=>"010100000",
  36616=>"101011011",
  36617=>"010001110",
  36618=>"100111111",
  36619=>"011000011",
  36620=>"101001111",
  36621=>"111111101",
  36622=>"101000000",
  36623=>"100110001",
  36624=>"110100001",
  36625=>"011101010",
  36626=>"100111011",
  36627=>"010110001",
  36628=>"001011000",
  36629=>"110000100",
  36630=>"101111100",
  36631=>"111111010",
  36632=>"011010011",
  36633=>"111000101",
  36634=>"111111100",
  36635=>"110010101",
  36636=>"011100000",
  36637=>"101010011",
  36638=>"000100111",
  36639=>"100001000",
  36640=>"100001111",
  36641=>"010011101",
  36642=>"011011001",
  36643=>"011100100",
  36644=>"101100101",
  36645=>"001001100",
  36646=>"101000011",
  36647=>"111110010",
  36648=>"000110110",
  36649=>"101001011",
  36650=>"101011000",
  36651=>"001001101",
  36652=>"000011101",
  36653=>"001011000",
  36654=>"100110000",
  36655=>"001001010",
  36656=>"011101011",
  36657=>"000011111",
  36658=>"111110001",
  36659=>"100011000",
  36660=>"001000011",
  36661=>"101000010",
  36662=>"111000111",
  36663=>"000101001",
  36664=>"000001010",
  36665=>"111000100",
  36666=>"111100010",
  36667=>"101110101",
  36668=>"110100111",
  36669=>"001000001",
  36670=>"000100010",
  36671=>"110001000",
  36672=>"011100111",
  36673=>"000010111",
  36674=>"101100101",
  36675=>"100000001",
  36676=>"011000110",
  36677=>"001010100",
  36678=>"000101100",
  36679=>"010000110",
  36680=>"001010111",
  36681=>"010001100",
  36682=>"010000101",
  36683=>"000101101",
  36684=>"101111011",
  36685=>"010000000",
  36686=>"010001001",
  36687=>"010110001",
  36688=>"110110110",
  36689=>"100100000",
  36690=>"110000001",
  36691=>"011101011",
  36692=>"111101101",
  36693=>"000000111",
  36694=>"011010001",
  36695=>"010101000",
  36696=>"100101010",
  36697=>"110111011",
  36698=>"110101001",
  36699=>"101010100",
  36700=>"000101010",
  36701=>"010100110",
  36702=>"111011001",
  36703=>"000000100",
  36704=>"100000011",
  36705=>"011001010",
  36706=>"010110000",
  36707=>"100101100",
  36708=>"001000101",
  36709=>"000000100",
  36710=>"101010110",
  36711=>"100111111",
  36712=>"010010100",
  36713=>"101101111",
  36714=>"110101001",
  36715=>"011100010",
  36716=>"101000000",
  36717=>"101001001",
  36718=>"110110011",
  36719=>"101010111",
  36720=>"110010000",
  36721=>"101100110",
  36722=>"111011011",
  36723=>"000101010",
  36724=>"011001000",
  36725=>"111110011",
  36726=>"101110111",
  36727=>"110110011",
  36728=>"010010000",
  36729=>"010010001",
  36730=>"000011011",
  36731=>"010100000",
  36732=>"001100011",
  36733=>"010011001",
  36734=>"100111111",
  36735=>"110011010",
  36736=>"011101000",
  36737=>"110011000",
  36738=>"010011001",
  36739=>"000010000",
  36740=>"111100011",
  36741=>"000101111",
  36742=>"111100111",
  36743=>"010101100",
  36744=>"111101110",
  36745=>"111101110",
  36746=>"111111110",
  36747=>"101101101",
  36748=>"110111110",
  36749=>"111110100",
  36750=>"010000111",
  36751=>"001111010",
  36752=>"100100110",
  36753=>"000110010",
  36754=>"010001100",
  36755=>"101110010",
  36756=>"110110000",
  36757=>"010100101",
  36758=>"001011011",
  36759=>"001101111",
  36760=>"010001011",
  36761=>"110100000",
  36762=>"001111001",
  36763=>"011101001",
  36764=>"100111011",
  36765=>"100101000",
  36766=>"001011111",
  36767=>"000011110",
  36768=>"010001011",
  36769=>"110111110",
  36770=>"111001111",
  36771=>"110111001",
  36772=>"110100111",
  36773=>"001000010",
  36774=>"110000010",
  36775=>"110000111",
  36776=>"100100111",
  36777=>"011010010",
  36778=>"010010100",
  36779=>"010111100",
  36780=>"101111000",
  36781=>"110111000",
  36782=>"010100111",
  36783=>"000001000",
  36784=>"100010011",
  36785=>"011101011",
  36786=>"111101110",
  36787=>"110011100",
  36788=>"110010000",
  36789=>"010011100",
  36790=>"001001101",
  36791=>"010111100",
  36792=>"011110110",
  36793=>"111110100",
  36794=>"110010000",
  36795=>"100011100",
  36796=>"000011111",
  36797=>"100101001",
  36798=>"111111001",
  36799=>"101100101",
  36800=>"010010110",
  36801=>"011011111",
  36802=>"111011001",
  36803=>"111001011",
  36804=>"000110001",
  36805=>"000111100",
  36806=>"011000001",
  36807=>"000111101",
  36808=>"110110100",
  36809=>"000010000",
  36810=>"100101111",
  36811=>"100100100",
  36812=>"100111011",
  36813=>"011111110",
  36814=>"110011000",
  36815=>"101001111",
  36816=>"101010111",
  36817=>"010100111",
  36818=>"011110001",
  36819=>"011101000",
  36820=>"100011100",
  36821=>"110100101",
  36822=>"101001101",
  36823=>"100100101",
  36824=>"100110110",
  36825=>"100111100",
  36826=>"011110011",
  36827=>"111010010",
  36828=>"011101101",
  36829=>"111111111",
  36830=>"110001000",
  36831=>"000011100",
  36832=>"101011011",
  36833=>"000100100",
  36834=>"100111111",
  36835=>"001111001",
  36836=>"111100010",
  36837=>"011001110",
  36838=>"001100010",
  36839=>"000001000",
  36840=>"010111001",
  36841=>"011110100",
  36842=>"110010111",
  36843=>"100111000",
  36844=>"011011110",
  36845=>"101011001",
  36846=>"001011001",
  36847=>"101110010",
  36848=>"011011111",
  36849=>"001001001",
  36850=>"011101010",
  36851=>"100100010",
  36852=>"011100110",
  36853=>"101101010",
  36854=>"000010101",
  36855=>"111000001",
  36856=>"010111001",
  36857=>"000000010",
  36858=>"111101001",
  36859=>"110010111",
  36860=>"101100011",
  36861=>"100011110",
  36862=>"011001111",
  36863=>"101101110",
  36864=>"111001000",
  36865=>"100010000",
  36866=>"100010110",
  36867=>"100101100",
  36868=>"111010010",
  36869=>"110000000",
  36870=>"000100100",
  36871=>"111000101",
  36872=>"010000000",
  36873=>"011100100",
  36874=>"100010100",
  36875=>"011101000",
  36876=>"111011010",
  36877=>"000010100",
  36878=>"101001111",
  36879=>"101110000",
  36880=>"101101011",
  36881=>"111001100",
  36882=>"101010100",
  36883=>"010100001",
  36884=>"011100111",
  36885=>"111110111",
  36886=>"110111110",
  36887=>"000001100",
  36888=>"011000000",
  36889=>"000011111",
  36890=>"010011101",
  36891=>"001001010",
  36892=>"101101010",
  36893=>"100111011",
  36894=>"101101100",
  36895=>"101111010",
  36896=>"011111011",
  36897=>"100000011",
  36898=>"110000110",
  36899=>"000000101",
  36900=>"000101111",
  36901=>"011000010",
  36902=>"001110011",
  36903=>"011110000",
  36904=>"111110010",
  36905=>"011101001",
  36906=>"101000001",
  36907=>"000101010",
  36908=>"000001010",
  36909=>"010100010",
  36910=>"111001110",
  36911=>"010110101",
  36912=>"110110101",
  36913=>"010010010",
  36914=>"011001111",
  36915=>"111010000",
  36916=>"111001111",
  36917=>"001000001",
  36918=>"100100010",
  36919=>"101001010",
  36920=>"101110000",
  36921=>"001100010",
  36922=>"101100000",
  36923=>"110001011",
  36924=>"011000000",
  36925=>"000001001",
  36926=>"000100100",
  36927=>"110010100",
  36928=>"000000101",
  36929=>"000000000",
  36930=>"111000010",
  36931=>"010010100",
  36932=>"100010101",
  36933=>"011001010",
  36934=>"101111100",
  36935=>"001011001",
  36936=>"111001010",
  36937=>"001001001",
  36938=>"100000110",
  36939=>"110010000",
  36940=>"100010101",
  36941=>"110111111",
  36942=>"011001110",
  36943=>"100001000",
  36944=>"110010101",
  36945=>"001100011",
  36946=>"100100100",
  36947=>"111101010",
  36948=>"111100110",
  36949=>"010100010",
  36950=>"111001000",
  36951=>"000001000",
  36952=>"011111111",
  36953=>"111011001",
  36954=>"101010010",
  36955=>"011010011",
  36956=>"000010101",
  36957=>"101100111",
  36958=>"011011111",
  36959=>"110010010",
  36960=>"110001000",
  36961=>"101110110",
  36962=>"011111101",
  36963=>"010011101",
  36964=>"010001000",
  36965=>"111111110",
  36966=>"001010011",
  36967=>"000011010",
  36968=>"111100101",
  36969=>"110111000",
  36970=>"011110111",
  36971=>"101010111",
  36972=>"110001101",
  36973=>"110101110",
  36974=>"000000000",
  36975=>"100010111",
  36976=>"111010000",
  36977=>"000000111",
  36978=>"101100011",
  36979=>"010101010",
  36980=>"100100011",
  36981=>"110001001",
  36982=>"000001111",
  36983=>"001111110",
  36984=>"111100001",
  36985=>"111011011",
  36986=>"011011100",
  36987=>"100101110",
  36988=>"100010001",
  36989=>"111010011",
  36990=>"111000010",
  36991=>"001010101",
  36992=>"100110100",
  36993=>"100000010",
  36994=>"110101100",
  36995=>"100111011",
  36996=>"100110000",
  36997=>"001101111",
  36998=>"110010110",
  36999=>"001000100",
  37000=>"000000001",
  37001=>"111000110",
  37002=>"110001110",
  37003=>"110011000",
  37004=>"000100100",
  37005=>"111111110",
  37006=>"110110011",
  37007=>"000101000",
  37008=>"110111111",
  37009=>"001101000",
  37010=>"001010000",
  37011=>"111010010",
  37012=>"111100000",
  37013=>"100111111",
  37014=>"100001001",
  37015=>"100110111",
  37016=>"011100011",
  37017=>"000100000",
  37018=>"100110111",
  37019=>"000011001",
  37020=>"001110011",
  37021=>"100100000",
  37022=>"111011101",
  37023=>"011011001",
  37024=>"111001001",
  37025=>"001100011",
  37026=>"000001010",
  37027=>"001111001",
  37028=>"111100010",
  37029=>"100100111",
  37030=>"001111101",
  37031=>"011111000",
  37032=>"111111100",
  37033=>"001011010",
  37034=>"001010001",
  37035=>"010001001",
  37036=>"000010010",
  37037=>"000001010",
  37038=>"111111100",
  37039=>"011011101",
  37040=>"100101001",
  37041=>"111100111",
  37042=>"100111001",
  37043=>"010000111",
  37044=>"000011101",
  37045=>"100100100",
  37046=>"010101010",
  37047=>"011111110",
  37048=>"101001110",
  37049=>"011001001",
  37050=>"110010101",
  37051=>"101010100",
  37052=>"101000001",
  37053=>"010111011",
  37054=>"010000110",
  37055=>"011111011",
  37056=>"001001000",
  37057=>"101111100",
  37058=>"100111110",
  37059=>"100010010",
  37060=>"000011101",
  37061=>"001110110",
  37062=>"000100010",
  37063=>"001100111",
  37064=>"101001011",
  37065=>"110001000",
  37066=>"000010000",
  37067=>"000011111",
  37068=>"010110010",
  37069=>"000001100",
  37070=>"000111111",
  37071=>"010110011",
  37072=>"100100000",
  37073=>"100000101",
  37074=>"010000000",
  37075=>"000110110",
  37076=>"010011111",
  37077=>"101111011",
  37078=>"000000000",
  37079=>"100101010",
  37080=>"101100111",
  37081=>"001001000",
  37082=>"010001110",
  37083=>"011010001",
  37084=>"001011100",
  37085=>"111010101",
  37086=>"010000001",
  37087=>"000000110",
  37088=>"000101000",
  37089=>"001011101",
  37090=>"100111001",
  37091=>"111100101",
  37092=>"100011101",
  37093=>"010010110",
  37094=>"110000101",
  37095=>"001100101",
  37096=>"000011001",
  37097=>"100010111",
  37098=>"010001111",
  37099=>"011101101",
  37100=>"110100111",
  37101=>"001111011",
  37102=>"111110011",
  37103=>"111100101",
  37104=>"001000001",
  37105=>"111101100",
  37106=>"000101111",
  37107=>"011011110",
  37108=>"110110011",
  37109=>"101001000",
  37110=>"000101101",
  37111=>"010010100",
  37112=>"010111100",
  37113=>"111101101",
  37114=>"110100001",
  37115=>"110010011",
  37116=>"100101001",
  37117=>"001001000",
  37118=>"010010110",
  37119=>"101100110",
  37120=>"100010011",
  37121=>"111100011",
  37122=>"011001001",
  37123=>"011000101",
  37124=>"010111100",
  37125=>"111011001",
  37126=>"111111001",
  37127=>"100000101",
  37128=>"000101111",
  37129=>"001100100",
  37130=>"011101010",
  37131=>"010101101",
  37132=>"110010000",
  37133=>"111111010",
  37134=>"100010011",
  37135=>"110101111",
  37136=>"100011111",
  37137=>"011111011",
  37138=>"101110110",
  37139=>"011000000",
  37140=>"001111001",
  37141=>"111101110",
  37142=>"010101001",
  37143=>"100100100",
  37144=>"011000101",
  37145=>"000101111",
  37146=>"001000110",
  37147=>"000010000",
  37148=>"010000101",
  37149=>"011100100",
  37150=>"110001011",
  37151=>"101101010",
  37152=>"010110111",
  37153=>"111011010",
  37154=>"110100001",
  37155=>"111010010",
  37156=>"001000100",
  37157=>"010110101",
  37158=>"010110110",
  37159=>"100101100",
  37160=>"001001111",
  37161=>"010010111",
  37162=>"100011000",
  37163=>"111100000",
  37164=>"010011001",
  37165=>"000001100",
  37166=>"001101111",
  37167=>"111011011",
  37168=>"001001101",
  37169=>"000111111",
  37170=>"000101001",
  37171=>"001110000",
  37172=>"110100100",
  37173=>"011111001",
  37174=>"000001001",
  37175=>"011100000",
  37176=>"101100000",
  37177=>"000011010",
  37178=>"010101100",
  37179=>"001101000",
  37180=>"111010001",
  37181=>"000000101",
  37182=>"010101111",
  37183=>"100101001",
  37184=>"111011110",
  37185=>"101010000",
  37186=>"110100100",
  37187=>"111000111",
  37188=>"101011110",
  37189=>"000100111",
  37190=>"100000100",
  37191=>"101100001",
  37192=>"111111011",
  37193=>"001110100",
  37194=>"001111011",
  37195=>"010011111",
  37196=>"010000010",
  37197=>"110111001",
  37198=>"000111111",
  37199=>"100111001",
  37200=>"111100010",
  37201=>"001000001",
  37202=>"100001110",
  37203=>"001000000",
  37204=>"010001000",
  37205=>"000101010",
  37206=>"101000111",
  37207=>"000101110",
  37208=>"110101011",
  37209=>"000011000",
  37210=>"010000011",
  37211=>"010000000",
  37212=>"010000110",
  37213=>"110010100",
  37214=>"110111010",
  37215=>"101001011",
  37216=>"011010111",
  37217=>"110101000",
  37218=>"001010111",
  37219=>"001010101",
  37220=>"100110110",
  37221=>"010111011",
  37222=>"001111011",
  37223=>"111001001",
  37224=>"001010101",
  37225=>"001100001",
  37226=>"111000011",
  37227=>"000110000",
  37228=>"010011010",
  37229=>"000011100",
  37230=>"101100101",
  37231=>"011101010",
  37232=>"100110010",
  37233=>"010000001",
  37234=>"001011100",
  37235=>"010101100",
  37236=>"011000111",
  37237=>"111011010",
  37238=>"101010011",
  37239=>"010110000",
  37240=>"011110001",
  37241=>"010000010",
  37242=>"101001101",
  37243=>"101101010",
  37244=>"001000111",
  37245=>"011101111",
  37246=>"100111011",
  37247=>"111000110",
  37248=>"100011100",
  37249=>"001100010",
  37250=>"101100101",
  37251=>"110001011",
  37252=>"011000001",
  37253=>"000101001",
  37254=>"110001100",
  37255=>"010011101",
  37256=>"011101101",
  37257=>"001110101",
  37258=>"110001000",
  37259=>"001000001",
  37260=>"001000000",
  37261=>"100001001",
  37262=>"110000101",
  37263=>"000011000",
  37264=>"111010100",
  37265=>"001101111",
  37266=>"101000110",
  37267=>"111010111",
  37268=>"100010101",
  37269=>"001100101",
  37270=>"110001111",
  37271=>"110100100",
  37272=>"000101110",
  37273=>"100100101",
  37274=>"110001010",
  37275=>"111011001",
  37276=>"001010010",
  37277=>"110001100",
  37278=>"011110011",
  37279=>"000011111",
  37280=>"101110101",
  37281=>"110101111",
  37282=>"000000001",
  37283=>"100100100",
  37284=>"000011010",
  37285=>"010110001",
  37286=>"110000101",
  37287=>"001011111",
  37288=>"101100100",
  37289=>"001100111",
  37290=>"001010101",
  37291=>"111101000",
  37292=>"110011101",
  37293=>"100011001",
  37294=>"111111011",
  37295=>"000001100",
  37296=>"111110110",
  37297=>"100100110",
  37298=>"011110100",
  37299=>"001001000",
  37300=>"110110100",
  37301=>"110011110",
  37302=>"100011100",
  37303=>"010100111",
  37304=>"110010010",
  37305=>"101100000",
  37306=>"000000000",
  37307=>"100101100",
  37308=>"110100100",
  37309=>"001010111",
  37310=>"100100010",
  37311=>"110010000",
  37312=>"100000100",
  37313=>"010011000",
  37314=>"101000110",
  37315=>"110110011",
  37316=>"001011010",
  37317=>"101110101",
  37318=>"010100000",
  37319=>"001100100",
  37320=>"100010010",
  37321=>"110000100",
  37322=>"101001100",
  37323=>"100100000",
  37324=>"110010110",
  37325=>"111011000",
  37326=>"001100001",
  37327=>"100110000",
  37328=>"010101000",
  37329=>"100011001",
  37330=>"000011111",
  37331=>"000011000",
  37332=>"001111111",
  37333=>"111100110",
  37334=>"000110011",
  37335=>"001011010",
  37336=>"010110011",
  37337=>"110110111",
  37338=>"111111001",
  37339=>"100000111",
  37340=>"000111101",
  37341=>"111110000",
  37342=>"000101010",
  37343=>"010010110",
  37344=>"110110100",
  37345=>"010011110",
  37346=>"000011011",
  37347=>"110100011",
  37348=>"111100100",
  37349=>"110101010",
  37350=>"110101000",
  37351=>"000111101",
  37352=>"010100001",
  37353=>"100101010",
  37354=>"100000000",
  37355=>"001010101",
  37356=>"111100101",
  37357=>"000101100",
  37358=>"011110000",
  37359=>"111000001",
  37360=>"010110001",
  37361=>"000001011",
  37362=>"101111000",
  37363=>"111010110",
  37364=>"110010101",
  37365=>"000000000",
  37366=>"011001110",
  37367=>"101111101",
  37368=>"101110100",
  37369=>"001101000",
  37370=>"111101101",
  37371=>"110010001",
  37372=>"001110111",
  37373=>"000011010",
  37374=>"000010000",
  37375=>"000000000",
  37376=>"100011100",
  37377=>"010111001",
  37378=>"001011101",
  37379=>"010000001",
  37380=>"100111101",
  37381=>"001110111",
  37382=>"110001010",
  37383=>"111011001",
  37384=>"011100101",
  37385=>"011001111",
  37386=>"100110011",
  37387=>"000101100",
  37388=>"000001110",
  37389=>"000100101",
  37390=>"001110000",
  37391=>"100100000",
  37392=>"001001111",
  37393=>"011111111",
  37394=>"110010111",
  37395=>"110111101",
  37396=>"110011010",
  37397=>"110001111",
  37398=>"100111010",
  37399=>"101111001",
  37400=>"010101111",
  37401=>"010110100",
  37402=>"011010100",
  37403=>"000011100",
  37404=>"011001110",
  37405=>"011000000",
  37406=>"000101111",
  37407=>"111001111",
  37408=>"101001111",
  37409=>"010000111",
  37410=>"100000000",
  37411=>"111001110",
  37412=>"111011111",
  37413=>"100101011",
  37414=>"010101010",
  37415=>"010001001",
  37416=>"111110001",
  37417=>"100110111",
  37418=>"111000000",
  37419=>"111111000",
  37420=>"100001111",
  37421=>"110111011",
  37422=>"000101111",
  37423=>"111101011",
  37424=>"101000011",
  37425=>"101001101",
  37426=>"101000100",
  37427=>"001000011",
  37428=>"001011001",
  37429=>"000000001",
  37430=>"101010100",
  37431=>"000110000",
  37432=>"101100000",
  37433=>"111110110",
  37434=>"010100010",
  37435=>"100101110",
  37436=>"100010100",
  37437=>"101101101",
  37438=>"101111011",
  37439=>"001001101",
  37440=>"111110110",
  37441=>"000110010",
  37442=>"001000000",
  37443=>"010100010",
  37444=>"000000101",
  37445=>"011111001",
  37446=>"001000110",
  37447=>"100010000",
  37448=>"011100010",
  37449=>"100011011",
  37450=>"001101100",
  37451=>"100000101",
  37452=>"110011010",
  37453=>"110101110",
  37454=>"011011110",
  37455=>"011110011",
  37456=>"110001101",
  37457=>"001110000",
  37458=>"111001111",
  37459=>"100010001",
  37460=>"110101100",
  37461=>"001111001",
  37462=>"101101001",
  37463=>"101101100",
  37464=>"010100010",
  37465=>"000111010",
  37466=>"000011000",
  37467=>"110100010",
  37468=>"001101001",
  37469=>"001000101",
  37470=>"100100111",
  37471=>"010001001",
  37472=>"001100110",
  37473=>"000000110",
  37474=>"010010101",
  37475=>"000000111",
  37476=>"100011001",
  37477=>"111111100",
  37478=>"100111101",
  37479=>"111010110",
  37480=>"011011100",
  37481=>"001011100",
  37482=>"000000111",
  37483=>"101111110",
  37484=>"000110000",
  37485=>"100001111",
  37486=>"101101010",
  37487=>"110011101",
  37488=>"001101110",
  37489=>"101100000",
  37490=>"100001010",
  37491=>"001110001",
  37492=>"111101111",
  37493=>"101000001",
  37494=>"110011110",
  37495=>"101110111",
  37496=>"000010000",
  37497=>"101001100",
  37498=>"011111001",
  37499=>"011100000",
  37500=>"000000000",
  37501=>"001000000",
  37502=>"010101101",
  37503=>"100111101",
  37504=>"001101010",
  37505=>"110111110",
  37506=>"101001110",
  37507=>"010000111",
  37508=>"101110100",
  37509=>"100000001",
  37510=>"001111001",
  37511=>"111101001",
  37512=>"000111101",
  37513=>"010001111",
  37514=>"001111010",
  37515=>"100000010",
  37516=>"010010010",
  37517=>"001000000",
  37518=>"101011000",
  37519=>"011101000",
  37520=>"011010000",
  37521=>"011011011",
  37522=>"000010010",
  37523=>"101100110",
  37524=>"101010100",
  37525=>"100110100",
  37526=>"000000111",
  37527=>"000001110",
  37528=>"000001010",
  37529=>"111010100",
  37530=>"100101000",
  37531=>"101100000",
  37532=>"110010100",
  37533=>"010010111",
  37534=>"011001011",
  37535=>"000110100",
  37536=>"100100010",
  37537=>"001000110",
  37538=>"100100010",
  37539=>"010010001",
  37540=>"110101000",
  37541=>"000110001",
  37542=>"101111010",
  37543=>"001010000",
  37544=>"111001001",
  37545=>"001110101",
  37546=>"011100000",
  37547=>"001101001",
  37548=>"110010100",
  37549=>"001110100",
  37550=>"111111100",
  37551=>"001001010",
  37552=>"000000010",
  37553=>"000010111",
  37554=>"100001010",
  37555=>"100001010",
  37556=>"101101011",
  37557=>"011011011",
  37558=>"100010001",
  37559=>"001011100",
  37560=>"000011100",
  37561=>"100000111",
  37562=>"011010011",
  37563=>"010001001",
  37564=>"100011011",
  37565=>"010011011",
  37566=>"011010001",
  37567=>"100100011",
  37568=>"110111101",
  37569=>"101101000",
  37570=>"111111101",
  37571=>"001011100",
  37572=>"000011101",
  37573=>"000001111",
  37574=>"111001101",
  37575=>"010000000",
  37576=>"110101000",
  37577=>"101111110",
  37578=>"111000110",
  37579=>"111101001",
  37580=>"000001000",
  37581=>"001010100",
  37582=>"110101100",
  37583=>"011001111",
  37584=>"010110000",
  37585=>"110111100",
  37586=>"111100010",
  37587=>"000100000",
  37588=>"110100101",
  37589=>"000010001",
  37590=>"111000001",
  37591=>"100111111",
  37592=>"100110101",
  37593=>"010001000",
  37594=>"110001011",
  37595=>"110101100",
  37596=>"101101011",
  37597=>"110000100",
  37598=>"110001100",
  37599=>"101101111",
  37600=>"100010100",
  37601=>"110111010",
  37602=>"100010111",
  37603=>"010100110",
  37604=>"001110110",
  37605=>"001011101",
  37606=>"010010101",
  37607=>"000110000",
  37608=>"010100110",
  37609=>"011100111",
  37610=>"010111100",
  37611=>"011101101",
  37612=>"100011000",
  37613=>"000001001",
  37614=>"000101001",
  37615=>"111110010",
  37616=>"001110011",
  37617=>"001110100",
  37618=>"000000000",
  37619=>"111011101",
  37620=>"010101110",
  37621=>"111000111",
  37622=>"001011100",
  37623=>"101000100",
  37624=>"111010001",
  37625=>"011111001",
  37626=>"010110101",
  37627=>"001100000",
  37628=>"011010010",
  37629=>"000110100",
  37630=>"010101011",
  37631=>"110001000",
  37632=>"110010010",
  37633=>"011111001",
  37634=>"111100010",
  37635=>"101001000",
  37636=>"110001001",
  37637=>"001100011",
  37638=>"101001011",
  37639=>"100011000",
  37640=>"100000001",
  37641=>"111101011",
  37642=>"000010000",
  37643=>"000001110",
  37644=>"000000101",
  37645=>"010010010",
  37646=>"100001010",
  37647=>"010000001",
  37648=>"011100010",
  37649=>"100110111",
  37650=>"111100000",
  37651=>"110000110",
  37652=>"000010010",
  37653=>"000011111",
  37654=>"110000000",
  37655=>"001000010",
  37656=>"001010000",
  37657=>"011010001",
  37658=>"000001000",
  37659=>"000010010",
  37660=>"010000000",
  37661=>"101001100",
  37662=>"100100100",
  37663=>"011011101",
  37664=>"100010100",
  37665=>"110101111",
  37666=>"000100011",
  37667=>"010000010",
  37668=>"000100101",
  37669=>"101100001",
  37670=>"000100110",
  37671=>"010110001",
  37672=>"101011100",
  37673=>"000101000",
  37674=>"101110010",
  37675=>"110001011",
  37676=>"100111011",
  37677=>"100111110",
  37678=>"111101011",
  37679=>"000001101",
  37680=>"000000000",
  37681=>"001101100",
  37682=>"000110000",
  37683=>"111000000",
  37684=>"111011010",
  37685=>"110010110",
  37686=>"110101011",
  37687=>"000001100",
  37688=>"101100000",
  37689=>"101110101",
  37690=>"000000010",
  37691=>"010001000",
  37692=>"101010101",
  37693=>"111000001",
  37694=>"001000000",
  37695=>"011111011",
  37696=>"011100110",
  37697=>"101111000",
  37698=>"101010111",
  37699=>"001000110",
  37700=>"010110000",
  37701=>"010111011",
  37702=>"000001001",
  37703=>"001101100",
  37704=>"101110001",
  37705=>"000110000",
  37706=>"010010111",
  37707=>"001000101",
  37708=>"001110010",
  37709=>"001110010",
  37710=>"010000000",
  37711=>"000001001",
  37712=>"111101000",
  37713=>"000111011",
  37714=>"000001010",
  37715=>"111101010",
  37716=>"000100001",
  37717=>"101111011",
  37718=>"100000010",
  37719=>"011100110",
  37720=>"011011011",
  37721=>"010110000",
  37722=>"010111000",
  37723=>"101101110",
  37724=>"011011111",
  37725=>"110011000",
  37726=>"011010001",
  37727=>"110000011",
  37728=>"100011000",
  37729=>"001101011",
  37730=>"110010000",
  37731=>"111001101",
  37732=>"111010101",
  37733=>"110000000",
  37734=>"110101111",
  37735=>"010001001",
  37736=>"000110001",
  37737=>"110100010",
  37738=>"100111001",
  37739=>"001111111",
  37740=>"111001100",
  37741=>"000001001",
  37742=>"101110111",
  37743=>"010001010",
  37744=>"100011010",
  37745=>"101101110",
  37746=>"101000111",
  37747=>"010001101",
  37748=>"000000000",
  37749=>"000110000",
  37750=>"000010011",
  37751=>"100000101",
  37752=>"011010111",
  37753=>"010101100",
  37754=>"000000010",
  37755=>"000000000",
  37756=>"001000010",
  37757=>"111000010",
  37758=>"001110010",
  37759=>"011011101",
  37760=>"001111011",
  37761=>"010110100",
  37762=>"001101000",
  37763=>"101101100",
  37764=>"101101010",
  37765=>"111110000",
  37766=>"001100111",
  37767=>"001100010",
  37768=>"101111111",
  37769=>"000101111",
  37770=>"100111011",
  37771=>"101011001",
  37772=>"000100000",
  37773=>"110011111",
  37774=>"000011110",
  37775=>"101100101",
  37776=>"110010111",
  37777=>"101111111",
  37778=>"000111011",
  37779=>"110011111",
  37780=>"000001010",
  37781=>"100010110",
  37782=>"111101010",
  37783=>"100010100",
  37784=>"000111100",
  37785=>"001001000",
  37786=>"100101111",
  37787=>"001000000",
  37788=>"100001011",
  37789=>"111000000",
  37790=>"001101100",
  37791=>"110110001",
  37792=>"100000000",
  37793=>"011101001",
  37794=>"111111010",
  37795=>"000001111",
  37796=>"010000101",
  37797=>"111101000",
  37798=>"101110001",
  37799=>"110000011",
  37800=>"000001010",
  37801=>"110111111",
  37802=>"011110001",
  37803=>"010111111",
  37804=>"111001000",
  37805=>"101001101",
  37806=>"000001001",
  37807=>"000000000",
  37808=>"101000010",
  37809=>"111111111",
  37810=>"001010100",
  37811=>"100010010",
  37812=>"000111111",
  37813=>"101010011",
  37814=>"011111011",
  37815=>"011011111",
  37816=>"111101011",
  37817=>"001110100",
  37818=>"110111001",
  37819=>"101000010",
  37820=>"110011010",
  37821=>"111000111",
  37822=>"010011110",
  37823=>"101101111",
  37824=>"111110010",
  37825=>"010000100",
  37826=>"010000011",
  37827=>"100011100",
  37828=>"010010110",
  37829=>"011010100",
  37830=>"011100011",
  37831=>"010111001",
  37832=>"010001100",
  37833=>"001100000",
  37834=>"011011111",
  37835=>"111001101",
  37836=>"110011001",
  37837=>"010000010",
  37838=>"100010010",
  37839=>"011000011",
  37840=>"010101010",
  37841=>"111110101",
  37842=>"000010111",
  37843=>"100100100",
  37844=>"000001011",
  37845=>"011000101",
  37846=>"101011101",
  37847=>"111111001",
  37848=>"000100100",
  37849=>"001001111",
  37850=>"001011101",
  37851=>"011010100",
  37852=>"001111010",
  37853=>"111111010",
  37854=>"111010000",
  37855=>"101000001",
  37856=>"001000111",
  37857=>"111110101",
  37858=>"100100111",
  37859=>"111000001",
  37860=>"010000111",
  37861=>"000100001",
  37862=>"010010100",
  37863=>"000100010",
  37864=>"000000000",
  37865=>"101110101",
  37866=>"000110011",
  37867=>"011101101",
  37868=>"010110001",
  37869=>"100100100",
  37870=>"000100000",
  37871=>"111111100",
  37872=>"010011000",
  37873=>"000000101",
  37874=>"001001001",
  37875=>"000000111",
  37876=>"010010011",
  37877=>"110011000",
  37878=>"110111101",
  37879=>"101100010",
  37880=>"100100111",
  37881=>"111010100",
  37882=>"101101000",
  37883=>"100011001",
  37884=>"000010100",
  37885=>"001110001",
  37886=>"001001101",
  37887=>"010000100",
  37888=>"111111001",
  37889=>"000101011",
  37890=>"000111011",
  37891=>"110111010",
  37892=>"001000111",
  37893=>"001010010",
  37894=>"100100111",
  37895=>"101001110",
  37896=>"010010101",
  37897=>"001000010",
  37898=>"110100011",
  37899=>"111110110",
  37900=>"011011101",
  37901=>"101101111",
  37902=>"011010000",
  37903=>"101001111",
  37904=>"101011010",
  37905=>"111001000",
  37906=>"010001001",
  37907=>"000100010",
  37908=>"010001011",
  37909=>"110000110",
  37910=>"001001110",
  37911=>"100000000",
  37912=>"000000101",
  37913=>"110001001",
  37914=>"111010101",
  37915=>"111011001",
  37916=>"110000000",
  37917=>"111110010",
  37918=>"000001001",
  37919=>"111101100",
  37920=>"111000101",
  37921=>"001000111",
  37922=>"101110000",
  37923=>"000001100",
  37924=>"000000011",
  37925=>"010000110",
  37926=>"111011111",
  37927=>"110000101",
  37928=>"000010111",
  37929=>"001011011",
  37930=>"110101101",
  37931=>"000101111",
  37932=>"000000011",
  37933=>"111010111",
  37934=>"011011111",
  37935=>"000110011",
  37936=>"001001101",
  37937=>"110111101",
  37938=>"011011111",
  37939=>"111000000",
  37940=>"011110001",
  37941=>"100111011",
  37942=>"101000010",
  37943=>"010011011",
  37944=>"011010011",
  37945=>"000010001",
  37946=>"000011101",
  37947=>"001100001",
  37948=>"100001101",
  37949=>"001101100",
  37950=>"110000011",
  37951=>"111010100",
  37952=>"011101010",
  37953=>"001100110",
  37954=>"010101001",
  37955=>"101011111",
  37956=>"000000110",
  37957=>"010100101",
  37958=>"010001110",
  37959=>"100110000",
  37960=>"100010000",
  37961=>"100110100",
  37962=>"000101110",
  37963=>"100001101",
  37964=>"110110001",
  37965=>"110001000",
  37966=>"000001100",
  37967=>"011001000",
  37968=>"010100000",
  37969=>"001001100",
  37970=>"100100000",
  37971=>"110100011",
  37972=>"000100010",
  37973=>"001101010",
  37974=>"000110110",
  37975=>"001101011",
  37976=>"111111101",
  37977=>"100110000",
  37978=>"100100001",
  37979=>"111111010",
  37980=>"011100011",
  37981=>"101100101",
  37982=>"011100000",
  37983=>"011111101",
  37984=>"011011000",
  37985=>"011110111",
  37986=>"111110111",
  37987=>"101000111",
  37988=>"000000101",
  37989=>"010100100",
  37990=>"111110001",
  37991=>"010010001",
  37992=>"111101000",
  37993=>"101100100",
  37994=>"100001111",
  37995=>"001011001",
  37996=>"100000100",
  37997=>"101101010",
  37998=>"111001001",
  37999=>"100101100",
  38000=>"010011011",
  38001=>"010011101",
  38002=>"101000010",
  38003=>"011011111",
  38004=>"111110011",
  38005=>"011110110",
  38006=>"110111111",
  38007=>"000001100",
  38008=>"010001100",
  38009=>"000001010",
  38010=>"001011111",
  38011=>"000000000",
  38012=>"001100001",
  38013=>"010100001",
  38014=>"111110000",
  38015=>"011001000",
  38016=>"001010100",
  38017=>"101101111",
  38018=>"111011110",
  38019=>"110101001",
  38020=>"101000100",
  38021=>"001101111",
  38022=>"011001110",
  38023=>"111110111",
  38024=>"100110011",
  38025=>"001111100",
  38026=>"100010011",
  38027=>"000111001",
  38028=>"000011100",
  38029=>"111101011",
  38030=>"010000011",
  38031=>"110001100",
  38032=>"001010101",
  38033=>"011101001",
  38034=>"100010000",
  38035=>"111010100",
  38036=>"001011111",
  38037=>"100010100",
  38038=>"110001111",
  38039=>"001001010",
  38040=>"101010100",
  38041=>"000001000",
  38042=>"011100111",
  38043=>"110011101",
  38044=>"001000110",
  38045=>"100100101",
  38046=>"101011110",
  38047=>"111010011",
  38048=>"001101101",
  38049=>"111110101",
  38050=>"001110110",
  38051=>"010001101",
  38052=>"101011110",
  38053=>"100101101",
  38054=>"000000001",
  38055=>"001000000",
  38056=>"001001111",
  38057=>"110111111",
  38058=>"100001011",
  38059=>"011011100",
  38060=>"101011110",
  38061=>"100100111",
  38062=>"010101101",
  38063=>"101101101",
  38064=>"010010101",
  38065=>"010100110",
  38066=>"111001101",
  38067=>"101010101",
  38068=>"100101001",
  38069=>"011000001",
  38070=>"011001010",
  38071=>"101100010",
  38072=>"101111101",
  38073=>"000001000",
  38074=>"101001100",
  38075=>"000000011",
  38076=>"001010001",
  38077=>"000000101",
  38078=>"101100110",
  38079=>"011100001",
  38080=>"110011011",
  38081=>"011000000",
  38082=>"001011101",
  38083=>"110001000",
  38084=>"100110101",
  38085=>"100101111",
  38086=>"111101101",
  38087=>"110111001",
  38088=>"101011011",
  38089=>"111100101",
  38090=>"000111101",
  38091=>"010000101",
  38092=>"111110001",
  38093=>"100000000",
  38094=>"011001001",
  38095=>"011010000",
  38096=>"101111110",
  38097=>"000001000",
  38098=>"001100111",
  38099=>"101000111",
  38100=>"011011111",
  38101=>"110100000",
  38102=>"001000000",
  38103=>"001111110",
  38104=>"100100111",
  38105=>"010001100",
  38106=>"001001000",
  38107=>"111100100",
  38108=>"010011101",
  38109=>"100000101",
  38110=>"111101000",
  38111=>"100011010",
  38112=>"100001111",
  38113=>"000000111",
  38114=>"100000000",
  38115=>"101011101",
  38116=>"100111101",
  38117=>"001101100",
  38118=>"000000011",
  38119=>"000101110",
  38120=>"011011000",
  38121=>"000011000",
  38122=>"011010111",
  38123=>"000101011",
  38124=>"001000100",
  38125=>"000010001",
  38126=>"110100111",
  38127=>"001101110",
  38128=>"110011001",
  38129=>"001011001",
  38130=>"100111000",
  38131=>"100101101",
  38132=>"111100011",
  38133=>"100101000",
  38134=>"111001010",
  38135=>"011111101",
  38136=>"000000011",
  38137=>"101111100",
  38138=>"000100001",
  38139=>"010101001",
  38140=>"101101101",
  38141=>"011110110",
  38142=>"111111111",
  38143=>"001110111",
  38144=>"001010011",
  38145=>"100010110",
  38146=>"111000010",
  38147=>"011101110",
  38148=>"111011001",
  38149=>"010100010",
  38150=>"001110110",
  38151=>"000001111",
  38152=>"101111000",
  38153=>"010000110",
  38154=>"001011011",
  38155=>"110101001",
  38156=>"100101111",
  38157=>"011011010",
  38158=>"101010101",
  38159=>"011010000",
  38160=>"001011010",
  38161=>"010110100",
  38162=>"101100111",
  38163=>"100010011",
  38164=>"100110000",
  38165=>"110111111",
  38166=>"001110111",
  38167=>"010000101",
  38168=>"110101001",
  38169=>"110110110",
  38170=>"111111011",
  38171=>"000001000",
  38172=>"011110110",
  38173=>"011001100",
  38174=>"101111110",
  38175=>"101101101",
  38176=>"010010000",
  38177=>"011001010",
  38178=>"100100010",
  38179=>"010110100",
  38180=>"100010110",
  38181=>"101110100",
  38182=>"011011110",
  38183=>"011111110",
  38184=>"110000100",
  38185=>"101001010",
  38186=>"110101111",
  38187=>"111100011",
  38188=>"011000010",
  38189=>"111000110",
  38190=>"011000111",
  38191=>"010001000",
  38192=>"010100011",
  38193=>"111111000",
  38194=>"101011011",
  38195=>"010001010",
  38196=>"000000100",
  38197=>"000001001",
  38198=>"100010111",
  38199=>"010100101",
  38200=>"001001111",
  38201=>"100100011",
  38202=>"010001111",
  38203=>"000100111",
  38204=>"101000010",
  38205=>"101111001",
  38206=>"111110011",
  38207=>"111111110",
  38208=>"001100010",
  38209=>"000001110",
  38210=>"000110110",
  38211=>"001011001",
  38212=>"000111111",
  38213=>"111010011",
  38214=>"101001010",
  38215=>"111100100",
  38216=>"010011110",
  38217=>"100110101",
  38218=>"001001111",
  38219=>"000010011",
  38220=>"011111110",
  38221=>"000010110",
  38222=>"010010001",
  38223=>"011111010",
  38224=>"011110010",
  38225=>"100111110",
  38226=>"011010110",
  38227=>"000100111",
  38228=>"101001010",
  38229=>"011101001",
  38230=>"100110111",
  38231=>"100101101",
  38232=>"011010011",
  38233=>"111010011",
  38234=>"100001101",
  38235=>"000001111",
  38236=>"000110001",
  38237=>"010001110",
  38238=>"010010001",
  38239=>"000010100",
  38240=>"111110011",
  38241=>"010000101",
  38242=>"000101111",
  38243=>"101000111",
  38244=>"001100010",
  38245=>"001011011",
  38246=>"000111101",
  38247=>"101101000",
  38248=>"101010110",
  38249=>"101101001",
  38250=>"110100010",
  38251=>"001011010",
  38252=>"000000010",
  38253=>"100110111",
  38254=>"100011001",
  38255=>"000111101",
  38256=>"001001011",
  38257=>"110100010",
  38258=>"110010000",
  38259=>"100101110",
  38260=>"110010110",
  38261=>"011011101",
  38262=>"100100011",
  38263=>"100100110",
  38264=>"111110100",
  38265=>"010010011",
  38266=>"110011110",
  38267=>"101100011",
  38268=>"101100100",
  38269=>"011100011",
  38270=>"000001111",
  38271=>"101101111",
  38272=>"010010100",
  38273=>"000110011",
  38274=>"100111001",
  38275=>"001000010",
  38276=>"001101000",
  38277=>"101000001",
  38278=>"010110111",
  38279=>"100100001",
  38280=>"000010111",
  38281=>"011111111",
  38282=>"010010001",
  38283=>"010011010",
  38284=>"110111000",
  38285=>"011011111",
  38286=>"001001001",
  38287=>"100000100",
  38288=>"111010000",
  38289=>"001001100",
  38290=>"010001111",
  38291=>"011011111",
  38292=>"001100101",
  38293=>"011001100",
  38294=>"000100101",
  38295=>"101001000",
  38296=>"010100101",
  38297=>"001001000",
  38298=>"001001110",
  38299=>"111001011",
  38300=>"101011011",
  38301=>"000100011",
  38302=>"100000000",
  38303=>"110110111",
  38304=>"101101100",
  38305=>"000101011",
  38306=>"010100111",
  38307=>"001011100",
  38308=>"110011000",
  38309=>"111110111",
  38310=>"011001011",
  38311=>"111000111",
  38312=>"010000000",
  38313=>"100001010",
  38314=>"001001101",
  38315=>"110010001",
  38316=>"011110110",
  38317=>"000011000",
  38318=>"001000101",
  38319=>"100101110",
  38320=>"101000111",
  38321=>"010101011",
  38322=>"010011010",
  38323=>"001111100",
  38324=>"001001000",
  38325=>"001010010",
  38326=>"111111111",
  38327=>"011010010",
  38328=>"001110001",
  38329=>"100100000",
  38330=>"111101000",
  38331=>"010111111",
  38332=>"110000110",
  38333=>"010010000",
  38334=>"110000111",
  38335=>"010111110",
  38336=>"111111001",
  38337=>"010011111",
  38338=>"111101101",
  38339=>"111010010",
  38340=>"010111001",
  38341=>"000010000",
  38342=>"000000000",
  38343=>"110101011",
  38344=>"010110010",
  38345=>"011100001",
  38346=>"000000001",
  38347=>"011010010",
  38348=>"010101000",
  38349=>"000001000",
  38350=>"010001111",
  38351=>"001011000",
  38352=>"010100010",
  38353=>"010000110",
  38354=>"011111011",
  38355=>"010001110",
  38356=>"110110101",
  38357=>"011100111",
  38358=>"101100110",
  38359=>"101101101",
  38360=>"101011001",
  38361=>"100011101",
  38362=>"001111001",
  38363=>"010111100",
  38364=>"100001100",
  38365=>"001101010",
  38366=>"000001001",
  38367=>"011100110",
  38368=>"000101100",
  38369=>"111111110",
  38370=>"110001100",
  38371=>"011000101",
  38372=>"111100100",
  38373=>"010111101",
  38374=>"100000001",
  38375=>"011101100",
  38376=>"000110100",
  38377=>"000101001",
  38378=>"000011110",
  38379=>"101111001",
  38380=>"001100001",
  38381=>"110000000",
  38382=>"000111001",
  38383=>"011100111",
  38384=>"110001110",
  38385=>"011101101",
  38386=>"110011001",
  38387=>"011110100",
  38388=>"110110011",
  38389=>"100001111",
  38390=>"010001111",
  38391=>"011100010",
  38392=>"111010001",
  38393=>"000110001",
  38394=>"000101000",
  38395=>"101101101",
  38396=>"000010111",
  38397=>"110010010",
  38398=>"010000010",
  38399=>"011110011",
  38400=>"011011010",
  38401=>"001111011",
  38402=>"001000000",
  38403=>"001000001",
  38404=>"101101001",
  38405=>"010101101",
  38406=>"110011000",
  38407=>"111111011",
  38408=>"111101000",
  38409=>"110101101",
  38410=>"110101110",
  38411=>"001111101",
  38412=>"101101111",
  38413=>"010101010",
  38414=>"101110100",
  38415=>"111100100",
  38416=>"001001001",
  38417=>"001010010",
  38418=>"011101011",
  38419=>"001011010",
  38420=>"001001101",
  38421=>"010010010",
  38422=>"010100011",
  38423=>"000101011",
  38424=>"100011101",
  38425=>"100000001",
  38426=>"011001010",
  38427=>"111001110",
  38428=>"111110111",
  38429=>"000111101",
  38430=>"011100111",
  38431=>"011000110",
  38432=>"011000010",
  38433=>"011110111",
  38434=>"000101111",
  38435=>"101101101",
  38436=>"011010111",
  38437=>"110100101",
  38438=>"110011000",
  38439=>"100000101",
  38440=>"110110000",
  38441=>"111000001",
  38442=>"010001110",
  38443=>"100100000",
  38444=>"001110010",
  38445=>"101010101",
  38446=>"010001000",
  38447=>"100110000",
  38448=>"100110100",
  38449=>"010000001",
  38450=>"000101101",
  38451=>"111100101",
  38452=>"001101000",
  38453=>"010011101",
  38454=>"001001001",
  38455=>"010010011",
  38456=>"110110010",
  38457=>"100010001",
  38458=>"101101011",
  38459=>"110001000",
  38460=>"100011101",
  38461=>"011101110",
  38462=>"011101011",
  38463=>"100000100",
  38464=>"010111011",
  38465=>"011101100",
  38466=>"000011111",
  38467=>"100010000",
  38468=>"011101101",
  38469=>"111100001",
  38470=>"101111011",
  38471=>"000110111",
  38472=>"000110111",
  38473=>"010011110",
  38474=>"001011000",
  38475=>"111011111",
  38476=>"000010010",
  38477=>"000100000",
  38478=>"000011000",
  38479=>"110101001",
  38480=>"010101111",
  38481=>"000000010",
  38482=>"010111000",
  38483=>"101010000",
  38484=>"000000011",
  38485=>"000111001",
  38486=>"001100011",
  38487=>"000110010",
  38488=>"011100001",
  38489=>"101000001",
  38490=>"001101001",
  38491=>"110110111",
  38492=>"010010001",
  38493=>"100101000",
  38494=>"001101001",
  38495=>"001110110",
  38496=>"101111100",
  38497=>"111110001",
  38498=>"000010101",
  38499=>"001100011",
  38500=>"010100011",
  38501=>"110110011",
  38502=>"000010000",
  38503=>"000111000",
  38504=>"110110101",
  38505=>"000101010",
  38506=>"010110011",
  38507=>"100111100",
  38508=>"001111010",
  38509=>"110001101",
  38510=>"001001001",
  38511=>"100111100",
  38512=>"101001111",
  38513=>"111000110",
  38514=>"000100001",
  38515=>"100001000",
  38516=>"101011011",
  38517=>"001101001",
  38518=>"101111101",
  38519=>"100110100",
  38520=>"010001111",
  38521=>"111101111",
  38522=>"111100101",
  38523=>"011100100",
  38524=>"101001000",
  38525=>"000011010",
  38526=>"001000100",
  38527=>"111111100",
  38528=>"001000100",
  38529=>"111110011",
  38530=>"001011100",
  38531=>"100010111",
  38532=>"010111100",
  38533=>"100100001",
  38534=>"011111011",
  38535=>"111100011",
  38536=>"011110000",
  38537=>"000010000",
  38538=>"001000011",
  38539=>"110110111",
  38540=>"100011010",
  38541=>"110100101",
  38542=>"011110010",
  38543=>"001001000",
  38544=>"010111101",
  38545=>"011000011",
  38546=>"100111101",
  38547=>"100111000",
  38548=>"101101001",
  38549=>"111110011",
  38550=>"101110111",
  38551=>"110000001",
  38552=>"001101111",
  38553=>"100001010",
  38554=>"110011110",
  38555=>"000100110",
  38556=>"101001111",
  38557=>"011101110",
  38558=>"001010111",
  38559=>"011101011",
  38560=>"111010101",
  38561=>"010101110",
  38562=>"011111110",
  38563=>"011001000",
  38564=>"101001001",
  38565=>"001010010",
  38566=>"101100111",
  38567=>"001001001",
  38568=>"010110100",
  38569=>"101000101",
  38570=>"010101000",
  38571=>"110111010",
  38572=>"111111100",
  38573=>"000110001",
  38574=>"111111000",
  38575=>"011000001",
  38576=>"010000111",
  38577=>"100110001",
  38578=>"110011000",
  38579=>"011011011",
  38580=>"001101111",
  38581=>"010101001",
  38582=>"101010110",
  38583=>"101110001",
  38584=>"011101101",
  38585=>"100001100",
  38586=>"000010001",
  38587=>"111011111",
  38588=>"101100100",
  38589=>"001011010",
  38590=>"101001011",
  38591=>"110101010",
  38592=>"110010101",
  38593=>"010111011",
  38594=>"010100001",
  38595=>"011000000",
  38596=>"100000001",
  38597=>"001001000",
  38598=>"010110000",
  38599=>"100100001",
  38600=>"100000011",
  38601=>"110001001",
  38602=>"001111100",
  38603=>"010101101",
  38604=>"001001001",
  38605=>"011110110",
  38606=>"011011110",
  38607=>"010111111",
  38608=>"001100110",
  38609=>"001001010",
  38610=>"101000000",
  38611=>"011010010",
  38612=>"010111101",
  38613=>"001001000",
  38614=>"000000001",
  38615=>"001101110",
  38616=>"000101011",
  38617=>"110110110",
  38618=>"101000000",
  38619=>"000111110",
  38620=>"101101101",
  38621=>"001000011",
  38622=>"000110110",
  38623=>"111010000",
  38624=>"011000111",
  38625=>"001010000",
  38626=>"110100111",
  38627=>"010010101",
  38628=>"001111110",
  38629=>"100010111",
  38630=>"100100010",
  38631=>"110110110",
  38632=>"101101001",
  38633=>"001011001",
  38634=>"111110100",
  38635=>"001000011",
  38636=>"001101011",
  38637=>"111101000",
  38638=>"111110100",
  38639=>"101100101",
  38640=>"100000101",
  38641=>"000100010",
  38642=>"000001010",
  38643=>"000000011",
  38644=>"011111011",
  38645=>"100111001",
  38646=>"001000001",
  38647=>"101000000",
  38648=>"111001100",
  38649=>"010111001",
  38650=>"001100111",
  38651=>"101110100",
  38652=>"010001111",
  38653=>"011010100",
  38654=>"101010010",
  38655=>"000100000",
  38656=>"100110011",
  38657=>"010010100",
  38658=>"111111000",
  38659=>"001000111",
  38660=>"101010110",
  38661=>"101011111",
  38662=>"110000101",
  38663=>"011110111",
  38664=>"000101101",
  38665=>"100100101",
  38666=>"000000100",
  38667=>"110101001",
  38668=>"101000100",
  38669=>"110001111",
  38670=>"010110110",
  38671=>"010111100",
  38672=>"000100000",
  38673=>"101110100",
  38674=>"110111011",
  38675=>"001000110",
  38676=>"001011011",
  38677=>"100001001",
  38678=>"011110000",
  38679=>"100100100",
  38680=>"001000111",
  38681=>"100001001",
  38682=>"111110001",
  38683=>"111111001",
  38684=>"001101000",
  38685=>"110001011",
  38686=>"110000010",
  38687=>"010111000",
  38688=>"000001001",
  38689=>"101011101",
  38690=>"001000000",
  38691=>"111111101",
  38692=>"111010111",
  38693=>"001000001",
  38694=>"101010100",
  38695=>"011101110",
  38696=>"110101001",
  38697=>"110010101",
  38698=>"010000101",
  38699=>"110011001",
  38700=>"110100001",
  38701=>"101001111",
  38702=>"001101010",
  38703=>"111000000",
  38704=>"001111100",
  38705=>"111100100",
  38706=>"101001101",
  38707=>"110010101",
  38708=>"110111000",
  38709=>"100111111",
  38710=>"000100001",
  38711=>"111101101",
  38712=>"100100010",
  38713=>"011101001",
  38714=>"110000110",
  38715=>"000001011",
  38716=>"111111110",
  38717=>"000100111",
  38718=>"100111011",
  38719=>"110110100",
  38720=>"000000101",
  38721=>"110001010",
  38722=>"100000111",
  38723=>"010110101",
  38724=>"001100010",
  38725=>"000110101",
  38726=>"101100001",
  38727=>"000101001",
  38728=>"100011011",
  38729=>"100010001",
  38730=>"000011010",
  38731=>"100101001",
  38732=>"001001000",
  38733=>"111110000",
  38734=>"110101001",
  38735=>"011110000",
  38736=>"001000000",
  38737=>"100001010",
  38738=>"101000101",
  38739=>"011011100",
  38740=>"010001000",
  38741=>"011001100",
  38742=>"101100111",
  38743=>"100110010",
  38744=>"000100000",
  38745=>"001000111",
  38746=>"011100001",
  38747=>"011101001",
  38748=>"000110010",
  38749=>"110111110",
  38750=>"100100000",
  38751=>"000100011",
  38752=>"000110010",
  38753=>"100101011",
  38754=>"001110110",
  38755=>"101001011",
  38756=>"100111011",
  38757=>"101110111",
  38758=>"100001111",
  38759=>"111001111",
  38760=>"000101000",
  38761=>"111110110",
  38762=>"010101110",
  38763=>"001101000",
  38764=>"010100101",
  38765=>"100101111",
  38766=>"100101011",
  38767=>"000011110",
  38768=>"101001101",
  38769=>"001011001",
  38770=>"011000011",
  38771=>"101111101",
  38772=>"100111011",
  38773=>"110101100",
  38774=>"110100000",
  38775=>"100101111",
  38776=>"010011110",
  38777=>"001100100",
  38778=>"001000100",
  38779=>"001101011",
  38780=>"000111000",
  38781=>"101100001",
  38782=>"111001100",
  38783=>"101010111",
  38784=>"001110111",
  38785=>"101001001",
  38786=>"000010010",
  38787=>"001011111",
  38788=>"101000010",
  38789=>"001101010",
  38790=>"011101101",
  38791=>"111010000",
  38792=>"010111011",
  38793=>"110100100",
  38794=>"111111101",
  38795=>"101000011",
  38796=>"001101110",
  38797=>"110010001",
  38798=>"111011110",
  38799=>"100010100",
  38800=>"100101000",
  38801=>"011000100",
  38802=>"100011001",
  38803=>"111000000",
  38804=>"011010010",
  38805=>"111011001",
  38806=>"011100110",
  38807=>"100010001",
  38808=>"111111011",
  38809=>"100010001",
  38810=>"101100111",
  38811=>"010001001",
  38812=>"100111010",
  38813=>"011010100",
  38814=>"011010001",
  38815=>"001111001",
  38816=>"101011011",
  38817=>"011100100",
  38818=>"100110111",
  38819=>"010111101",
  38820=>"000110000",
  38821=>"111010011",
  38822=>"101111100",
  38823=>"100011101",
  38824=>"111011011",
  38825=>"000011111",
  38826=>"001011010",
  38827=>"001001100",
  38828=>"110010110",
  38829=>"101111001",
  38830=>"000101011",
  38831=>"000100101",
  38832=>"001000001",
  38833=>"011100011",
  38834=>"011110110",
  38835=>"011011100",
  38836=>"110011010",
  38837=>"110111010",
  38838=>"000110000",
  38839=>"111111000",
  38840=>"001011000",
  38841=>"100000100",
  38842=>"000101000",
  38843=>"001100001",
  38844=>"110011100",
  38845=>"010110100",
  38846=>"100001100",
  38847=>"101001000",
  38848=>"110100100",
  38849=>"011110011",
  38850=>"010001100",
  38851=>"011101101",
  38852=>"100001100",
  38853=>"100001000",
  38854=>"101001111",
  38855=>"000000001",
  38856=>"101110000",
  38857=>"000110111",
  38858=>"100100111",
  38859=>"001111011",
  38860=>"010011000",
  38861=>"111010110",
  38862=>"110010001",
  38863=>"010001001",
  38864=>"010000011",
  38865=>"011110110",
  38866=>"011100001",
  38867=>"010100101",
  38868=>"100110110",
  38869=>"111011101",
  38870=>"111010000",
  38871=>"110111101",
  38872=>"000001010",
  38873=>"111101010",
  38874=>"110100010",
  38875=>"011110001",
  38876=>"001111111",
  38877=>"110101011",
  38878=>"101111000",
  38879=>"011011101",
  38880=>"100010000",
  38881=>"100101001",
  38882=>"100110011",
  38883=>"011100111",
  38884=>"011011111",
  38885=>"000010010",
  38886=>"000001000",
  38887=>"101000011",
  38888=>"101100100",
  38889=>"011010011",
  38890=>"010110011",
  38891=>"111011000",
  38892=>"101111011",
  38893=>"000000011",
  38894=>"110010101",
  38895=>"100110001",
  38896=>"101001111",
  38897=>"101010110",
  38898=>"110001100",
  38899=>"100011101",
  38900=>"110111101",
  38901=>"011110101",
  38902=>"110100110",
  38903=>"110000110",
  38904=>"110010111",
  38905=>"101011101",
  38906=>"001111100",
  38907=>"001111111",
  38908=>"101110101",
  38909=>"000010000",
  38910=>"100101111",
  38911=>"001000001",
  38912=>"110101100",
  38913=>"000000001",
  38914=>"110100111",
  38915=>"101101001",
  38916=>"110001010",
  38917=>"110100100",
  38918=>"000011100",
  38919=>"110010110",
  38920=>"110110001",
  38921=>"101001001",
  38922=>"101000101",
  38923=>"100010010",
  38924=>"110000111",
  38925=>"110101011",
  38926=>"100011101",
  38927=>"110000000",
  38928=>"101101111",
  38929=>"110001000",
  38930=>"111111111",
  38931=>"100000010",
  38932=>"011100111",
  38933=>"010111101",
  38934=>"110111101",
  38935=>"101010111",
  38936=>"110000011",
  38937=>"000000111",
  38938=>"100001000",
  38939=>"101111111",
  38940=>"000101011",
  38941=>"000011001",
  38942=>"011011000",
  38943=>"100100001",
  38944=>"100100010",
  38945=>"101000010",
  38946=>"100000000",
  38947=>"101000111",
  38948=>"011010011",
  38949=>"101100001",
  38950=>"111110111",
  38951=>"101010101",
  38952=>"101001011",
  38953=>"100111100",
  38954=>"110011101",
  38955=>"011100111",
  38956=>"111110110",
  38957=>"100101011",
  38958=>"101000011",
  38959=>"010000001",
  38960=>"101010010",
  38961=>"011101111",
  38962=>"101010110",
  38963=>"010101110",
  38964=>"100101000",
  38965=>"010010000",
  38966=>"000000001",
  38967=>"110011011",
  38968=>"000011111",
  38969=>"101000010",
  38970=>"101101001",
  38971=>"100000110",
  38972=>"110000011",
  38973=>"111111101",
  38974=>"100000111",
  38975=>"001000001",
  38976=>"110100001",
  38977=>"001010000",
  38978=>"110000011",
  38979=>"010000100",
  38980=>"101011011",
  38981=>"011100011",
  38982=>"111000111",
  38983=>"000101000",
  38984=>"001011100",
  38985=>"011001010",
  38986=>"011010100",
  38987=>"011101011",
  38988=>"010111110",
  38989=>"011001000",
  38990=>"011011000",
  38991=>"101001011",
  38992=>"101110111",
  38993=>"101100110",
  38994=>"100010011",
  38995=>"011110011",
  38996=>"100111110",
  38997=>"111110011",
  38998=>"111011100",
  38999=>"001100100",
  39000=>"010101110",
  39001=>"100011110",
  39002=>"011010011",
  39003=>"001110100",
  39004=>"010000011",
  39005=>"101011110",
  39006=>"110110000",
  39007=>"001111010",
  39008=>"101010010",
  39009=>"111000011",
  39010=>"100110100",
  39011=>"000000010",
  39012=>"010011010",
  39013=>"110110111",
  39014=>"000011101",
  39015=>"100010010",
  39016=>"001001110",
  39017=>"111111101",
  39018=>"000111001",
  39019=>"100110111",
  39020=>"110010101",
  39021=>"110010110",
  39022=>"100011010",
  39023=>"100001000",
  39024=>"100110000",
  39025=>"011100010",
  39026=>"000011001",
  39027=>"000010111",
  39028=>"111001000",
  39029=>"010010110",
  39030=>"011010000",
  39031=>"001001000",
  39032=>"000100100",
  39033=>"111111010",
  39034=>"101111111",
  39035=>"011110011",
  39036=>"000010010",
  39037=>"110000101",
  39038=>"110000010",
  39039=>"011101101",
  39040=>"011001001",
  39041=>"100011100",
  39042=>"000001101",
  39043=>"100011100",
  39044=>"010000010",
  39045=>"000011010",
  39046=>"010111101",
  39047=>"110100001",
  39048=>"100001010",
  39049=>"000010101",
  39050=>"101110100",
  39051=>"100001001",
  39052=>"000101110",
  39053=>"111101010",
  39054=>"111010010",
  39055=>"111110001",
  39056=>"000101010",
  39057=>"010111100",
  39058=>"000100010",
  39059=>"001101011",
  39060=>"000010010",
  39061=>"000011111",
  39062=>"101011100",
  39063=>"001110010",
  39064=>"001000101",
  39065=>"110011010",
  39066=>"100100101",
  39067=>"000010100",
  39068=>"011000010",
  39069=>"110010101",
  39070=>"100001100",
  39071=>"000000011",
  39072=>"111010000",
  39073=>"010010101",
  39074=>"000100010",
  39075=>"000001101",
  39076=>"101111101",
  39077=>"101001110",
  39078=>"110000000",
  39079=>"110011110",
  39080=>"100111101",
  39081=>"101110100",
  39082=>"010000111",
  39083=>"111101010",
  39084=>"111001001",
  39085=>"110110111",
  39086=>"100101001",
  39087=>"101001010",
  39088=>"111000101",
  39089=>"111100101",
  39090=>"101010000",
  39091=>"101100010",
  39092=>"110011100",
  39093=>"110011111",
  39094=>"111001001",
  39095=>"101110111",
  39096=>"110000000",
  39097=>"000101000",
  39098=>"100101011",
  39099=>"011110111",
  39100=>"101100010",
  39101=>"011011001",
  39102=>"001110000",
  39103=>"111000001",
  39104=>"000100011",
  39105=>"000011111",
  39106=>"000111011",
  39107=>"010100011",
  39108=>"011001001",
  39109=>"010100101",
  39110=>"111100101",
  39111=>"011110110",
  39112=>"100000100",
  39113=>"111101000",
  39114=>"110011110",
  39115=>"000010111",
  39116=>"001111010",
  39117=>"010011101",
  39118=>"000000010",
  39119=>"111110000",
  39120=>"111111111",
  39121=>"100110010",
  39122=>"100101001",
  39123=>"101000011",
  39124=>"111101111",
  39125=>"101010100",
  39126=>"111010010",
  39127=>"110011100",
  39128=>"100110000",
  39129=>"100110111",
  39130=>"011001111",
  39131=>"101101111",
  39132=>"010000101",
  39133=>"111101000",
  39134=>"101000000",
  39135=>"011111000",
  39136=>"000100010",
  39137=>"011010111",
  39138=>"000001111",
  39139=>"100110001",
  39140=>"111001001",
  39141=>"001001010",
  39142=>"010101100",
  39143=>"010001010",
  39144=>"110001100",
  39145=>"011110011",
  39146=>"010101110",
  39147=>"001111111",
  39148=>"100011101",
  39149=>"010010000",
  39150=>"100111101",
  39151=>"001001000",
  39152=>"001110100",
  39153=>"101101101",
  39154=>"011000100",
  39155=>"001100100",
  39156=>"110010000",
  39157=>"111100001",
  39158=>"011101100",
  39159=>"110010001",
  39160=>"001101011",
  39161=>"110100111",
  39162=>"101001100",
  39163=>"100010011",
  39164=>"100110110",
  39165=>"011110111",
  39166=>"001111100",
  39167=>"100001110",
  39168=>"010101111",
  39169=>"110010101",
  39170=>"001110100",
  39171=>"110100000",
  39172=>"010111111",
  39173=>"100111101",
  39174=>"011100000",
  39175=>"001101110",
  39176=>"000001110",
  39177=>"001000101",
  39178=>"001000111",
  39179=>"011100110",
  39180=>"000010111",
  39181=>"001111100",
  39182=>"110011100",
  39183=>"100011010",
  39184=>"010110110",
  39185=>"100101010",
  39186=>"001001100",
  39187=>"101011011",
  39188=>"100110101",
  39189=>"110110010",
  39190=>"111110110",
  39191=>"001110011",
  39192=>"110010001",
  39193=>"000100101",
  39194=>"110001101",
  39195=>"010000100",
  39196=>"101001110",
  39197=>"110000110",
  39198=>"111010110",
  39199=>"101000000",
  39200=>"100111100",
  39201=>"101011011",
  39202=>"110111110",
  39203=>"100011000",
  39204=>"010110110",
  39205=>"010001100",
  39206=>"111110001",
  39207=>"100111011",
  39208=>"100100110",
  39209=>"110110110",
  39210=>"010101001",
  39211=>"010000100",
  39212=>"101000001",
  39213=>"100101100",
  39214=>"100000001",
  39215=>"110001101",
  39216=>"011100000",
  39217=>"110110010",
  39218=>"010000011",
  39219=>"010010010",
  39220=>"011001000",
  39221=>"100001001",
  39222=>"111101100",
  39223=>"001101111",
  39224=>"000101101",
  39225=>"100111110",
  39226=>"110110000",
  39227=>"011110011",
  39228=>"001101011",
  39229=>"010011000",
  39230=>"011010010",
  39231=>"001001101",
  39232=>"101111111",
  39233=>"010010000",
  39234=>"100100010",
  39235=>"010000101",
  39236=>"111110000",
  39237=>"001001010",
  39238=>"100101001",
  39239=>"110011001",
  39240=>"100110101",
  39241=>"011100111",
  39242=>"011001010",
  39243=>"110111111",
  39244=>"001111001",
  39245=>"100000001",
  39246=>"111011000",
  39247=>"001101100",
  39248=>"010001110",
  39249=>"101100001",
  39250=>"111000100",
  39251=>"111100111",
  39252=>"001101010",
  39253=>"001110101",
  39254=>"011101000",
  39255=>"111101011",
  39256=>"010001101",
  39257=>"001101011",
  39258=>"000010100",
  39259=>"110010100",
  39260=>"000100001",
  39261=>"110100101",
  39262=>"110001001",
  39263=>"010010101",
  39264=>"010101011",
  39265=>"000011100",
  39266=>"000010000",
  39267=>"110100100",
  39268=>"101100110",
  39269=>"100111000",
  39270=>"110110000",
  39271=>"010000011",
  39272=>"110101100",
  39273=>"000010110",
  39274=>"111111011",
  39275=>"101010101",
  39276=>"011111101",
  39277=>"000001100",
  39278=>"000010000",
  39279=>"011100110",
  39280=>"000000010",
  39281=>"001011001",
  39282=>"111001011",
  39283=>"100111000",
  39284=>"110100110",
  39285=>"001000000",
  39286=>"111101001",
  39287=>"111010011",
  39288=>"001011111",
  39289=>"010111001",
  39290=>"011110110",
  39291=>"100111000",
  39292=>"100110001",
  39293=>"110101101",
  39294=>"011111111",
  39295=>"111011000",
  39296=>"111011100",
  39297=>"000110000",
  39298=>"101001100",
  39299=>"101111010",
  39300=>"001010110",
  39301=>"000011101",
  39302=>"000110111",
  39303=>"011000001",
  39304=>"101101000",
  39305=>"001011001",
  39306=>"010010000",
  39307=>"011011101",
  39308=>"000110011",
  39309=>"000110000",
  39310=>"101110111",
  39311=>"011010011",
  39312=>"001001100",
  39313=>"110001110",
  39314=>"110110011",
  39315=>"101001010",
  39316=>"111010110",
  39317=>"000111010",
  39318=>"010010111",
  39319=>"101110001",
  39320=>"110110100",
  39321=>"010110111",
  39322=>"011001100",
  39323=>"011010101",
  39324=>"010100111",
  39325=>"011111010",
  39326=>"111110001",
  39327=>"011001110",
  39328=>"111110000",
  39329=>"011011001",
  39330=>"100001101",
  39331=>"011001000",
  39332=>"100011111",
  39333=>"001010101",
  39334=>"011011000",
  39335=>"110001000",
  39336=>"001011001",
  39337=>"011100100",
  39338=>"000100011",
  39339=>"100000000",
  39340=>"000110110",
  39341=>"001110010",
  39342=>"011111110",
  39343=>"011100110",
  39344=>"111011111",
  39345=>"111000011",
  39346=>"111001011",
  39347=>"001000100",
  39348=>"110111011",
  39349=>"011111001",
  39350=>"000111111",
  39351=>"111111101",
  39352=>"101111001",
  39353=>"001110001",
  39354=>"101011000",
  39355=>"010111111",
  39356=>"101101000",
  39357=>"011100011",
  39358=>"111101010",
  39359=>"000100000",
  39360=>"011110001",
  39361=>"010100000",
  39362=>"011000010",
  39363=>"111001011",
  39364=>"011011000",
  39365=>"011101101",
  39366=>"111100010",
  39367=>"010100100",
  39368=>"111101111",
  39369=>"000011110",
  39370=>"001101101",
  39371=>"100011100",
  39372=>"001010010",
  39373=>"011011010",
  39374=>"100110111",
  39375=>"110100101",
  39376=>"111110110",
  39377=>"001010111",
  39378=>"001010011",
  39379=>"100111110",
  39380=>"000110001",
  39381=>"010000001",
  39382=>"100001101",
  39383=>"000010001",
  39384=>"011011001",
  39385=>"000001111",
  39386=>"101000000",
  39387=>"000001111",
  39388=>"100111101",
  39389=>"001001101",
  39390=>"000010100",
  39391=>"100110000",
  39392=>"100101001",
  39393=>"100111001",
  39394=>"101001000",
  39395=>"001101110",
  39396=>"001001100",
  39397=>"011111111",
  39398=>"011001010",
  39399=>"001010110",
  39400=>"111010001",
  39401=>"010110100",
  39402=>"000011110",
  39403=>"110001101",
  39404=>"100100100",
  39405=>"110001011",
  39406=>"100000111",
  39407=>"000100110",
  39408=>"001000001",
  39409=>"011110010",
  39410=>"101010001",
  39411=>"110011101",
  39412=>"111100010",
  39413=>"000110111",
  39414=>"100010110",
  39415=>"101001011",
  39416=>"100011000",
  39417=>"010010001",
  39418=>"101011010",
  39419=>"100010111",
  39420=>"000101111",
  39421=>"011010101",
  39422=>"001101011",
  39423=>"001011011",
  39424=>"011110010",
  39425=>"100001011",
  39426=>"110001011",
  39427=>"111100110",
  39428=>"101000110",
  39429=>"010110010",
  39430=>"111111011",
  39431=>"011010000",
  39432=>"111001001",
  39433=>"001101110",
  39434=>"110110000",
  39435=>"010100000",
  39436=>"100110111",
  39437=>"001101110",
  39438=>"101110011",
  39439=>"000100111",
  39440=>"010100111",
  39441=>"010111111",
  39442=>"000000010",
  39443=>"010011011",
  39444=>"001100010",
  39445=>"010100110",
  39446=>"110000000",
  39447=>"111111011",
  39448=>"111011001",
  39449=>"000100000",
  39450=>"001000101",
  39451=>"010000101",
  39452=>"000110000",
  39453=>"001110010",
  39454=>"101010110",
  39455=>"101110110",
  39456=>"001100011",
  39457=>"000111001",
  39458=>"011000000",
  39459=>"111001110",
  39460=>"110100011",
  39461=>"101101010",
  39462=>"000000000",
  39463=>"100100110",
  39464=>"010010101",
  39465=>"001111000",
  39466=>"000101011",
  39467=>"110000000",
  39468=>"110100001",
  39469=>"000010110",
  39470=>"000110010",
  39471=>"100100011",
  39472=>"001000000",
  39473=>"000100110",
  39474=>"000010001",
  39475=>"100001010",
  39476=>"011101010",
  39477=>"010010011",
  39478=>"000111001",
  39479=>"010101000",
  39480=>"000011000",
  39481=>"010011111",
  39482=>"111001111",
  39483=>"101001001",
  39484=>"001001111",
  39485=>"110010000",
  39486=>"010000010",
  39487=>"011110100",
  39488=>"111110110",
  39489=>"110001010",
  39490=>"111111001",
  39491=>"101100001",
  39492=>"110010000",
  39493=>"010100011",
  39494=>"100010001",
  39495=>"101001110",
  39496=>"110011101",
  39497=>"111111001",
  39498=>"110001111",
  39499=>"100100111",
  39500=>"010010001",
  39501=>"101100101",
  39502=>"101111111",
  39503=>"001000011",
  39504=>"010011111",
  39505=>"001010101",
  39506=>"111111111",
  39507=>"100000001",
  39508=>"000111101",
  39509=>"100101010",
  39510=>"001111000",
  39511=>"101100010",
  39512=>"110111111",
  39513=>"010111011",
  39514=>"000000000",
  39515=>"000001100",
  39516=>"100010101",
  39517=>"101010001",
  39518=>"000100010",
  39519=>"011100101",
  39520=>"100101101",
  39521=>"111101001",
  39522=>"000000100",
  39523=>"111110100",
  39524=>"000100110",
  39525=>"010011111",
  39526=>"101111000",
  39527=>"100010111",
  39528=>"110001101",
  39529=>"010000000",
  39530=>"011111101",
  39531=>"100010000",
  39532=>"010100111",
  39533=>"011010101",
  39534=>"110010000",
  39535=>"001101111",
  39536=>"110000101",
  39537=>"000111001",
  39538=>"101010110",
  39539=>"010000110",
  39540=>"101101101",
  39541=>"100000000",
  39542=>"101110111",
  39543=>"100110101",
  39544=>"000110101",
  39545=>"110101010",
  39546=>"101011001",
  39547=>"001100101",
  39548=>"000010101",
  39549=>"010001010",
  39550=>"011110111",
  39551=>"100100100",
  39552=>"001010011",
  39553=>"011111110",
  39554=>"111000000",
  39555=>"100001100",
  39556=>"001101111",
  39557=>"011001111",
  39558=>"111110001",
  39559=>"000001001",
  39560=>"110110000",
  39561=>"011111011",
  39562=>"001001000",
  39563=>"110010100",
  39564=>"100000110",
  39565=>"111001000",
  39566=>"001011000",
  39567=>"000101100",
  39568=>"000001010",
  39569=>"110010010",
  39570=>"000111001",
  39571=>"010001001",
  39572=>"100101100",
  39573=>"111100001",
  39574=>"011111101",
  39575=>"001010001",
  39576=>"101011011",
  39577=>"001101000",
  39578=>"010110100",
  39579=>"101101001",
  39580=>"101001000",
  39581=>"100110001",
  39582=>"111110000",
  39583=>"111100011",
  39584=>"001010011",
  39585=>"011111001",
  39586=>"101000101",
  39587=>"000101011",
  39588=>"100010001",
  39589=>"100000001",
  39590=>"101100011",
  39591=>"100010101",
  39592=>"110001011",
  39593=>"101000000",
  39594=>"100011101",
  39595=>"011000001",
  39596=>"111001010",
  39597=>"000110100",
  39598=>"101100100",
  39599=>"100001100",
  39600=>"101111001",
  39601=>"011101000",
  39602=>"011100010",
  39603=>"010001000",
  39604=>"100010011",
  39605=>"011100111",
  39606=>"100000010",
  39607=>"011111101",
  39608=>"000010010",
  39609=>"110010011",
  39610=>"001100000",
  39611=>"000000110",
  39612=>"110011111",
  39613=>"101101010",
  39614=>"100111111",
  39615=>"000100101",
  39616=>"111001110",
  39617=>"001010000",
  39618=>"000011101",
  39619=>"001110111",
  39620=>"000001010",
  39621=>"010101111",
  39622=>"010000101",
  39623=>"001111000",
  39624=>"111101000",
  39625=>"010011001",
  39626=>"001001000",
  39627=>"101010011",
  39628=>"000100111",
  39629=>"010000001",
  39630=>"111000111",
  39631=>"011001101",
  39632=>"010101010",
  39633=>"001010100",
  39634=>"110111000",
  39635=>"101110001",
  39636=>"011011010",
  39637=>"010000101",
  39638=>"001100101",
  39639=>"011111111",
  39640=>"011100010",
  39641=>"100101100",
  39642=>"111110111",
  39643=>"101111000",
  39644=>"100111001",
  39645=>"011000000",
  39646=>"000010011",
  39647=>"000010111",
  39648=>"001101110",
  39649=>"101111101",
  39650=>"010010010",
  39651=>"000001001",
  39652=>"101000101",
  39653=>"100011110",
  39654=>"000011101",
  39655=>"000001110",
  39656=>"101101011",
  39657=>"000010100",
  39658=>"000001111",
  39659=>"000001001",
  39660=>"000001110",
  39661=>"010100001",
  39662=>"100111100",
  39663=>"000010101",
  39664=>"001010100",
  39665=>"001100001",
  39666=>"100101010",
  39667=>"101101000",
  39668=>"111110000",
  39669=>"001111010",
  39670=>"101111000",
  39671=>"001011010",
  39672=>"000001111",
  39673=>"101011100",
  39674=>"101011101",
  39675=>"101001101",
  39676=>"011000100",
  39677=>"101100101",
  39678=>"110010011",
  39679=>"000001100",
  39680=>"100011001",
  39681=>"001001010",
  39682=>"000000101",
  39683=>"000000110",
  39684=>"011110110",
  39685=>"100010011",
  39686=>"100000111",
  39687=>"011010010",
  39688=>"010000011",
  39689=>"100011001",
  39690=>"111101011",
  39691=>"010111010",
  39692=>"001011101",
  39693=>"001011101",
  39694=>"101110111",
  39695=>"111000010",
  39696=>"010101000",
  39697=>"001000110",
  39698=>"111110111",
  39699=>"100001010",
  39700=>"101101100",
  39701=>"101100010",
  39702=>"110110110",
  39703=>"110110110",
  39704=>"001011001",
  39705=>"101000100",
  39706=>"011111110",
  39707=>"011100100",
  39708=>"011000110",
  39709=>"011110001",
  39710=>"011000000",
  39711=>"110101110",
  39712=>"101100110",
  39713=>"010111010",
  39714=>"110100100",
  39715=>"001111010",
  39716=>"101111001",
  39717=>"111101010",
  39718=>"101011001",
  39719=>"000001000",
  39720=>"101100100",
  39721=>"000000000",
  39722=>"000100011",
  39723=>"110010000",
  39724=>"101100010",
  39725=>"101101110",
  39726=>"011011011",
  39727=>"100010111",
  39728=>"110001101",
  39729=>"011101100",
  39730=>"110100111",
  39731=>"000100011",
  39732=>"001111111",
  39733=>"000011000",
  39734=>"101001110",
  39735=>"101000001",
  39736=>"110101001",
  39737=>"110010110",
  39738=>"100111101",
  39739=>"101111010",
  39740=>"111111110",
  39741=>"000001101",
  39742=>"111110100",
  39743=>"001100100",
  39744=>"011100001",
  39745=>"001101100",
  39746=>"111101110",
  39747=>"010000000",
  39748=>"101101100",
  39749=>"010111011",
  39750=>"001010001",
  39751=>"001101000",
  39752=>"010010110",
  39753=>"011011100",
  39754=>"010111010",
  39755=>"000101011",
  39756=>"000100110",
  39757=>"110001011",
  39758=>"000000111",
  39759=>"000010001",
  39760=>"111110110",
  39761=>"100011101",
  39762=>"100000110",
  39763=>"011110110",
  39764=>"110000010",
  39765=>"100100010",
  39766=>"111110000",
  39767=>"001001000",
  39768=>"101000111",
  39769=>"010001001",
  39770=>"100100110",
  39771=>"000001001",
  39772=>"101011110",
  39773=>"100011100",
  39774=>"111000110",
  39775=>"101111001",
  39776=>"110000111",
  39777=>"010000001",
  39778=>"010111110",
  39779=>"110011011",
  39780=>"100111111",
  39781=>"011111100",
  39782=>"000111101",
  39783=>"110001110",
  39784=>"010111101",
  39785=>"101110000",
  39786=>"100001001",
  39787=>"111000011",
  39788=>"000100100",
  39789=>"100101011",
  39790=>"111011110",
  39791=>"001110100",
  39792=>"000010110",
  39793=>"011111110",
  39794=>"110111110",
  39795=>"100011010",
  39796=>"101011110",
  39797=>"101011101",
  39798=>"000111001",
  39799=>"100101100",
  39800=>"001101011",
  39801=>"000111001",
  39802=>"011100001",
  39803=>"110101110",
  39804=>"001001101",
  39805=>"001101111",
  39806=>"111111110",
  39807=>"011010000",
  39808=>"110001001",
  39809=>"111110000",
  39810=>"001010000",
  39811=>"000100101",
  39812=>"011000110",
  39813=>"000111001",
  39814=>"101010100",
  39815=>"001110001",
  39816=>"111000111",
  39817=>"101011011",
  39818=>"111011001",
  39819=>"001001111",
  39820=>"111111101",
  39821=>"111010101",
  39822=>"000001010",
  39823=>"010001111",
  39824=>"110100001",
  39825=>"101010001",
  39826=>"000000000",
  39827=>"000001000",
  39828=>"011011000",
  39829=>"000011110",
  39830=>"101001110",
  39831=>"011110010",
  39832=>"010001100",
  39833=>"110110101",
  39834=>"011000110",
  39835=>"000000100",
  39836=>"000010100",
  39837=>"011001110",
  39838=>"101111101",
  39839=>"011011100",
  39840=>"000011110",
  39841=>"101110111",
  39842=>"011011100",
  39843=>"111010001",
  39844=>"011000100",
  39845=>"011001110",
  39846=>"000100110",
  39847=>"010001000",
  39848=>"000010010",
  39849=>"001010000",
  39850=>"100110110",
  39851=>"101000111",
  39852=>"010101000",
  39853=>"010101000",
  39854=>"010110011",
  39855=>"000010000",
  39856=>"001000101",
  39857=>"001111100",
  39858=>"010101100",
  39859=>"011111100",
  39860=>"100011000",
  39861=>"111000010",
  39862=>"111000111",
  39863=>"100100000",
  39864=>"100100000",
  39865=>"010001101",
  39866=>"101101101",
  39867=>"101110011",
  39868=>"001100101",
  39869=>"110110111",
  39870=>"010011011",
  39871=>"111000110",
  39872=>"010111111",
  39873=>"010111001",
  39874=>"000010110",
  39875=>"110011011",
  39876=>"111110110",
  39877=>"000100000",
  39878=>"001001100",
  39879=>"001001110",
  39880=>"101110100",
  39881=>"011011000",
  39882=>"110000111",
  39883=>"000110101",
  39884=>"000100111",
  39885=>"100110110",
  39886=>"011101011",
  39887=>"100110111",
  39888=>"101111011",
  39889=>"011010110",
  39890=>"100110101",
  39891=>"000001000",
  39892=>"110101000",
  39893=>"110010000",
  39894=>"000011011",
  39895=>"000101111",
  39896=>"000110000",
  39897=>"001000101",
  39898=>"011011001",
  39899=>"001011001",
  39900=>"111000100",
  39901=>"111101011",
  39902=>"000000111",
  39903=>"111010011",
  39904=>"001111100",
  39905=>"110010110",
  39906=>"110010001",
  39907=>"010010011",
  39908=>"100001011",
  39909=>"001110101",
  39910=>"011111000",
  39911=>"101000111",
  39912=>"000011100",
  39913=>"010011101",
  39914=>"111011111",
  39915=>"100001111",
  39916=>"100010111",
  39917=>"010101000",
  39918=>"111101001",
  39919=>"001111001",
  39920=>"010011011",
  39921=>"010011011",
  39922=>"010001101",
  39923=>"000011001",
  39924=>"000000011",
  39925=>"011111011",
  39926=>"011110100",
  39927=>"100110111",
  39928=>"011110111",
  39929=>"001100110",
  39930=>"110101010",
  39931=>"001011001",
  39932=>"011001011",
  39933=>"111000100",
  39934=>"000111010",
  39935=>"001001111",
  39936=>"111100111",
  39937=>"001110111",
  39938=>"001011100",
  39939=>"001111110",
  39940=>"011111101",
  39941=>"110101001",
  39942=>"011001000",
  39943=>"110101111",
  39944=>"110011100",
  39945=>"000110100",
  39946=>"111110010",
  39947=>"110111110",
  39948=>"000111111",
  39949=>"000101010",
  39950=>"011011100",
  39951=>"111000110",
  39952=>"011110100",
  39953=>"010100010",
  39954=>"010010010",
  39955=>"100000001",
  39956=>"000111011",
  39957=>"001000111",
  39958=>"011101101",
  39959=>"010100000",
  39960=>"110100010",
  39961=>"010011101",
  39962=>"000000100",
  39963=>"101001010",
  39964=>"110001001",
  39965=>"000110011",
  39966=>"000100011",
  39967=>"100010010",
  39968=>"000001000",
  39969=>"110011100",
  39970=>"001101001",
  39971=>"011111110",
  39972=>"110101010",
  39973=>"101110111",
  39974=>"111010100",
  39975=>"000010111",
  39976=>"001110111",
  39977=>"000101001",
  39978=>"111000001",
  39979=>"111001111",
  39980=>"111000100",
  39981=>"010010010",
  39982=>"001010011",
  39983=>"000110001",
  39984=>"100011101",
  39985=>"101101111",
  39986=>"110001100",
  39987=>"100010000",
  39988=>"100110111",
  39989=>"010111000",
  39990=>"111001011",
  39991=>"000110110",
  39992=>"001001100",
  39993=>"010110111",
  39994=>"001011100",
  39995=>"011011111",
  39996=>"001111010",
  39997=>"111110001",
  39998=>"011111111",
  39999=>"010101101",
  40000=>"010001001",
  40001=>"000101111",
  40002=>"100100011",
  40003=>"100101011",
  40004=>"000001000",
  40005=>"000100011",
  40006=>"110011000",
  40007=>"001010010",
  40008=>"101000110",
  40009=>"101011110",
  40010=>"001000001",
  40011=>"111110110",
  40012=>"100000101",
  40013=>"111101010",
  40014=>"101011011",
  40015=>"011011010",
  40016=>"100000111",
  40017=>"100011010",
  40018=>"101000011",
  40019=>"001010000",
  40020=>"101000001",
  40021=>"001000001",
  40022=>"110111010",
  40023=>"011101111",
  40024=>"110011111",
  40025=>"000000110",
  40026=>"001110011",
  40027=>"101011000",
  40028=>"110101001",
  40029=>"010001010",
  40030=>"000011110",
  40031=>"001000111",
  40032=>"010111100",
  40033=>"000000101",
  40034=>"011101010",
  40035=>"111001001",
  40036=>"011110000",
  40037=>"100100111",
  40038=>"101100000",
  40039=>"010100011",
  40040=>"100100001",
  40041=>"110101001",
  40042=>"110011000",
  40043=>"010010111",
  40044=>"110010100",
  40045=>"010000011",
  40046=>"100110111",
  40047=>"011100110",
  40048=>"100111000",
  40049=>"001011100",
  40050=>"000100011",
  40051=>"111011100",
  40052=>"001110011",
  40053=>"110110110",
  40054=>"010011011",
  40055=>"010100010",
  40056=>"011001000",
  40057=>"111101100",
  40058=>"110111111",
  40059=>"011001001",
  40060=>"111101011",
  40061=>"110111111",
  40062=>"101111111",
  40063=>"100011010",
  40064=>"011111010",
  40065=>"111100101",
  40066=>"111101111",
  40067=>"101001000",
  40068=>"100101100",
  40069=>"111110101",
  40070=>"111010101",
  40071=>"101100100",
  40072=>"111011010",
  40073=>"001010000",
  40074=>"100011001",
  40075=>"000101011",
  40076=>"110100000",
  40077=>"111110000",
  40078=>"100101110",
  40079=>"111010000",
  40080=>"011111010",
  40081=>"010110001",
  40082=>"100000101",
  40083=>"111110100",
  40084=>"010001111",
  40085=>"010111111",
  40086=>"001001001",
  40087=>"011001101",
  40088=>"111010010",
  40089=>"101001101",
  40090=>"000011010",
  40091=>"101110110",
  40092=>"001010000",
  40093=>"101010010",
  40094=>"001000001",
  40095=>"011010000",
  40096=>"000100100",
  40097=>"010100100",
  40098=>"000010000",
  40099=>"001001101",
  40100=>"110101111",
  40101=>"000011101",
  40102=>"001001100",
  40103=>"110100100",
  40104=>"100101000",
  40105=>"000100011",
  40106=>"110101000",
  40107=>"111111011",
  40108=>"110010101",
  40109=>"001100111",
  40110=>"101001111",
  40111=>"011011000",
  40112=>"010001001",
  40113=>"101011010",
  40114=>"111011010",
  40115=>"110110000",
  40116=>"101011000",
  40117=>"100001100",
  40118=>"000010111",
  40119=>"101010100",
  40120=>"010110010",
  40121=>"011110000",
  40122=>"001011001",
  40123=>"000011100",
  40124=>"110010010",
  40125=>"000010010",
  40126=>"101111110",
  40127=>"101000110",
  40128=>"111110011",
  40129=>"001100010",
  40130=>"010000111",
  40131=>"010001001",
  40132=>"011011001",
  40133=>"010010100",
  40134=>"000101011",
  40135=>"111001001",
  40136=>"100000110",
  40137=>"100011001",
  40138=>"101000111",
  40139=>"111101010",
  40140=>"001000101",
  40141=>"010100001",
  40142=>"100001011",
  40143=>"110010000",
  40144=>"011010011",
  40145=>"100000010",
  40146=>"110111111",
  40147=>"011101101",
  40148=>"000100101",
  40149=>"010000001",
  40150=>"011101100",
  40151=>"000011010",
  40152=>"100000110",
  40153=>"100100111",
  40154=>"000011111",
  40155=>"100100011",
  40156=>"101001111",
  40157=>"001000000",
  40158=>"010110111",
  40159=>"000011110",
  40160=>"000101110",
  40161=>"110110000",
  40162=>"100010011",
  40163=>"000011000",
  40164=>"111000100",
  40165=>"001110100",
  40166=>"101110100",
  40167=>"101101100",
  40168=>"000111111",
  40169=>"001000110",
  40170=>"110000000",
  40171=>"111010111",
  40172=>"000001010",
  40173=>"111111101",
  40174=>"001100100",
  40175=>"111000000",
  40176=>"010001010",
  40177=>"110101001",
  40178=>"110110100",
  40179=>"111111101",
  40180=>"001000101",
  40181=>"001010000",
  40182=>"100000101",
  40183=>"000000101",
  40184=>"010011110",
  40185=>"001000100",
  40186=>"101111010",
  40187=>"000010100",
  40188=>"110100110",
  40189=>"111011100",
  40190=>"110111111",
  40191=>"111111110",
  40192=>"011100000",
  40193=>"000010001",
  40194=>"010011101",
  40195=>"111111000",
  40196=>"001011111",
  40197=>"101111010",
  40198=>"100001111",
  40199=>"000001010",
  40200=>"010101010",
  40201=>"011111101",
  40202=>"100111000",
  40203=>"111010110",
  40204=>"000100100",
  40205=>"010111001",
  40206=>"100100111",
  40207=>"111101111",
  40208=>"011001010",
  40209=>"011110101",
  40210=>"001000111",
  40211=>"001100000",
  40212=>"110101111",
  40213=>"010100110",
  40214=>"111011100",
  40215=>"011111101",
  40216=>"101000011",
  40217=>"110101011",
  40218=>"010001010",
  40219=>"101111001",
  40220=>"111000011",
  40221=>"000011010",
  40222=>"001110000",
  40223=>"000110000",
  40224=>"001011000",
  40225=>"010100110",
  40226=>"001000101",
  40227=>"100000100",
  40228=>"111001111",
  40229=>"111011100",
  40230=>"110111111",
  40231=>"011000010",
  40232=>"100101011",
  40233=>"001011000",
  40234=>"001101011",
  40235=>"111001001",
  40236=>"010111001",
  40237=>"111010001",
  40238=>"010111110",
  40239=>"001010110",
  40240=>"001000000",
  40241=>"100010000",
  40242=>"011110010",
  40243=>"101011111",
  40244=>"000010010",
  40245=>"101101111",
  40246=>"000001100",
  40247=>"101100010",
  40248=>"110010010",
  40249=>"010101001",
  40250=>"100100111",
  40251=>"001011011",
  40252=>"001101001",
  40253=>"100100101",
  40254=>"001101100",
  40255=>"110001000",
  40256=>"101001010",
  40257=>"110100010",
  40258=>"100001100",
  40259=>"000101001",
  40260=>"011011111",
  40261=>"000011000",
  40262=>"010000000",
  40263=>"000000101",
  40264=>"010000000",
  40265=>"001001100",
  40266=>"000000110",
  40267=>"111010110",
  40268=>"000010001",
  40269=>"000000011",
  40270=>"100011101",
  40271=>"011010001",
  40272=>"110110011",
  40273=>"100000100",
  40274=>"101000000",
  40275=>"111010110",
  40276=>"100000100",
  40277=>"100001011",
  40278=>"110101011",
  40279=>"100101101",
  40280=>"000000000",
  40281=>"100110111",
  40282=>"100001111",
  40283=>"000010011",
  40284=>"110010110",
  40285=>"000101011",
  40286=>"110010101",
  40287=>"000100010",
  40288=>"111110111",
  40289=>"111001111",
  40290=>"100111011",
  40291=>"111100100",
  40292=>"101010111",
  40293=>"001000110",
  40294=>"011001100",
  40295=>"001101000",
  40296=>"110101011",
  40297=>"111111111",
  40298=>"111000010",
  40299=>"001111011",
  40300=>"101110011",
  40301=>"110110100",
  40302=>"101011101",
  40303=>"000001101",
  40304=>"100100010",
  40305=>"001001010",
  40306=>"011000100",
  40307=>"000111011",
  40308=>"000111000",
  40309=>"001000010",
  40310=>"001111001",
  40311=>"110101001",
  40312=>"001000010",
  40313=>"100000001",
  40314=>"000111011",
  40315=>"111010001",
  40316=>"011111100",
  40317=>"000010000",
  40318=>"001001011",
  40319=>"010001110",
  40320=>"010001000",
  40321=>"011000000",
  40322=>"000110110",
  40323=>"110000100",
  40324=>"111010101",
  40325=>"011110111",
  40326=>"111000001",
  40327=>"011011010",
  40328=>"110011101",
  40329=>"111110010",
  40330=>"111001010",
  40331=>"111101110",
  40332=>"100000110",
  40333=>"100001101",
  40334=>"110100100",
  40335=>"011100000",
  40336=>"001111100",
  40337=>"000011000",
  40338=>"001100100",
  40339=>"101001001",
  40340=>"011001100",
  40341=>"111000001",
  40342=>"101100101",
  40343=>"001100111",
  40344=>"011101101",
  40345=>"011110100",
  40346=>"110001111",
  40347=>"000110010",
  40348=>"111110111",
  40349=>"100001001",
  40350=>"001100011",
  40351=>"111110010",
  40352=>"001000000",
  40353=>"010011101",
  40354=>"111101001",
  40355=>"100001100",
  40356=>"110011110",
  40357=>"010110011",
  40358=>"101011100",
  40359=>"101111100",
  40360=>"110111111",
  40361=>"100010101",
  40362=>"000010000",
  40363=>"000101110",
  40364=>"100010011",
  40365=>"001010001",
  40366=>"000010000",
  40367=>"010100110",
  40368=>"010011010",
  40369=>"000000000",
  40370=>"101000010",
  40371=>"111000011",
  40372=>"111111010",
  40373=>"101110000",
  40374=>"010110010",
  40375=>"001010010",
  40376=>"111010010",
  40377=>"000110101",
  40378=>"110110010",
  40379=>"001011100",
  40380=>"100101100",
  40381=>"111011100",
  40382=>"001101111",
  40383=>"000110111",
  40384=>"101101111",
  40385=>"010011001",
  40386=>"011001011",
  40387=>"101000011",
  40388=>"010111011",
  40389=>"100101001",
  40390=>"010110101",
  40391=>"100001000",
  40392=>"010001001",
  40393=>"010110011",
  40394=>"111000111",
  40395=>"100001100",
  40396=>"010110000",
  40397=>"101010001",
  40398=>"110100101",
  40399=>"110011110",
  40400=>"101111101",
  40401=>"111001110",
  40402=>"010110011",
  40403=>"100000110",
  40404=>"100000111",
  40405=>"011010110",
  40406=>"110000001",
  40407=>"101100110",
  40408=>"001100100",
  40409=>"011010010",
  40410=>"010100000",
  40411=>"110110110",
  40412=>"001010110",
  40413=>"001111100",
  40414=>"001011011",
  40415=>"000101010",
  40416=>"100111100",
  40417=>"111101111",
  40418=>"000011110",
  40419=>"000111100",
  40420=>"101010010",
  40421=>"110110100",
  40422=>"111101011",
  40423=>"110100000",
  40424=>"101110100",
  40425=>"000111011",
  40426=>"111100001",
  40427=>"110111100",
  40428=>"000000110",
  40429=>"101111101",
  40430=>"110101111",
  40431=>"010010000",
  40432=>"001001000",
  40433=>"111111101",
  40434=>"101110100",
  40435=>"111101001",
  40436=>"100001011",
  40437=>"111001110",
  40438=>"000100110",
  40439=>"001000000",
  40440=>"100001001",
  40441=>"001110011",
  40442=>"100110110",
  40443=>"111010000",
  40444=>"100111001",
  40445=>"010001100",
  40446=>"010101101",
  40447=>"111010111",
  40448=>"100001101",
  40449=>"100111101",
  40450=>"100101010",
  40451=>"000001010",
  40452=>"000010011",
  40453=>"111111111",
  40454=>"100001001",
  40455=>"000010110",
  40456=>"111110101",
  40457=>"101001000",
  40458=>"111010111",
  40459=>"001111001",
  40460=>"001001011",
  40461=>"100011111",
  40462=>"100110110",
  40463=>"000110011",
  40464=>"000000000",
  40465=>"011110111",
  40466=>"001011000",
  40467=>"100011111",
  40468=>"101011100",
  40469=>"101100011",
  40470=>"000000101",
  40471=>"001110101",
  40472=>"011111110",
  40473=>"110010000",
  40474=>"101100110",
  40475=>"100010101",
  40476=>"110000011",
  40477=>"111001011",
  40478=>"001001000",
  40479=>"011011110",
  40480=>"010000001",
  40481=>"101000101",
  40482=>"110000000",
  40483=>"111011011",
  40484=>"110011010",
  40485=>"011101111",
  40486=>"101010001",
  40487=>"100111100",
  40488=>"010011010",
  40489=>"100110010",
  40490=>"010011000",
  40491=>"011101110",
  40492=>"110100000",
  40493=>"000100101",
  40494=>"111101101",
  40495=>"010111110",
  40496=>"011011000",
  40497=>"000010110",
  40498=>"000010101",
  40499=>"100101011",
  40500=>"000011111",
  40501=>"000000000",
  40502=>"100101100",
  40503=>"111101011",
  40504=>"000111111",
  40505=>"100100011",
  40506=>"010001001",
  40507=>"100000101",
  40508=>"011110010",
  40509=>"011111101",
  40510=>"101000111",
  40511=>"101101100",
  40512=>"101111101",
  40513=>"000000010",
  40514=>"000000111",
  40515=>"010101100",
  40516=>"101110110",
  40517=>"011101101",
  40518=>"001110011",
  40519=>"110100101",
  40520=>"000101000",
  40521=>"000001001",
  40522=>"100110111",
  40523=>"001000100",
  40524=>"111101010",
  40525=>"100000100",
  40526=>"011100100",
  40527=>"100110100",
  40528=>"001001011",
  40529=>"000110000",
  40530=>"100100010",
  40531=>"000010001",
  40532=>"010001000",
  40533=>"011000000",
  40534=>"010001100",
  40535=>"101000100",
  40536=>"101010111",
  40537=>"000111111",
  40538=>"000101111",
  40539=>"000001100",
  40540=>"000101010",
  40541=>"100111010",
  40542=>"000001111",
  40543=>"011111010",
  40544=>"111010000",
  40545=>"010101100",
  40546=>"001010010",
  40547=>"111010010",
  40548=>"111101011",
  40549=>"000011010",
  40550=>"011010000",
  40551=>"101111011",
  40552=>"110001000",
  40553=>"001011000",
  40554=>"000100101",
  40555=>"001100000",
  40556=>"111010101",
  40557=>"000011100",
  40558=>"110111011",
  40559=>"111011101",
  40560=>"111110001",
  40561=>"010011001",
  40562=>"111000001",
  40563=>"001001000",
  40564=>"001100001",
  40565=>"111110101",
  40566=>"011000000",
  40567=>"100001101",
  40568=>"001101110",
  40569=>"000110000",
  40570=>"101111000",
  40571=>"000001101",
  40572=>"010110000",
  40573=>"110010110",
  40574=>"010000101",
  40575=>"101011110",
  40576=>"001011000",
  40577=>"011100111",
  40578=>"010101111",
  40579=>"000111110",
  40580=>"001110111",
  40581=>"000110110",
  40582=>"001100011",
  40583=>"111010011",
  40584=>"110011110",
  40585=>"010110010",
  40586=>"111101111",
  40587=>"111100000",
  40588=>"111100101",
  40589=>"000011111",
  40590=>"000101111",
  40591=>"010111000",
  40592=>"110001111",
  40593=>"010100000",
  40594=>"010010000",
  40595=>"000110101",
  40596=>"110000000",
  40597=>"100000000",
  40598=>"111111001",
  40599=>"101111101",
  40600=>"101000100",
  40601=>"011010000",
  40602=>"011111100",
  40603=>"111111010",
  40604=>"011110101",
  40605=>"000110011",
  40606=>"111000111",
  40607=>"001000000",
  40608=>"001000011",
  40609=>"100010100",
  40610=>"001000010",
  40611=>"101010111",
  40612=>"011001100",
  40613=>"100010000",
  40614=>"000100101",
  40615=>"000000000",
  40616=>"001010111",
  40617=>"110010010",
  40618=>"101010101",
  40619=>"011000011",
  40620=>"101001101",
  40621=>"110000010",
  40622=>"010110100",
  40623=>"100101001",
  40624=>"100100100",
  40625=>"110001100",
  40626=>"000010011",
  40627=>"000101010",
  40628=>"000000100",
  40629=>"010111001",
  40630=>"010000011",
  40631=>"000000111",
  40632=>"111011101",
  40633=>"110000010",
  40634=>"101000110",
  40635=>"100101010",
  40636=>"000101100",
  40637=>"101001000",
  40638=>"010011101",
  40639=>"110010011",
  40640=>"001010110",
  40641=>"111110010",
  40642=>"100000000",
  40643=>"111010001",
  40644=>"001011111",
  40645=>"010011111",
  40646=>"000000110",
  40647=>"110000000",
  40648=>"101101010",
  40649=>"010110000",
  40650=>"000000110",
  40651=>"110110001",
  40652=>"000001001",
  40653=>"111011111",
  40654=>"101100010",
  40655=>"110111100",
  40656=>"111110100",
  40657=>"111000000",
  40658=>"110101110",
  40659=>"010110101",
  40660=>"111101101",
  40661=>"000111110",
  40662=>"011101100",
  40663=>"110100001",
  40664=>"101001110",
  40665=>"110111100",
  40666=>"000001110",
  40667=>"101010010",
  40668=>"010001001",
  40669=>"110110101",
  40670=>"000101111",
  40671=>"110011101",
  40672=>"000001110",
  40673=>"100111010",
  40674=>"100000100",
  40675=>"010011011",
  40676=>"111000100",
  40677=>"100001011",
  40678=>"001001110",
  40679=>"111010101",
  40680=>"101110010",
  40681=>"001111100",
  40682=>"001011001",
  40683=>"111101111",
  40684=>"011101010",
  40685=>"111111101",
  40686=>"011001100",
  40687=>"101110000",
  40688=>"000101111",
  40689=>"110001100",
  40690=>"000111010",
  40691=>"101101101",
  40692=>"101011101",
  40693=>"111011101",
  40694=>"001111001",
  40695=>"110000010",
  40696=>"100100001",
  40697=>"011101010",
  40698=>"100010101",
  40699=>"110111001",
  40700=>"001101101",
  40701=>"001110000",
  40702=>"010101000",
  40703=>"111111111",
  40704=>"100110000",
  40705=>"111110111",
  40706=>"110101010",
  40707=>"101100111",
  40708=>"000001000",
  40709=>"000011010",
  40710=>"100000011",
  40711=>"001011001",
  40712=>"101010011",
  40713=>"000100101",
  40714=>"110001100",
  40715=>"000111101",
  40716=>"111111011",
  40717=>"100011100",
  40718=>"110100000",
  40719=>"111110100",
  40720=>"111010010",
  40721=>"010101110",
  40722=>"010011101",
  40723=>"100111011",
  40724=>"101110010",
  40725=>"000010010",
  40726=>"010110110",
  40727=>"000010010",
  40728=>"110011001",
  40729=>"001001100",
  40730=>"000000010",
  40731=>"000000110",
  40732=>"010011011",
  40733=>"101011000",
  40734=>"110010000",
  40735=>"110011101",
  40736=>"101110111",
  40737=>"101011010",
  40738=>"101011000",
  40739=>"110010010",
  40740=>"001010001",
  40741=>"101000101",
  40742=>"101001111",
  40743=>"011000010",
  40744=>"010001011",
  40745=>"000101001",
  40746=>"000000000",
  40747=>"001111111",
  40748=>"011011011",
  40749=>"111010101",
  40750=>"011100011",
  40751=>"111101000",
  40752=>"101101011",
  40753=>"110011000",
  40754=>"000000100",
  40755=>"011101100",
  40756=>"111100110",
  40757=>"111100000",
  40758=>"111010111",
  40759=>"110111100",
  40760=>"001011111",
  40761=>"000101011",
  40762=>"000000010",
  40763=>"011111001",
  40764=>"100111111",
  40765=>"010100010",
  40766=>"100010001",
  40767=>"000100101",
  40768=>"010011000",
  40769=>"101010000",
  40770=>"111110111",
  40771=>"000001000",
  40772=>"001000101",
  40773=>"010000101",
  40774=>"010101111",
  40775=>"010111111",
  40776=>"110101111",
  40777=>"000010111",
  40778=>"101011100",
  40779=>"010001011",
  40780=>"010011000",
  40781=>"011100111",
  40782=>"000001110",
  40783=>"110010111",
  40784=>"110001011",
  40785=>"000000011",
  40786=>"000010101",
  40787=>"101100111",
  40788=>"010111011",
  40789=>"001000110",
  40790=>"100101011",
  40791=>"110011011",
  40792=>"110000010",
  40793=>"111100001",
  40794=>"110101000",
  40795=>"101101110",
  40796=>"101111101",
  40797=>"100001001",
  40798=>"110001011",
  40799=>"000100100",
  40800=>"010011010",
  40801=>"001100000",
  40802=>"001000001",
  40803=>"111100010",
  40804=>"001100000",
  40805=>"101110110",
  40806=>"110110011",
  40807=>"110110101",
  40808=>"111000100",
  40809=>"111011100",
  40810=>"111110010",
  40811=>"111010111",
  40812=>"001100000",
  40813=>"110110000",
  40814=>"111100001",
  40815=>"101111110",
  40816=>"000010110",
  40817=>"000001110",
  40818=>"001100011",
  40819=>"000010110",
  40820=>"000100100",
  40821=>"100011000",
  40822=>"011110000",
  40823=>"110001010",
  40824=>"111010110",
  40825=>"111100100",
  40826=>"100000000",
  40827=>"001101000",
  40828=>"100011000",
  40829=>"100111011",
  40830=>"010011011",
  40831=>"010010001",
  40832=>"001010110",
  40833=>"000001111",
  40834=>"000000011",
  40835=>"011010110",
  40836=>"000010000",
  40837=>"000010011",
  40838=>"011010000",
  40839=>"010110101",
  40840=>"111000001",
  40841=>"100000010",
  40842=>"110000010",
  40843=>"100000000",
  40844=>"100001001",
  40845=>"000010101",
  40846=>"110111011",
  40847=>"000010001",
  40848=>"101101011",
  40849=>"110111001",
  40850=>"100110100",
  40851=>"000100101",
  40852=>"111110101",
  40853=>"100001000",
  40854=>"110101101",
  40855=>"010101110",
  40856=>"101110101",
  40857=>"000100001",
  40858=>"111100100",
  40859=>"010011110",
  40860=>"100011010",
  40861=>"100000010",
  40862=>"111000000",
  40863=>"001000000",
  40864=>"110100110",
  40865=>"100011100",
  40866=>"010110010",
  40867=>"011100101",
  40868=>"001001100",
  40869=>"001001110",
  40870=>"111000000",
  40871=>"101101101",
  40872=>"010100111",
  40873=>"110010101",
  40874=>"111011001",
  40875=>"100110001",
  40876=>"110000101",
  40877=>"100101010",
  40878=>"011001100",
  40879=>"001110110",
  40880=>"111101100",
  40881=>"111111101",
  40882=>"010110001",
  40883=>"001000111",
  40884=>"111100101",
  40885=>"011001000",
  40886=>"010010111",
  40887=>"110000000",
  40888=>"101010010",
  40889=>"110100111",
  40890=>"001100011",
  40891=>"010000101",
  40892=>"011111111",
  40893=>"110100110",
  40894=>"101101101",
  40895=>"100101000",
  40896=>"100000110",
  40897=>"011101100",
  40898=>"010010000",
  40899=>"111001101",
  40900=>"010101000",
  40901=>"010000001",
  40902=>"000110011",
  40903=>"111110011",
  40904=>"101001001",
  40905=>"010000111",
  40906=>"011100101",
  40907=>"001111110",
  40908=>"000010100",
  40909=>"011011110",
  40910=>"100110010",
  40911=>"000011100",
  40912=>"110000100",
  40913=>"011010101",
  40914=>"100111010",
  40915=>"101101101",
  40916=>"001011000",
  40917=>"000010111",
  40918=>"111001010",
  40919=>"010010001",
  40920=>"100011010",
  40921=>"000011101",
  40922=>"001000100",
  40923=>"000001010",
  40924=>"010100111",
  40925=>"100011011",
  40926=>"110011101",
  40927=>"011101111",
  40928=>"111101011",
  40929=>"101110100",
  40930=>"010000010",
  40931=>"100000000",
  40932=>"100100000",
  40933=>"100100011",
  40934=>"010111001",
  40935=>"001000111",
  40936=>"000000111",
  40937=>"101111100",
  40938=>"000100111",
  40939=>"011010000",
  40940=>"111111111",
  40941=>"011100001",
  40942=>"101000010",
  40943=>"000001010",
  40944=>"000110011",
  40945=>"101011111",
  40946=>"010011011",
  40947=>"011000110",
  40948=>"001111101",
  40949=>"100001001",
  40950=>"010101111",
  40951=>"101111111",
  40952=>"101111110",
  40953=>"101111101",
  40954=>"010111010",
  40955=>"010111100",
  40956=>"100100011",
  40957=>"000111000",
  40958=>"110001010",
  40959=>"110111100",
  40960=>"010101101",
  40961=>"100000000",
  40962=>"010010101",
  40963=>"100100000",
  40964=>"000001101",
  40965=>"100010011",
  40966=>"011101000",
  40967=>"010111101",
  40968=>"011101011",
  40969=>"000101110",
  40970=>"100001011",
  40971=>"001100100",
  40972=>"011111110",
  40973=>"111100011",
  40974=>"001101100",
  40975=>"110000111",
  40976=>"100000001",
  40977=>"111011111",
  40978=>"100001110",
  40979=>"001000001",
  40980=>"010001100",
  40981=>"110110111",
  40982=>"001110000",
  40983=>"001111001",
  40984=>"101111110",
  40985=>"011110110",
  40986=>"100001101",
  40987=>"000000011",
  40988=>"001100100",
  40989=>"110010011",
  40990=>"011001100",
  40991=>"110101000",
  40992=>"010010111",
  40993=>"011110101",
  40994=>"111111001",
  40995=>"001001111",
  40996=>"111000010",
  40997=>"111000101",
  40998=>"001000011",
  40999=>"011000010",
  41000=>"011100011",
  41001=>"111100001",
  41002=>"111101001",
  41003=>"011100011",
  41004=>"000111101",
  41005=>"100100010",
  41006=>"001000101",
  41007=>"001111011",
  41008=>"001001101",
  41009=>"101110011",
  41010=>"110111010",
  41011=>"001100000",
  41012=>"010011100",
  41013=>"000000010",
  41014=>"100000100",
  41015=>"111001110",
  41016=>"010011100",
  41017=>"010010011",
  41018=>"011110000",
  41019=>"010011111",
  41020=>"100011010",
  41021=>"100110000",
  41022=>"010110001",
  41023=>"001010001",
  41024=>"111110111",
  41025=>"011000000",
  41026=>"001101101",
  41027=>"001110101",
  41028=>"100100100",
  41029=>"010101101",
  41030=>"100001001",
  41031=>"110011011",
  41032=>"100101100",
  41033=>"110000110",
  41034=>"110010100",
  41035=>"111001010",
  41036=>"011001011",
  41037=>"100100001",
  41038=>"000111011",
  41039=>"011100000",
  41040=>"011001000",
  41041=>"101111100",
  41042=>"000110000",
  41043=>"001000111",
  41044=>"101111101",
  41045=>"111010011",
  41046=>"110111100",
  41047=>"000111010",
  41048=>"000111000",
  41049=>"000011111",
  41050=>"110010010",
  41051=>"110101001",
  41052=>"011111101",
  41053=>"101111010",
  41054=>"101011010",
  41055=>"100001101",
  41056=>"001011111",
  41057=>"100001001",
  41058=>"101111100",
  41059=>"010000100",
  41060=>"111001010",
  41061=>"010100000",
  41062=>"000010011",
  41063=>"110010110",
  41064=>"111110011",
  41065=>"110110001",
  41066=>"000000010",
  41067=>"011000100",
  41068=>"001011000",
  41069=>"111100011",
  41070=>"100101000",
  41071=>"000101000",
  41072=>"111001101",
  41073=>"101111111",
  41074=>"111011100",
  41075=>"001101100",
  41076=>"010010100",
  41077=>"000100100",
  41078=>"111111001",
  41079=>"100110111",
  41080=>"010101110",
  41081=>"110000110",
  41082=>"101101111",
  41083=>"111100010",
  41084=>"100100000",
  41085=>"101110000",
  41086=>"101011100",
  41087=>"111110100",
  41088=>"111111111",
  41089=>"101100101",
  41090=>"010111000",
  41091=>"011111110",
  41092=>"000000010",
  41093=>"011001010",
  41094=>"101011110",
  41095=>"001100110",
  41096=>"010101010",
  41097=>"100011100",
  41098=>"010000101",
  41099=>"100000000",
  41100=>"011010000",
  41101=>"100001111",
  41102=>"000100000",
  41103=>"011011100",
  41104=>"011010000",
  41105=>"111110111",
  41106=>"010100000",
  41107=>"010110100",
  41108=>"110110100",
  41109=>"101100001",
  41110=>"011001110",
  41111=>"110110001",
  41112=>"110111000",
  41113=>"100011000",
  41114=>"100001001",
  41115=>"000001010",
  41116=>"111100011",
  41117=>"101001000",
  41118=>"110011010",
  41119=>"001001101",
  41120=>"101100110",
  41121=>"000010001",
  41122=>"111111011",
  41123=>"110110111",
  41124=>"011010100",
  41125=>"010001110",
  41126=>"100100000",
  41127=>"100100110",
  41128=>"010010000",
  41129=>"011100000",
  41130=>"110111000",
  41131=>"111000010",
  41132=>"000010001",
  41133=>"110011101",
  41134=>"011111011",
  41135=>"000100000",
  41136=>"000000110",
  41137=>"001010000",
  41138=>"110100111",
  41139=>"101111011",
  41140=>"100110101",
  41141=>"101110111",
  41142=>"000010101",
  41143=>"001000000",
  41144=>"010000010",
  41145=>"101011111",
  41146=>"011001111",
  41147=>"011011111",
  41148=>"111000000",
  41149=>"000000001",
  41150=>"101111111",
  41151=>"000101100",
  41152=>"001000100",
  41153=>"100000000",
  41154=>"111110010",
  41155=>"000010010",
  41156=>"011110100",
  41157=>"001010011",
  41158=>"100001110",
  41159=>"000000001",
  41160=>"010001000",
  41161=>"111101100",
  41162=>"100000111",
  41163=>"100010011",
  41164=>"101011001",
  41165=>"000101111",
  41166=>"001000111",
  41167=>"011111111",
  41168=>"010001111",
  41169=>"000111000",
  41170=>"001001111",
  41171=>"000100010",
  41172=>"100100010",
  41173=>"100110110",
  41174=>"100011110",
  41175=>"011111110",
  41176=>"111100001",
  41177=>"001100001",
  41178=>"101100100",
  41179=>"110111110",
  41180=>"101001001",
  41181=>"000001100",
  41182=>"010000000",
  41183=>"011101111",
  41184=>"010010010",
  41185=>"111110101",
  41186=>"001010111",
  41187=>"101000100",
  41188=>"101011001",
  41189=>"110101101",
  41190=>"000010110",
  41191=>"011101100",
  41192=>"100000110",
  41193=>"000110010",
  41194=>"000101100",
  41195=>"011110000",
  41196=>"001111110",
  41197=>"001110010",
  41198=>"001000010",
  41199=>"101111000",
  41200=>"000001101",
  41201=>"111001110",
  41202=>"001110110",
  41203=>"100001100",
  41204=>"101001101",
  41205=>"100011001",
  41206=>"110110010",
  41207=>"011000010",
  41208=>"100001110",
  41209=>"110001111",
  41210=>"110010000",
  41211=>"001000111",
  41212=>"010010011",
  41213=>"001100000",
  41214=>"010111010",
  41215=>"110001100",
  41216=>"010111001",
  41217=>"110101010",
  41218=>"011000010",
  41219=>"011111011",
  41220=>"110101110",
  41221=>"101101011",
  41222=>"101001000",
  41223=>"111101101",
  41224=>"101111001",
  41225=>"000001010",
  41226=>"011010011",
  41227=>"001010101",
  41228=>"110101011",
  41229=>"000010100",
  41230=>"010000101",
  41231=>"000111110",
  41232=>"010011000",
  41233=>"101101000",
  41234=>"000001000",
  41235=>"001111111",
  41236=>"000101111",
  41237=>"000111010",
  41238=>"010111010",
  41239=>"001110011",
  41240=>"100111000",
  41241=>"100100010",
  41242=>"101010000",
  41243=>"111110111",
  41244=>"111000001",
  41245=>"111100101",
  41246=>"000001111",
  41247=>"010001110",
  41248=>"011000100",
  41249=>"100101100",
  41250=>"111011011",
  41251=>"000110011",
  41252=>"110100001",
  41253=>"111000111",
  41254=>"010110000",
  41255=>"001101100",
  41256=>"000101100",
  41257=>"001001101",
  41258=>"101110100",
  41259=>"001010100",
  41260=>"001110110",
  41261=>"111010111",
  41262=>"000111001",
  41263=>"110111100",
  41264=>"100010000",
  41265=>"001000000",
  41266=>"010110111",
  41267=>"111000010",
  41268=>"110000001",
  41269=>"001011100",
  41270=>"100011000",
  41271=>"110111111",
  41272=>"110110010",
  41273=>"110111101",
  41274=>"111101100",
  41275=>"111101010",
  41276=>"000000100",
  41277=>"110001000",
  41278=>"110110101",
  41279=>"001001110",
  41280=>"111111111",
  41281=>"111101011",
  41282=>"101010100",
  41283=>"110100011",
  41284=>"100111111",
  41285=>"001100111",
  41286=>"011101111",
  41287=>"100101100",
  41288=>"100101101",
  41289=>"100001011",
  41290=>"111100110",
  41291=>"001011110",
  41292=>"001011110",
  41293=>"000011001",
  41294=>"001000100",
  41295=>"100101110",
  41296=>"000110111",
  41297=>"001111011",
  41298=>"110101000",
  41299=>"011000111",
  41300=>"011101111",
  41301=>"111111001",
  41302=>"101101100",
  41303=>"110101010",
  41304=>"011011010",
  41305=>"000011010",
  41306=>"111010000",
  41307=>"010010010",
  41308=>"100100010",
  41309=>"110011110",
  41310=>"010110101",
  41311=>"101011110",
  41312=>"111110100",
  41313=>"111101011",
  41314=>"000000100",
  41315=>"011100110",
  41316=>"000000010",
  41317=>"001011010",
  41318=>"010000001",
  41319=>"101111111",
  41320=>"101110111",
  41321=>"001101110",
  41322=>"010101001",
  41323=>"011110011",
  41324=>"101111100",
  41325=>"000010101",
  41326=>"001001111",
  41327=>"000001111",
  41328=>"110111010",
  41329=>"010111011",
  41330=>"010111001",
  41331=>"000011110",
  41332=>"011010111",
  41333=>"100010111",
  41334=>"011101000",
  41335=>"110001101",
  41336=>"111011000",
  41337=>"111001111",
  41338=>"110110010",
  41339=>"101100110",
  41340=>"010100110",
  41341=>"110000101",
  41342=>"001100010",
  41343=>"001011110",
  41344=>"001010010",
  41345=>"110010011",
  41346=>"111010001",
  41347=>"000100011",
  41348=>"001111001",
  41349=>"101001001",
  41350=>"000111011",
  41351=>"000011000",
  41352=>"011010100",
  41353=>"111111111",
  41354=>"010000110",
  41355=>"001100101",
  41356=>"110110110",
  41357=>"010110011",
  41358=>"101010101",
  41359=>"101111111",
  41360=>"001000100",
  41361=>"011000110",
  41362=>"000101001",
  41363=>"101101010",
  41364=>"101110000",
  41365=>"000000101",
  41366=>"000011001",
  41367=>"001011001",
  41368=>"011100110",
  41369=>"001011101",
  41370=>"000100010",
  41371=>"111011000",
  41372=>"101111000",
  41373=>"011111010",
  41374=>"000111000",
  41375=>"111111100",
  41376=>"000110110",
  41377=>"110110100",
  41378=>"110011000",
  41379=>"010100000",
  41380=>"011000000",
  41381=>"100000101",
  41382=>"000000000",
  41383=>"001001110",
  41384=>"001000100",
  41385=>"001111000",
  41386=>"010110101",
  41387=>"010100000",
  41388=>"011001011",
  41389=>"110101010",
  41390=>"111111001",
  41391=>"001101011",
  41392=>"011001001",
  41393=>"000011011",
  41394=>"011011010",
  41395=>"100111010",
  41396=>"011111000",
  41397=>"010101001",
  41398=>"000000001",
  41399=>"010110100",
  41400=>"001000100",
  41401=>"010011001",
  41402=>"110011110",
  41403=>"101111111",
  41404=>"101110100",
  41405=>"110101111",
  41406=>"001100000",
  41407=>"111011101",
  41408=>"010001010",
  41409=>"001000000",
  41410=>"110011101",
  41411=>"010001001",
  41412=>"010001000",
  41413=>"111111111",
  41414=>"001000101",
  41415=>"011001011",
  41416=>"001110010",
  41417=>"001000110",
  41418=>"001111011",
  41419=>"001101010",
  41420=>"000001010",
  41421=>"011100110",
  41422=>"000010100",
  41423=>"110000101",
  41424=>"001000101",
  41425=>"110011100",
  41426=>"111011111",
  41427=>"100110010",
  41428=>"110111101",
  41429=>"110010001",
  41430=>"111110111",
  41431=>"011010110",
  41432=>"111000110",
  41433=>"110011011",
  41434=>"010001110",
  41435=>"000001110",
  41436=>"100110010",
  41437=>"001110111",
  41438=>"100011011",
  41439=>"000101001",
  41440=>"000011000",
  41441=>"101010110",
  41442=>"000001100",
  41443=>"100001110",
  41444=>"011001101",
  41445=>"001111110",
  41446=>"100001000",
  41447=>"011111101",
  41448=>"000000110",
  41449=>"001000111",
  41450=>"011001011",
  41451=>"111111001",
  41452=>"010011110",
  41453=>"011101110",
  41454=>"101000110",
  41455=>"110000110",
  41456=>"110011111",
  41457=>"100110110",
  41458=>"010010100",
  41459=>"011011011",
  41460=>"110110101",
  41461=>"011111100",
  41462=>"110010101",
  41463=>"101000011",
  41464=>"010011011",
  41465=>"110110000",
  41466=>"111111010",
  41467=>"100110101",
  41468=>"101110110",
  41469=>"000000101",
  41470=>"011101010",
  41471=>"111001101",
  41472=>"100101011",
  41473=>"100111011",
  41474=>"111100111",
  41475=>"111000000",
  41476=>"110100000",
  41477=>"100001010",
  41478=>"111001011",
  41479=>"011111110",
  41480=>"010001010",
  41481=>"011001000",
  41482=>"010110110",
  41483=>"101100010",
  41484=>"011011011",
  41485=>"101100000",
  41486=>"101111010",
  41487=>"001101101",
  41488=>"001000001",
  41489=>"010111111",
  41490=>"011001101",
  41491=>"101110000",
  41492=>"101110001",
  41493=>"000011101",
  41494=>"000010001",
  41495=>"010110111",
  41496=>"000101101",
  41497=>"100110110",
  41498=>"010100000",
  41499=>"111111110",
  41500=>"010100010",
  41501=>"111110010",
  41502=>"010100010",
  41503=>"001011011",
  41504=>"011000100",
  41505=>"001010101",
  41506=>"011010000",
  41507=>"111101100",
  41508=>"000010100",
  41509=>"000001111",
  41510=>"001010010",
  41511=>"111010011",
  41512=>"100011010",
  41513=>"010110110",
  41514=>"101000001",
  41515=>"010011010",
  41516=>"000101111",
  41517=>"000100111",
  41518=>"111111100",
  41519=>"101111101",
  41520=>"111010110",
  41521=>"101000010",
  41522=>"110111100",
  41523=>"011011111",
  41524=>"000000110",
  41525=>"001001000",
  41526=>"010101110",
  41527=>"110011011",
  41528=>"001100111",
  41529=>"101111101",
  41530=>"000110111",
  41531=>"100111000",
  41532=>"100001011",
  41533=>"111111000",
  41534=>"000101010",
  41535=>"001101100",
  41536=>"101101010",
  41537=>"111110010",
  41538=>"011000100",
  41539=>"011111111",
  41540=>"111100100",
  41541=>"101101101",
  41542=>"100000110",
  41543=>"101110010",
  41544=>"001100011",
  41545=>"010000111",
  41546=>"000010000",
  41547=>"010101111",
  41548=>"010100101",
  41549=>"100000010",
  41550=>"111000001",
  41551=>"111110010",
  41552=>"001101111",
  41553=>"010010000",
  41554=>"111011000",
  41555=>"001010010",
  41556=>"001001101",
  41557=>"001010101",
  41558=>"001000011",
  41559=>"100001000",
  41560=>"111101011",
  41561=>"101011011",
  41562=>"100111101",
  41563=>"100101011",
  41564=>"000111000",
  41565=>"101110001",
  41566=>"101110100",
  41567=>"111111011",
  41568=>"101111100",
  41569=>"111111001",
  41570=>"010111011",
  41571=>"010100001",
  41572=>"000011000",
  41573=>"111110100",
  41574=>"011110111",
  41575=>"111101111",
  41576=>"110011010",
  41577=>"100001110",
  41578=>"110100100",
  41579=>"101011110",
  41580=>"000000101",
  41581=>"100101110",
  41582=>"000010110",
  41583=>"100100111",
  41584=>"010100000",
  41585=>"111010001",
  41586=>"101110101",
  41587=>"000000000",
  41588=>"100010010",
  41589=>"000011110",
  41590=>"110111110",
  41591=>"000000101",
  41592=>"100001111",
  41593=>"100101011",
  41594=>"111110000",
  41595=>"110110011",
  41596=>"011101101",
  41597=>"100100000",
  41598=>"111100100",
  41599=>"000000101",
  41600=>"101010010",
  41601=>"111100110",
  41602=>"000010010",
  41603=>"010010100",
  41604=>"011001010",
  41605=>"011111100",
  41606=>"000001100",
  41607=>"001100110",
  41608=>"011000000",
  41609=>"101011010",
  41610=>"001001100",
  41611=>"111000111",
  41612=>"000101110",
  41613=>"010110011",
  41614=>"101101101",
  41615=>"001011100",
  41616=>"010001110",
  41617=>"101000000",
  41618=>"111100011",
  41619=>"010011101",
  41620=>"001000011",
  41621=>"101001011",
  41622=>"011010000",
  41623=>"010001111",
  41624=>"101011100",
  41625=>"001011111",
  41626=>"011011101",
  41627=>"111001101",
  41628=>"111110101",
  41629=>"000100110",
  41630=>"010001110",
  41631=>"111010101",
  41632=>"010100011",
  41633=>"010011100",
  41634=>"111111110",
  41635=>"100100000",
  41636=>"000011001",
  41637=>"011001010",
  41638=>"001000011",
  41639=>"100111100",
  41640=>"110000111",
  41641=>"100101100",
  41642=>"110110001",
  41643=>"100110110",
  41644=>"110101001",
  41645=>"011010011",
  41646=>"110010001",
  41647=>"011110111",
  41648=>"010001001",
  41649=>"101110110",
  41650=>"101101010",
  41651=>"001011010",
  41652=>"001001110",
  41653=>"010100001",
  41654=>"000110101",
  41655=>"001001001",
  41656=>"001110101",
  41657=>"001100010",
  41658=>"010001111",
  41659=>"110111110",
  41660=>"101101110",
  41661=>"100010010",
  41662=>"110001111",
  41663=>"000111011",
  41664=>"101110111",
  41665=>"000111100",
  41666=>"111100010",
  41667=>"101111111",
  41668=>"111001111",
  41669=>"111111110",
  41670=>"100100111",
  41671=>"010010110",
  41672=>"111001010",
  41673=>"110100100",
  41674=>"010101000",
  41675=>"010001011",
  41676=>"011111111",
  41677=>"010110000",
  41678=>"010110101",
  41679=>"000000001",
  41680=>"100111011",
  41681=>"010001111",
  41682=>"110011101",
  41683=>"100110111",
  41684=>"100001111",
  41685=>"000000010",
  41686=>"110111101",
  41687=>"011011100",
  41688=>"011100010",
  41689=>"010000101",
  41690=>"001001110",
  41691=>"111101111",
  41692=>"100011100",
  41693=>"111001000",
  41694=>"100001010",
  41695=>"111000000",
  41696=>"000110111",
  41697=>"011110110",
  41698=>"010001010",
  41699=>"101110100",
  41700=>"010001000",
  41701=>"110111111",
  41702=>"000001010",
  41703=>"010101110",
  41704=>"100001001",
  41705=>"010101001",
  41706=>"111101101",
  41707=>"010010001",
  41708=>"010100101",
  41709=>"110000001",
  41710=>"110010000",
  41711=>"001101101",
  41712=>"100111000",
  41713=>"000110000",
  41714=>"100001100",
  41715=>"000000010",
  41716=>"010000100",
  41717=>"010011110",
  41718=>"000011101",
  41719=>"011011101",
  41720=>"010110111",
  41721=>"100111111",
  41722=>"011000111",
  41723=>"000000110",
  41724=>"110010101",
  41725=>"111001101",
  41726=>"010001010",
  41727=>"000011101",
  41728=>"100111110",
  41729=>"010000101",
  41730=>"001011111",
  41731=>"001000011",
  41732=>"101011011",
  41733=>"001100000",
  41734=>"000110110",
  41735=>"110111011",
  41736=>"100001001",
  41737=>"011000100",
  41738=>"101011001",
  41739=>"100001010",
  41740=>"111010001",
  41741=>"101111110",
  41742=>"001000100",
  41743=>"101010110",
  41744=>"001011101",
  41745=>"100011111",
  41746=>"110100100",
  41747=>"001000101",
  41748=>"011010111",
  41749=>"100000000",
  41750=>"111111100",
  41751=>"111100111",
  41752=>"011001010",
  41753=>"110011011",
  41754=>"101001111",
  41755=>"000110011",
  41756=>"010000001",
  41757=>"010111011",
  41758=>"101101001",
  41759=>"011010011",
  41760=>"000000000",
  41761=>"111111101",
  41762=>"000001100",
  41763=>"110000000",
  41764=>"001001100",
  41765=>"010001000",
  41766=>"111011110",
  41767=>"010111110",
  41768=>"010100000",
  41769=>"100000100",
  41770=>"110100000",
  41771=>"101011100",
  41772=>"110100001",
  41773=>"000100001",
  41774=>"001111001",
  41775=>"011010110",
  41776=>"001010001",
  41777=>"111000110",
  41778=>"011001111",
  41779=>"100100011",
  41780=>"000111101",
  41781=>"101010111",
  41782=>"110000111",
  41783=>"101001101",
  41784=>"101101001",
  41785=>"100000111",
  41786=>"111101010",
  41787=>"111000010",
  41788=>"100011101",
  41789=>"010011100",
  41790=>"100011001",
  41791=>"001001011",
  41792=>"101011100",
  41793=>"110110100",
  41794=>"000001010",
  41795=>"011111100",
  41796=>"110110000",
  41797=>"100000010",
  41798=>"011010011",
  41799=>"010101011",
  41800=>"001111000",
  41801=>"001001110",
  41802=>"011100010",
  41803=>"010100010",
  41804=>"011010010",
  41805=>"110011111",
  41806=>"010010111",
  41807=>"111000111",
  41808=>"111011110",
  41809=>"010010100",
  41810=>"011111011",
  41811=>"010010101",
  41812=>"101010010",
  41813=>"010110011",
  41814=>"111001110",
  41815=>"110111011",
  41816=>"100110001",
  41817=>"011001111",
  41818=>"110101001",
  41819=>"010110010",
  41820=>"001000100",
  41821=>"111101101",
  41822=>"001000100",
  41823=>"000000101",
  41824=>"100111101",
  41825=>"101110010",
  41826=>"111001100",
  41827=>"100111100",
  41828=>"111011101",
  41829=>"110001100",
  41830=>"110100000",
  41831=>"111001110",
  41832=>"000111001",
  41833=>"000011110",
  41834=>"010100111",
  41835=>"100110010",
  41836=>"100100010",
  41837=>"111001101",
  41838=>"011111111",
  41839=>"110010011",
  41840=>"111110111",
  41841=>"011011110",
  41842=>"000001101",
  41843=>"010100101",
  41844=>"011100101",
  41845=>"000110111",
  41846=>"100011110",
  41847=>"001111101",
  41848=>"101101000",
  41849=>"010101010",
  41850=>"011010111",
  41851=>"001101100",
  41852=>"110010101",
  41853=>"011001111",
  41854=>"010111010",
  41855=>"010101001",
  41856=>"010101100",
  41857=>"000010000",
  41858=>"001001001",
  41859=>"000110101",
  41860=>"110111001",
  41861=>"001000001",
  41862=>"011000000",
  41863=>"110010100",
  41864=>"010001000",
  41865=>"011100111",
  41866=>"010100101",
  41867=>"000010000",
  41868=>"011111001",
  41869=>"011110010",
  41870=>"111111110",
  41871=>"101001110",
  41872=>"110011111",
  41873=>"110000111",
  41874=>"100011100",
  41875=>"000111111",
  41876=>"000001000",
  41877=>"001001100",
  41878=>"101111100",
  41879=>"110101000",
  41880=>"111010010",
  41881=>"000100001",
  41882=>"111011110",
  41883=>"001101010",
  41884=>"011101110",
  41885=>"000000000",
  41886=>"101011000",
  41887=>"111000011",
  41888=>"111101111",
  41889=>"110000011",
  41890=>"111110010",
  41891=>"111000100",
  41892=>"101000001",
  41893=>"100110001",
  41894=>"010010010",
  41895=>"110001010",
  41896=>"000001011",
  41897=>"000000110",
  41898=>"010111010",
  41899=>"011000110",
  41900=>"110110011",
  41901=>"011010111",
  41902=>"011011100",
  41903=>"111011000",
  41904=>"101101011",
  41905=>"010011111",
  41906=>"111111011",
  41907=>"111111110",
  41908=>"010101001",
  41909=>"100110111",
  41910=>"010110001",
  41911=>"001010101",
  41912=>"110001010",
  41913=>"100011000",
  41914=>"111110011",
  41915=>"100011000",
  41916=>"110001011",
  41917=>"111111111",
  41918=>"111100110",
  41919=>"010101110",
  41920=>"011010000",
  41921=>"101010001",
  41922=>"110101110",
  41923=>"101110100",
  41924=>"011000100",
  41925=>"011100011",
  41926=>"110101000",
  41927=>"101001010",
  41928=>"001001100",
  41929=>"000101000",
  41930=>"010010110",
  41931=>"111000001",
  41932=>"100111010",
  41933=>"101100011",
  41934=>"010110110",
  41935=>"111010101",
  41936=>"001101001",
  41937=>"101110010",
  41938=>"111101000",
  41939=>"101111101",
  41940=>"000100100",
  41941=>"001000010",
  41942=>"101001000",
  41943=>"011010111",
  41944=>"000111011",
  41945=>"111110111",
  41946=>"011110110",
  41947=>"100110001",
  41948=>"110000101",
  41949=>"110000011",
  41950=>"101000000",
  41951=>"110000100",
  41952=>"101101011",
  41953=>"011110110",
  41954=>"111101011",
  41955=>"010111001",
  41956=>"100100000",
  41957=>"111111111",
  41958=>"010001110",
  41959=>"000000101",
  41960=>"000011111",
  41961=>"000010101",
  41962=>"010001100",
  41963=>"010001001",
  41964=>"000111010",
  41965=>"111110000",
  41966=>"011000100",
  41967=>"001101000",
  41968=>"100011111",
  41969=>"100000100",
  41970=>"010011010",
  41971=>"010111011",
  41972=>"110011111",
  41973=>"010110001",
  41974=>"011011000",
  41975=>"010011111",
  41976=>"111111000",
  41977=>"001001010",
  41978=>"101110111",
  41979=>"101001000",
  41980=>"000110001",
  41981=>"000111010",
  41982=>"110101001",
  41983=>"001010001",
  41984=>"100100000",
  41985=>"100001110",
  41986=>"000100001",
  41987=>"111111100",
  41988=>"010111111",
  41989=>"001111100",
  41990=>"001011000",
  41991=>"001000100",
  41992=>"111011100",
  41993=>"101101111",
  41994=>"011101111",
  41995=>"000111110",
  41996=>"000101000",
  41997=>"110010100",
  41998=>"101100011",
  41999=>"111001111",
  42000=>"110111010",
  42001=>"111001011",
  42002=>"001001111",
  42003=>"000001010",
  42004=>"000001100",
  42005=>"011011110",
  42006=>"110011011",
  42007=>"011111010",
  42008=>"100000111",
  42009=>"101101000",
  42010=>"010100101",
  42011=>"000101000",
  42012=>"001101100",
  42013=>"111111011",
  42014=>"011000010",
  42015=>"011000000",
  42016=>"011000100",
  42017=>"001011011",
  42018=>"001101101",
  42019=>"001101000",
  42020=>"000000010",
  42021=>"001110111",
  42022=>"010011000",
  42023=>"011001000",
  42024=>"111000111",
  42025=>"000001011",
  42026=>"001000100",
  42027=>"110111011",
  42028=>"011010101",
  42029=>"100111010",
  42030=>"100010010",
  42031=>"101110110",
  42032=>"110101001",
  42033=>"010110010",
  42034=>"011011010",
  42035=>"100000101",
  42036=>"101010001",
  42037=>"100110100",
  42038=>"001100011",
  42039=>"011010001",
  42040=>"000000011",
  42041=>"001000010",
  42042=>"101101010",
  42043=>"000001000",
  42044=>"100111101",
  42045=>"011011000",
  42046=>"000010110",
  42047=>"101110110",
  42048=>"100000110",
  42049=>"000110000",
  42050=>"000100000",
  42051=>"011010100",
  42052=>"101011011",
  42053=>"111000110",
  42054=>"000000011",
  42055=>"010101100",
  42056=>"000010000",
  42057=>"110101011",
  42058=>"101011111",
  42059=>"000011000",
  42060=>"101001101",
  42061=>"111111101",
  42062=>"010111001",
  42063=>"011000100",
  42064=>"010011111",
  42065=>"101101110",
  42066=>"100001000",
  42067=>"001100110",
  42068=>"111000010",
  42069=>"101000110",
  42070=>"011111011",
  42071=>"011000011",
  42072=>"000111111",
  42073=>"110111001",
  42074=>"101110101",
  42075=>"000110101",
  42076=>"011110110",
  42077=>"110111011",
  42078=>"001110000",
  42079=>"100100110",
  42080=>"111111100",
  42081=>"000110001",
  42082=>"101110010",
  42083=>"101001100",
  42084=>"010010011",
  42085=>"100010000",
  42086=>"011011000",
  42087=>"110010100",
  42088=>"101111101",
  42089=>"100000110",
  42090=>"000011101",
  42091=>"111110000",
  42092=>"010111010",
  42093=>"010110100",
  42094=>"100110011",
  42095=>"101111011",
  42096=>"110000010",
  42097=>"010111000",
  42098=>"000110100",
  42099=>"101110010",
  42100=>"001111010",
  42101=>"100111110",
  42102=>"001001110",
  42103=>"000100010",
  42104=>"010011101",
  42105=>"110111110",
  42106=>"110110111",
  42107=>"000000100",
  42108=>"000011111",
  42109=>"111000011",
  42110=>"010010101",
  42111=>"011000111",
  42112=>"000000100",
  42113=>"110111111",
  42114=>"001100011",
  42115=>"101110000",
  42116=>"000010000",
  42117=>"000010101",
  42118=>"111011101",
  42119=>"111111001",
  42120=>"110001000",
  42121=>"101111010",
  42122=>"110110111",
  42123=>"110011000",
  42124=>"010101111",
  42125=>"010011001",
  42126=>"010000001",
  42127=>"010010010",
  42128=>"011000001",
  42129=>"010011111",
  42130=>"101101111",
  42131=>"110100001",
  42132=>"011001011",
  42133=>"101010000",
  42134=>"111011101",
  42135=>"000110111",
  42136=>"110100111",
  42137=>"100111100",
  42138=>"110010000",
  42139=>"001101000",
  42140=>"110101000",
  42141=>"001011010",
  42142=>"100101100",
  42143=>"000111110",
  42144=>"001111010",
  42145=>"011101000",
  42146=>"110111000",
  42147=>"000011111",
  42148=>"110110111",
  42149=>"111111010",
  42150=>"111110010",
  42151=>"111000100",
  42152=>"111111100",
  42153=>"101010011",
  42154=>"001101110",
  42155=>"000000011",
  42156=>"101000100",
  42157=>"000010101",
  42158=>"001100000",
  42159=>"011010110",
  42160=>"010011000",
  42161=>"010111111",
  42162=>"100000101",
  42163=>"001000100",
  42164=>"001001000",
  42165=>"101111111",
  42166=>"111101100",
  42167=>"011110111",
  42168=>"010011101",
  42169=>"010110111",
  42170=>"001111000",
  42171=>"011001100",
  42172=>"110011101",
  42173=>"010101010",
  42174=>"101011111",
  42175=>"000100100",
  42176=>"100001111",
  42177=>"010111100",
  42178=>"011000010",
  42179=>"100000001",
  42180=>"000010110",
  42181=>"100111110",
  42182=>"100101001",
  42183=>"110010101",
  42184=>"100110101",
  42185=>"101001010",
  42186=>"100111101",
  42187=>"111001000",
  42188=>"110010110",
  42189=>"110110100",
  42190=>"110110001",
  42191=>"011100101",
  42192=>"010010111",
  42193=>"010110101",
  42194=>"101000100",
  42195=>"101101110",
  42196=>"001101100",
  42197=>"000111100",
  42198=>"011111101",
  42199=>"000000000",
  42200=>"001001101",
  42201=>"110010101",
  42202=>"110001101",
  42203=>"010000011",
  42204=>"001001001",
  42205=>"010010110",
  42206=>"101111010",
  42207=>"011110000",
  42208=>"001101000",
  42209=>"011111111",
  42210=>"111101011",
  42211=>"000101010",
  42212=>"111110110",
  42213=>"101000110",
  42214=>"100011100",
  42215=>"101100010",
  42216=>"111100000",
  42217=>"101011100",
  42218=>"110111000",
  42219=>"011001011",
  42220=>"001011001",
  42221=>"001111000",
  42222=>"010010110",
  42223=>"010000110",
  42224=>"110001111",
  42225=>"110110010",
  42226=>"011001100",
  42227=>"101111001",
  42228=>"100110100",
  42229=>"100010011",
  42230=>"111100101",
  42231=>"001101011",
  42232=>"100100000",
  42233=>"000000101",
  42234=>"110101110",
  42235=>"101010011",
  42236=>"100101100",
  42237=>"111111101",
  42238=>"011011110",
  42239=>"000010011",
  42240=>"010101100",
  42241=>"110010111",
  42242=>"011101101",
  42243=>"010110000",
  42244=>"100010111",
  42245=>"110000010",
  42246=>"111001111",
  42247=>"001010101",
  42248=>"111101111",
  42249=>"010010001",
  42250=>"101101000",
  42251=>"010010101",
  42252=>"000100011",
  42253=>"100010010",
  42254=>"100010101",
  42255=>"101001010",
  42256=>"100100111",
  42257=>"110110010",
  42258=>"100000000",
  42259=>"111001011",
  42260=>"001000000",
  42261=>"011100101",
  42262=>"110001110",
  42263=>"111100001",
  42264=>"101000011",
  42265=>"001001101",
  42266=>"100101110",
  42267=>"101111010",
  42268=>"111000010",
  42269=>"100101100",
  42270=>"010110010",
  42271=>"101111001",
  42272=>"000111100",
  42273=>"110100110",
  42274=>"001011001",
  42275=>"101011001",
  42276=>"000011110",
  42277=>"010010000",
  42278=>"101100001",
  42279=>"011110001",
  42280=>"001001011",
  42281=>"110110001",
  42282=>"001000000",
  42283=>"000000001",
  42284=>"110010101",
  42285=>"000100111",
  42286=>"001000110",
  42287=>"111001110",
  42288=>"101111110",
  42289=>"010010001",
  42290=>"001110111",
  42291=>"000111010",
  42292=>"010111110",
  42293=>"001101111",
  42294=>"110000100",
  42295=>"110111111",
  42296=>"100100000",
  42297=>"011000000",
  42298=>"100000111",
  42299=>"110000101",
  42300=>"011100000",
  42301=>"110111101",
  42302=>"111100011",
  42303=>"101111011",
  42304=>"100011000",
  42305=>"110010000",
  42306=>"000000010",
  42307=>"111101111",
  42308=>"011111001",
  42309=>"100011000",
  42310=>"101001010",
  42311=>"111101100",
  42312=>"000100100",
  42313=>"110000011",
  42314=>"111010001",
  42315=>"111000110",
  42316=>"011010110",
  42317=>"000100001",
  42318=>"100000010",
  42319=>"000000100",
  42320=>"101000100",
  42321=>"110101110",
  42322=>"111000111",
  42323=>"110111101",
  42324=>"111100011",
  42325=>"010010010",
  42326=>"110101010",
  42327=>"110111000",
  42328=>"000000010",
  42329=>"010101100",
  42330=>"111101100",
  42331=>"100001000",
  42332=>"111011100",
  42333=>"101111111",
  42334=>"010001011",
  42335=>"000010001",
  42336=>"011000011",
  42337=>"100111110",
  42338=>"000000000",
  42339=>"000010101",
  42340=>"011101010",
  42341=>"100100100",
  42342=>"111000100",
  42343=>"101000000",
  42344=>"001000000",
  42345=>"111111011",
  42346=>"110010110",
  42347=>"010001000",
  42348=>"100011000",
  42349=>"111111010",
  42350=>"010100010",
  42351=>"101111000",
  42352=>"001101101",
  42353=>"000000110",
  42354=>"001011011",
  42355=>"111000110",
  42356=>"100100011",
  42357=>"011111111",
  42358=>"000010010",
  42359=>"011101000",
  42360=>"101110110",
  42361=>"100010100",
  42362=>"100111100",
  42363=>"010101101",
  42364=>"010100111",
  42365=>"101100111",
  42366=>"110001100",
  42367=>"011100111",
  42368=>"011111111",
  42369=>"001000100",
  42370=>"111110011",
  42371=>"110111100",
  42372=>"100111011",
  42373=>"001001100",
  42374=>"011000111",
  42375=>"010111101",
  42376=>"011010011",
  42377=>"001100111",
  42378=>"011001110",
  42379=>"111011100",
  42380=>"101110001",
  42381=>"100000000",
  42382=>"111000000",
  42383=>"000000001",
  42384=>"010000111",
  42385=>"101100101",
  42386=>"110110000",
  42387=>"001100011",
  42388=>"001101001",
  42389=>"000110010",
  42390=>"010100011",
  42391=>"100110100",
  42392=>"011011011",
  42393=>"111101111",
  42394=>"010101010",
  42395=>"010100110",
  42396=>"000010010",
  42397=>"100111111",
  42398=>"010000111",
  42399=>"100000000",
  42400=>"010010100",
  42401=>"100111010",
  42402=>"000111011",
  42403=>"110001010",
  42404=>"011111110",
  42405=>"010001100",
  42406=>"001011001",
  42407=>"101110011",
  42408=>"101011111",
  42409=>"001011011",
  42410=>"010001001",
  42411=>"000001110",
  42412=>"000001100",
  42413=>"110110001",
  42414=>"100101000",
  42415=>"000010001",
  42416=>"001110110",
  42417=>"010110110",
  42418=>"101101111",
  42419=>"011011101",
  42420=>"001100100",
  42421=>"011000000",
  42422=>"100100000",
  42423=>"000111101",
  42424=>"111001010",
  42425=>"011011110",
  42426=>"111100001",
  42427=>"111111100",
  42428=>"111111010",
  42429=>"000100100",
  42430=>"011111100",
  42431=>"111100011",
  42432=>"001100100",
  42433=>"001000101",
  42434=>"111001111",
  42435=>"001001011",
  42436=>"110111100",
  42437=>"000110111",
  42438=>"011101111",
  42439=>"000100000",
  42440=>"100000000",
  42441=>"110010110",
  42442=>"101010001",
  42443=>"011011110",
  42444=>"010000110",
  42445=>"111010001",
  42446=>"010010100",
  42447=>"010111000",
  42448=>"011010010",
  42449=>"110110100",
  42450=>"100001110",
  42451=>"111100011",
  42452=>"001101110",
  42453=>"000000000",
  42454=>"001111000",
  42455=>"010000111",
  42456=>"000010111",
  42457=>"100111111",
  42458=>"101011111",
  42459=>"110000101",
  42460=>"001110010",
  42461=>"110110111",
  42462=>"001110001",
  42463=>"010000111",
  42464=>"101000001",
  42465=>"111001000",
  42466=>"101011010",
  42467=>"110110011",
  42468=>"100100010",
  42469=>"101111110",
  42470=>"000101010",
  42471=>"010011001",
  42472=>"001001110",
  42473=>"110110111",
  42474=>"111010001",
  42475=>"100110000",
  42476=>"000010110",
  42477=>"111011000",
  42478=>"110111100",
  42479=>"010111101",
  42480=>"011100001",
  42481=>"110111010",
  42482=>"110001111",
  42483=>"100111100",
  42484=>"101000100",
  42485=>"000001011",
  42486=>"100101110",
  42487=>"000111001",
  42488=>"011000101",
  42489=>"001000110",
  42490=>"010000001",
  42491=>"001011011",
  42492=>"111111101",
  42493=>"111001010",
  42494=>"010000001",
  42495=>"110000001",
  42496=>"010001010",
  42497=>"000000011",
  42498=>"110011011",
  42499=>"001001000",
  42500=>"010010001",
  42501=>"111001010",
  42502=>"001111111",
  42503=>"000000010",
  42504=>"110101011",
  42505=>"111111110",
  42506=>"010001001",
  42507=>"011001100",
  42508=>"001001000",
  42509=>"110001001",
  42510=>"110111100",
  42511=>"111101100",
  42512=>"110110111",
  42513=>"100111111",
  42514=>"000101010",
  42515=>"011010111",
  42516=>"100000110",
  42517=>"001110110",
  42518=>"110101001",
  42519=>"101010000",
  42520=>"111010010",
  42521=>"001001001",
  42522=>"010000100",
  42523=>"101011110",
  42524=>"000001110",
  42525=>"000101010",
  42526=>"011111011",
  42527=>"101011010",
  42528=>"010000101",
  42529=>"101111100",
  42530=>"001000011",
  42531=>"011101101",
  42532=>"101111000",
  42533=>"111101010",
  42534=>"101001011",
  42535=>"000000111",
  42536=>"100000101",
  42537=>"111001110",
  42538=>"011110010",
  42539=>"001000110",
  42540=>"000100001",
  42541=>"000001000",
  42542=>"000110000",
  42543=>"101100011",
  42544=>"000110100",
  42545=>"100001110",
  42546=>"101011100",
  42547=>"111010011",
  42548=>"111000111",
  42549=>"001101101",
  42550=>"110111101",
  42551=>"100110010",
  42552=>"110011111",
  42553=>"101111110",
  42554=>"101110001",
  42555=>"001110100",
  42556=>"001000111",
  42557=>"001101111",
  42558=>"110010010",
  42559=>"110100000",
  42560=>"010001101",
  42561=>"110010100",
  42562=>"111101011",
  42563=>"100011010",
  42564=>"110000111",
  42565=>"101100111",
  42566=>"010001000",
  42567=>"000001110",
  42568=>"010000000",
  42569=>"100000010",
  42570=>"111000001",
  42571=>"010001011",
  42572=>"110010010",
  42573=>"011110111",
  42574=>"111011000",
  42575=>"011011010",
  42576=>"100110111",
  42577=>"101001011",
  42578=>"100000010",
  42579=>"101000011",
  42580=>"001011100",
  42581=>"101000101",
  42582=>"100101101",
  42583=>"100110010",
  42584=>"110111101",
  42585=>"100011110",
  42586=>"000101011",
  42587=>"000000101",
  42588=>"010011111",
  42589=>"000110001",
  42590=>"000111101",
  42591=>"001111010",
  42592=>"111010100",
  42593=>"000101000",
  42594=>"011100101",
  42595=>"101100101",
  42596=>"011000111",
  42597=>"000011010",
  42598=>"000100010",
  42599=>"001001001",
  42600=>"000000010",
  42601=>"010001111",
  42602=>"110101001",
  42603=>"011101011",
  42604=>"100010010",
  42605=>"000010110",
  42606=>"001000000",
  42607=>"001100011",
  42608=>"100001001",
  42609=>"111101000",
  42610=>"100110100",
  42611=>"010100001",
  42612=>"000000100",
  42613=>"000101100",
  42614=>"001100101",
  42615=>"110101100",
  42616=>"100011000",
  42617=>"100011011",
  42618=>"110111001",
  42619=>"000001000",
  42620=>"101101010",
  42621=>"110100011",
  42622=>"110100111",
  42623=>"101001100",
  42624=>"101001101",
  42625=>"101011011",
  42626=>"011110010",
  42627=>"111101110",
  42628=>"000110100",
  42629=>"101011011",
  42630=>"000000101",
  42631=>"111111111",
  42632=>"001000110",
  42633=>"001001100",
  42634=>"111100000",
  42635=>"100000011",
  42636=>"001000000",
  42637=>"100001001",
  42638=>"001100101",
  42639=>"110011000",
  42640=>"001101000",
  42641=>"010101011",
  42642=>"100000000",
  42643=>"010011111",
  42644=>"010100110",
  42645=>"001010010",
  42646=>"101101001",
  42647=>"011110000",
  42648=>"010000001",
  42649=>"010100001",
  42650=>"010110011",
  42651=>"111001010",
  42652=>"001011111",
  42653=>"010001001",
  42654=>"111010111",
  42655=>"100011100",
  42656=>"011001000",
  42657=>"010100001",
  42658=>"011101000",
  42659=>"001100101",
  42660=>"010110111",
  42661=>"010111110",
  42662=>"000101000",
  42663=>"001000110",
  42664=>"010111101",
  42665=>"111111000",
  42666=>"110001111",
  42667=>"000100101",
  42668=>"001000110",
  42669=>"101110101",
  42670=>"100111110",
  42671=>"101010100",
  42672=>"000110010",
  42673=>"010110100",
  42674=>"111011111",
  42675=>"000000110",
  42676=>"010001110",
  42677=>"011011110",
  42678=>"011011000",
  42679=>"110000010",
  42680=>"100000110",
  42681=>"110101011",
  42682=>"000001100",
  42683=>"001000111",
  42684=>"011100111",
  42685=>"010011001",
  42686=>"000000110",
  42687=>"011100110",
  42688=>"011111011",
  42689=>"110010110",
  42690=>"110001101",
  42691=>"001011001",
  42692=>"100111100",
  42693=>"010101101",
  42694=>"100111010",
  42695=>"100001111",
  42696=>"000100000",
  42697=>"001110111",
  42698=>"111101110",
  42699=>"000001000",
  42700=>"100110000",
  42701=>"101011111",
  42702=>"100100001",
  42703=>"110000101",
  42704=>"001000101",
  42705=>"100011111",
  42706=>"000001000",
  42707=>"010011000",
  42708=>"001010111",
  42709=>"000111111",
  42710=>"100111101",
  42711=>"100100111",
  42712=>"100101001",
  42713=>"100111000",
  42714=>"001000100",
  42715=>"111110100",
  42716=>"110001111",
  42717=>"110001000",
  42718=>"011111100",
  42719=>"000001111",
  42720=>"000100011",
  42721=>"001101110",
  42722=>"001011100",
  42723=>"001110011",
  42724=>"101101110",
  42725=>"010110000",
  42726=>"001000001",
  42727=>"011000111",
  42728=>"101100110",
  42729=>"011101011",
  42730=>"011000001",
  42731=>"010100001",
  42732=>"000100000",
  42733=>"000100100",
  42734=>"011110100",
  42735=>"000100100",
  42736=>"111011010",
  42737=>"001101000",
  42738=>"001100100",
  42739=>"010111000",
  42740=>"000010001",
  42741=>"111110011",
  42742=>"011011100",
  42743=>"011111111",
  42744=>"000001101",
  42745=>"101010100",
  42746=>"011100000",
  42747=>"000001001",
  42748=>"100101111",
  42749=>"001111010",
  42750=>"110001001",
  42751=>"100101010",
  42752=>"010111101",
  42753=>"111101100",
  42754=>"011000010",
  42755=>"100001000",
  42756=>"001110111",
  42757=>"011101011",
  42758=>"001100011",
  42759=>"100110001",
  42760=>"011101110",
  42761=>"001010011",
  42762=>"011011000",
  42763=>"100010010",
  42764=>"000111010",
  42765=>"001110001",
  42766=>"111000000",
  42767=>"001000010",
  42768=>"011000000",
  42769=>"000001000",
  42770=>"100111110",
  42771=>"101000111",
  42772=>"011001101",
  42773=>"110101010",
  42774=>"010011010",
  42775=>"011001101",
  42776=>"110110110",
  42777=>"110111000",
  42778=>"100010110",
  42779=>"111111101",
  42780=>"000010010",
  42781=>"000001100",
  42782=>"101110001",
  42783=>"000100100",
  42784=>"011001110",
  42785=>"000100011",
  42786=>"100010001",
  42787=>"100001100",
  42788=>"101110010",
  42789=>"000000010",
  42790=>"010100100",
  42791=>"101100100",
  42792=>"111111110",
  42793=>"111100001",
  42794=>"111111111",
  42795=>"010011010",
  42796=>"001101001",
  42797=>"000110111",
  42798=>"010011010",
  42799=>"100000011",
  42800=>"101000101",
  42801=>"010100001",
  42802=>"111001000",
  42803=>"011100111",
  42804=>"101011101",
  42805=>"001000011",
  42806=>"110101100",
  42807=>"111111110",
  42808=>"111111001",
  42809=>"000010011",
  42810=>"001000111",
  42811=>"111110101",
  42812=>"111111111",
  42813=>"000000111",
  42814=>"010010110",
  42815=>"100110101",
  42816=>"111011110",
  42817=>"011000110",
  42818=>"000101000",
  42819=>"011000100",
  42820=>"100000100",
  42821=>"011000111",
  42822=>"100000010",
  42823=>"110010000",
  42824=>"011101100",
  42825=>"111100011",
  42826=>"000101001",
  42827=>"101011011",
  42828=>"010000010",
  42829=>"001100000",
  42830=>"100001000",
  42831=>"110011000",
  42832=>"000110001",
  42833=>"101100111",
  42834=>"010101011",
  42835=>"011110101",
  42836=>"000111110",
  42837=>"001111110",
  42838=>"111011000",
  42839=>"101001110",
  42840=>"111111101",
  42841=>"100110100",
  42842=>"010000111",
  42843=>"000001110",
  42844=>"000111010",
  42845=>"001010010",
  42846=>"100010101",
  42847=>"000001111",
  42848=>"000111010",
  42849=>"001100110",
  42850=>"000000011",
  42851=>"010001111",
  42852=>"000011101",
  42853=>"010101000",
  42854=>"100100100",
  42855=>"100101110",
  42856=>"000010101",
  42857=>"110110001",
  42858=>"000100111",
  42859=>"011001001",
  42860=>"111110100",
  42861=>"101111100",
  42862=>"000101011",
  42863=>"010110100",
  42864=>"111010100",
  42865=>"000100101",
  42866=>"100101101",
  42867=>"111011011",
  42868=>"010000010",
  42869=>"110100000",
  42870=>"100100010",
  42871=>"110001000",
  42872=>"110110001",
  42873=>"100110100",
  42874=>"001011001",
  42875=>"010100001",
  42876=>"100110100",
  42877=>"100110110",
  42878=>"100001010",
  42879=>"100001111",
  42880=>"000010010",
  42881=>"111100011",
  42882=>"110000010",
  42883=>"011110100",
  42884=>"011001001",
  42885=>"001101000",
  42886=>"110111111",
  42887=>"100011000",
  42888=>"100111111",
  42889=>"000010011",
  42890=>"001100111",
  42891=>"101100010",
  42892=>"001011111",
  42893=>"100101100",
  42894=>"001010111",
  42895=>"010011011",
  42896=>"000011011",
  42897=>"010100000",
  42898=>"100001000",
  42899=>"011000100",
  42900=>"010000110",
  42901=>"110001011",
  42902=>"001011001",
  42903=>"101000011",
  42904=>"000000100",
  42905=>"011111101",
  42906=>"000101000",
  42907=>"001110100",
  42908=>"111010010",
  42909=>"000101001",
  42910=>"111100111",
  42911=>"111110000",
  42912=>"000110001",
  42913=>"101111101",
  42914=>"111100101",
  42915=>"111100111",
  42916=>"001110011",
  42917=>"001101101",
  42918=>"110001011",
  42919=>"111011001",
  42920=>"011001100",
  42921=>"000010000",
  42922=>"010001100",
  42923=>"101111111",
  42924=>"001100000",
  42925=>"011110110",
  42926=>"001100001",
  42927=>"000101001",
  42928=>"101100001",
  42929=>"000111111",
  42930=>"011001110",
  42931=>"001100111",
  42932=>"111110111",
  42933=>"110001011",
  42934=>"001100000",
  42935=>"110000010",
  42936=>"010111111",
  42937=>"100101101",
  42938=>"110001001",
  42939=>"011111110",
  42940=>"111110010",
  42941=>"101101111",
  42942=>"000010010",
  42943=>"000100110",
  42944=>"101000011",
  42945=>"110101011",
  42946=>"011001000",
  42947=>"000101110",
  42948=>"111011010",
  42949=>"011110001",
  42950=>"000010010",
  42951=>"101001010",
  42952=>"011011011",
  42953=>"101000101",
  42954=>"011000000",
  42955=>"111001011",
  42956=>"110011101",
  42957=>"010001001",
  42958=>"111111111",
  42959=>"001110001",
  42960=>"001001011",
  42961=>"010100101",
  42962=>"010000110",
  42963=>"100010101",
  42964=>"110110110",
  42965=>"001100100",
  42966=>"000101110",
  42967=>"001001111",
  42968=>"110110000",
  42969=>"101011101",
  42970=>"011100101",
  42971=>"000000000",
  42972=>"001100101",
  42973=>"111000000",
  42974=>"100011110",
  42975=>"010011110",
  42976=>"100111001",
  42977=>"011101110",
  42978=>"101100010",
  42979=>"100110000",
  42980=>"100011001",
  42981=>"111001000",
  42982=>"001000000",
  42983=>"000100101",
  42984=>"000100010",
  42985=>"011010111",
  42986=>"011000001",
  42987=>"010101100",
  42988=>"110110101",
  42989=>"100001011",
  42990=>"111010110",
  42991=>"111011001",
  42992=>"011111101",
  42993=>"100100110",
  42994=>"010001000",
  42995=>"111010110",
  42996=>"010000011",
  42997=>"111110101",
  42998=>"100111011",
  42999=>"110101000",
  43000=>"110111001",
  43001=>"011001011",
  43002=>"001110010",
  43003=>"011111100",
  43004=>"000101011",
  43005=>"101100000",
  43006=>"101011000",
  43007=>"100011000",
  43008=>"000000110",
  43009=>"000011101",
  43010=>"111000110",
  43011=>"010011011",
  43012=>"111110010",
  43013=>"010101100",
  43014=>"001011111",
  43015=>"001000000",
  43016=>"011111110",
  43017=>"101001011",
  43018=>"001010111",
  43019=>"001001011",
  43020=>"100101000",
  43021=>"101110101",
  43022=>"001101000",
  43023=>"001001011",
  43024=>"001001001",
  43025=>"000000000",
  43026=>"010011010",
  43027=>"101000011",
  43028=>"011101010",
  43029=>"100101011",
  43030=>"011011010",
  43031=>"001101000",
  43032=>"001011000",
  43033=>"001110010",
  43034=>"110100100",
  43035=>"010001000",
  43036=>"011000111",
  43037=>"011101100",
  43038=>"110100000",
  43039=>"111011101",
  43040=>"010001110",
  43041=>"100100010",
  43042=>"001001000",
  43043=>"100000101",
  43044=>"001111010",
  43045=>"110000110",
  43046=>"111101001",
  43047=>"100010001",
  43048=>"101010001",
  43049=>"010101001",
  43050=>"010110101",
  43051=>"000101101",
  43052=>"101011001",
  43053=>"010110011",
  43054=>"111011110",
  43055=>"100010101",
  43056=>"010010111",
  43057=>"111110110",
  43058=>"101101111",
  43059=>"010100001",
  43060=>"001001000",
  43061=>"010100011",
  43062=>"011011011",
  43063=>"100001110",
  43064=>"010101100",
  43065=>"000011011",
  43066=>"100111001",
  43067=>"000010001",
  43068=>"111100000",
  43069=>"111110100",
  43070=>"110010111",
  43071=>"110010010",
  43072=>"011000011",
  43073=>"110101010",
  43074=>"011001000",
  43075=>"011100011",
  43076=>"001001000",
  43077=>"011010111",
  43078=>"010001000",
  43079=>"000010010",
  43080=>"101100000",
  43081=>"111010000",
  43082=>"000011101",
  43083=>"000000111",
  43084=>"100001011",
  43085=>"000111000",
  43086=>"011100010",
  43087=>"100011010",
  43088=>"010001001",
  43089=>"101001010",
  43090=>"111010101",
  43091=>"010110000",
  43092=>"100000010",
  43093=>"010100000",
  43094=>"010001001",
  43095=>"001100000",
  43096=>"010000011",
  43097=>"001011110",
  43098=>"000010000",
  43099=>"011001001",
  43100=>"000111000",
  43101=>"001010010",
  43102=>"111010111",
  43103=>"011000110",
  43104=>"001001000",
  43105=>"100110000",
  43106=>"110000010",
  43107=>"000111101",
  43108=>"010000000",
  43109=>"000000000",
  43110=>"000011101",
  43111=>"100010101",
  43112=>"010100001",
  43113=>"011010101",
  43114=>"100010100",
  43115=>"001111101",
  43116=>"010100101",
  43117=>"010100010",
  43118=>"110110001",
  43119=>"111110010",
  43120=>"011000101",
  43121=>"011010001",
  43122=>"110111010",
  43123=>"011010101",
  43124=>"011110011",
  43125=>"100001111",
  43126=>"001101111",
  43127=>"001000001",
  43128=>"100110101",
  43129=>"010110111",
  43130=>"000000101",
  43131=>"100000110",
  43132=>"010101101",
  43133=>"000110010",
  43134=>"100111100",
  43135=>"010011000",
  43136=>"000000000",
  43137=>"011100010",
  43138=>"010111101",
  43139=>"101110001",
  43140=>"111001001",
  43141=>"111110101",
  43142=>"101001011",
  43143=>"000100110",
  43144=>"100011101",
  43145=>"100101111",
  43146=>"001101000",
  43147=>"110110110",
  43148=>"000001001",
  43149=>"001101100",
  43150=>"101111101",
  43151=>"010001110",
  43152=>"010001111",
  43153=>"110100011",
  43154=>"011101011",
  43155=>"100010110",
  43156=>"010001000",
  43157=>"111010001",
  43158=>"000001000",
  43159=>"100000101",
  43160=>"110100010",
  43161=>"101000101",
  43162=>"010100010",
  43163=>"100001010",
  43164=>"101001001",
  43165=>"000010000",
  43166=>"101000101",
  43167=>"111111010",
  43168=>"011001000",
  43169=>"111100110",
  43170=>"101010010",
  43171=>"000001110",
  43172=>"010110110",
  43173=>"000101111",
  43174=>"010010100",
  43175=>"111101000",
  43176=>"010110011",
  43177=>"100110000",
  43178=>"100110101",
  43179=>"011111101",
  43180=>"100000000",
  43181=>"110100000",
  43182=>"011100111",
  43183=>"000001010",
  43184=>"110100011",
  43185=>"011101001",
  43186=>"000011111",
  43187=>"011001001",
  43188=>"101111001",
  43189=>"010100001",
  43190=>"111100001",
  43191=>"010110100",
  43192=>"001000100",
  43193=>"100110010",
  43194=>"111111110",
  43195=>"011011100",
  43196=>"010010100",
  43197=>"011111001",
  43198=>"110001011",
  43199=>"110011001",
  43200=>"110110001",
  43201=>"110000010",
  43202=>"011011010",
  43203=>"000110000",
  43204=>"011000001",
  43205=>"110011011",
  43206=>"101101000",
  43207=>"101010000",
  43208=>"011100001",
  43209=>"001101111",
  43210=>"001010001",
  43211=>"100111000",
  43212=>"101111001",
  43213=>"011110101",
  43214=>"000010010",
  43215=>"000011100",
  43216=>"110110001",
  43217=>"001111011",
  43218=>"101101011",
  43219=>"100001100",
  43220=>"101000100",
  43221=>"101111010",
  43222=>"011110110",
  43223=>"001111101",
  43224=>"001001001",
  43225=>"001110001",
  43226=>"011110000",
  43227=>"000101001",
  43228=>"011010101",
  43229=>"001011000",
  43230=>"111011100",
  43231=>"100010000",
  43232=>"100001010",
  43233=>"010101011",
  43234=>"010010101",
  43235=>"110000011",
  43236=>"000010100",
  43237=>"001100010",
  43238=>"000000111",
  43239=>"010011100",
  43240=>"010101101",
  43241=>"100101011",
  43242=>"111011111",
  43243=>"001000110",
  43244=>"000000101",
  43245=>"000010001",
  43246=>"110101001",
  43247=>"101110010",
  43248=>"110111011",
  43249=>"101010000",
  43250=>"111100100",
  43251=>"100001011",
  43252=>"111001001",
  43253=>"011100111",
  43254=>"101001100",
  43255=>"111111101",
  43256=>"000011011",
  43257=>"111000111",
  43258=>"110111000",
  43259=>"000001001",
  43260=>"000100101",
  43261=>"110100110",
  43262=>"111111110",
  43263=>"000000110",
  43264=>"110010100",
  43265=>"010011100",
  43266=>"111100000",
  43267=>"011010111",
  43268=>"101101010",
  43269=>"101001110",
  43270=>"010100111",
  43271=>"100011010",
  43272=>"010111011",
  43273=>"110110000",
  43274=>"111101010",
  43275=>"001101110",
  43276=>"000101101",
  43277=>"100001111",
  43278=>"111001100",
  43279=>"000000010",
  43280=>"010011111",
  43281=>"011001110",
  43282=>"110110110",
  43283=>"011000100",
  43284=>"111101001",
  43285=>"001110110",
  43286=>"111000000",
  43287=>"101101010",
  43288=>"101101011",
  43289=>"110000000",
  43290=>"011000000",
  43291=>"000000110",
  43292=>"000111000",
  43293=>"110111100",
  43294=>"110011011",
  43295=>"001101001",
  43296=>"001000100",
  43297=>"010111010",
  43298=>"000111111",
  43299=>"110101010",
  43300=>"100110001",
  43301=>"011110111",
  43302=>"000000111",
  43303=>"110110011",
  43304=>"010000111",
  43305=>"011110100",
  43306=>"011101110",
  43307=>"100100000",
  43308=>"000001101",
  43309=>"001000010",
  43310=>"000101101",
  43311=>"100011011",
  43312=>"010110100",
  43313=>"110001010",
  43314=>"111011010",
  43315=>"100010000",
  43316=>"110110100",
  43317=>"001101010",
  43318=>"010111000",
  43319=>"111001100",
  43320=>"100101101",
  43321=>"111110001",
  43322=>"110001110",
  43323=>"010000100",
  43324=>"101110001",
  43325=>"110001110",
  43326=>"001000101",
  43327=>"001101000",
  43328=>"001101011",
  43329=>"101011101",
  43330=>"001111100",
  43331=>"100101101",
  43332=>"000100001",
  43333=>"101111001",
  43334=>"111011001",
  43335=>"101101101",
  43336=>"000100111",
  43337=>"111011010",
  43338=>"011111110",
  43339=>"000000000",
  43340=>"001110110",
  43341=>"001101001",
  43342=>"010001000",
  43343=>"111101101",
  43344=>"010101001",
  43345=>"011111001",
  43346=>"111101001",
  43347=>"000000110",
  43348=>"101001011",
  43349=>"111011011",
  43350=>"100100110",
  43351=>"100010010",
  43352=>"010000000",
  43353=>"101100110",
  43354=>"111110010",
  43355=>"111011101",
  43356=>"100111101",
  43357=>"111101100",
  43358=>"010001110",
  43359=>"110100100",
  43360=>"110111100",
  43361=>"000111110",
  43362=>"001110101",
  43363=>"001000110",
  43364=>"110011101",
  43365=>"000101111",
  43366=>"011100111",
  43367=>"111101101",
  43368=>"010000111",
  43369=>"000000100",
  43370=>"001100010",
  43371=>"010100010",
  43372=>"111000000",
  43373=>"101111000",
  43374=>"001001111",
  43375=>"011001001",
  43376=>"001000111",
  43377=>"101000011",
  43378=>"110111010",
  43379=>"111111001",
  43380=>"101011000",
  43381=>"010011100",
  43382=>"010010001",
  43383=>"110100110",
  43384=>"011101110",
  43385=>"001100000",
  43386=>"000001010",
  43387=>"101011010",
  43388=>"101101100",
  43389=>"001001010",
  43390=>"001100000",
  43391=>"011000000",
  43392=>"010111000",
  43393=>"001011001",
  43394=>"110111001",
  43395=>"001101010",
  43396=>"110101101",
  43397=>"010001011",
  43398=>"111101100",
  43399=>"001001100",
  43400=>"111010101",
  43401=>"101001010",
  43402=>"000010001",
  43403=>"011000110",
  43404=>"010001011",
  43405=>"011001010",
  43406=>"100111010",
  43407=>"010110000",
  43408=>"100100111",
  43409=>"000010010",
  43410=>"010001101",
  43411=>"101110101",
  43412=>"000100000",
  43413=>"001111101",
  43414=>"101101111",
  43415=>"100000000",
  43416=>"101110111",
  43417=>"011100100",
  43418=>"110000110",
  43419=>"110000100",
  43420=>"111011010",
  43421=>"010000111",
  43422=>"011010011",
  43423=>"001001011",
  43424=>"010010101",
  43425=>"111100101",
  43426=>"011110100",
  43427=>"110010100",
  43428=>"010110100",
  43429=>"101100000",
  43430=>"011010100",
  43431=>"100000001",
  43432=>"110010011",
  43433=>"100001101",
  43434=>"001101000",
  43435=>"010000100",
  43436=>"001000100",
  43437=>"000110110",
  43438=>"110111000",
  43439=>"101111110",
  43440=>"000011010",
  43441=>"110001000",
  43442=>"011110111",
  43443=>"001110000",
  43444=>"110111110",
  43445=>"101010001",
  43446=>"010001111",
  43447=>"001111110",
  43448=>"100100000",
  43449=>"110011000",
  43450=>"010100100",
  43451=>"101100110",
  43452=>"001110100",
  43453=>"110000000",
  43454=>"000001001",
  43455=>"101100100",
  43456=>"100010011",
  43457=>"101000001",
  43458=>"000111111",
  43459=>"100100001",
  43460=>"001001000",
  43461=>"010111110",
  43462=>"001000100",
  43463=>"100111010",
  43464=>"111100111",
  43465=>"011100110",
  43466=>"100101010",
  43467=>"100111001",
  43468=>"000010000",
  43469=>"001010110",
  43470=>"000101000",
  43471=>"101010101",
  43472=>"100010111",
  43473=>"100111010",
  43474=>"101000010",
  43475=>"010111111",
  43476=>"110101001",
  43477=>"001011001",
  43478=>"001000111",
  43479=>"110011100",
  43480=>"110010100",
  43481=>"000010000",
  43482=>"101001110",
  43483=>"101110101",
  43484=>"000010110",
  43485=>"010100110",
  43486=>"101011101",
  43487=>"100100011",
  43488=>"111101111",
  43489=>"101001101",
  43490=>"110010110",
  43491=>"111100010",
  43492=>"100101101",
  43493=>"110010100",
  43494=>"100011100",
  43495=>"100001010",
  43496=>"011100010",
  43497=>"010001010",
  43498=>"010110101",
  43499=>"000101100",
  43500=>"010011100",
  43501=>"110000010",
  43502=>"110011010",
  43503=>"001100110",
  43504=>"110000100",
  43505=>"100011001",
  43506=>"110011100",
  43507=>"000001101",
  43508=>"110010000",
  43509=>"100001101",
  43510=>"100101111",
  43511=>"110111111",
  43512=>"111110000",
  43513=>"001100000",
  43514=>"000110101",
  43515=>"111011010",
  43516=>"011000110",
  43517=>"101101101",
  43518=>"110111001",
  43519=>"110100100",
  43520=>"000101001",
  43521=>"101101111",
  43522=>"101010111",
  43523=>"110110010",
  43524=>"111010001",
  43525=>"001111100",
  43526=>"010101001",
  43527=>"111101111",
  43528=>"000100000",
  43529=>"010010101",
  43530=>"010011110",
  43531=>"101111100",
  43532=>"010101011",
  43533=>"000000000",
  43534=>"001000010",
  43535=>"111000111",
  43536=>"110000001",
  43537=>"110100110",
  43538=>"010111010",
  43539=>"111011011",
  43540=>"100011000",
  43541=>"100001011",
  43542=>"100000010",
  43543=>"100110111",
  43544=>"100110101",
  43545=>"111101010",
  43546=>"010010001",
  43547=>"101011011",
  43548=>"011000110",
  43549=>"000101110",
  43550=>"101001010",
  43551=>"010001000",
  43552=>"010000011",
  43553=>"110001100",
  43554=>"001100111",
  43555=>"011100100",
  43556=>"111100100",
  43557=>"000111010",
  43558=>"110001110",
  43559=>"010110000",
  43560=>"000111000",
  43561=>"010111110",
  43562=>"000011100",
  43563=>"101001011",
  43564=>"100001110",
  43565=>"101100011",
  43566=>"001001000",
  43567=>"000000011",
  43568=>"100100101",
  43569=>"000101111",
  43570=>"101101110",
  43571=>"011100111",
  43572=>"011011000",
  43573=>"001110111",
  43574=>"011000011",
  43575=>"111101001",
  43576=>"011011011",
  43577=>"000110000",
  43578=>"110111001",
  43579=>"000011011",
  43580=>"010011111",
  43581=>"100011000",
  43582=>"111110101",
  43583=>"111010110",
  43584=>"001000000",
  43585=>"001100100",
  43586=>"000011101",
  43587=>"011001011",
  43588=>"000001010",
  43589=>"100110010",
  43590=>"000101000",
  43591=>"010000011",
  43592=>"111100011",
  43593=>"100101011",
  43594=>"100000110",
  43595=>"101111011",
  43596=>"011100000",
  43597=>"100100011",
  43598=>"011100000",
  43599=>"001011110",
  43600=>"100011011",
  43601=>"111101110",
  43602=>"100101000",
  43603=>"000000000",
  43604=>"001011111",
  43605=>"010000011",
  43606=>"100000101",
  43607=>"111110011",
  43608=>"101010011",
  43609=>"101111100",
  43610=>"011110000",
  43611=>"110000010",
  43612=>"101001001",
  43613=>"100010101",
  43614=>"110011011",
  43615=>"100001000",
  43616=>"110100000",
  43617=>"001100000",
  43618=>"110110010",
  43619=>"011010110",
  43620=>"111111101",
  43621=>"001010011",
  43622=>"001100110",
  43623=>"000001101",
  43624=>"110010111",
  43625=>"111101001",
  43626=>"111111000",
  43627=>"100111100",
  43628=>"000011110",
  43629=>"110011111",
  43630=>"100110101",
  43631=>"101101001",
  43632=>"111000001",
  43633=>"000010000",
  43634=>"111001000",
  43635=>"000000100",
  43636=>"011011001",
  43637=>"000011100",
  43638=>"100110011",
  43639=>"001100000",
  43640=>"011100000",
  43641=>"000111110",
  43642=>"111101011",
  43643=>"111001101",
  43644=>"001000110",
  43645=>"011101111",
  43646=>"000000100",
  43647=>"000011110",
  43648=>"000011100",
  43649=>"100111111",
  43650=>"000110110",
  43651=>"000101110",
  43652=>"010101100",
  43653=>"001100101",
  43654=>"011100110",
  43655=>"110111101",
  43656=>"011011011",
  43657=>"000000110",
  43658=>"010100010",
  43659=>"011110000",
  43660=>"111110000",
  43661=>"000101010",
  43662=>"011110010",
  43663=>"010010111",
  43664=>"010100110",
  43665=>"111100110",
  43666=>"111001101",
  43667=>"101101111",
  43668=>"101000011",
  43669=>"101100100",
  43670=>"111010000",
  43671=>"110011001",
  43672=>"101110011",
  43673=>"111001001",
  43674=>"000100110",
  43675=>"110110111",
  43676=>"100011111",
  43677=>"111000110",
  43678=>"111111010",
  43679=>"000110011",
  43680=>"011101111",
  43681=>"101001000",
  43682=>"101001001",
  43683=>"111111010",
  43684=>"101100101",
  43685=>"010110111",
  43686=>"100000010",
  43687=>"111110100",
  43688=>"101111100",
  43689=>"001110000",
  43690=>"100100111",
  43691=>"100100010",
  43692=>"100001100",
  43693=>"011100000",
  43694=>"000010000",
  43695=>"000001100",
  43696=>"000100111",
  43697=>"010000101",
  43698=>"001101001",
  43699=>"000010010",
  43700=>"000001010",
  43701=>"011001001",
  43702=>"100100100",
  43703=>"101010010",
  43704=>"000111101",
  43705=>"000010111",
  43706=>"111111110",
  43707=>"100111000",
  43708=>"000010000",
  43709=>"010001010",
  43710=>"100010010",
  43711=>"100000000",
  43712=>"000111100",
  43713=>"101100000",
  43714=>"101101100",
  43715=>"110101111",
  43716=>"110111001",
  43717=>"101100110",
  43718=>"111110100",
  43719=>"110010001",
  43720=>"110001101",
  43721=>"011110000",
  43722=>"100011111",
  43723=>"000011000",
  43724=>"000000111",
  43725=>"101101001",
  43726=>"101101101",
  43727=>"110110011",
  43728=>"001101011",
  43729=>"000010100",
  43730=>"101010110",
  43731=>"011010110",
  43732=>"100110010",
  43733=>"001101111",
  43734=>"101100100",
  43735=>"000000100",
  43736=>"001010110",
  43737=>"110001001",
  43738=>"000101101",
  43739=>"001000001",
  43740=>"101000110",
  43741=>"010100101",
  43742=>"100000011",
  43743=>"100011001",
  43744=>"010001000",
  43745=>"100000011",
  43746=>"100111000",
  43747=>"101001011",
  43748=>"011011110",
  43749=>"100000101",
  43750=>"001010010",
  43751=>"100110111",
  43752=>"001100011",
  43753=>"101001001",
  43754=>"001101110",
  43755=>"011010110",
  43756=>"000110111",
  43757=>"011000110",
  43758=>"111110101",
  43759=>"101101101",
  43760=>"110100000",
  43761=>"000101001",
  43762=>"001011000",
  43763=>"010111000",
  43764=>"111111100",
  43765=>"110100001",
  43766=>"000011011",
  43767=>"011001110",
  43768=>"011010101",
  43769=>"111110110",
  43770=>"001001111",
  43771=>"101100011",
  43772=>"111000010",
  43773=>"010100001",
  43774=>"100001101",
  43775=>"011110100",
  43776=>"011100111",
  43777=>"101101111",
  43778=>"001011000",
  43779=>"001010101",
  43780=>"011111110",
  43781=>"001110101",
  43782=>"100010100",
  43783=>"011100110",
  43784=>"001110010",
  43785=>"010001001",
  43786=>"101111010",
  43787=>"101010100",
  43788=>"000001100",
  43789=>"111101111",
  43790=>"101111110",
  43791=>"011010100",
  43792=>"001100010",
  43793=>"000100011",
  43794=>"001101010",
  43795=>"111001101",
  43796=>"011000010",
  43797=>"001010001",
  43798=>"110000100",
  43799=>"100100000",
  43800=>"000000000",
  43801=>"011000110",
  43802=>"111011101",
  43803=>"111101111",
  43804=>"000000111",
  43805=>"011001110",
  43806=>"100010000",
  43807=>"100101010",
  43808=>"011010001",
  43809=>"100110011",
  43810=>"000110111",
  43811=>"110100011",
  43812=>"111010111",
  43813=>"011101011",
  43814=>"011000111",
  43815=>"100111111",
  43816=>"100100000",
  43817=>"100111001",
  43818=>"011011001",
  43819=>"010101111",
  43820=>"110011011",
  43821=>"111101110",
  43822=>"000011110",
  43823=>"001001101",
  43824=>"000100010",
  43825=>"001010010",
  43826=>"000011001",
  43827=>"100001101",
  43828=>"110011000",
  43829=>"110001111",
  43830=>"011000011",
  43831=>"101000110",
  43832=>"001110101",
  43833=>"100110000",
  43834=>"001000100",
  43835=>"100110001",
  43836=>"001101011",
  43837=>"010000000",
  43838=>"101010000",
  43839=>"011011010",
  43840=>"101000111",
  43841=>"100001000",
  43842=>"001000101",
  43843=>"110110000",
  43844=>"110111111",
  43845=>"011101110",
  43846=>"100001101",
  43847=>"111010101",
  43848=>"001111101",
  43849=>"110111100",
  43850=>"000000111",
  43851=>"010000101",
  43852=>"011111000",
  43853=>"010011100",
  43854=>"010110111",
  43855=>"111011010",
  43856=>"101100010",
  43857=>"000001101",
  43858=>"001110101",
  43859=>"110000001",
  43860=>"110111111",
  43861=>"111111011",
  43862=>"010010110",
  43863=>"000111000",
  43864=>"000000000",
  43865=>"011011100",
  43866=>"110000010",
  43867=>"111000110",
  43868=>"110101100",
  43869=>"010100101",
  43870=>"010000011",
  43871=>"000000100",
  43872=>"100010110",
  43873=>"001010100",
  43874=>"000000111",
  43875=>"100011111",
  43876=>"100000110",
  43877=>"010100000",
  43878=>"000000100",
  43879=>"111110111",
  43880=>"010000000",
  43881=>"011010110",
  43882=>"001101000",
  43883=>"100000100",
  43884=>"010110100",
  43885=>"100010101",
  43886=>"000111101",
  43887=>"100011001",
  43888=>"000010010",
  43889=>"111011101",
  43890=>"001000001",
  43891=>"010100001",
  43892=>"101101110",
  43893=>"101101101",
  43894=>"100011001",
  43895=>"110101000",
  43896=>"001001111",
  43897=>"100001110",
  43898=>"011011101",
  43899=>"110111001",
  43900=>"100111101",
  43901=>"001000010",
  43902=>"010000100",
  43903=>"100000110",
  43904=>"101111101",
  43905=>"111101100",
  43906=>"000000110",
  43907=>"010000110",
  43908=>"011000010",
  43909=>"100100100",
  43910=>"000100110",
  43911=>"000001101",
  43912=>"011001100",
  43913=>"101000000",
  43914=>"011100111",
  43915=>"100101000",
  43916=>"101001110",
  43917=>"110010010",
  43918=>"111001011",
  43919=>"111111011",
  43920=>"011010100",
  43921=>"111001101",
  43922=>"100110010",
  43923=>"100101111",
  43924=>"100001001",
  43925=>"101101111",
  43926=>"001001000",
  43927=>"011110010",
  43928=>"101010010",
  43929=>"100100010",
  43930=>"000110001",
  43931=>"010101011",
  43932=>"010000011",
  43933=>"101100010",
  43934=>"011000010",
  43935=>"001101001",
  43936=>"001110110",
  43937=>"000010110",
  43938=>"000110111",
  43939=>"100110110",
  43940=>"011010001",
  43941=>"100100011",
  43942=>"000101111",
  43943=>"011010000",
  43944=>"011001000",
  43945=>"101101101",
  43946=>"101101111",
  43947=>"011000101",
  43948=>"110100111",
  43949=>"111101110",
  43950=>"011101001",
  43951=>"100101101",
  43952=>"011100111",
  43953=>"111111011",
  43954=>"101100111",
  43955=>"011010101",
  43956=>"001010111",
  43957=>"000001011",
  43958=>"111010100",
  43959=>"001101101",
  43960=>"111001111",
  43961=>"110011011",
  43962=>"011011010",
  43963=>"101100010",
  43964=>"100101011",
  43965=>"010100111",
  43966=>"110110011",
  43967=>"110011000",
  43968=>"011011111",
  43969=>"100000100",
  43970=>"001101011",
  43971=>"010000001",
  43972=>"010010110",
  43973=>"100100001",
  43974=>"011111001",
  43975=>"000100011",
  43976=>"000100101",
  43977=>"000011101",
  43978=>"111100101",
  43979=>"110100010",
  43980=>"111010001",
  43981=>"000100111",
  43982=>"000011101",
  43983=>"010101011",
  43984=>"011111011",
  43985=>"000110101",
  43986=>"000000101",
  43987=>"100011011",
  43988=>"010001111",
  43989=>"100111110",
  43990=>"100010100",
  43991=>"101001111",
  43992=>"110001000",
  43993=>"111110001",
  43994=>"111100000",
  43995=>"001110111",
  43996=>"101101101",
  43997=>"111101111",
  43998=>"110110011",
  43999=>"001010010",
  44000=>"101100110",
  44001=>"010001011",
  44002=>"000010100",
  44003=>"100000011",
  44004=>"001010000",
  44005=>"000001001",
  44006=>"101000010",
  44007=>"101111011",
  44008=>"101000111",
  44009=>"100010001",
  44010=>"000000010",
  44011=>"000010011",
  44012=>"010111001",
  44013=>"111001100",
  44014=>"000110100",
  44015=>"001111011",
  44016=>"111000110",
  44017=>"100111111",
  44018=>"000000100",
  44019=>"001101000",
  44020=>"101010111",
  44021=>"010001000",
  44022=>"110101110",
  44023=>"100101001",
  44024=>"111000110",
  44025=>"001111111",
  44026=>"110101111",
  44027=>"000001000",
  44028=>"101101111",
  44029=>"110000100",
  44030=>"111101100",
  44031=>"111111000",
  44032=>"000101000",
  44033=>"111001110",
  44034=>"111111010",
  44035=>"001001001",
  44036=>"011010110",
  44037=>"010011011",
  44038=>"110110111",
  44039=>"100101110",
  44040=>"010000010",
  44041=>"010111101",
  44042=>"001111110",
  44043=>"111011001",
  44044=>"111111111",
  44045=>"100110001",
  44046=>"001011111",
  44047=>"011011100",
  44048=>"001010000",
  44049=>"111010100",
  44050=>"010001111",
  44051=>"101110111",
  44052=>"111000100",
  44053=>"100010000",
  44054=>"001100101",
  44055=>"101110011",
  44056=>"010101100",
  44057=>"111011000",
  44058=>"101011111",
  44059=>"010100110",
  44060=>"111100011",
  44061=>"010000111",
  44062=>"011110011",
  44063=>"010100101",
  44064=>"110110111",
  44065=>"010000101",
  44066=>"000110110",
  44067=>"101010001",
  44068=>"101000001",
  44069=>"101101101",
  44070=>"010001100",
  44071=>"010100101",
  44072=>"100110100",
  44073=>"010100010",
  44074=>"000011110",
  44075=>"101101100",
  44076=>"001111100",
  44077=>"011010101",
  44078=>"100100001",
  44079=>"001000111",
  44080=>"110010011",
  44081=>"010011010",
  44082=>"100000010",
  44083=>"000101011",
  44084=>"010011001",
  44085=>"101101000",
  44086=>"111000110",
  44087=>"001000000",
  44088=>"000111111",
  44089=>"010011000",
  44090=>"010000000",
  44091=>"110011111",
  44092=>"000110000",
  44093=>"001001011",
  44094=>"001011111",
  44095=>"000101111",
  44096=>"111111000",
  44097=>"100000001",
  44098=>"001100001",
  44099=>"100010010",
  44100=>"010011101",
  44101=>"111100111",
  44102=>"111011100",
  44103=>"001011111",
  44104=>"101001011",
  44105=>"000110111",
  44106=>"011010001",
  44107=>"011010100",
  44108=>"100010100",
  44109=>"001000010",
  44110=>"000010111",
  44111=>"011000111",
  44112=>"111011011",
  44113=>"111101111",
  44114=>"101010001",
  44115=>"011000110",
  44116=>"010000111",
  44117=>"100111101",
  44118=>"011100101",
  44119=>"011010100",
  44120=>"001110100",
  44121=>"111001101",
  44122=>"110111001",
  44123=>"110000111",
  44124=>"010010110",
  44125=>"000011111",
  44126=>"001001001",
  44127=>"011010011",
  44128=>"000000110",
  44129=>"111001000",
  44130=>"010001110",
  44131=>"010100101",
  44132=>"011010001",
  44133=>"110000001",
  44134=>"000000111",
  44135=>"111011000",
  44136=>"001101011",
  44137=>"100000111",
  44138=>"010100110",
  44139=>"000101101",
  44140=>"011001110",
  44141=>"111010100",
  44142=>"110001000",
  44143=>"010100011",
  44144=>"000001100",
  44145=>"001100001",
  44146=>"111111011",
  44147=>"000101100",
  44148=>"101101000",
  44149=>"101001010",
  44150=>"100111001",
  44151=>"110000111",
  44152=>"010100110",
  44153=>"010100101",
  44154=>"001001101",
  44155=>"011001010",
  44156=>"001101110",
  44157=>"010100111",
  44158=>"011010111",
  44159=>"011000010",
  44160=>"111010011",
  44161=>"101011011",
  44162=>"111010111",
  44163=>"100010100",
  44164=>"110011011",
  44165=>"110001110",
  44166=>"010110010",
  44167=>"110101100",
  44168=>"100100000",
  44169=>"000001100",
  44170=>"100100010",
  44171=>"110001000",
  44172=>"001110011",
  44173=>"011000100",
  44174=>"100010000",
  44175=>"101011111",
  44176=>"010111100",
  44177=>"110010110",
  44178=>"100001000",
  44179=>"101101010",
  44180=>"001010010",
  44181=>"011000100",
  44182=>"011011001",
  44183=>"111110000",
  44184=>"111111100",
  44185=>"011000101",
  44186=>"110001111",
  44187=>"001100000",
  44188=>"000110010",
  44189=>"101001101",
  44190=>"101001100",
  44191=>"100100011",
  44192=>"010100110",
  44193=>"011101010",
  44194=>"000010111",
  44195=>"010001100",
  44196=>"101100010",
  44197=>"111100011",
  44198=>"101011110",
  44199=>"100110101",
  44200=>"101001001",
  44201=>"011001110",
  44202=>"001110111",
  44203=>"000111100",
  44204=>"001000101",
  44205=>"010100010",
  44206=>"001011111",
  44207=>"111001111",
  44208=>"001101110",
  44209=>"001010001",
  44210=>"110001100",
  44211=>"101011000",
  44212=>"000001111",
  44213=>"110010101",
  44214=>"000100001",
  44215=>"000110000",
  44216=>"010010101",
  44217=>"011111101",
  44218=>"010110011",
  44219=>"101101011",
  44220=>"010110101",
  44221=>"001001101",
  44222=>"111111100",
  44223=>"100111100",
  44224=>"001011011",
  44225=>"101000000",
  44226=>"111010001",
  44227=>"101001101",
  44228=>"000101100",
  44229=>"110110101",
  44230=>"111010110",
  44231=>"111110101",
  44232=>"011111100",
  44233=>"011110111",
  44234=>"111001010",
  44235=>"000100010",
  44236=>"011111010",
  44237=>"111010101",
  44238=>"000110010",
  44239=>"111011000",
  44240=>"100110111",
  44241=>"110000000",
  44242=>"010001000",
  44243=>"111001001",
  44244=>"001010001",
  44245=>"100011110",
  44246=>"101110101",
  44247=>"111000111",
  44248=>"000000001",
  44249=>"101011111",
  44250=>"001110111",
  44251=>"110110011",
  44252=>"000100000",
  44253=>"011000111",
  44254=>"001100000",
  44255=>"100011000",
  44256=>"111110111",
  44257=>"101111111",
  44258=>"010111111",
  44259=>"111000101",
  44260=>"010111000",
  44261=>"011011101",
  44262=>"011011010",
  44263=>"110011010",
  44264=>"101001111",
  44265=>"110101101",
  44266=>"110100010",
  44267=>"100010010",
  44268=>"110011001",
  44269=>"000010110",
  44270=>"110010000",
  44271=>"110000000",
  44272=>"110100000",
  44273=>"010110010",
  44274=>"100010011",
  44275=>"100111010",
  44276=>"110110011",
  44277=>"011000010",
  44278=>"111010001",
  44279=>"011010111",
  44280=>"001111110",
  44281=>"011001010",
  44282=>"001011111",
  44283=>"111011011",
  44284=>"110111100",
  44285=>"000000100",
  44286=>"100110001",
  44287=>"011100100",
  44288=>"110011001",
  44289=>"001101110",
  44290=>"011010100",
  44291=>"000000100",
  44292=>"101101111",
  44293=>"110110011",
  44294=>"110111011",
  44295=>"101100000",
  44296=>"110010101",
  44297=>"011001100",
  44298=>"110101101",
  44299=>"101111011",
  44300=>"010000001",
  44301=>"110101010",
  44302=>"110100000",
  44303=>"000100001",
  44304=>"100001100",
  44305=>"000111001",
  44306=>"001010110",
  44307=>"001010010",
  44308=>"000011100",
  44309=>"111000010",
  44310=>"110110111",
  44311=>"000101110",
  44312=>"010101111",
  44313=>"101000000",
  44314=>"010000001",
  44315=>"001110100",
  44316=>"000010101",
  44317=>"010011010",
  44318=>"011011111",
  44319=>"111001111",
  44320=>"001000010",
  44321=>"010101000",
  44322=>"110011000",
  44323=>"011100110",
  44324=>"010101111",
  44325=>"010110111",
  44326=>"000001000",
  44327=>"001111101",
  44328=>"111010110",
  44329=>"101100110",
  44330=>"111101111",
  44331=>"001010100",
  44332=>"001001010",
  44333=>"010101001",
  44334=>"011100001",
  44335=>"000111101",
  44336=>"011100101",
  44337=>"011011001",
  44338=>"010001010",
  44339=>"001010101",
  44340=>"001110000",
  44341=>"101000100",
  44342=>"010100000",
  44343=>"000101111",
  44344=>"000001010",
  44345=>"011100101",
  44346=>"010110110",
  44347=>"110110100",
  44348=>"000011110",
  44349=>"110011001",
  44350=>"000111100",
  44351=>"100000111",
  44352=>"011000000",
  44353=>"011111011",
  44354=>"101001100",
  44355=>"011101000",
  44356=>"011000000",
  44357=>"101100110",
  44358=>"000000010",
  44359=>"011111111",
  44360=>"010010000",
  44361=>"010010111",
  44362=>"010101111",
  44363=>"000000010",
  44364=>"100000000",
  44365=>"111010100",
  44366=>"100011000",
  44367=>"110100010",
  44368=>"101101110",
  44369=>"011111101",
  44370=>"111110111",
  44371=>"001010000",
  44372=>"100100001",
  44373=>"010100101",
  44374=>"101101010",
  44375=>"001101000",
  44376=>"010010111",
  44377=>"111110001",
  44378=>"011001110",
  44379=>"100111111",
  44380=>"001100101",
  44381=>"010111000",
  44382=>"000010011",
  44383=>"001110001",
  44384=>"000001001",
  44385=>"011110101",
  44386=>"000011011",
  44387=>"000001110",
  44388=>"010000010",
  44389=>"010000011",
  44390=>"010111100",
  44391=>"111101001",
  44392=>"001110101",
  44393=>"010000101",
  44394=>"001110001",
  44395=>"101110001",
  44396=>"010010001",
  44397=>"010100110",
  44398=>"000111100",
  44399=>"110100001",
  44400=>"000101100",
  44401=>"010010000",
  44402=>"011110100",
  44403=>"110100100",
  44404=>"110011000",
  44405=>"011011110",
  44406=>"100001100",
  44407=>"100100000",
  44408=>"100110010",
  44409=>"111011010",
  44410=>"110100001",
  44411=>"001111101",
  44412=>"101100000",
  44413=>"000001111",
  44414=>"000110000",
  44415=>"011001001",
  44416=>"000110110",
  44417=>"000000110",
  44418=>"100001010",
  44419=>"110101111",
  44420=>"100011001",
  44421=>"101101101",
  44422=>"111000110",
  44423=>"110001000",
  44424=>"100101010",
  44425=>"110110011",
  44426=>"100011001",
  44427=>"101000000",
  44428=>"010010101",
  44429=>"110101111",
  44430=>"011010011",
  44431=>"100001000",
  44432=>"001100011",
  44433=>"110001000",
  44434=>"110010011",
  44435=>"000000100",
  44436=>"011011001",
  44437=>"000110011",
  44438=>"001001010",
  44439=>"011100100",
  44440=>"000110010",
  44441=>"001010101",
  44442=>"100111011",
  44443=>"110110011",
  44444=>"110101001",
  44445=>"101011111",
  44446=>"000101101",
  44447=>"000110001",
  44448=>"111100000",
  44449=>"011100000",
  44450=>"110010111",
  44451=>"011010000",
  44452=>"111111110",
  44453=>"110011000",
  44454=>"110011000",
  44455=>"111010010",
  44456=>"111001110",
  44457=>"010100110",
  44458=>"111011110",
  44459=>"011110100",
  44460=>"111110111",
  44461=>"101011110",
  44462=>"010110100",
  44463=>"110111000",
  44464=>"010010100",
  44465=>"010110010",
  44466=>"001010010",
  44467=>"011100110",
  44468=>"010001101",
  44469=>"111111011",
  44470=>"100101010",
  44471=>"011110000",
  44472=>"011110001",
  44473=>"001111000",
  44474=>"000000010",
  44475=>"011000111",
  44476=>"101110010",
  44477=>"011010010",
  44478=>"110010100",
  44479=>"010011110",
  44480=>"011001100",
  44481=>"010101110",
  44482=>"010010110",
  44483=>"111111100",
  44484=>"010010000",
  44485=>"001111100",
  44486=>"010000000",
  44487=>"110000010",
  44488=>"011010001",
  44489=>"110000111",
  44490=>"010000100",
  44491=>"100010110",
  44492=>"110010110",
  44493=>"011011000",
  44494=>"010111011",
  44495=>"100100010",
  44496=>"010111101",
  44497=>"001011110",
  44498=>"110011110",
  44499=>"010010000",
  44500=>"010101111",
  44501=>"000100110",
  44502=>"111000010",
  44503=>"110000100",
  44504=>"011111001",
  44505=>"101100000",
  44506=>"111101000",
  44507=>"010001011",
  44508=>"100101011",
  44509=>"101010110",
  44510=>"111010000",
  44511=>"010111000",
  44512=>"100110101",
  44513=>"100110011",
  44514=>"000101100",
  44515=>"011101001",
  44516=>"011101011",
  44517=>"001011000",
  44518=>"011100001",
  44519=>"000001101",
  44520=>"111111111",
  44521=>"000110001",
  44522=>"101101110",
  44523=>"011100111",
  44524=>"001101010",
  44525=>"100110000",
  44526=>"011000110",
  44527=>"001111010",
  44528=>"010110100",
  44529=>"111010100",
  44530=>"101101101",
  44531=>"000110100",
  44532=>"110010111",
  44533=>"110000110",
  44534=>"111000111",
  44535=>"100100111",
  44536=>"000111001",
  44537=>"001111001",
  44538=>"000011000",
  44539=>"101001101",
  44540=>"101010001",
  44541=>"100000110",
  44542=>"100111011",
  44543=>"000000011",
  44544=>"011010001",
  44545=>"101011110",
  44546=>"011011011",
  44547=>"010000000",
  44548=>"010011000",
  44549=>"000101000",
  44550=>"110100010",
  44551=>"111100000",
  44552=>"111001110",
  44553=>"001011010",
  44554=>"101001010",
  44555=>"100100111",
  44556=>"000111111",
  44557=>"000001001",
  44558=>"001011101",
  44559=>"011111010",
  44560=>"100000110",
  44561=>"011011100",
  44562=>"110101011",
  44563=>"100010001",
  44564=>"110000110",
  44565=>"100101111",
  44566=>"100010000",
  44567=>"100001100",
  44568=>"001000100",
  44569=>"010100110",
  44570=>"001011000",
  44571=>"000100010",
  44572=>"000000000",
  44573=>"100010110",
  44574=>"101111110",
  44575=>"010010101",
  44576=>"110111010",
  44577=>"100110001",
  44578=>"101011101",
  44579=>"011101010",
  44580=>"101110000",
  44581=>"010101110",
  44582=>"000100101",
  44583=>"001011011",
  44584=>"110101000",
  44585=>"010110011",
  44586=>"011011101",
  44587=>"101011010",
  44588=>"000100110",
  44589=>"111000100",
  44590=>"110100100",
  44591=>"110110001",
  44592=>"010000001",
  44593=>"001001000",
  44594=>"101010111",
  44595=>"110111111",
  44596=>"010100111",
  44597=>"011011101",
  44598=>"011011011",
  44599=>"110111101",
  44600=>"001100110",
  44601=>"100101010",
  44602=>"101111010",
  44603=>"101111000",
  44604=>"101100111",
  44605=>"101101111",
  44606=>"010111011",
  44607=>"010011001",
  44608=>"011001101",
  44609=>"110000000",
  44610=>"100011100",
  44611=>"001010111",
  44612=>"011000111",
  44613=>"100011100",
  44614=>"001000001",
  44615=>"101010111",
  44616=>"001001001",
  44617=>"000100101",
  44618=>"110100011",
  44619=>"100010001",
  44620=>"110110101",
  44621=>"011000001",
  44622=>"101010000",
  44623=>"100001110",
  44624=>"010000001",
  44625=>"101101011",
  44626=>"010111101",
  44627=>"011011001",
  44628=>"001010111",
  44629=>"111001110",
  44630=>"100110101",
  44631=>"010100100",
  44632=>"010000010",
  44633=>"101101001",
  44634=>"111101101",
  44635=>"110110000",
  44636=>"011000001",
  44637=>"001111001",
  44638=>"111011001",
  44639=>"110101111",
  44640=>"111100011",
  44641=>"000000011",
  44642=>"110101111",
  44643=>"001000111",
  44644=>"001001010",
  44645=>"111011101",
  44646=>"111000000",
  44647=>"101000111",
  44648=>"110100011",
  44649=>"110110000",
  44650=>"111111000",
  44651=>"111001100",
  44652=>"100101001",
  44653=>"011100010",
  44654=>"010100111",
  44655=>"111110001",
  44656=>"101011001",
  44657=>"011000010",
  44658=>"111000101",
  44659=>"000100111",
  44660=>"010011011",
  44661=>"101100101",
  44662=>"111111110",
  44663=>"011001111",
  44664=>"001010010",
  44665=>"001010111",
  44666=>"010110000",
  44667=>"001011101",
  44668=>"000010111",
  44669=>"100101011",
  44670=>"000001010",
  44671=>"001110001",
  44672=>"101000000",
  44673=>"101000111",
  44674=>"000101100",
  44675=>"110101001",
  44676=>"010110010",
  44677=>"101010101",
  44678=>"011011100",
  44679=>"111001001",
  44680=>"101010111",
  44681=>"001001010",
  44682=>"001010100",
  44683=>"010000001",
  44684=>"011111010",
  44685=>"010011000",
  44686=>"100001011",
  44687=>"010010001",
  44688=>"011101110",
  44689=>"001101001",
  44690=>"010001101",
  44691=>"011001011",
  44692=>"011101000",
  44693=>"111110001",
  44694=>"010101110",
  44695=>"011001101",
  44696=>"100101101",
  44697=>"001101101",
  44698=>"110100100",
  44699=>"000011110",
  44700=>"110100101",
  44701=>"001111101",
  44702=>"000000110",
  44703=>"100101101",
  44704=>"010100001",
  44705=>"010100111",
  44706=>"001101110",
  44707=>"010010110",
  44708=>"101101101",
  44709=>"000000001",
  44710=>"010000111",
  44711=>"000110001",
  44712=>"111010000",
  44713=>"100000111",
  44714=>"000110100",
  44715=>"001010000",
  44716=>"001111100",
  44717=>"000111000",
  44718=>"100001110",
  44719=>"111111001",
  44720=>"001010111",
  44721=>"011101100",
  44722=>"100011101",
  44723=>"110001010",
  44724=>"001110101",
  44725=>"100111010",
  44726=>"011101111",
  44727=>"111101001",
  44728=>"011001001",
  44729=>"001100010",
  44730=>"110111110",
  44731=>"010100000",
  44732=>"000111011",
  44733=>"000100101",
  44734=>"101010111",
  44735=>"100000100",
  44736=>"011100011",
  44737=>"101001101",
  44738=>"000110100",
  44739=>"010110111",
  44740=>"101010000",
  44741=>"001011101",
  44742=>"001000000",
  44743=>"011111111",
  44744=>"100111000",
  44745=>"010111110",
  44746=>"000010011",
  44747=>"001111011",
  44748=>"000100001",
  44749=>"111100011",
  44750=>"000001000",
  44751=>"000010001",
  44752=>"011001110",
  44753=>"110101000",
  44754=>"011110110",
  44755=>"000101101",
  44756=>"001100110",
  44757=>"000100010",
  44758=>"111111010",
  44759=>"100110101",
  44760=>"100111011",
  44761=>"000010010",
  44762=>"111110011",
  44763=>"100001010",
  44764=>"000111001",
  44765=>"100100100",
  44766=>"101100100",
  44767=>"011011011",
  44768=>"011100000",
  44769=>"010011001",
  44770=>"000110110",
  44771=>"001111100",
  44772=>"100110001",
  44773=>"110101000",
  44774=>"010001100",
  44775=>"110111010",
  44776=>"011110100",
  44777=>"111110001",
  44778=>"111111000",
  44779=>"010111001",
  44780=>"000001001",
  44781=>"111001000",
  44782=>"011110100",
  44783=>"101110111",
  44784=>"110001001",
  44785=>"111011110",
  44786=>"111111011",
  44787=>"011111011",
  44788=>"101101001",
  44789=>"100001110",
  44790=>"011101100",
  44791=>"000010100",
  44792=>"000101001",
  44793=>"110100110",
  44794=>"110110000",
  44795=>"100100001",
  44796=>"101000110",
  44797=>"100101011",
  44798=>"101111000",
  44799=>"011001110",
  44800=>"101101101",
  44801=>"100010011",
  44802=>"011010111",
  44803=>"110101111",
  44804=>"101000000",
  44805=>"001001010",
  44806=>"010111011",
  44807=>"100111100",
  44808=>"110101110",
  44809=>"010101100",
  44810=>"101000110",
  44811=>"111100010",
  44812=>"000000011",
  44813=>"000101100",
  44814=>"000111011",
  44815=>"011110000",
  44816=>"011001110",
  44817=>"000111101",
  44818=>"000010010",
  44819=>"110000100",
  44820=>"101011000",
  44821=>"100011101",
  44822=>"110101000",
  44823=>"000010000",
  44824=>"101101011",
  44825=>"011100100",
  44826=>"001000101",
  44827=>"010000101",
  44828=>"101011001",
  44829=>"011101110",
  44830=>"111100111",
  44831=>"001100111",
  44832=>"011100000",
  44833=>"010111101",
  44834=>"100001010",
  44835=>"001101111",
  44836=>"100010001",
  44837=>"110110101",
  44838=>"110111111",
  44839=>"100111001",
  44840=>"000100111",
  44841=>"011000101",
  44842=>"000111111",
  44843=>"101011000",
  44844=>"001001010",
  44845=>"000000100",
  44846=>"011111011",
  44847=>"001010000",
  44848=>"100010011",
  44849=>"110010111",
  44850=>"111011010",
  44851=>"000110010",
  44852=>"100001111",
  44853=>"100011101",
  44854=>"001101101",
  44855=>"001011110",
  44856=>"000010000",
  44857=>"011101111",
  44858=>"110000111",
  44859=>"111110010",
  44860=>"000100000",
  44861=>"111100110",
  44862=>"100101010",
  44863=>"000010111",
  44864=>"101111100",
  44865=>"000101001",
  44866=>"111001001",
  44867=>"110010010",
  44868=>"001111110",
  44869=>"110100110",
  44870=>"111110001",
  44871=>"011111011",
  44872=>"010001000",
  44873=>"111111000",
  44874=>"010000111",
  44875=>"011010101",
  44876=>"001110001",
  44877=>"001010110",
  44878=>"110101011",
  44879=>"101000000",
  44880=>"101001011",
  44881=>"011110111",
  44882=>"100010011",
  44883=>"011000111",
  44884=>"111001111",
  44885=>"111001001",
  44886=>"110111110",
  44887=>"111100110",
  44888=>"000111000",
  44889=>"101000111",
  44890=>"001001011",
  44891=>"100000000",
  44892=>"010000111",
  44893=>"101111011",
  44894=>"111111011",
  44895=>"011011011",
  44896=>"100101011",
  44897=>"100111010",
  44898=>"011110110",
  44899=>"100001011",
  44900=>"010110110",
  44901=>"111000110",
  44902=>"111110110",
  44903=>"011101011",
  44904=>"010000010",
  44905=>"110100110",
  44906=>"100110010",
  44907=>"011101110",
  44908=>"110001110",
  44909=>"101000011",
  44910=>"101100110",
  44911=>"010111111",
  44912=>"100101001",
  44913=>"111101011",
  44914=>"101111110",
  44915=>"010001000",
  44916=>"011011101",
  44917=>"110110011",
  44918=>"100010011",
  44919=>"000010011",
  44920=>"110101111",
  44921=>"010011100",
  44922=>"000010000",
  44923=>"010011111",
  44924=>"000010010",
  44925=>"110011111",
  44926=>"000010000",
  44927=>"010111001",
  44928=>"011000011",
  44929=>"001111111",
  44930=>"001000110",
  44931=>"110001110",
  44932=>"100110111",
  44933=>"010100111",
  44934=>"011011101",
  44935=>"101000011",
  44936=>"000000101",
  44937=>"001001110",
  44938=>"000000101",
  44939=>"100111011",
  44940=>"010011101",
  44941=>"010111001",
  44942=>"111011110",
  44943=>"110101101",
  44944=>"011000000",
  44945=>"110000110",
  44946=>"100011111",
  44947=>"000000110",
  44948=>"010111010",
  44949=>"110110110",
  44950=>"111100100",
  44951=>"011100101",
  44952=>"101110111",
  44953=>"010010001",
  44954=>"000101111",
  44955=>"100010110",
  44956=>"010011000",
  44957=>"101110010",
  44958=>"100110100",
  44959=>"011000000",
  44960=>"010111000",
  44961=>"101100100",
  44962=>"110100000",
  44963=>"000110101",
  44964=>"000111110",
  44965=>"010010100",
  44966=>"000110011",
  44967=>"000000011",
  44968=>"010011101",
  44969=>"001000001",
  44970=>"001011111",
  44971=>"101101011",
  44972=>"001110111",
  44973=>"110100001",
  44974=>"000000111",
  44975=>"101001001",
  44976=>"010010000",
  44977=>"110001100",
  44978=>"000010101",
  44979=>"111001000",
  44980=>"111101111",
  44981=>"101110101",
  44982=>"010111111",
  44983=>"000111100",
  44984=>"001010010",
  44985=>"010010001",
  44986=>"011001010",
  44987=>"000000100",
  44988=>"010011101",
  44989=>"000100000",
  44990=>"111011010",
  44991=>"111000110",
  44992=>"100011110",
  44993=>"101001001",
  44994=>"100000110",
  44995=>"010101011",
  44996=>"000100100",
  44997=>"110101000",
  44998=>"101011001",
  44999=>"010000111",
  45000=>"111100101",
  45001=>"101100111",
  45002=>"011111011",
  45003=>"001110101",
  45004=>"011101111",
  45005=>"111001011",
  45006=>"011100101",
  45007=>"001001010",
  45008=>"110001011",
  45009=>"111001011",
  45010=>"010000100",
  45011=>"100101100",
  45012=>"101101111",
  45013=>"001011011",
  45014=>"010100000",
  45015=>"011000000",
  45016=>"010010011",
  45017=>"101110111",
  45018=>"001101010",
  45019=>"101010010",
  45020=>"100000010",
  45021=>"111111010",
  45022=>"100010111",
  45023=>"111000010",
  45024=>"011011011",
  45025=>"001011101",
  45026=>"110110111",
  45027=>"110100101",
  45028=>"011011011",
  45029=>"010100000",
  45030=>"001111011",
  45031=>"000111001",
  45032=>"111010001",
  45033=>"000110110",
  45034=>"011010001",
  45035=>"010111100",
  45036=>"001010001",
  45037=>"101010110",
  45038=>"001101100",
  45039=>"001010010",
  45040=>"011000101",
  45041=>"101100101",
  45042=>"111000011",
  45043=>"011100001",
  45044=>"011000000",
  45045=>"000100111",
  45046=>"111000000",
  45047=>"010100111",
  45048=>"111000111",
  45049=>"111100001",
  45050=>"100000001",
  45051=>"110011110",
  45052=>"001000111",
  45053=>"001110101",
  45054=>"101011110",
  45055=>"011111011",
  45056=>"101101100",
  45057=>"111101010",
  45058=>"101010100",
  45059=>"101000010",
  45060=>"111000101",
  45061=>"100100101",
  45062=>"011000000",
  45063=>"000101000",
  45064=>"101011110",
  45065=>"100110001",
  45066=>"001100000",
  45067=>"000101011",
  45068=>"100101010",
  45069=>"011001000",
  45070=>"000101010",
  45071=>"001110110",
  45072=>"111001100",
  45073=>"000111000",
  45074=>"110010001",
  45075=>"001011011",
  45076=>"110100010",
  45077=>"110011011",
  45078=>"011000011",
  45079=>"001000100",
  45080=>"110110011",
  45081=>"011100100",
  45082=>"001100111",
  45083=>"011110011",
  45084=>"001100000",
  45085=>"101000010",
  45086=>"110010010",
  45087=>"110110010",
  45088=>"101011101",
  45089=>"100000100",
  45090=>"011001101",
  45091=>"110011010",
  45092=>"011110011",
  45093=>"110110101",
  45094=>"110010110",
  45095=>"101001010",
  45096=>"100011010",
  45097=>"001011110",
  45098=>"101001110",
  45099=>"000100010",
  45100=>"100001001",
  45101=>"011010011",
  45102=>"110000001",
  45103=>"101101001",
  45104=>"010110100",
  45105=>"101001101",
  45106=>"010101101",
  45107=>"001010010",
  45108=>"101101111",
  45109=>"000000001",
  45110=>"011100101",
  45111=>"011011100",
  45112=>"101101000",
  45113=>"000100100",
  45114=>"111111000",
  45115=>"000001111",
  45116=>"110100001",
  45117=>"001100010",
  45118=>"101101000",
  45119=>"101101001",
  45120=>"101000011",
  45121=>"001101010",
  45122=>"101100000",
  45123=>"010101111",
  45124=>"011011111",
  45125=>"111000100",
  45126=>"111010011",
  45127=>"000100101",
  45128=>"001001100",
  45129=>"010110011",
  45130=>"000000000",
  45131=>"000010010",
  45132=>"011010000",
  45133=>"010100101",
  45134=>"101110110",
  45135=>"110000101",
  45136=>"000110001",
  45137=>"101011000",
  45138=>"110110010",
  45139=>"011010111",
  45140=>"010000110",
  45141=>"111111100",
  45142=>"101000110",
  45143=>"001000001",
  45144=>"101001110",
  45145=>"011000010",
  45146=>"100011110",
  45147=>"101111110",
  45148=>"110001111",
  45149=>"100101101",
  45150=>"100010110",
  45151=>"111001001",
  45152=>"000100010",
  45153=>"011111011",
  45154=>"110101100",
  45155=>"011110110",
  45156=>"011001010",
  45157=>"100011010",
  45158=>"001111001",
  45159=>"000100110",
  45160=>"010010101",
  45161=>"110011000",
  45162=>"010001000",
  45163=>"110100100",
  45164=>"000001101",
  45165=>"000100001",
  45166=>"111001101",
  45167=>"100101101",
  45168=>"010001010",
  45169=>"010110100",
  45170=>"111001101",
  45171=>"001011001",
  45172=>"001010000",
  45173=>"100010111",
  45174=>"000010010",
  45175=>"100100110",
  45176=>"101011111",
  45177=>"110111110",
  45178=>"011010000",
  45179=>"110100110",
  45180=>"100001101",
  45181=>"011000000",
  45182=>"011100101",
  45183=>"101110010",
  45184=>"001011111",
  45185=>"001011101",
  45186=>"000110010",
  45187=>"001000101",
  45188=>"001000011",
  45189=>"101000101",
  45190=>"011001011",
  45191=>"000000001",
  45192=>"101011110",
  45193=>"001111010",
  45194=>"001010000",
  45195=>"111111011",
  45196=>"110101100",
  45197=>"010001000",
  45198=>"100000101",
  45199=>"110101010",
  45200=>"111011111",
  45201=>"011010011",
  45202=>"010100000",
  45203=>"101011001",
  45204=>"101001011",
  45205=>"110100001",
  45206=>"001000010",
  45207=>"110000001",
  45208=>"011110001",
  45209=>"011011101",
  45210=>"011010101",
  45211=>"100101010",
  45212=>"111001001",
  45213=>"100101000",
  45214=>"101111100",
  45215=>"010001110",
  45216=>"111011100",
  45217=>"111001011",
  45218=>"100010000",
  45219=>"010010001",
  45220=>"100001000",
  45221=>"111110110",
  45222=>"100000011",
  45223=>"110011001",
  45224=>"000001110",
  45225=>"010010100",
  45226=>"110100001",
  45227=>"111111110",
  45228=>"111001010",
  45229=>"110001011",
  45230=>"010011101",
  45231=>"100100100",
  45232=>"000010111",
  45233=>"000010010",
  45234=>"011010010",
  45235=>"001110101",
  45236=>"001101010",
  45237=>"000101010",
  45238=>"010100110",
  45239=>"011001100",
  45240=>"100010000",
  45241=>"110110101",
  45242=>"010000011",
  45243=>"111000000",
  45244=>"000101110",
  45245=>"001010101",
  45246=>"000111100",
  45247=>"101000001",
  45248=>"001100111",
  45249=>"101111101",
  45250=>"001110010",
  45251=>"101011010",
  45252=>"111001110",
  45253=>"000101010",
  45254=>"000101111",
  45255=>"111101101",
  45256=>"111000110",
  45257=>"000111011",
  45258=>"000110000",
  45259=>"010111110",
  45260=>"110100010",
  45261=>"101101101",
  45262=>"000101111",
  45263=>"101010010",
  45264=>"000111000",
  45265=>"001010011",
  45266=>"010100111",
  45267=>"110111000",
  45268=>"111001100",
  45269=>"100111100",
  45270=>"101000111",
  45271=>"010001011",
  45272=>"100001010",
  45273=>"011000100",
  45274=>"111110101",
  45275=>"111100100",
  45276=>"110011111",
  45277=>"010000100",
  45278=>"001011100",
  45279=>"111000000",
  45280=>"100101100",
  45281=>"001011110",
  45282=>"000001101",
  45283=>"001010110",
  45284=>"111111110",
  45285=>"101010011",
  45286=>"111101011",
  45287=>"111111111",
  45288=>"010101100",
  45289=>"100011100",
  45290=>"011000000",
  45291=>"111010110",
  45292=>"011011000",
  45293=>"101111011",
  45294=>"100110110",
  45295=>"111111111",
  45296=>"110101100",
  45297=>"111100101",
  45298=>"011110001",
  45299=>"110000101",
  45300=>"001111001",
  45301=>"110011001",
  45302=>"011011010",
  45303=>"001111101",
  45304=>"011001011",
  45305=>"011000001",
  45306=>"101000101",
  45307=>"110000000",
  45308=>"100010110",
  45309=>"010010111",
  45310=>"111001011",
  45311=>"110011110",
  45312=>"010001101",
  45313=>"101110001",
  45314=>"011101000",
  45315=>"010110110",
  45316=>"110001110",
  45317=>"011011110",
  45318=>"111001010",
  45319=>"011000101",
  45320=>"001100111",
  45321=>"110101001",
  45322=>"001011000",
  45323=>"101011010",
  45324=>"011111110",
  45325=>"110101100",
  45326=>"001001100",
  45327=>"110111111",
  45328=>"000000010",
  45329=>"000010100",
  45330=>"001010011",
  45331=>"010101111",
  45332=>"001000110",
  45333=>"100100101",
  45334=>"111110001",
  45335=>"001101110",
  45336=>"001000001",
  45337=>"110111000",
  45338=>"100000101",
  45339=>"100101100",
  45340=>"000111110",
  45341=>"110001010",
  45342=>"011010101",
  45343=>"001001101",
  45344=>"010111100",
  45345=>"100011011",
  45346=>"001010100",
  45347=>"000100111",
  45348=>"111010010",
  45349=>"001100110",
  45350=>"101111010",
  45351=>"011010010",
  45352=>"111111100",
  45353=>"110111000",
  45354=>"110101110",
  45355=>"000011011",
  45356=>"000100111",
  45357=>"100000001",
  45358=>"010101111",
  45359=>"100001001",
  45360=>"011001010",
  45361=>"010001010",
  45362=>"001000110",
  45363=>"000000001",
  45364=>"110100001",
  45365=>"111010101",
  45366=>"001011101",
  45367=>"000011110",
  45368=>"110111011",
  45369=>"110010000",
  45370=>"100100100",
  45371=>"110110011",
  45372=>"011111101",
  45373=>"001010000",
  45374=>"101101101",
  45375=>"100000001",
  45376=>"001100111",
  45377=>"100011000",
  45378=>"100110101",
  45379=>"111011000",
  45380=>"001000100",
  45381=>"111101101",
  45382=>"011011001",
  45383=>"110001001",
  45384=>"000011011",
  45385=>"101001011",
  45386=>"100101101",
  45387=>"000010000",
  45388=>"101111100",
  45389=>"110001011",
  45390=>"111100101",
  45391=>"100100110",
  45392=>"110101001",
  45393=>"111111101",
  45394=>"111110111",
  45395=>"100100010",
  45396=>"000001010",
  45397=>"101101110",
  45398=>"110001101",
  45399=>"101111110",
  45400=>"010100011",
  45401=>"100011100",
  45402=>"011110100",
  45403=>"010110100",
  45404=>"010110000",
  45405=>"010010011",
  45406=>"001011100",
  45407=>"000101101",
  45408=>"001000110",
  45409=>"111000011",
  45410=>"110011000",
  45411=>"000101111",
  45412=>"101001111",
  45413=>"101110001",
  45414=>"110011010",
  45415=>"010000100",
  45416=>"101101001",
  45417=>"100001101",
  45418=>"011110110",
  45419=>"001100000",
  45420=>"011011001",
  45421=>"011101111",
  45422=>"000011111",
  45423=>"101000110",
  45424=>"111010011",
  45425=>"110111011",
  45426=>"000101111",
  45427=>"111100010",
  45428=>"010000010",
  45429=>"001000101",
  45430=>"000100011",
  45431=>"101000011",
  45432=>"111101100",
  45433=>"110011111",
  45434=>"001101000",
  45435=>"110110101",
  45436=>"100110100",
  45437=>"001000110",
  45438=>"111010110",
  45439=>"011011011",
  45440=>"110101111",
  45441=>"010100000",
  45442=>"100111000",
  45443=>"010001000",
  45444=>"100000100",
  45445=>"000000000",
  45446=>"000111010",
  45447=>"011011101",
  45448=>"101000011",
  45449=>"100100001",
  45450=>"000000111",
  45451=>"100000111",
  45452=>"100000101",
  45453=>"100001010",
  45454=>"111100111",
  45455=>"000011000",
  45456=>"010001011",
  45457=>"001000001",
  45458=>"100001100",
  45459=>"111100001",
  45460=>"111110010",
  45461=>"111111111",
  45462=>"010110011",
  45463=>"110010011",
  45464=>"000110001",
  45465=>"101000111",
  45466=>"100000111",
  45467=>"110100010",
  45468=>"011001010",
  45469=>"001101111",
  45470=>"011010000",
  45471=>"001110011",
  45472=>"010001011",
  45473=>"011010111",
  45474=>"100001010",
  45475=>"000010010",
  45476=>"010001110",
  45477=>"100000000",
  45478=>"100010010",
  45479=>"001111100",
  45480=>"100110001",
  45481=>"001100010",
  45482=>"110111100",
  45483=>"100011001",
  45484=>"110101101",
  45485=>"100100001",
  45486=>"101100001",
  45487=>"011010001",
  45488=>"111001000",
  45489=>"011101101",
  45490=>"010000101",
  45491=>"011101001",
  45492=>"010011010",
  45493=>"111110010",
  45494=>"001101111",
  45495=>"001000010",
  45496=>"011110111",
  45497=>"011101100",
  45498=>"000000011",
  45499=>"110100110",
  45500=>"100111111",
  45501=>"001110001",
  45502=>"110010100",
  45503=>"011011101",
  45504=>"110001000",
  45505=>"001011000",
  45506=>"001000010",
  45507=>"100001111",
  45508=>"110000000",
  45509=>"110000111",
  45510=>"001010100",
  45511=>"000000000",
  45512=>"011100011",
  45513=>"101001001",
  45514=>"001001101",
  45515=>"100011100",
  45516=>"001001010",
  45517=>"111011000",
  45518=>"100111110",
  45519=>"111110001",
  45520=>"100100111",
  45521=>"110111000",
  45522=>"101001011",
  45523=>"101010110",
  45524=>"101101011",
  45525=>"111110100",
  45526=>"000001100",
  45527=>"110100100",
  45528=>"000110110",
  45529=>"000011111",
  45530=>"110110111",
  45531=>"001110010",
  45532=>"010011101",
  45533=>"001010001",
  45534=>"101011011",
  45535=>"010010101",
  45536=>"110101000",
  45537=>"101110011",
  45538=>"110101011",
  45539=>"001100010",
  45540=>"101011100",
  45541=>"110111100",
  45542=>"001000100",
  45543=>"000000000",
  45544=>"101010001",
  45545=>"011011100",
  45546=>"010001010",
  45547=>"111001111",
  45548=>"111001010",
  45549=>"000000110",
  45550=>"100101000",
  45551=>"000111100",
  45552=>"001000111",
  45553=>"000111111",
  45554=>"100000000",
  45555=>"001101010",
  45556=>"011111011",
  45557=>"100101110",
  45558=>"011101110",
  45559=>"101111111",
  45560=>"110001111",
  45561=>"010100110",
  45562=>"111101100",
  45563=>"001110100",
  45564=>"111100111",
  45565=>"100010001",
  45566=>"100100100",
  45567=>"100011100",
  45568=>"110010010",
  45569=>"101011010",
  45570=>"100101000",
  45571=>"000000001",
  45572=>"001111101",
  45573=>"010110011",
  45574=>"111011111",
  45575=>"110111001",
  45576=>"011101000",
  45577=>"100001111",
  45578=>"001000001",
  45579=>"010100111",
  45580=>"101111101",
  45581=>"111001001",
  45582=>"011010111",
  45583=>"101011010",
  45584=>"010100111",
  45585=>"110100000",
  45586=>"111010001",
  45587=>"101010111",
  45588=>"001111000",
  45589=>"000000010",
  45590=>"010011111",
  45591=>"010011010",
  45592=>"101100011",
  45593=>"110110011",
  45594=>"011101101",
  45595=>"100001111",
  45596=>"000100011",
  45597=>"011011111",
  45598=>"011100000",
  45599=>"100111111",
  45600=>"000110100",
  45601=>"011000101",
  45602=>"100000001",
  45603=>"100001101",
  45604=>"001011110",
  45605=>"000101010",
  45606=>"011010011",
  45607=>"010010000",
  45608=>"001000101",
  45609=>"100110011",
  45610=>"111001011",
  45611=>"010110000",
  45612=>"100101011",
  45613=>"100100100",
  45614=>"001100010",
  45615=>"000101001",
  45616=>"011100010",
  45617=>"011111010",
  45618=>"111100011",
  45619=>"110001011",
  45620=>"001110000",
  45621=>"011001101",
  45622=>"000000111",
  45623=>"100101000",
  45624=>"101100101",
  45625=>"000001111",
  45626=>"011111101",
  45627=>"011011010",
  45628=>"000011000",
  45629=>"110101101",
  45630=>"101101011",
  45631=>"010001010",
  45632=>"001101101",
  45633=>"111000001",
  45634=>"011111110",
  45635=>"001010100",
  45636=>"000010000",
  45637=>"001011000",
  45638=>"110101110",
  45639=>"101111001",
  45640=>"100111101",
  45641=>"001010011",
  45642=>"000101001",
  45643=>"001011111",
  45644=>"000101010",
  45645=>"001100010",
  45646=>"011101101",
  45647=>"010101010",
  45648=>"101011000",
  45649=>"011111001",
  45650=>"100110111",
  45651=>"110101000",
  45652=>"011110110",
  45653=>"011001001",
  45654=>"100110100",
  45655=>"110111011",
  45656=>"100010111",
  45657=>"101100111",
  45658=>"010101100",
  45659=>"100001110",
  45660=>"000001011",
  45661=>"111010011",
  45662=>"000111101",
  45663=>"010111001",
  45664=>"101110010",
  45665=>"111101110",
  45666=>"001001100",
  45667=>"000001110",
  45668=>"000000110",
  45669=>"110000110",
  45670=>"000110001",
  45671=>"001101111",
  45672=>"111000001",
  45673=>"111000001",
  45674=>"110110001",
  45675=>"100100100",
  45676=>"001011100",
  45677=>"101100111",
  45678=>"100000100",
  45679=>"011001000",
  45680=>"000101010",
  45681=>"001100111",
  45682=>"110010100",
  45683=>"001101010",
  45684=>"011001001",
  45685=>"111011111",
  45686=>"110010111",
  45687=>"000100110",
  45688=>"001011000",
  45689=>"111010101",
  45690=>"011111010",
  45691=>"000000111",
  45692=>"010110001",
  45693=>"010011010",
  45694=>"111000101",
  45695=>"100110100",
  45696=>"010010000",
  45697=>"101001011",
  45698=>"101000110",
  45699=>"011010100",
  45700=>"011010000",
  45701=>"111001010",
  45702=>"001111111",
  45703=>"010110010",
  45704=>"011000011",
  45705=>"001001001",
  45706=>"000101110",
  45707=>"011110001",
  45708=>"110011100",
  45709=>"000100100",
  45710=>"110111111",
  45711=>"101100000",
  45712=>"110100001",
  45713=>"100011001",
  45714=>"010101101",
  45715=>"011001000",
  45716=>"100000000",
  45717=>"101000101",
  45718=>"011010001",
  45719=>"101000001",
  45720=>"100010100",
  45721=>"010100000",
  45722=>"001101100",
  45723=>"011111011",
  45724=>"001000101",
  45725=>"011010100",
  45726=>"100100101",
  45727=>"001110010",
  45728=>"101010000",
  45729=>"000010111",
  45730=>"000010110",
  45731=>"100011000",
  45732=>"001001111",
  45733=>"110111011",
  45734=>"010000110",
  45735=>"000101000",
  45736=>"010100110",
  45737=>"101000110",
  45738=>"000000100",
  45739=>"010011001",
  45740=>"101101011",
  45741=>"100000010",
  45742=>"010100100",
  45743=>"111101011",
  45744=>"101001100",
  45745=>"100100101",
  45746=>"011010101",
  45747=>"000010000",
  45748=>"000011100",
  45749=>"010010101",
  45750=>"010100100",
  45751=>"001000110",
  45752=>"001110100",
  45753=>"010000001",
  45754=>"111001101",
  45755=>"001110100",
  45756=>"100010111",
  45757=>"001010111",
  45758=>"111100011",
  45759=>"101100001",
  45760=>"010100110",
  45761=>"000111000",
  45762=>"111000001",
  45763=>"000011000",
  45764=>"111010011",
  45765=>"000011011",
  45766=>"000110111",
  45767=>"110010010",
  45768=>"001001111",
  45769=>"010010010",
  45770=>"111111100",
  45771=>"000011001",
  45772=>"110000100",
  45773=>"010001011",
  45774=>"011110001",
  45775=>"100101001",
  45776=>"000110101",
  45777=>"000010110",
  45778=>"000010010",
  45779=>"011100011",
  45780=>"011110001",
  45781=>"101101111",
  45782=>"010110011",
  45783=>"011000110",
  45784=>"100100111",
  45785=>"011100011",
  45786=>"100001001",
  45787=>"001100000",
  45788=>"110110110",
  45789=>"100010001",
  45790=>"110101010",
  45791=>"011100000",
  45792=>"111011111",
  45793=>"011000110",
  45794=>"110100001",
  45795=>"111100111",
  45796=>"101000011",
  45797=>"000011010",
  45798=>"000010110",
  45799=>"001110111",
  45800=>"100011011",
  45801=>"000010100",
  45802=>"111000011",
  45803=>"001011100",
  45804=>"000101011",
  45805=>"101001111",
  45806=>"001111011",
  45807=>"001010110",
  45808=>"111010111",
  45809=>"110010111",
  45810=>"110111110",
  45811=>"101011110",
  45812=>"110001001",
  45813=>"010001101",
  45814=>"010111111",
  45815=>"000100100",
  45816=>"111001000",
  45817=>"010011110",
  45818=>"001101000",
  45819=>"001010000",
  45820=>"011010110",
  45821=>"001111110",
  45822=>"100100010",
  45823=>"010101001",
  45824=>"110000101",
  45825=>"111111001",
  45826=>"000110011",
  45827=>"101001000",
  45828=>"000010111",
  45829=>"110001101",
  45830=>"100001110",
  45831=>"111111011",
  45832=>"110001100",
  45833=>"010010100",
  45834=>"110111001",
  45835=>"001010001",
  45836=>"000010011",
  45837=>"100011110",
  45838=>"111000100",
  45839=>"011111000",
  45840=>"010011001",
  45841=>"000100000",
  45842=>"111111111",
  45843=>"111011100",
  45844=>"000000010",
  45845=>"100001000",
  45846=>"110001100",
  45847=>"101111110",
  45848=>"001000000",
  45849=>"111010011",
  45850=>"010100010",
  45851=>"011010000",
  45852=>"111110100",
  45853=>"101011010",
  45854=>"011001001",
  45855=>"100011110",
  45856=>"000010011",
  45857=>"110100110",
  45858=>"101110101",
  45859=>"011001100",
  45860=>"110111010",
  45861=>"100001101",
  45862=>"111100000",
  45863=>"101011010",
  45864=>"011010111",
  45865=>"101011101",
  45866=>"000000000",
  45867=>"111111100",
  45868=>"001110110",
  45869=>"000001110",
  45870=>"101110111",
  45871=>"101101101",
  45872=>"001010111",
  45873=>"100110110",
  45874=>"101100101",
  45875=>"000000101",
  45876=>"011100001",
  45877=>"111010000",
  45878=>"111001011",
  45879=>"100101110",
  45880=>"101110000",
  45881=>"101011111",
  45882=>"000011101",
  45883=>"010001011",
  45884=>"101110001",
  45885=>"011100100",
  45886=>"011100011",
  45887=>"110100111",
  45888=>"101100111",
  45889=>"110010000",
  45890=>"101001100",
  45891=>"010110100",
  45892=>"110001111",
  45893=>"101000000",
  45894=>"100000000",
  45895=>"011100111",
  45896=>"010011111",
  45897=>"110111110",
  45898=>"010000111",
  45899=>"001000001",
  45900=>"001000101",
  45901=>"010000110",
  45902=>"110111001",
  45903=>"101011000",
  45904=>"100000110",
  45905=>"011101101",
  45906=>"001100010",
  45907=>"000111100",
  45908=>"110011001",
  45909=>"000001000",
  45910=>"001110101",
  45911=>"111111111",
  45912=>"100110110",
  45913=>"001100001",
  45914=>"011001000",
  45915=>"000011100",
  45916=>"101000011",
  45917=>"101011000",
  45918=>"000011111",
  45919=>"001111010",
  45920=>"000010101",
  45921=>"110111100",
  45922=>"000010110",
  45923=>"100011001",
  45924=>"101111100",
  45925=>"000001101",
  45926=>"000101111",
  45927=>"011111100",
  45928=>"001111111",
  45929=>"111010101",
  45930=>"110000001",
  45931=>"010100011",
  45932=>"001001001",
  45933=>"101111101",
  45934=>"100111100",
  45935=>"011110100",
  45936=>"110000110",
  45937=>"110111100",
  45938=>"111101101",
  45939=>"011110111",
  45940=>"110101010",
  45941=>"100110010",
  45942=>"000100011",
  45943=>"111001101",
  45944=>"001010110",
  45945=>"111010110",
  45946=>"000111011",
  45947=>"101111101",
  45948=>"010001011",
  45949=>"110011010",
  45950=>"100111010",
  45951=>"010010011",
  45952=>"001011110",
  45953=>"001001111",
  45954=>"001110011",
  45955=>"001010011",
  45956=>"100001111",
  45957=>"111101011",
  45958=>"000011000",
  45959=>"000001000",
  45960=>"110101011",
  45961=>"101011101",
  45962=>"010101010",
  45963=>"111111000",
  45964=>"000100100",
  45965=>"101011100",
  45966=>"110000001",
  45967=>"001000000",
  45968=>"001011001",
  45969=>"100011001",
  45970=>"000101100",
  45971=>"100111001",
  45972=>"011110111",
  45973=>"011001111",
  45974=>"010001101",
  45975=>"010111110",
  45976=>"000110000",
  45977=>"010011101",
  45978=>"011100100",
  45979=>"101101011",
  45980=>"011010010",
  45981=>"001010001",
  45982=>"100110000",
  45983=>"010110100",
  45984=>"111010101",
  45985=>"011001000",
  45986=>"101111010",
  45987=>"100001001",
  45988=>"100001010",
  45989=>"100011011",
  45990=>"111001000",
  45991=>"111000100",
  45992=>"000101111",
  45993=>"000001100",
  45994=>"100010110",
  45995=>"111110011",
  45996=>"100010000",
  45997=>"001101000",
  45998=>"000111001",
  45999=>"001101101",
  46000=>"110000010",
  46001=>"101011101",
  46002=>"100111001",
  46003=>"010110000",
  46004=>"100101100",
  46005=>"000111110",
  46006=>"011011011",
  46007=>"011101111",
  46008=>"000011100",
  46009=>"001100101",
  46010=>"011110110",
  46011=>"000000101",
  46012=>"000110011",
  46013=>"101000000",
  46014=>"011000010",
  46015=>"101101100",
  46016=>"000110001",
  46017=>"000110101",
  46018=>"110101101",
  46019=>"001100110",
  46020=>"000001010",
  46021=>"101101001",
  46022=>"110000000",
  46023=>"010000100",
  46024=>"110011001",
  46025=>"111100111",
  46026=>"001101011",
  46027=>"010100011",
  46028=>"100111010",
  46029=>"101001010",
  46030=>"111100111",
  46031=>"100110100",
  46032=>"101100110",
  46033=>"111011001",
  46034=>"000001011",
  46035=>"110010000",
  46036=>"100110111",
  46037=>"010011010",
  46038=>"100100001",
  46039=>"100001010",
  46040=>"010000001",
  46041=>"000100000",
  46042=>"011000000",
  46043=>"101011111",
  46044=>"100011110",
  46045=>"110100100",
  46046=>"111110111",
  46047=>"000101010",
  46048=>"100011011",
  46049=>"100111000",
  46050=>"000001001",
  46051=>"001001001",
  46052=>"001011011",
  46053=>"100011011",
  46054=>"000001110",
  46055=>"001001111",
  46056=>"110000101",
  46057=>"010001001",
  46058=>"010001001",
  46059=>"011101110",
  46060=>"111011111",
  46061=>"001111001",
  46062=>"111111000",
  46063=>"011011011",
  46064=>"100011010",
  46065=>"101100111",
  46066=>"000001110",
  46067=>"110011100",
  46068=>"100010110",
  46069=>"010001010",
  46070=>"101001010",
  46071=>"111001001",
  46072=>"100010110",
  46073=>"011010010",
  46074=>"000111001",
  46075=>"100000011",
  46076=>"101110101",
  46077=>"011111101",
  46078=>"011011010",
  46079=>"110000001",
  46080=>"001101010",
  46081=>"001000011",
  46082=>"111111000",
  46083=>"001011001",
  46084=>"000100001",
  46085=>"011101010",
  46086=>"011001111",
  46087=>"001110101",
  46088=>"010011101",
  46089=>"101101011",
  46090=>"100001101",
  46091=>"010101000",
  46092=>"100111100",
  46093=>"011000011",
  46094=>"001111001",
  46095=>"101101110",
  46096=>"011011001",
  46097=>"100010011",
  46098=>"111100000",
  46099=>"111100000",
  46100=>"011100110",
  46101=>"000110110",
  46102=>"011010000",
  46103=>"100000111",
  46104=>"011011100",
  46105=>"000110011",
  46106=>"000100100",
  46107=>"000100001",
  46108=>"001101110",
  46109=>"000010000",
  46110=>"101100011",
  46111=>"001000110",
  46112=>"010101001",
  46113=>"101001010",
  46114=>"010101101",
  46115=>"111001101",
  46116=>"110001101",
  46117=>"111111011",
  46118=>"111111011",
  46119=>"010001001",
  46120=>"000111010",
  46121=>"111111100",
  46122=>"110111111",
  46123=>"001101101",
  46124=>"000010000",
  46125=>"100000011",
  46126=>"101011000",
  46127=>"001110101",
  46128=>"000000000",
  46129=>"000001000",
  46130=>"010011010",
  46131=>"111111110",
  46132=>"100001111",
  46133=>"000001001",
  46134=>"101010101",
  46135=>"110101011",
  46136=>"100001000",
  46137=>"100010010",
  46138=>"010111011",
  46139=>"111001010",
  46140=>"100100000",
  46141=>"110111111",
  46142=>"110001100",
  46143=>"000011110",
  46144=>"001000000",
  46145=>"100111010",
  46146=>"011010101",
  46147=>"110101110",
  46148=>"011011100",
  46149=>"010110101",
  46150=>"010101100",
  46151=>"111111101",
  46152=>"010101000",
  46153=>"000000001",
  46154=>"010001011",
  46155=>"010001111",
  46156=>"000111010",
  46157=>"110011101",
  46158=>"101001011",
  46159=>"111110101",
  46160=>"000001001",
  46161=>"001110000",
  46162=>"010011000",
  46163=>"011000000",
  46164=>"011000111",
  46165=>"100001010",
  46166=>"110000110",
  46167=>"001101001",
  46168=>"001010001",
  46169=>"111000101",
  46170=>"100000111",
  46171=>"111010000",
  46172=>"000110011",
  46173=>"101000100",
  46174=>"011001111",
  46175=>"101101101",
  46176=>"001100111",
  46177=>"110011001",
  46178=>"101111001",
  46179=>"010101011",
  46180=>"001100010",
  46181=>"111010000",
  46182=>"000000100",
  46183=>"111000100",
  46184=>"000011100",
  46185=>"001010111",
  46186=>"110011001",
  46187=>"111101011",
  46188=>"101001111",
  46189=>"000101001",
  46190=>"111111111",
  46191=>"110010110",
  46192=>"111111111",
  46193=>"010111011",
  46194=>"101111111",
  46195=>"010010000",
  46196=>"011010000",
  46197=>"111011000",
  46198=>"000111011",
  46199=>"000011011",
  46200=>"100111001",
  46201=>"101000000",
  46202=>"001110101",
  46203=>"110001010",
  46204=>"100001010",
  46205=>"110101100",
  46206=>"111110010",
  46207=>"110011100",
  46208=>"111111010",
  46209=>"000000001",
  46210=>"100010101",
  46211=>"110100010",
  46212=>"001001010",
  46213=>"100010000",
  46214=>"110100100",
  46215=>"010000001",
  46216=>"111101100",
  46217=>"011101110",
  46218=>"111000000",
  46219=>"100010100",
  46220=>"111011101",
  46221=>"101001101",
  46222=>"011110010",
  46223=>"011100111",
  46224=>"000000001",
  46225=>"010111101",
  46226=>"100010110",
  46227=>"111011001",
  46228=>"011101101",
  46229=>"111010011",
  46230=>"101000010",
  46231=>"000001110",
  46232=>"000000110",
  46233=>"010101111",
  46234=>"110100000",
  46235=>"000010010",
  46236=>"111111011",
  46237=>"100000101",
  46238=>"000100010",
  46239=>"010100100",
  46240=>"110001011",
  46241=>"110011101",
  46242=>"111101111",
  46243=>"100011011",
  46244=>"001010001",
  46245=>"111110010",
  46246=>"100001101",
  46247=>"001001101",
  46248=>"011011001",
  46249=>"011000011",
  46250=>"101001101",
  46251=>"011001010",
  46252=>"001011111",
  46253=>"001111111",
  46254=>"000101100",
  46255=>"110011110",
  46256=>"011010101",
  46257=>"010010010",
  46258=>"101000101",
  46259=>"001001000",
  46260=>"001011111",
  46261=>"111011100",
  46262=>"111100110",
  46263=>"011100000",
  46264=>"000010011",
  46265=>"111101100",
  46266=>"011101001",
  46267=>"011111011",
  46268=>"001010111",
  46269=>"111111110",
  46270=>"000011110",
  46271=>"010101100",
  46272=>"100011011",
  46273=>"001000101",
  46274=>"111000000",
  46275=>"011011010",
  46276=>"100100010",
  46277=>"001010001",
  46278=>"111000111",
  46279=>"000001111",
  46280=>"011101000",
  46281=>"100010001",
  46282=>"000000011",
  46283=>"110110000",
  46284=>"101101011",
  46285=>"011101000",
  46286=>"000001110",
  46287=>"101000100",
  46288=>"001000001",
  46289=>"001010101",
  46290=>"101011100",
  46291=>"010000000",
  46292=>"110011000",
  46293=>"110000000",
  46294=>"101011011",
  46295=>"000000000",
  46296=>"100110001",
  46297=>"101100101",
  46298=>"100111001",
  46299=>"001000110",
  46300=>"010110111",
  46301=>"011111000",
  46302=>"111000010",
  46303=>"011001111",
  46304=>"111101001",
  46305=>"010110000",
  46306=>"000010000",
  46307=>"001111101",
  46308=>"000111101",
  46309=>"111000011",
  46310=>"101011000",
  46311=>"010111011",
  46312=>"110011110",
  46313=>"001000101",
  46314=>"111110110",
  46315=>"001000000",
  46316=>"011010010",
  46317=>"011000010",
  46318=>"011100011",
  46319=>"111110111",
  46320=>"101110011",
  46321=>"010100101",
  46322=>"001001010",
  46323=>"101000001",
  46324=>"001000111",
  46325=>"000000111",
  46326=>"001110101",
  46327=>"000011111",
  46328=>"001000101",
  46329=>"010110001",
  46330=>"111100011",
  46331=>"000011100",
  46332=>"110011011",
  46333=>"000011011",
  46334=>"011110100",
  46335=>"010000110",
  46336=>"101010000",
  46337=>"000010000",
  46338=>"010011110",
  46339=>"010000010",
  46340=>"010101110",
  46341=>"111010011",
  46342=>"100100101",
  46343=>"000100101",
  46344=>"000000000",
  46345=>"101010011",
  46346=>"011000001",
  46347=>"100010100",
  46348=>"110111001",
  46349=>"101011011",
  46350=>"100010000",
  46351=>"111001100",
  46352=>"001111010",
  46353=>"101111101",
  46354=>"111001101",
  46355=>"100000101",
  46356=>"111111100",
  46357=>"101111010",
  46358=>"111111100",
  46359=>"100110111",
  46360=>"110101011",
  46361=>"000101010",
  46362=>"110111000",
  46363=>"000101010",
  46364=>"111000110",
  46365=>"001111010",
  46366=>"110101100",
  46367=>"111011001",
  46368=>"000001010",
  46369=>"000010000",
  46370=>"101001111",
  46371=>"011000110",
  46372=>"110110010",
  46373=>"011111000",
  46374=>"011101110",
  46375=>"110000000",
  46376=>"100010110",
  46377=>"100110111",
  46378=>"000000000",
  46379=>"010010010",
  46380=>"110001100",
  46381=>"001010100",
  46382=>"111111110",
  46383=>"000101110",
  46384=>"100101011",
  46385=>"110101011",
  46386=>"111110001",
  46387=>"100011000",
  46388=>"010101001",
  46389=>"101001000",
  46390=>"000100001",
  46391=>"111010011",
  46392=>"001110110",
  46393=>"011001100",
  46394=>"100111100",
  46395=>"001111100",
  46396=>"101001101",
  46397=>"100100100",
  46398=>"101110111",
  46399=>"000010000",
  46400=>"000010011",
  46401=>"000000101",
  46402=>"110110100",
  46403=>"110011111",
  46404=>"101111000",
  46405=>"110011101",
  46406=>"000000110",
  46407=>"100011101",
  46408=>"110100111",
  46409=>"100101111",
  46410=>"010000100",
  46411=>"001011000",
  46412=>"101110110",
  46413=>"010111100",
  46414=>"011111000",
  46415=>"110011100",
  46416=>"010000110",
  46417=>"011000010",
  46418=>"111110010",
  46419=>"110110100",
  46420=>"110001101",
  46421=>"011100000",
  46422=>"111101111",
  46423=>"111011011",
  46424=>"100001000",
  46425=>"100101111",
  46426=>"010100110",
  46427=>"011000000",
  46428=>"011000000",
  46429=>"010100001",
  46430=>"010000001",
  46431=>"111001111",
  46432=>"000111101",
  46433=>"110111110",
  46434=>"110000011",
  46435=>"100100010",
  46436=>"110101111",
  46437=>"111111010",
  46438=>"100000111",
  46439=>"011010111",
  46440=>"011010011",
  46441=>"111101101",
  46442=>"101000010",
  46443=>"101011000",
  46444=>"101000110",
  46445=>"000101001",
  46446=>"110000010",
  46447=>"010101011",
  46448=>"111010000",
  46449=>"111010001",
  46450=>"110010011",
  46451=>"001000110",
  46452=>"001010000",
  46453=>"010110010",
  46454=>"111110110",
  46455=>"100101101",
  46456=>"001000000",
  46457=>"010010011",
  46458=>"010001111",
  46459=>"100000011",
  46460=>"110000000",
  46461=>"010001110",
  46462=>"111001110",
  46463=>"111011110",
  46464=>"111100111",
  46465=>"010100100",
  46466=>"011011000",
  46467=>"010000101",
  46468=>"000100001",
  46469=>"010110101",
  46470=>"001110111",
  46471=>"110010111",
  46472=>"001100100",
  46473=>"111100111",
  46474=>"001001001",
  46475=>"011111000",
  46476=>"101001111",
  46477=>"110010000",
  46478=>"011110001",
  46479=>"000110011",
  46480=>"101110111",
  46481=>"010000010",
  46482=>"001001011",
  46483=>"000011100",
  46484=>"110110000",
  46485=>"111110010",
  46486=>"100110110",
  46487=>"000100101",
  46488=>"110101111",
  46489=>"111011000",
  46490=>"010000111",
  46491=>"000100001",
  46492=>"010110110",
  46493=>"000000000",
  46494=>"110011000",
  46495=>"110010001",
  46496=>"111101101",
  46497=>"000100100",
  46498=>"110100001",
  46499=>"001011000",
  46500=>"100101110",
  46501=>"000101100",
  46502=>"011110001",
  46503=>"000001011",
  46504=>"111111110",
  46505=>"111011111",
  46506=>"100101001",
  46507=>"001101001",
  46508=>"101000000",
  46509=>"001001110",
  46510=>"001011100",
  46511=>"111111111",
  46512=>"101111101",
  46513=>"111111111",
  46514=>"011101111",
  46515=>"100101110",
  46516=>"100011000",
  46517=>"100001010",
  46518=>"111000000",
  46519=>"010011000",
  46520=>"000100101",
  46521=>"111001010",
  46522=>"011000111",
  46523=>"100000110",
  46524=>"011011000",
  46525=>"101001111",
  46526=>"010010001",
  46527=>"011101101",
  46528=>"101000111",
  46529=>"110011111",
  46530=>"011101111",
  46531=>"110101111",
  46532=>"100011011",
  46533=>"000000101",
  46534=>"111101100",
  46535=>"111111101",
  46536=>"001101010",
  46537=>"101100011",
  46538=>"011011110",
  46539=>"000111010",
  46540=>"001011111",
  46541=>"011111100",
  46542=>"000000010",
  46543=>"111011001",
  46544=>"101100000",
  46545=>"111011000",
  46546=>"001101111",
  46547=>"001101010",
  46548=>"011110011",
  46549=>"010010011",
  46550=>"101011011",
  46551=>"111001101",
  46552=>"110110001",
  46553=>"010100000",
  46554=>"011101011",
  46555=>"000110101",
  46556=>"100011001",
  46557=>"110110110",
  46558=>"000000111",
  46559=>"000100110",
  46560=>"101110010",
  46561=>"011001010",
  46562=>"101110111",
  46563=>"000000110",
  46564=>"011011101",
  46565=>"110110110",
  46566=>"001100110",
  46567=>"110100101",
  46568=>"000101110",
  46569=>"010011100",
  46570=>"010111110",
  46571=>"011111001",
  46572=>"101100111",
  46573=>"001111111",
  46574=>"000011100",
  46575=>"110000111",
  46576=>"100001011",
  46577=>"110011100",
  46578=>"100111110",
  46579=>"101110111",
  46580=>"101010100",
  46581=>"000000110",
  46582=>"101001011",
  46583=>"010000000",
  46584=>"110101110",
  46585=>"011100000",
  46586=>"111011100",
  46587=>"000010000",
  46588=>"000011000",
  46589=>"011100000",
  46590=>"001011011",
  46591=>"001111111",
  46592=>"000110000",
  46593=>"110001100",
  46594=>"110010100",
  46595=>"111100111",
  46596=>"000101101",
  46597=>"000110101",
  46598=>"010000010",
  46599=>"110010100",
  46600=>"000101101",
  46601=>"100110110",
  46602=>"000010000",
  46603=>"110010111",
  46604=>"100111010",
  46605=>"111010000",
  46606=>"111101110",
  46607=>"111011111",
  46608=>"110101100",
  46609=>"010000100",
  46610=>"101001010",
  46611=>"101001011",
  46612=>"010000001",
  46613=>"000011110",
  46614=>"011001001",
  46615=>"111011111",
  46616=>"100000110",
  46617=>"001100000",
  46618=>"001011001",
  46619=>"101111110",
  46620=>"010000100",
  46621=>"001001011",
  46622=>"110010010",
  46623=>"001010001",
  46624=>"101101110",
  46625=>"011011111",
  46626=>"111101111",
  46627=>"001010110",
  46628=>"000010001",
  46629=>"010100000",
  46630=>"000011101",
  46631=>"011001111",
  46632=>"011000011",
  46633=>"000101010",
  46634=>"100100010",
  46635=>"101011000",
  46636=>"000000011",
  46637=>"010011100",
  46638=>"001100000",
  46639=>"000000100",
  46640=>"110000100",
  46641=>"000101010",
  46642=>"100010110",
  46643=>"101010101",
  46644=>"100110010",
  46645=>"010001111",
  46646=>"000100000",
  46647=>"101011110",
  46648=>"110011010",
  46649=>"011111100",
  46650=>"100000110",
  46651=>"000111001",
  46652=>"110111111",
  46653=>"001000101",
  46654=>"010000000",
  46655=>"000110011",
  46656=>"100101110",
  46657=>"000100100",
  46658=>"000001011",
  46659=>"111011110",
  46660=>"000101001",
  46661=>"111110000",
  46662=>"001001011",
  46663=>"010000001",
  46664=>"101111000",
  46665=>"010011010",
  46666=>"010011100",
  46667=>"000101100",
  46668=>"001111001",
  46669=>"111100000",
  46670=>"110000111",
  46671=>"010111111",
  46672=>"010111000",
  46673=>"110110010",
  46674=>"010000011",
  46675=>"000110110",
  46676=>"111010001",
  46677=>"101011011",
  46678=>"111001111",
  46679=>"010010110",
  46680=>"001110111",
  46681=>"101111101",
  46682=>"111100110",
  46683=>"011110110",
  46684=>"000000110",
  46685=>"110000100",
  46686=>"101101101",
  46687=>"100001001",
  46688=>"001100101",
  46689=>"110000001",
  46690=>"000001100",
  46691=>"111000110",
  46692=>"000000011",
  46693=>"110100000",
  46694=>"101110111",
  46695=>"111001100",
  46696=>"111111100",
  46697=>"101111011",
  46698=>"100000001",
  46699=>"011011000",
  46700=>"111011101",
  46701=>"100100000",
  46702=>"111011010",
  46703=>"011010101",
  46704=>"111100100",
  46705=>"001100110",
  46706=>"001001011",
  46707=>"011000011",
  46708=>"101110101",
  46709=>"010010010",
  46710=>"010111101",
  46711=>"011101000",
  46712=>"011111010",
  46713=>"101100110",
  46714=>"111110010",
  46715=>"100110010",
  46716=>"110000010",
  46717=>"110001001",
  46718=>"100001111",
  46719=>"110111101",
  46720=>"010010100",
  46721=>"010000100",
  46722=>"101101100",
  46723=>"101101000",
  46724=>"011000000",
  46725=>"000001000",
  46726=>"001101100",
  46727=>"010110001",
  46728=>"110101010",
  46729=>"001101110",
  46730=>"000011100",
  46731=>"011011011",
  46732=>"100111000",
  46733=>"011111011",
  46734=>"111001000",
  46735=>"101100000",
  46736=>"110001111",
  46737=>"110000010",
  46738=>"111010110",
  46739=>"010010110",
  46740=>"111011100",
  46741=>"001101001",
  46742=>"000101011",
  46743=>"111101111",
  46744=>"010001011",
  46745=>"100110111",
  46746=>"011001000",
  46747=>"111001111",
  46748=>"011010001",
  46749=>"111010011",
  46750=>"100010010",
  46751=>"110111110",
  46752=>"110100010",
  46753=>"010010011",
  46754=>"111010001",
  46755=>"110110001",
  46756=>"110110101",
  46757=>"101101010",
  46758=>"111011010",
  46759=>"110011111",
  46760=>"100001010",
  46761=>"111000101",
  46762=>"001111000",
  46763=>"111001001",
  46764=>"111101001",
  46765=>"100110010",
  46766=>"000000010",
  46767=>"011011111",
  46768=>"001000110",
  46769=>"001011100",
  46770=>"000101111",
  46771=>"100101001",
  46772=>"001000010",
  46773=>"110001010",
  46774=>"011111000",
  46775=>"100100111",
  46776=>"110010100",
  46777=>"101100100",
  46778=>"111011001",
  46779=>"010000110",
  46780=>"110101100",
  46781=>"010111010",
  46782=>"000100001",
  46783=>"100010110",
  46784=>"000010101",
  46785=>"001111100",
  46786=>"011111111",
  46787=>"000101111",
  46788=>"010001110",
  46789=>"111110111",
  46790=>"000110101",
  46791=>"000001001",
  46792=>"101000100",
  46793=>"111010011",
  46794=>"011101000",
  46795=>"111111110",
  46796=>"001010010",
  46797=>"001101100",
  46798=>"000100001",
  46799=>"010010010",
  46800=>"110100101",
  46801=>"010101011",
  46802=>"001100110",
  46803=>"010000001",
  46804=>"111000000",
  46805=>"011111111",
  46806=>"001010111",
  46807=>"011111010",
  46808=>"100001111",
  46809=>"001000011",
  46810=>"111010000",
  46811=>"010111100",
  46812=>"101100100",
  46813=>"100001101",
  46814=>"111111100",
  46815=>"000110110",
  46816=>"101010000",
  46817=>"111011101",
  46818=>"111011111",
  46819=>"010111011",
  46820=>"000101000",
  46821=>"101000110",
  46822=>"000001111",
  46823=>"111000010",
  46824=>"010110101",
  46825=>"101111010",
  46826=>"101000111",
  46827=>"100111010",
  46828=>"001001001",
  46829=>"001011101",
  46830=>"000101101",
  46831=>"000010100",
  46832=>"100001001",
  46833=>"100100001",
  46834=>"010101011",
  46835=>"101000011",
  46836=>"110101100",
  46837=>"110010111",
  46838=>"110111111",
  46839=>"100110001",
  46840=>"100001111",
  46841=>"010010111",
  46842=>"001001011",
  46843=>"101001001",
  46844=>"001101000",
  46845=>"011100000",
  46846=>"010001001",
  46847=>"010010111",
  46848=>"001000000",
  46849=>"111010100",
  46850=>"011010001",
  46851=>"011001110",
  46852=>"000100011",
  46853=>"000101011",
  46854=>"001011010",
  46855=>"000011101",
  46856=>"111000101",
  46857=>"111101010",
  46858=>"001000001",
  46859=>"100110111",
  46860=>"110101110",
  46861=>"010110110",
  46862=>"101111101",
  46863=>"010100110",
  46864=>"111110110",
  46865=>"101000011",
  46866=>"110110101",
  46867=>"100111011",
  46868=>"001001011",
  46869=>"011010011",
  46870=>"110100011",
  46871=>"100101010",
  46872=>"001000111",
  46873=>"100100011",
  46874=>"001011000",
  46875=>"010110011",
  46876=>"010011100",
  46877=>"000010110",
  46878=>"111011000",
  46879=>"100010011",
  46880=>"010111110",
  46881=>"110001100",
  46882=>"010101000",
  46883=>"111001011",
  46884=>"000100101",
  46885=>"000100011",
  46886=>"110000100",
  46887=>"001110101",
  46888=>"010101010",
  46889=>"010100000",
  46890=>"101011000",
  46891=>"100100100",
  46892=>"011001100",
  46893=>"010111001",
  46894=>"001000010",
  46895=>"001010001",
  46896=>"100101011",
  46897=>"001000010",
  46898=>"111100101",
  46899=>"000000010",
  46900=>"000100101",
  46901=>"010110001",
  46902=>"101110110",
  46903=>"110010010",
  46904=>"101000101",
  46905=>"101000000",
  46906=>"000010111",
  46907=>"101011101",
  46908=>"111000100",
  46909=>"101011001",
  46910=>"001001101",
  46911=>"100101000",
  46912=>"011101011",
  46913=>"000000110",
  46914=>"111101111",
  46915=>"110100111",
  46916=>"100100101",
  46917=>"111000100",
  46918=>"010000010",
  46919=>"110010101",
  46920=>"111110111",
  46921=>"001010111",
  46922=>"111001000",
  46923=>"011111100",
  46924=>"110010000",
  46925=>"011011010",
  46926=>"000110100",
  46927=>"001101111",
  46928=>"111000111",
  46929=>"111100011",
  46930=>"000111100",
  46931=>"010011010",
  46932=>"010000000",
  46933=>"000001010",
  46934=>"101011001",
  46935=>"000010101",
  46936=>"001000110",
  46937=>"110011010",
  46938=>"100101010",
  46939=>"101101100",
  46940=>"111000001",
  46941=>"001000100",
  46942=>"001110001",
  46943=>"101111011",
  46944=>"100101110",
  46945=>"100110011",
  46946=>"101100011",
  46947=>"011101000",
  46948=>"011000110",
  46949=>"000110110",
  46950=>"110110011",
  46951=>"101000111",
  46952=>"001001001",
  46953=>"000110101",
  46954=>"001001001",
  46955=>"001110111",
  46956=>"000000001",
  46957=>"100111001",
  46958=>"110101010",
  46959=>"111001000",
  46960=>"001011011",
  46961=>"110011101",
  46962=>"011010011",
  46963=>"101011011",
  46964=>"000111100",
  46965=>"111101100",
  46966=>"100110110",
  46967=>"010000010",
  46968=>"011011001",
  46969=>"010101110",
  46970=>"111101101",
  46971=>"001100011",
  46972=>"001111001",
  46973=>"001011001",
  46974=>"101100111",
  46975=>"000100100",
  46976=>"000001010",
  46977=>"111001001",
  46978=>"011111011",
  46979=>"101110011",
  46980=>"100001110",
  46981=>"101110110",
  46982=>"101100111",
  46983=>"101110000",
  46984=>"000010001",
  46985=>"110011001",
  46986=>"010110111",
  46987=>"010111000",
  46988=>"101110101",
  46989=>"010001111",
  46990=>"011100000",
  46991=>"100001101",
  46992=>"111000001",
  46993=>"000100011",
  46994=>"111101001",
  46995=>"111111111",
  46996=>"011011111",
  46997=>"110000011",
  46998=>"010011010",
  46999=>"101111001",
  47000=>"110011110",
  47001=>"111100100",
  47002=>"010111011",
  47003=>"011111000",
  47004=>"010110101",
  47005=>"000010101",
  47006=>"010010001",
  47007=>"111000100",
  47008=>"101000111",
  47009=>"110100111",
  47010=>"110100111",
  47011=>"001101110",
  47012=>"101111101",
  47013=>"010010011",
  47014=>"001111101",
  47015=>"111110111",
  47016=>"011001001",
  47017=>"101111110",
  47018=>"000010001",
  47019=>"010100100",
  47020=>"101100011",
  47021=>"111011010",
  47022=>"111011111",
  47023=>"001100010",
  47024=>"110011010",
  47025=>"101000111",
  47026=>"000101001",
  47027=>"000000111",
  47028=>"101011110",
  47029=>"011110000",
  47030=>"110011100",
  47031=>"101111111",
  47032=>"001110110",
  47033=>"111011111",
  47034=>"110110101",
  47035=>"111100101",
  47036=>"010010000",
  47037=>"010010011",
  47038=>"000000001",
  47039=>"111011101",
  47040=>"101001001",
  47041=>"010101110",
  47042=>"001110000",
  47043=>"000101110",
  47044=>"110010011",
  47045=>"011010011",
  47046=>"100101001",
  47047=>"010000100",
  47048=>"010100111",
  47049=>"100110011",
  47050=>"010000001",
  47051=>"001101101",
  47052=>"111111010",
  47053=>"110111111",
  47054=>"110000011",
  47055=>"101110110",
  47056=>"011110100",
  47057=>"110000110",
  47058=>"011110000",
  47059=>"111101010",
  47060=>"000100011",
  47061=>"000001000",
  47062=>"000100000",
  47063=>"010010100",
  47064=>"000110000",
  47065=>"000111100",
  47066=>"110111100",
  47067=>"011010011",
  47068=>"111110010",
  47069=>"100110111",
  47070=>"001000100",
  47071=>"000100111",
  47072=>"000011010",
  47073=>"110001111",
  47074=>"111010010",
  47075=>"101001101",
  47076=>"111101101",
  47077=>"000000100",
  47078=>"011000001",
  47079=>"100111100",
  47080=>"000001111",
  47081=>"000011011",
  47082=>"010011010",
  47083=>"001001110",
  47084=>"011010001",
  47085=>"000010110",
  47086=>"011011010",
  47087=>"111100100",
  47088=>"010011100",
  47089=>"100101101",
  47090=>"001010010",
  47091=>"101101001",
  47092=>"101000001",
  47093=>"011011100",
  47094=>"000111110",
  47095=>"010110010",
  47096=>"111110011",
  47097=>"011110111",
  47098=>"101110100",
  47099=>"000110100",
  47100=>"001010000",
  47101=>"000000100",
  47102=>"001011010",
  47103=>"100111110",
  47104=>"000001111",
  47105=>"010101111",
  47106=>"000100100",
  47107=>"100000111",
  47108=>"011000011",
  47109=>"001101101",
  47110=>"000010101",
  47111=>"111100000",
  47112=>"111111110",
  47113=>"100111101",
  47114=>"011011000",
  47115=>"011010001",
  47116=>"010001110",
  47117=>"100010100",
  47118=>"101001110",
  47119=>"010110000",
  47120=>"100111010",
  47121=>"110111011",
  47122=>"100011011",
  47123=>"100110010",
  47124=>"100010111",
  47125=>"001001001",
  47126=>"111001001",
  47127=>"110100011",
  47128=>"001111010",
  47129=>"001000110",
  47130=>"101110111",
  47131=>"111111011",
  47132=>"001001110",
  47133=>"000010011",
  47134=>"001000100",
  47135=>"010010101",
  47136=>"100001000",
  47137=>"011000100",
  47138=>"010000001",
  47139=>"100110110",
  47140=>"101001011",
  47141=>"001100000",
  47142=>"011011001",
  47143=>"101111110",
  47144=>"000101011",
  47145=>"000000101",
  47146=>"010000101",
  47147=>"110110010",
  47148=>"101100001",
  47149=>"111001001",
  47150=>"110011101",
  47151=>"101001000",
  47152=>"000110001",
  47153=>"100110100",
  47154=>"000001010",
  47155=>"010011100",
  47156=>"110011011",
  47157=>"000100100",
  47158=>"110111011",
  47159=>"100101011",
  47160=>"000111110",
  47161=>"000100101",
  47162=>"001011010",
  47163=>"001001111",
  47164=>"010011001",
  47165=>"111100101",
  47166=>"011010011",
  47167=>"100000110",
  47168=>"101110100",
  47169=>"000111010",
  47170=>"101111000",
  47171=>"100010000",
  47172=>"101110111",
  47173=>"101011010",
  47174=>"000010011",
  47175=>"100010001",
  47176=>"001001111",
  47177=>"011011001",
  47178=>"111001011",
  47179=>"001110100",
  47180=>"000010010",
  47181=>"010101111",
  47182=>"001111000",
  47183=>"011110001",
  47184=>"100110001",
  47185=>"111101101",
  47186=>"111101010",
  47187=>"000011111",
  47188=>"111110011",
  47189=>"000111101",
  47190=>"010111101",
  47191=>"110110010",
  47192=>"001010011",
  47193=>"000001011",
  47194=>"101001100",
  47195=>"010010101",
  47196=>"000000010",
  47197=>"000001010",
  47198=>"101000110",
  47199=>"100011110",
  47200=>"111111111",
  47201=>"011011000",
  47202=>"011101000",
  47203=>"100100101",
  47204=>"111010010",
  47205=>"001010101",
  47206=>"101010001",
  47207=>"000111000",
  47208=>"101001100",
  47209=>"101010011",
  47210=>"000000010",
  47211=>"100110000",
  47212=>"011111111",
  47213=>"101110110",
  47214=>"101111101",
  47215=>"001000001",
  47216=>"110011000",
  47217=>"010010010",
  47218=>"111010010",
  47219=>"111010101",
  47220=>"110000110",
  47221=>"001100110",
  47222=>"111001011",
  47223=>"100010100",
  47224=>"111101110",
  47225=>"011010010",
  47226=>"111100001",
  47227=>"010011010",
  47228=>"101000101",
  47229=>"100001101",
  47230=>"000100010",
  47231=>"011010010",
  47232=>"100001110",
  47233=>"010011110",
  47234=>"011011001",
  47235=>"000000111",
  47236=>"101101001",
  47237=>"110110100",
  47238=>"101001110",
  47239=>"101101000",
  47240=>"001100000",
  47241=>"000100011",
  47242=>"000000101",
  47243=>"111010110",
  47244=>"000011110",
  47245=>"011110111",
  47246=>"001100000",
  47247=>"001110010",
  47248=>"011110111",
  47249=>"110011111",
  47250=>"010100001",
  47251=>"111110100",
  47252=>"000000110",
  47253=>"010000011",
  47254=>"000010010",
  47255=>"000100111",
  47256=>"000110101",
  47257=>"111001011",
  47258=>"010011101",
  47259=>"110101001",
  47260=>"010011000",
  47261=>"100001110",
  47262=>"111111101",
  47263=>"111101101",
  47264=>"101111100",
  47265=>"101010111",
  47266=>"010001000",
  47267=>"100010010",
  47268=>"000100110",
  47269=>"000111111",
  47270=>"011100111",
  47271=>"010001110",
  47272=>"011111111",
  47273=>"001011111",
  47274=>"011011101",
  47275=>"110100011",
  47276=>"010101000",
  47277=>"100101110",
  47278=>"101010111",
  47279=>"110100101",
  47280=>"011100101",
  47281=>"110101000",
  47282=>"101001110",
  47283=>"000111100",
  47284=>"100111101",
  47285=>"010111001",
  47286=>"111110110",
  47287=>"101100101",
  47288=>"000010000",
  47289=>"000011010",
  47290=>"000101100",
  47291=>"110001110",
  47292=>"001111101",
  47293=>"100011001",
  47294=>"011101010",
  47295=>"111000010",
  47296=>"100110101",
  47297=>"110011000",
  47298=>"111001101",
  47299=>"010010100",
  47300=>"000111011",
  47301=>"101010011",
  47302=>"110001111",
  47303=>"110100101",
  47304=>"101001111",
  47305=>"001000001",
  47306=>"110101100",
  47307=>"101110001",
  47308=>"110111011",
  47309=>"110011110",
  47310=>"100101011",
  47311=>"101001111",
  47312=>"011011001",
  47313=>"111000100",
  47314=>"010100100",
  47315=>"011001100",
  47316=>"001100101",
  47317=>"100111111",
  47318=>"001010001",
  47319=>"000111011",
  47320=>"101101101",
  47321=>"100001001",
  47322=>"001001000",
  47323=>"111100110",
  47324=>"111011101",
  47325=>"010111000",
  47326=>"010011000",
  47327=>"011101001",
  47328=>"001000010",
  47329=>"001100111",
  47330=>"110100110",
  47331=>"101010001",
  47332=>"011111000",
  47333=>"010011010",
  47334=>"100100000",
  47335=>"100011100",
  47336=>"000110111",
  47337=>"101011001",
  47338=>"110111110",
  47339=>"000000001",
  47340=>"001100000",
  47341=>"001111010",
  47342=>"101000111",
  47343=>"101111001",
  47344=>"011010011",
  47345=>"010111010",
  47346=>"000101000",
  47347=>"011110100",
  47348=>"101100011",
  47349=>"001101110",
  47350=>"100000000",
  47351=>"111111001",
  47352=>"111110000",
  47353=>"000100111",
  47354=>"001011110",
  47355=>"100101001",
  47356=>"001010111",
  47357=>"001111001",
  47358=>"010000001",
  47359=>"001001011",
  47360=>"001000100",
  47361=>"110010101",
  47362=>"011011110",
  47363=>"000100100",
  47364=>"011011111",
  47365=>"100100010",
  47366=>"101100111",
  47367=>"101011010",
  47368=>"011010110",
  47369=>"010010110",
  47370=>"000001000",
  47371=>"110011000",
  47372=>"010000011",
  47373=>"111110010",
  47374=>"000011101",
  47375=>"001101110",
  47376=>"110101011",
  47377=>"000011101",
  47378=>"111101010",
  47379=>"011100110",
  47380=>"110001100",
  47381=>"000111000",
  47382=>"001100010",
  47383=>"001001111",
  47384=>"001000101",
  47385=>"000011001",
  47386=>"111111000",
  47387=>"001101111",
  47388=>"100110110",
  47389=>"111100000",
  47390=>"101111101",
  47391=>"010000001",
  47392=>"000110001",
  47393=>"111000101",
  47394=>"000011110",
  47395=>"101111011",
  47396=>"100001000",
  47397=>"110101100",
  47398=>"000010110",
  47399=>"111001011",
  47400=>"111011100",
  47401=>"010000000",
  47402=>"100100011",
  47403=>"110110111",
  47404=>"001101000",
  47405=>"111101111",
  47406=>"100000111",
  47407=>"111100110",
  47408=>"000111001",
  47409=>"111111010",
  47410=>"011000000",
  47411=>"000010110",
  47412=>"110010001",
  47413=>"011000010",
  47414=>"011001111",
  47415=>"101110000",
  47416=>"111010111",
  47417=>"000000100",
  47418=>"110111001",
  47419=>"111011101",
  47420=>"011111000",
  47421=>"110110001",
  47422=>"001100101",
  47423=>"110101011",
  47424=>"101001000",
  47425=>"100101011",
  47426=>"000001100",
  47427=>"010010111",
  47428=>"101100010",
  47429=>"010111100",
  47430=>"110100101",
  47431=>"000111111",
  47432=>"100000100",
  47433=>"010110010",
  47434=>"010011110",
  47435=>"110110100",
  47436=>"011001000",
  47437=>"000001111",
  47438=>"001010000",
  47439=>"000101000",
  47440=>"110000011",
  47441=>"010001101",
  47442=>"011011110",
  47443=>"000001000",
  47444=>"011000100",
  47445=>"010011001",
  47446=>"001010110",
  47447=>"011000011",
  47448=>"001100000",
  47449=>"001000010",
  47450=>"000111100",
  47451=>"011110011",
  47452=>"110001110",
  47453=>"011000011",
  47454=>"100100100",
  47455=>"001001110",
  47456=>"011011001",
  47457=>"011100011",
  47458=>"111111111",
  47459=>"000110110",
  47460=>"000000000",
  47461=>"101010010",
  47462=>"000101001",
  47463=>"101111001",
  47464=>"010001100",
  47465=>"111100010",
  47466=>"010000110",
  47467=>"000000110",
  47468=>"001000101",
  47469=>"111010110",
  47470=>"000010101",
  47471=>"001000010",
  47472=>"000010111",
  47473=>"110011001",
  47474=>"001001010",
  47475=>"011001011",
  47476=>"111100100",
  47477=>"100010101",
  47478=>"100100110",
  47479=>"000011101",
  47480=>"001010110",
  47481=>"000101110",
  47482=>"000010111",
  47483=>"001001111",
  47484=>"000001100",
  47485=>"100101100",
  47486=>"100111010",
  47487=>"110001110",
  47488=>"000110000",
  47489=>"100101110",
  47490=>"110100010",
  47491=>"101101000",
  47492=>"001110110",
  47493=>"110111000",
  47494=>"011110010",
  47495=>"110101001",
  47496=>"001011101",
  47497=>"011010000",
  47498=>"101111100",
  47499=>"000000011",
  47500=>"000101100",
  47501=>"100110111",
  47502=>"100101100",
  47503=>"110100111",
  47504=>"110011100",
  47505=>"100000111",
  47506=>"111101001",
  47507=>"001111111",
  47508=>"000100110",
  47509=>"010111100",
  47510=>"101101001",
  47511=>"111100111",
  47512=>"010000010",
  47513=>"011000001",
  47514=>"111101001",
  47515=>"101110011",
  47516=>"101100111",
  47517=>"111110101",
  47518=>"001110111",
  47519=>"001101000",
  47520=>"111011100",
  47521=>"011100101",
  47522=>"111111100",
  47523=>"000010011",
  47524=>"111010111",
  47525=>"101101000",
  47526=>"010111111",
  47527=>"111000111",
  47528=>"101100011",
  47529=>"111110010",
  47530=>"001110011",
  47531=>"110001000",
  47532=>"101001101",
  47533=>"000110001",
  47534=>"111111011",
  47535=>"010000000",
  47536=>"111111010",
  47537=>"010010001",
  47538=>"110110011",
  47539=>"111100000",
  47540=>"001111010",
  47541=>"101011000",
  47542=>"110100000",
  47543=>"011000010",
  47544=>"100000111",
  47545=>"010100010",
  47546=>"010000010",
  47547=>"110101111",
  47548=>"000011010",
  47549=>"111011100",
  47550=>"100000101",
  47551=>"001100101",
  47552=>"111000110",
  47553=>"111101010",
  47554=>"000100101",
  47555=>"101111010",
  47556=>"100110001",
  47557=>"011001100",
  47558=>"111000000",
  47559=>"000100110",
  47560=>"001000010",
  47561=>"000000001",
  47562=>"101000000",
  47563=>"100110111",
  47564=>"100000110",
  47565=>"001010111",
  47566=>"101011010",
  47567=>"100010010",
  47568=>"101011100",
  47569=>"111110101",
  47570=>"101101101",
  47571=>"110001001",
  47572=>"100101111",
  47573=>"100110010",
  47574=>"001101000",
  47575=>"001100100",
  47576=>"101110010",
  47577=>"101001110",
  47578=>"110111110",
  47579=>"111110100",
  47580=>"101101000",
  47581=>"001010110",
  47582=>"111100011",
  47583=>"000000001",
  47584=>"011001001",
  47585=>"000011011",
  47586=>"111000000",
  47587=>"100011001",
  47588=>"000111100",
  47589=>"001011101",
  47590=>"000100110",
  47591=>"110110110",
  47592=>"000010010",
  47593=>"110011111",
  47594=>"100110000",
  47595=>"010001101",
  47596=>"000000010",
  47597=>"101101001",
  47598=>"000010000",
  47599=>"000110111",
  47600=>"100001101",
  47601=>"101110101",
  47602=>"101100001",
  47603=>"111000111",
  47604=>"001001011",
  47605=>"001101101",
  47606=>"110101110",
  47607=>"001110110",
  47608=>"011010110",
  47609=>"111110100",
  47610=>"010010110",
  47611=>"111001001",
  47612=>"101010001",
  47613=>"110001001",
  47614=>"100010101",
  47615=>"101000110",
  47616=>"100100100",
  47617=>"111111011",
  47618=>"111001011",
  47619=>"010011001",
  47620=>"100010000",
  47621=>"011111010",
  47622=>"011111000",
  47623=>"110111010",
  47624=>"101111100",
  47625=>"111111110",
  47626=>"000000111",
  47627=>"000000010",
  47628=>"011100110",
  47629=>"111011101",
  47630=>"001010000",
  47631=>"000010001",
  47632=>"011010011",
  47633=>"000011010",
  47634=>"011110101",
  47635=>"100101011",
  47636=>"010001100",
  47637=>"001010001",
  47638=>"101011001",
  47639=>"101110000",
  47640=>"111101111",
  47641=>"110000000",
  47642=>"110101001",
  47643=>"111000101",
  47644=>"110001011",
  47645=>"110111001",
  47646=>"010111111",
  47647=>"111000111",
  47648=>"011011010",
  47649=>"111101110",
  47650=>"001000100",
  47651=>"000111010",
  47652=>"111000101",
  47653=>"100101111",
  47654=>"010100101",
  47655=>"100000101",
  47656=>"001011110",
  47657=>"010010110",
  47658=>"111110010",
  47659=>"010111110",
  47660=>"000110000",
  47661=>"110101000",
  47662=>"001100000",
  47663=>"100010010",
  47664=>"110001010",
  47665=>"000010001",
  47666=>"000000000",
  47667=>"100001010",
  47668=>"001001100",
  47669=>"011110011",
  47670=>"101011011",
  47671=>"000000001",
  47672=>"010101101",
  47673=>"111101011",
  47674=>"100110001",
  47675=>"101011110",
  47676=>"110000101",
  47677=>"000101101",
  47678=>"011001011",
  47679=>"011000010",
  47680=>"101100000",
  47681=>"011101010",
  47682=>"111110001",
  47683=>"111100000",
  47684=>"011101011",
  47685=>"010010110",
  47686=>"010101100",
  47687=>"101001110",
  47688=>"001000100",
  47689=>"101011101",
  47690=>"101110100",
  47691=>"100000011",
  47692=>"010100001",
  47693=>"110100110",
  47694=>"110001000",
  47695=>"100100101",
  47696=>"100101110",
  47697=>"000111010",
  47698=>"000101000",
  47699=>"000111001",
  47700=>"010010000",
  47701=>"100001111",
  47702=>"000110011",
  47703=>"001111111",
  47704=>"011110111",
  47705=>"000010010",
  47706=>"010011010",
  47707=>"100001100",
  47708=>"001111111",
  47709=>"111100010",
  47710=>"000010101",
  47711=>"010101010",
  47712=>"010011111",
  47713=>"110010011",
  47714=>"101001101",
  47715=>"000111111",
  47716=>"100001000",
  47717=>"110000101",
  47718=>"101000100",
  47719=>"111011010",
  47720=>"100101001",
  47721=>"000000001",
  47722=>"101011010",
  47723=>"011011010",
  47724=>"011101000",
  47725=>"001111011",
  47726=>"100000111",
  47727=>"111010010",
  47728=>"011001111",
  47729=>"000001001",
  47730=>"000010100",
  47731=>"011111001",
  47732=>"000011010",
  47733=>"100111111",
  47734=>"010110000",
  47735=>"011001000",
  47736=>"111111110",
  47737=>"011101011",
  47738=>"111011011",
  47739=>"000100011",
  47740=>"101100111",
  47741=>"011101111",
  47742=>"010011111",
  47743=>"011101100",
  47744=>"011100011",
  47745=>"001101100",
  47746=>"100101100",
  47747=>"100000001",
  47748=>"100000001",
  47749=>"100000001",
  47750=>"000100010",
  47751=>"111100011",
  47752=>"001001101",
  47753=>"010101100",
  47754=>"101010111",
  47755=>"110101001",
  47756=>"110111010",
  47757=>"010000010",
  47758=>"010110001",
  47759=>"011101001",
  47760=>"000010110",
  47761=>"000101000",
  47762=>"011111110",
  47763=>"010011100",
  47764=>"110100100",
  47765=>"101110110",
  47766=>"101111111",
  47767=>"011011010",
  47768=>"000110010",
  47769=>"111110011",
  47770=>"101010011",
  47771=>"000000000",
  47772=>"101101001",
  47773=>"000000010",
  47774=>"011011110",
  47775=>"000101110",
  47776=>"100011101",
  47777=>"100011100",
  47778=>"010101010",
  47779=>"101010100",
  47780=>"010111111",
  47781=>"001101101",
  47782=>"000001000",
  47783=>"010101111",
  47784=>"101010010",
  47785=>"100111000",
  47786=>"110000110",
  47787=>"010000100",
  47788=>"001000001",
  47789=>"100101001",
  47790=>"101010011",
  47791=>"010101010",
  47792=>"001110011",
  47793=>"100010001",
  47794=>"001010010",
  47795=>"000001001",
  47796=>"001001011",
  47797=>"011000011",
  47798=>"011010000",
  47799=>"101110010",
  47800=>"111100011",
  47801=>"111001010",
  47802=>"001101111",
  47803=>"110110000",
  47804=>"111001001",
  47805=>"101010100",
  47806=>"110000011",
  47807=>"000000010",
  47808=>"101111111",
  47809=>"110100100",
  47810=>"111111001",
  47811=>"101111000",
  47812=>"110001100",
  47813=>"010110110",
  47814=>"101011100",
  47815=>"001001111",
  47816=>"001000010",
  47817=>"010000100",
  47818=>"100101010",
  47819=>"000011000",
  47820=>"100001100",
  47821=>"101011001",
  47822=>"100111100",
  47823=>"001110101",
  47824=>"010010111",
  47825=>"111010110",
  47826=>"000000011",
  47827=>"010111100",
  47828=>"101111111",
  47829=>"011010000",
  47830=>"000011000",
  47831=>"111011010",
  47832=>"000101111",
  47833=>"011111100",
  47834=>"011001010",
  47835=>"111010111",
  47836=>"110100001",
  47837=>"010001110",
  47838=>"001001011",
  47839=>"010001110",
  47840=>"011111001",
  47841=>"110101100",
  47842=>"010110100",
  47843=>"100000101",
  47844=>"010000100",
  47845=>"111100111",
  47846=>"110010000",
  47847=>"100000000",
  47848=>"111010100",
  47849=>"010010010",
  47850=>"001000010",
  47851=>"101011100",
  47852=>"010000101",
  47853=>"100010001",
  47854=>"000101011",
  47855=>"100000111",
  47856=>"110111010",
  47857=>"101111100",
  47858=>"101100011",
  47859=>"100100111",
  47860=>"000011101",
  47861=>"101011110",
  47862=>"011010101",
  47863=>"110010100",
  47864=>"000000000",
  47865=>"101100111",
  47866=>"101000000",
  47867=>"111110010",
  47868=>"000011111",
  47869=>"000101100",
  47870=>"011110010",
  47871=>"110010101",
  47872=>"001101111",
  47873=>"000011000",
  47874=>"101110010",
  47875=>"000010100",
  47876=>"010001010",
  47877=>"010111110",
  47878=>"111110001",
  47879=>"011101010",
  47880=>"101101100",
  47881=>"001100000",
  47882=>"010000010",
  47883=>"110110001",
  47884=>"010000011",
  47885=>"100010010",
  47886=>"010110111",
  47887=>"100101110",
  47888=>"000010110",
  47889=>"000101001",
  47890=>"100011101",
  47891=>"101101111",
  47892=>"010011110",
  47893=>"001001111",
  47894=>"001110110",
  47895=>"010111001",
  47896=>"011010000",
  47897=>"001011111",
  47898=>"000001101",
  47899=>"100100001",
  47900=>"010001100",
  47901=>"101000110",
  47902=>"111001111",
  47903=>"100101111",
  47904=>"110100101",
  47905=>"001110011",
  47906=>"010100001",
  47907=>"111110001",
  47908=>"001101111",
  47909=>"111011111",
  47910=>"111101110",
  47911=>"110111011",
  47912=>"100010011",
  47913=>"000000100",
  47914=>"111110000",
  47915=>"110000110",
  47916=>"110101000",
  47917=>"111110001",
  47918=>"010110111",
  47919=>"010000100",
  47920=>"011010101",
  47921=>"000010011",
  47922=>"001011011",
  47923=>"100011001",
  47924=>"000101100",
  47925=>"001111100",
  47926=>"110100110",
  47927=>"110000011",
  47928=>"101100000",
  47929=>"101110101",
  47930=>"001110100",
  47931=>"100111110",
  47932=>"000100110",
  47933=>"010010100",
  47934=>"010111101",
  47935=>"011011101",
  47936=>"001111101",
  47937=>"000001011",
  47938=>"101001110",
  47939=>"001001010",
  47940=>"001011010",
  47941=>"111101110",
  47942=>"111101111",
  47943=>"000111110",
  47944=>"001101111",
  47945=>"000000101",
  47946=>"011111010",
  47947=>"100000110",
  47948=>"010010101",
  47949=>"001111100",
  47950=>"111011011",
  47951=>"100001011",
  47952=>"100100111",
  47953=>"100001000",
  47954=>"001101000",
  47955=>"001000011",
  47956=>"111010110",
  47957=>"101110010",
  47958=>"011000000",
  47959=>"000110110",
  47960=>"100010110",
  47961=>"100001110",
  47962=>"010010111",
  47963=>"111101101",
  47964=>"001011100",
  47965=>"000001001",
  47966=>"101101110",
  47967=>"000001110",
  47968=>"101001001",
  47969=>"010100011",
  47970=>"000011010",
  47971=>"010010001",
  47972=>"100100100",
  47973=>"010111010",
  47974=>"000010100",
  47975=>"000100101",
  47976=>"110011111",
  47977=>"101100001",
  47978=>"100101111",
  47979=>"011011000",
  47980=>"011101001",
  47981=>"010000100",
  47982=>"110000001",
  47983=>"110111111",
  47984=>"100011100",
  47985=>"000110000",
  47986=>"111000000",
  47987=>"010100111",
  47988=>"100000010",
  47989=>"100000110",
  47990=>"011100110",
  47991=>"010010010",
  47992=>"100000110",
  47993=>"100010110",
  47994=>"000111111",
  47995=>"010011110",
  47996=>"101100110",
  47997=>"111000011",
  47998=>"011110100",
  47999=>"110110001",
  48000=>"001000000",
  48001=>"000100011",
  48002=>"110001001",
  48003=>"110100010",
  48004=>"000111010",
  48005=>"011011010",
  48006=>"001110001",
  48007=>"110100010",
  48008=>"000001001",
  48009=>"111011101",
  48010=>"011101001",
  48011=>"110011011",
  48012=>"000111100",
  48013=>"001001111",
  48014=>"010111000",
  48015=>"110010110",
  48016=>"111001000",
  48017=>"101101101",
  48018=>"100110110",
  48019=>"101010010",
  48020=>"100011011",
  48021=>"100000000",
  48022=>"010011000",
  48023=>"100100110",
  48024=>"111110101",
  48025=>"000000100",
  48026=>"000111011",
  48027=>"000101100",
  48028=>"000101000",
  48029=>"100011101",
  48030=>"000001001",
  48031=>"110000010",
  48032=>"001111000",
  48033=>"111001100",
  48034=>"100100100",
  48035=>"110100110",
  48036=>"000110010",
  48037=>"100110110",
  48038=>"100001001",
  48039=>"110101000",
  48040=>"011000010",
  48041=>"111100010",
  48042=>"010110101",
  48043=>"011111101",
  48044=>"000011010",
  48045=>"101101100",
  48046=>"111010000",
  48047=>"110001111",
  48048=>"010010101",
  48049=>"101111001",
  48050=>"101000001",
  48051=>"100001001",
  48052=>"100010110",
  48053=>"001101100",
  48054=>"011101010",
  48055=>"101111101",
  48056=>"000010110",
  48057=>"110110010",
  48058=>"010010010",
  48059=>"110101011",
  48060=>"101110000",
  48061=>"011111100",
  48062=>"000001000",
  48063=>"001101010",
  48064=>"101110000",
  48065=>"010000100",
  48066=>"011000011",
  48067=>"101011110",
  48068=>"010100010",
  48069=>"001110010",
  48070=>"000111001",
  48071=>"010000010",
  48072=>"001000000",
  48073=>"001110010",
  48074=>"101001101",
  48075=>"110011100",
  48076=>"011111111",
  48077=>"001101111",
  48078=>"001010100",
  48079=>"011100011",
  48080=>"000111110",
  48081=>"001110100",
  48082=>"010000110",
  48083=>"100100011",
  48084=>"111101110",
  48085=>"010011011",
  48086=>"011110000",
  48087=>"110110000",
  48088=>"000000111",
  48089=>"010000010",
  48090=>"011110000",
  48091=>"010110011",
  48092=>"001111001",
  48093=>"100110000",
  48094=>"100011001",
  48095=>"000100100",
  48096=>"111011111",
  48097=>"101110011",
  48098=>"000001000",
  48099=>"110011011",
  48100=>"101011111",
  48101=>"000101000",
  48102=>"100100101",
  48103=>"111011011",
  48104=>"010000001",
  48105=>"101010101",
  48106=>"000001110",
  48107=>"010000000",
  48108=>"111001110",
  48109=>"100011100",
  48110=>"001111011",
  48111=>"110000101",
  48112=>"000101011",
  48113=>"000000101",
  48114=>"011010011",
  48115=>"110001110",
  48116=>"111110110",
  48117=>"001111110",
  48118=>"110111111",
  48119=>"100000111",
  48120=>"001000000",
  48121=>"000010001",
  48122=>"100001101",
  48123=>"101100111",
  48124=>"100101111",
  48125=>"110011101",
  48126=>"000001101",
  48127=>"111001100",
  48128=>"000010000",
  48129=>"110110000",
  48130=>"010010110",
  48131=>"101101010",
  48132=>"101100110",
  48133=>"010000110",
  48134=>"000011111",
  48135=>"111011111",
  48136=>"101101000",
  48137=>"001000100",
  48138=>"001000100",
  48139=>"110101001",
  48140=>"000000011",
  48141=>"101111011",
  48142=>"110101000",
  48143=>"111110100",
  48144=>"000011010",
  48145=>"011000001",
  48146=>"001000010",
  48147=>"000110110",
  48148=>"000000001",
  48149=>"111010011",
  48150=>"110101010",
  48151=>"000110000",
  48152=>"011000111",
  48153=>"011111111",
  48154=>"110001011",
  48155=>"000001101",
  48156=>"001000100",
  48157=>"111010011",
  48158=>"101111110",
  48159=>"011000100",
  48160=>"001010100",
  48161=>"000001011",
  48162=>"111000010",
  48163=>"001011110",
  48164=>"010101100",
  48165=>"101001110",
  48166=>"111000101",
  48167=>"010101011",
  48168=>"010001001",
  48169=>"100110111",
  48170=>"111001111",
  48171=>"001100100",
  48172=>"000000001",
  48173=>"111001111",
  48174=>"101101010",
  48175=>"111001100",
  48176=>"110000001",
  48177=>"110011000",
  48178=>"011001111",
  48179=>"101110000",
  48180=>"000110001",
  48181=>"000001000",
  48182=>"101111111",
  48183=>"101101000",
  48184=>"111111101",
  48185=>"100100110",
  48186=>"000110010",
  48187=>"111100000",
  48188=>"110001101",
  48189=>"011111001",
  48190=>"110111010",
  48191=>"010001110",
  48192=>"011011011",
  48193=>"010111001",
  48194=>"110101001",
  48195=>"001000110",
  48196=>"110000111",
  48197=>"100001000",
  48198=>"000001010",
  48199=>"001101101",
  48200=>"001110010",
  48201=>"100111000",
  48202=>"001010010",
  48203=>"101101100",
  48204=>"000101000",
  48205=>"010010110",
  48206=>"011010011",
  48207=>"000100101",
  48208=>"111110101",
  48209=>"001001010",
  48210=>"000001011",
  48211=>"011000100",
  48212=>"110110101",
  48213=>"101011100",
  48214=>"001011001",
  48215=>"011110011",
  48216=>"110010000",
  48217=>"100101111",
  48218=>"111011110",
  48219=>"001011001",
  48220=>"000100101",
  48221=>"111010110",
  48222=>"000110111",
  48223=>"010100110",
  48224=>"110000001",
  48225=>"001100100",
  48226=>"111111001",
  48227=>"101100011",
  48228=>"111100000",
  48229=>"011010011",
  48230=>"110101101",
  48231=>"001110111",
  48232=>"111010000",
  48233=>"110010111",
  48234=>"001001111",
  48235=>"010000110",
  48236=>"110100001",
  48237=>"010111000",
  48238=>"010001101",
  48239=>"101110110",
  48240=>"000110000",
  48241=>"100100100",
  48242=>"011000111",
  48243=>"010011000",
  48244=>"111010110",
  48245=>"111001011",
  48246=>"011010000",
  48247=>"010100111",
  48248=>"111111111",
  48249=>"001000000",
  48250=>"110001010",
  48251=>"101101001",
  48252=>"010001110",
  48253=>"011111101",
  48254=>"111000010",
  48255=>"100111000",
  48256=>"101010100",
  48257=>"010011110",
  48258=>"110111100",
  48259=>"101100101",
  48260=>"000001100",
  48261=>"100011001",
  48262=>"101100000",
  48263=>"111011001",
  48264=>"010111010",
  48265=>"111010110",
  48266=>"100010011",
  48267=>"100111111",
  48268=>"010000010",
  48269=>"111111000",
  48270=>"001001010",
  48271=>"001101010",
  48272=>"100111000",
  48273=>"011111111",
  48274=>"110111110",
  48275=>"010100101",
  48276=>"110010111",
  48277=>"001011111",
  48278=>"011000100",
  48279=>"100110100",
  48280=>"101111101",
  48281=>"111001110",
  48282=>"010000110",
  48283=>"111001101",
  48284=>"001001011",
  48285=>"111100010",
  48286=>"110101010",
  48287=>"101011000",
  48288=>"110110000",
  48289=>"111100011",
  48290=>"100001110",
  48291=>"001101110",
  48292=>"111000001",
  48293=>"000001101",
  48294=>"010001001",
  48295=>"100100101",
  48296=>"101011111",
  48297=>"011011001",
  48298=>"000001101",
  48299=>"111001111",
  48300=>"101111110",
  48301=>"010001001",
  48302=>"111011000",
  48303=>"001011100",
  48304=>"000110010",
  48305=>"001100100",
  48306=>"010010000",
  48307=>"001111110",
  48308=>"111010110",
  48309=>"011001000",
  48310=>"111110011",
  48311=>"101000000",
  48312=>"000001010",
  48313=>"101010100",
  48314=>"111001110",
  48315=>"011111101",
  48316=>"101101000",
  48317=>"111111100",
  48318=>"101101001",
  48319=>"110110000",
  48320=>"111100000",
  48321=>"001111100",
  48322=>"110000001",
  48323=>"000000101",
  48324=>"011111000",
  48325=>"000011110",
  48326=>"100111011",
  48327=>"001110101",
  48328=>"010101100",
  48329=>"110010101",
  48330=>"010111001",
  48331=>"100010100",
  48332=>"001100100",
  48333=>"010011011",
  48334=>"010111000",
  48335=>"011001101",
  48336=>"101101000",
  48337=>"111101000",
  48338=>"000100011",
  48339=>"011100110",
  48340=>"011111011",
  48341=>"010110111",
  48342=>"011111110",
  48343=>"101011011",
  48344=>"011110001",
  48345=>"000000100",
  48346=>"110110101",
  48347=>"001000101",
  48348=>"111111011",
  48349=>"011101001",
  48350=>"111100000",
  48351=>"011100011",
  48352=>"011101100",
  48353=>"110011001",
  48354=>"000000001",
  48355=>"111111110",
  48356=>"010011101",
  48357=>"001000111",
  48358=>"100110000",
  48359=>"111101000",
  48360=>"001111111",
  48361=>"111101101",
  48362=>"000000100",
  48363=>"001011100",
  48364=>"000011110",
  48365=>"110011110",
  48366=>"110001100",
  48367=>"101001111",
  48368=>"110100111",
  48369=>"101000100",
  48370=>"100001100",
  48371=>"111011101",
  48372=>"100111111",
  48373=>"010000100",
  48374=>"101111100",
  48375=>"000010110",
  48376=>"101000101",
  48377=>"101010111",
  48378=>"000010101",
  48379=>"010011001",
  48380=>"110000001",
  48381=>"000011001",
  48382=>"011000100",
  48383=>"011000000",
  48384=>"011010111",
  48385=>"111001001",
  48386=>"111000101",
  48387=>"100011010",
  48388=>"010001010",
  48389=>"010110110",
  48390=>"110010110",
  48391=>"110001001",
  48392=>"010010110",
  48393=>"100011010",
  48394=>"101101000",
  48395=>"101000101",
  48396=>"010011110",
  48397=>"000111111",
  48398=>"011000010",
  48399=>"000011100",
  48400=>"010100110",
  48401=>"100011001",
  48402=>"000010011",
  48403=>"100010000",
  48404=>"100111110",
  48405=>"100101110",
  48406=>"100100000",
  48407=>"111101001",
  48408=>"001101001",
  48409=>"100101111",
  48410=>"100110101",
  48411=>"011001100",
  48412=>"101011010",
  48413=>"010000111",
  48414=>"100011110",
  48415=>"110101000",
  48416=>"110001000",
  48417=>"110011110",
  48418=>"000001101",
  48419=>"110000111",
  48420=>"001111111",
  48421=>"010001111",
  48422=>"010011100",
  48423=>"011100110",
  48424=>"001100111",
  48425=>"000000010",
  48426=>"000100000",
  48427=>"111101110",
  48428=>"011111100",
  48429=>"101110001",
  48430=>"001001001",
  48431=>"011010110",
  48432=>"100110100",
  48433=>"011010100",
  48434=>"101001101",
  48435=>"100110010",
  48436=>"111010110",
  48437=>"110010011",
  48438=>"001000000",
  48439=>"001001000",
  48440=>"101000000",
  48441=>"101000000",
  48442=>"000111101",
  48443=>"000100111",
  48444=>"111000100",
  48445=>"110101010",
  48446=>"100001100",
  48447=>"101010011",
  48448=>"110110010",
  48449=>"111101011",
  48450=>"000001111",
  48451=>"001100001",
  48452=>"001010011",
  48453=>"110101100",
  48454=>"101011110",
  48455=>"010001111",
  48456=>"110000010",
  48457=>"111110111",
  48458=>"110111001",
  48459=>"110011110",
  48460=>"110010011",
  48461=>"111100001",
  48462=>"001000011",
  48463=>"000000101",
  48464=>"111010101",
  48465=>"101110011",
  48466=>"100101001",
  48467=>"010000111",
  48468=>"011101011",
  48469=>"100000111",
  48470=>"010000001",
  48471=>"000111110",
  48472=>"000110010",
  48473=>"100100111",
  48474=>"011100111",
  48475=>"100010010",
  48476=>"100010100",
  48477=>"011111111",
  48478=>"110011111",
  48479=>"001001000",
  48480=>"101101010",
  48481=>"101101100",
  48482=>"101101000",
  48483=>"000011010",
  48484=>"110111101",
  48485=>"000010000",
  48486=>"011001101",
  48487=>"101110010",
  48488=>"000010000",
  48489=>"001110000",
  48490=>"011100000",
  48491=>"101110000",
  48492=>"100000011",
  48493=>"101001100",
  48494=>"111101101",
  48495=>"001101101",
  48496=>"000001101",
  48497=>"111111011",
  48498=>"001101110",
  48499=>"111100000",
  48500=>"100010000",
  48501=>"111010101",
  48502=>"101011111",
  48503=>"100110011",
  48504=>"110111011",
  48505=>"110111011",
  48506=>"000000010",
  48507=>"001011010",
  48508=>"011111000",
  48509=>"000000110",
  48510=>"010000000",
  48511=>"111111111",
  48512=>"011010100",
  48513=>"001111111",
  48514=>"010111100",
  48515=>"010001000",
  48516=>"010011001",
  48517=>"101111100",
  48518=>"101001000",
  48519=>"000111001",
  48520=>"100100101",
  48521=>"000110111",
  48522=>"001000001",
  48523=>"000110001",
  48524=>"010000111",
  48525=>"001100000",
  48526=>"110100100",
  48527=>"000000110",
  48528=>"101100101",
  48529=>"110110000",
  48530=>"000001100",
  48531=>"011000010",
  48532=>"000111010",
  48533=>"011101010",
  48534=>"110111100",
  48535=>"101110000",
  48536=>"000101000",
  48537=>"100000000",
  48538=>"010001101",
  48539=>"010110001",
  48540=>"000101101",
  48541=>"111110010",
  48542=>"111100111",
  48543=>"000111000",
  48544=>"101010010",
  48545=>"010001110",
  48546=>"011101000",
  48547=>"111001111",
  48548=>"111001010",
  48549=>"001001101",
  48550=>"110101000",
  48551=>"001001100",
  48552=>"001000001",
  48553=>"111100101",
  48554=>"100011111",
  48555=>"111001110",
  48556=>"011110100",
  48557=>"000100000",
  48558=>"000111101",
  48559=>"111101100",
  48560=>"111011011",
  48561=>"010000010",
  48562=>"010100000",
  48563=>"100000010",
  48564=>"001000011",
  48565=>"011110110",
  48566=>"001100101",
  48567=>"011000101",
  48568=>"110111111",
  48569=>"010011111",
  48570=>"101111111",
  48571=>"010101001",
  48572=>"001101111",
  48573=>"000010001",
  48574=>"100111110",
  48575=>"010011010",
  48576=>"000101110",
  48577=>"011110001",
  48578=>"011101111",
  48579=>"010111110",
  48580=>"000100001",
  48581=>"110001000",
  48582=>"101010110",
  48583=>"111100111",
  48584=>"100111100",
  48585=>"111110101",
  48586=>"010100000",
  48587=>"000000010",
  48588=>"111011100",
  48589=>"100100111",
  48590=>"011001000",
  48591=>"001101100",
  48592=>"111111000",
  48593=>"101001001",
  48594=>"000000001",
  48595=>"100010111",
  48596=>"010000010",
  48597=>"111111101",
  48598=>"111001111",
  48599=>"001011110",
  48600=>"110011000",
  48601=>"111111110",
  48602=>"100011011",
  48603=>"101101000",
  48604=>"101101011",
  48605=>"111111000",
  48606=>"000100100",
  48607=>"001110000",
  48608=>"010101001",
  48609=>"111110100",
  48610=>"000111000",
  48611=>"101001001",
  48612=>"000111110",
  48613=>"101001100",
  48614=>"000111110",
  48615=>"010001011",
  48616=>"110010011",
  48617=>"011010110",
  48618=>"101111011",
  48619=>"001101110",
  48620=>"110111001",
  48621=>"101100001",
  48622=>"011010100",
  48623=>"100101011",
  48624=>"000011100",
  48625=>"010111110",
  48626=>"011101100",
  48627=>"100101010",
  48628=>"001000000",
  48629=>"000001000",
  48630=>"010111001",
  48631=>"100000100",
  48632=>"011111100",
  48633=>"000001111",
  48634=>"001011010",
  48635=>"011010101",
  48636=>"000010111",
  48637=>"100000100",
  48638=>"010111010",
  48639=>"000011101",
  48640=>"110010110",
  48641=>"001000101",
  48642=>"111110000",
  48643=>"011010011",
  48644=>"010000010",
  48645=>"000001001",
  48646=>"111111011",
  48647=>"100000110",
  48648=>"101100011",
  48649=>"110111101",
  48650=>"111101001",
  48651=>"101111110",
  48652=>"101101100",
  48653=>"101010100",
  48654=>"001001001",
  48655=>"011011001",
  48656=>"011111000",
  48657=>"010100110",
  48658=>"110010000",
  48659=>"111110000",
  48660=>"100110000",
  48661=>"001100010",
  48662=>"011110001",
  48663=>"101000001",
  48664=>"011011011",
  48665=>"110000111",
  48666=>"100101101",
  48667=>"111010000",
  48668=>"011000101",
  48669=>"101100110",
  48670=>"001010101",
  48671=>"000101000",
  48672=>"111111010",
  48673=>"001110010",
  48674=>"010011110",
  48675=>"000100000",
  48676=>"011000011",
  48677=>"010101011",
  48678=>"101011111",
  48679=>"000110100",
  48680=>"111101000",
  48681=>"001101001",
  48682=>"110100111",
  48683=>"100100111",
  48684=>"111110010",
  48685=>"101001011",
  48686=>"000001001",
  48687=>"001101100",
  48688=>"110001100",
  48689=>"101001101",
  48690=>"100000010",
  48691=>"101000000",
  48692=>"000011011",
  48693=>"110101111",
  48694=>"000111101",
  48695=>"111010001",
  48696=>"001001011",
  48697=>"111001000",
  48698=>"010101111",
  48699=>"011101101",
  48700=>"010000100",
  48701=>"010110011",
  48702=>"010110110",
  48703=>"011110000",
  48704=>"010000110",
  48705=>"111111110",
  48706=>"110111011",
  48707=>"001100010",
  48708=>"010110001",
  48709=>"111000100",
  48710=>"010100010",
  48711=>"010100111",
  48712=>"111111101",
  48713=>"110011011",
  48714=>"101000110",
  48715=>"101101101",
  48716=>"001001011",
  48717=>"000111011",
  48718=>"001110111",
  48719=>"101110011",
  48720=>"011111110",
  48721=>"101110010",
  48722=>"001001100",
  48723=>"000000110",
  48724=>"011101010",
  48725=>"011000011",
  48726=>"110010000",
  48727=>"010101110",
  48728=>"011111110",
  48729=>"011110100",
  48730=>"010100110",
  48731=>"001011010",
  48732=>"100010100",
  48733=>"000001010",
  48734=>"000101101",
  48735=>"110101010",
  48736=>"000011001",
  48737=>"011111111",
  48738=>"101110001",
  48739=>"110111011",
  48740=>"111110010",
  48741=>"101101010",
  48742=>"101010000",
  48743=>"110001010",
  48744=>"101100000",
  48745=>"011100010",
  48746=>"101001000",
  48747=>"110100101",
  48748=>"111111001",
  48749=>"101001001",
  48750=>"000111111",
  48751=>"011100100",
  48752=>"111111010",
  48753=>"100100100",
  48754=>"000001001",
  48755=>"100101101",
  48756=>"101111101",
  48757=>"000000110",
  48758=>"011001000",
  48759=>"110111000",
  48760=>"101100111",
  48761=>"100011100",
  48762=>"101100011",
  48763=>"110010011",
  48764=>"000101111",
  48765=>"110001101",
  48766=>"101101100",
  48767=>"100011101",
  48768=>"100001100",
  48769=>"010010001",
  48770=>"101000110",
  48771=>"101011010",
  48772=>"000110100",
  48773=>"000000100",
  48774=>"001000111",
  48775=>"111100111",
  48776=>"101110010",
  48777=>"111011000",
  48778=>"110011010",
  48779=>"000110111",
  48780=>"110000011",
  48781=>"010100111",
  48782=>"111111011",
  48783=>"010110111",
  48784=>"000000111",
  48785=>"000010101",
  48786=>"111000111",
  48787=>"101110000",
  48788=>"110101011",
  48789=>"000011001",
  48790=>"011010000",
  48791=>"011010111",
  48792=>"010111011",
  48793=>"111101100",
  48794=>"001001111",
  48795=>"000010111",
  48796=>"111110111",
  48797=>"001100000",
  48798=>"000110110",
  48799=>"011100011",
  48800=>"100000111",
  48801=>"101000001",
  48802=>"111001101",
  48803=>"011101000",
  48804=>"000110101",
  48805=>"101101101",
  48806=>"010000111",
  48807=>"111001001",
  48808=>"111010100",
  48809=>"001001011",
  48810=>"101101101",
  48811=>"101011001",
  48812=>"010100111",
  48813=>"000101111",
  48814=>"010101111",
  48815=>"111001001",
  48816=>"011101000",
  48817=>"101100101",
  48818=>"100010011",
  48819=>"111101111",
  48820=>"000011010",
  48821=>"111000111",
  48822=>"111110100",
  48823=>"110100110",
  48824=>"110110110",
  48825=>"110111011",
  48826=>"001101101",
  48827=>"110000101",
  48828=>"101010001",
  48829=>"011111001",
  48830=>"100101100",
  48831=>"111111011",
  48832=>"110001011",
  48833=>"110110100",
  48834=>"111010011",
  48835=>"110111001",
  48836=>"000110111",
  48837=>"011111011",
  48838=>"110110011",
  48839=>"101101111",
  48840=>"111100110",
  48841=>"001011011",
  48842=>"110010001",
  48843=>"001000111",
  48844=>"001011011",
  48845=>"101111000",
  48846=>"111011101",
  48847=>"111001001",
  48848=>"000001101",
  48849=>"101010100",
  48850=>"000010100",
  48851=>"101110110",
  48852=>"111011011",
  48853=>"111001100",
  48854=>"100001000",
  48855=>"110000000",
  48856=>"010001101",
  48857=>"110111010",
  48858=>"100000101",
  48859=>"110011001",
  48860=>"101011010",
  48861=>"100001001",
  48862=>"011111110",
  48863=>"100000001",
  48864=>"110011100",
  48865=>"111111010",
  48866=>"110000000",
  48867=>"111110100",
  48868=>"100100011",
  48869=>"101000011",
  48870=>"111111110",
  48871=>"011001110",
  48872=>"100111001",
  48873=>"100010010",
  48874=>"111010110",
  48875=>"111101111",
  48876=>"011000100",
  48877=>"100101001",
  48878=>"110101111",
  48879=>"110100001",
  48880=>"101110010",
  48881=>"101010101",
  48882=>"101011101",
  48883=>"000101111",
  48884=>"101001000",
  48885=>"111001111",
  48886=>"011110010",
  48887=>"000000100",
  48888=>"001010000",
  48889=>"101010000",
  48890=>"011001101",
  48891=>"000000010",
  48892=>"011111100",
  48893=>"001001011",
  48894=>"110110101",
  48895=>"000110010",
  48896=>"010010001",
  48897=>"100111001",
  48898=>"111000110",
  48899=>"110111001",
  48900=>"011010110",
  48901=>"110100000",
  48902=>"111011011",
  48903=>"110011001",
  48904=>"000011111",
  48905=>"111010110",
  48906=>"111000011",
  48907=>"111001001",
  48908=>"010000101",
  48909=>"101100010",
  48910=>"001011010",
  48911=>"000101001",
  48912=>"001010101",
  48913=>"100100101",
  48914=>"111111011",
  48915=>"010000000",
  48916=>"110110010",
  48917=>"011000001",
  48918=>"100100111",
  48919=>"001011111",
  48920=>"110111100",
  48921=>"000001110",
  48922=>"010100101",
  48923=>"111000000",
  48924=>"010001111",
  48925=>"101011001",
  48926=>"101111010",
  48927=>"001001111",
  48928=>"110001000",
  48929=>"011111110",
  48930=>"111101111",
  48931=>"011000110",
  48932=>"000000001",
  48933=>"110010101",
  48934=>"000100110",
  48935=>"100011001",
  48936=>"001001100",
  48937=>"101100101",
  48938=>"110011110",
  48939=>"100101111",
  48940=>"100100110",
  48941=>"111110110",
  48942=>"000100010",
  48943=>"111100100",
  48944=>"010011110",
  48945=>"100010111",
  48946=>"010011000",
  48947=>"010111101",
  48948=>"110111101",
  48949=>"010111001",
  48950=>"000010001",
  48951=>"000010001",
  48952=>"101101100",
  48953=>"101000101",
  48954=>"101111010",
  48955=>"001110100",
  48956=>"111001011",
  48957=>"000100100",
  48958=>"101001101",
  48959=>"100001101",
  48960=>"111011011",
  48961=>"100111111",
  48962=>"110010111",
  48963=>"010001111",
  48964=>"010000000",
  48965=>"110101010",
  48966=>"001110001",
  48967=>"100011010",
  48968=>"101001000",
  48969=>"010110010",
  48970=>"011011000",
  48971=>"010101000",
  48972=>"001110101",
  48973=>"001110010",
  48974=>"100001100",
  48975=>"010010011",
  48976=>"101000111",
  48977=>"111011000",
  48978=>"010011101",
  48979=>"100110101",
  48980=>"110110110",
  48981=>"000001001",
  48982=>"000101111",
  48983=>"011111110",
  48984=>"011001101",
  48985=>"100001001",
  48986=>"011010101",
  48987=>"000010101",
  48988=>"101101110",
  48989=>"000001111",
  48990=>"010011110",
  48991=>"011110001",
  48992=>"110100001",
  48993=>"001110001",
  48994=>"111011011",
  48995=>"000111010",
  48996=>"011010011",
  48997=>"010000110",
  48998=>"011011011",
  48999=>"001011101",
  49000=>"000010011",
  49001=>"101010011",
  49002=>"101100000",
  49003=>"000101010",
  49004=>"011010101",
  49005=>"011111100",
  49006=>"101010011",
  49007=>"010001001",
  49008=>"010010011",
  49009=>"001000110",
  49010=>"011110100",
  49011=>"101111101",
  49012=>"000101010",
  49013=>"111110011",
  49014=>"110010101",
  49015=>"100001100",
  49016=>"110101101",
  49017=>"001010000",
  49018=>"011011110",
  49019=>"010001001",
  49020=>"011010100",
  49021=>"110110001",
  49022=>"011010011",
  49023=>"001010111",
  49024=>"010000110",
  49025=>"100101100",
  49026=>"110011110",
  49027=>"010111101",
  49028=>"001101111",
  49029=>"000101000",
  49030=>"100100001",
  49031=>"101101001",
  49032=>"011111101",
  49033=>"101001000",
  49034=>"000100111",
  49035=>"101001110",
  49036=>"111110011",
  49037=>"101110000",
  49038=>"000010011",
  49039=>"101101010",
  49040=>"011000000",
  49041=>"000111000",
  49042=>"000010111",
  49043=>"101110011",
  49044=>"110101001",
  49045=>"111001011",
  49046=>"011000111",
  49047=>"111110101",
  49048=>"010101000",
  49049=>"101010100",
  49050=>"101111101",
  49051=>"011000001",
  49052=>"001010100",
  49053=>"010111110",
  49054=>"000100110",
  49055=>"000101101",
  49056=>"101101111",
  49057=>"100101000",
  49058=>"111110000",
  49059=>"111101101",
  49060=>"010000101",
  49061=>"011011010",
  49062=>"000100101",
  49063=>"000101101",
  49064=>"010111001",
  49065=>"000110101",
  49066=>"100000100",
  49067=>"000001111",
  49068=>"000101010",
  49069=>"011101010",
  49070=>"010010000",
  49071=>"000101001",
  49072=>"111010111",
  49073=>"101110010",
  49074=>"011011010",
  49075=>"111101111",
  49076=>"111001000",
  49077=>"101111111",
  49078=>"000100101",
  49079=>"001010111",
  49080=>"101111111",
  49081=>"000011101",
  49082=>"100100001",
  49083=>"101001101",
  49084=>"110100100",
  49085=>"010111000",
  49086=>"011111011",
  49087=>"010110000",
  49088=>"010110011",
  49089=>"010000111",
  49090=>"101001000",
  49091=>"101111111",
  49092=>"010100010",
  49093=>"110010101",
  49094=>"111101101",
  49095=>"011111000",
  49096=>"001010000",
  49097=>"100000001",
  49098=>"111000011",
  49099=>"001000010",
  49100=>"011000111",
  49101=>"110011100",
  49102=>"000100111",
  49103=>"010101010",
  49104=>"010010011",
  49105=>"111100111",
  49106=>"010000001",
  49107=>"011000001",
  49108=>"011001011",
  49109=>"000000000",
  49110=>"001111011",
  49111=>"101110001",
  49112=>"111100001",
  49113=>"110110110",
  49114=>"011110001",
  49115=>"000101111",
  49116=>"101111101",
  49117=>"010010001",
  49118=>"011010011",
  49119=>"101101110",
  49120=>"110000110",
  49121=>"110000000",
  49122=>"110001111",
  49123=>"110111011",
  49124=>"010000110",
  49125=>"011110000",
  49126=>"101011000",
  49127=>"010101001",
  49128=>"001000000",
  49129=>"111101110",
  49130=>"111110110",
  49131=>"000000000",
  49132=>"000111111",
  49133=>"000010010",
  49134=>"110000010",
  49135=>"110101011",
  49136=>"100101001",
  49137=>"100101110",
  49138=>"101101000",
  49139=>"001111011",
  49140=>"111001110",
  49141=>"111110100",
  49142=>"000000010",
  49143=>"011111101",
  49144=>"000010011",
  49145=>"001010000",
  49146=>"010011000",
  49147=>"100110011",
  49148=>"011001111",
  49149=>"000100111",
  49150=>"010000011",
  49151=>"100100001",
  49152=>"000100110",
  49153=>"010011011",
  49154=>"100010111",
  49155=>"011110111",
  49156=>"000110011",
  49157=>"001111000",
  49158=>"100000010",
  49159=>"011000100",
  49160=>"100100110",
  49161=>"101111111",
  49162=>"101100111",
  49163=>"100001001",
  49164=>"111001101",
  49165=>"000110011",
  49166=>"100001100",
  49167=>"111000000",
  49168=>"011111011",
  49169=>"000011101",
  49170=>"111101001",
  49171=>"111101111",
  49172=>"010000100",
  49173=>"110010000",
  49174=>"111011001",
  49175=>"111110100",
  49176=>"010010111",
  49177=>"011101001",
  49178=>"110010101",
  49179=>"001101010",
  49180=>"100111010",
  49181=>"011010100",
  49182=>"010000001",
  49183=>"010110100",
  49184=>"001010000",
  49185=>"100111010",
  49186=>"111111101",
  49187=>"000010100",
  49188=>"100011010",
  49189=>"011111010",
  49190=>"110110101",
  49191=>"110010100",
  49192=>"011011001",
  49193=>"101101100",
  49194=>"010010110",
  49195=>"100011111",
  49196=>"000001100",
  49197=>"110101011",
  49198=>"000101101",
  49199=>"111000101",
  49200=>"000110111",
  49201=>"110000001",
  49202=>"001011010",
  49203=>"110111000",
  49204=>"001111000",
  49205=>"111011000",
  49206=>"000001010",
  49207=>"011111101",
  49208=>"000101000",
  49209=>"111111111",
  49210=>"000101111",
  49211=>"100110101",
  49212=>"100001111",
  49213=>"011001110",
  49214=>"010000010",
  49215=>"110001011",
  49216=>"001110110",
  49217=>"000011110",
  49218=>"000011101",
  49219=>"101110011",
  49220=>"011011101",
  49221=>"000001110",
  49222=>"011100100",
  49223=>"100011100",
  49224=>"011000111",
  49225=>"001111110",
  49226=>"101001000",
  49227=>"101011011",
  49228=>"010001100",
  49229=>"011100000",
  49230=>"111001111",
  49231=>"011000101",
  49232=>"101000110",
  49233=>"111011111",
  49234=>"011000101",
  49235=>"010010110",
  49236=>"110000001",
  49237=>"101101011",
  49238=>"110011000",
  49239=>"101001001",
  49240=>"110101110",
  49241=>"010000001",
  49242=>"010000010",
  49243=>"110111000",
  49244=>"111000110",
  49245=>"100100011",
  49246=>"100010111",
  49247=>"010001110",
  49248=>"101101010",
  49249=>"000100110",
  49250=>"101100101",
  49251=>"001001011",
  49252=>"010101110",
  49253=>"011001110",
  49254=>"111011101",
  49255=>"111110001",
  49256=>"100001100",
  49257=>"100011101",
  49258=>"110100111",
  49259=>"111011010",
  49260=>"011111001",
  49261=>"111011100",
  49262=>"100001001",
  49263=>"010001111",
  49264=>"101010000",
  49265=>"010111101",
  49266=>"100101100",
  49267=>"001010001",
  49268=>"110100111",
  49269=>"111010000",
  49270=>"001011101",
  49271=>"000000111",
  49272=>"111100111",
  49273=>"100011100",
  49274=>"000011101",
  49275=>"110100000",
  49276=>"011010011",
  49277=>"110111000",
  49278=>"010011000",
  49279=>"101100110",
  49280=>"100100010",
  49281=>"000100111",
  49282=>"110110011",
  49283=>"101001000",
  49284=>"100001101",
  49285=>"100100101",
  49286=>"000100000",
  49287=>"110100011",
  49288=>"101101011",
  49289=>"010011010",
  49290=>"001000111",
  49291=>"111011011",
  49292=>"011001101",
  49293=>"100110101",
  49294=>"011110100",
  49295=>"011101011",
  49296=>"111000101",
  49297=>"011111010",
  49298=>"100100101",
  49299=>"111000010",
  49300=>"100001001",
  49301=>"000000001",
  49302=>"011000111",
  49303=>"100010001",
  49304=>"010111001",
  49305=>"111011100",
  49306=>"001100000",
  49307=>"110110110",
  49308=>"111000010",
  49309=>"110111001",
  49310=>"110001101",
  49311=>"100010111",
  49312=>"000011000",
  49313=>"000001000",
  49314=>"110011100",
  49315=>"000100001",
  49316=>"110001101",
  49317=>"010111011",
  49318=>"111001110",
  49319=>"110110100",
  49320=>"000110111",
  49321=>"111011001",
  49322=>"111111111",
  49323=>"010111000",
  49324=>"111110100",
  49325=>"010001111",
  49326=>"110101101",
  49327=>"000011110",
  49328=>"101001011",
  49329=>"000100100",
  49330=>"100011111",
  49331=>"100000100",
  49332=>"010001101",
  49333=>"111010010",
  49334=>"111000001",
  49335=>"010001000",
  49336=>"000100101",
  49337=>"001001011",
  49338=>"101010011",
  49339=>"111001001",
  49340=>"000101010",
  49341=>"111000101",
  49342=>"001101000",
  49343=>"111111111",
  49344=>"101100001",
  49345=>"111001101",
  49346=>"101001111",
  49347=>"010001111",
  49348=>"101011011",
  49349=>"011010010",
  49350=>"111001101",
  49351=>"000100100",
  49352=>"111011010",
  49353=>"010101011",
  49354=>"000100000",
  49355=>"100110101",
  49356=>"001010100",
  49357=>"011010101",
  49358=>"011101000",
  49359=>"001101011",
  49360=>"111101100",
  49361=>"011100011",
  49362=>"110110010",
  49363=>"000111001",
  49364=>"000100000",
  49365=>"111111011",
  49366=>"110011010",
  49367=>"000001110",
  49368=>"100110100",
  49369=>"110000100",
  49370=>"010000011",
  49371=>"100011010",
  49372=>"110001110",
  49373=>"000010100",
  49374=>"101000001",
  49375=>"101111000",
  49376=>"111010100",
  49377=>"111011101",
  49378=>"100110110",
  49379=>"010010010",
  49380=>"011001101",
  49381=>"001001001",
  49382=>"111001101",
  49383=>"011110010",
  49384=>"111011010",
  49385=>"001000110",
  49386=>"001010111",
  49387=>"101000100",
  49388=>"110111010",
  49389=>"111000101",
  49390=>"010101111",
  49391=>"001100110",
  49392=>"101010010",
  49393=>"011111010",
  49394=>"001110000",
  49395=>"100110100",
  49396=>"001110000",
  49397=>"001100111",
  49398=>"110100100",
  49399=>"101011101",
  49400=>"000001011",
  49401=>"010001111",
  49402=>"111111010",
  49403=>"101111000",
  49404=>"010101001",
  49405=>"111110111",
  49406=>"011100001",
  49407=>"100001010",
  49408=>"100010011",
  49409=>"101010000",
  49410=>"001001000",
  49411=>"001000111",
  49412=>"110100001",
  49413=>"001100111",
  49414=>"010010010",
  49415=>"001001110",
  49416=>"000110101",
  49417=>"000001000",
  49418=>"010000001",
  49419=>"101001011",
  49420=>"110110101",
  49421=>"100000010",
  49422=>"110100000",
  49423=>"010010000",
  49424=>"101101100",
  49425=>"011000001",
  49426=>"010100101",
  49427=>"000001110",
  49428=>"110111100",
  49429=>"011010011",
  49430=>"101101010",
  49431=>"011001111",
  49432=>"001010000",
  49433=>"000110001",
  49434=>"011010101",
  49435=>"010101101",
  49436=>"010001111",
  49437=>"000000100",
  49438=>"100111100",
  49439=>"010010100",
  49440=>"110010101",
  49441=>"110100011",
  49442=>"000010000",
  49443=>"001110010",
  49444=>"000100111",
  49445=>"001000001",
  49446=>"110100001",
  49447=>"001010000",
  49448=>"100011111",
  49449=>"100110011",
  49450=>"011000010",
  49451=>"000110001",
  49452=>"100111110",
  49453=>"111101100",
  49454=>"101000111",
  49455=>"100100011",
  49456=>"101101011",
  49457=>"010001001",
  49458=>"011011011",
  49459=>"001010000",
  49460=>"100001010",
  49461=>"100110010",
  49462=>"000111011",
  49463=>"100110001",
  49464=>"100100000",
  49465=>"100100001",
  49466=>"111001001",
  49467=>"111111011",
  49468=>"111010011",
  49469=>"001001110",
  49470=>"101101010",
  49471=>"101001000",
  49472=>"001100111",
  49473=>"011000010",
  49474=>"100000100",
  49475=>"010111110",
  49476=>"001000101",
  49477=>"111010010",
  49478=>"100000100",
  49479=>"011001000",
  49480=>"101000111",
  49481=>"110000111",
  49482=>"101001101",
  49483=>"001110011",
  49484=>"011111110",
  49485=>"011111011",
  49486=>"000111111",
  49487=>"010100111",
  49488=>"011010011",
  49489=>"001001011",
  49490=>"010110100",
  49491=>"010110101",
  49492=>"100010100",
  49493=>"110110111",
  49494=>"100011110",
  49495=>"101011111",
  49496=>"010010101",
  49497=>"000101100",
  49498=>"111001101",
  49499=>"001100010",
  49500=>"010011011",
  49501=>"001011101",
  49502=>"111000110",
  49503=>"011010100",
  49504=>"001010110",
  49505=>"010110110",
  49506=>"011011101",
  49507=>"011100001",
  49508=>"000010000",
  49509=>"101100100",
  49510=>"100000001",
  49511=>"111110001",
  49512=>"000001001",
  49513=>"110110001",
  49514=>"010001011",
  49515=>"010000010",
  49516=>"000100000",
  49517=>"111011010",
  49518=>"101000001",
  49519=>"011110010",
  49520=>"110101001",
  49521=>"011001010",
  49522=>"111010100",
  49523=>"111011101",
  49524=>"101011001",
  49525=>"101110000",
  49526=>"010010001",
  49527=>"110111111",
  49528=>"010010000",
  49529=>"010010100",
  49530=>"011111001",
  49531=>"010110110",
  49532=>"000011111",
  49533=>"110111110",
  49534=>"111110010",
  49535=>"110001000",
  49536=>"100001010",
  49537=>"001010101",
  49538=>"101000001",
  49539=>"100011011",
  49540=>"101101011",
  49541=>"101000000",
  49542=>"101101011",
  49543=>"111001101",
  49544=>"010001011",
  49545=>"111110111",
  49546=>"001101101",
  49547=>"001111110",
  49548=>"001111101",
  49549=>"000111101",
  49550=>"100101100",
  49551=>"100100100",
  49552=>"101101100",
  49553=>"011001000",
  49554=>"011011100",
  49555=>"100111110",
  49556=>"100110100",
  49557=>"110010101",
  49558=>"111111111",
  49559=>"100010000",
  49560=>"101110011",
  49561=>"110101110",
  49562=>"000111100",
  49563=>"001110001",
  49564=>"001011011",
  49565=>"100100000",
  49566=>"100010100",
  49567=>"110111110",
  49568=>"101100101",
  49569=>"111000001",
  49570=>"010000000",
  49571=>"001001000",
  49572=>"111111101",
  49573=>"110011100",
  49574=>"010111110",
  49575=>"001100000",
  49576=>"110100111",
  49577=>"111111111",
  49578=>"101011100",
  49579=>"010001100",
  49580=>"011100000",
  49581=>"011101111",
  49582=>"000011100",
  49583=>"101100011",
  49584=>"111101010",
  49585=>"101101100",
  49586=>"111001111",
  49587=>"011000101",
  49588=>"110110011",
  49589=>"110001111",
  49590=>"101110010",
  49591=>"111001010",
  49592=>"110110101",
  49593=>"001000100",
  49594=>"111011010",
  49595=>"101011011",
  49596=>"100110111",
  49597=>"111111111",
  49598=>"001111101",
  49599=>"000001000",
  49600=>"100010011",
  49601=>"011101011",
  49602=>"001110001",
  49603=>"011111011",
  49604=>"010000110",
  49605=>"101100110",
  49606=>"001100101",
  49607=>"000000110",
  49608=>"011001001",
  49609=>"101100100",
  49610=>"011101111",
  49611=>"100111111",
  49612=>"100111101",
  49613=>"101000011",
  49614=>"100101100",
  49615=>"011011100",
  49616=>"110011101",
  49617=>"001000011",
  49618=>"101101110",
  49619=>"111001110",
  49620=>"110110001",
  49621=>"100001110",
  49622=>"110001110",
  49623=>"010101001",
  49624=>"111001100",
  49625=>"100111101",
  49626=>"100011001",
  49627=>"000100110",
  49628=>"100111101",
  49629=>"101101000",
  49630=>"111010010",
  49631=>"001100011",
  49632=>"110100000",
  49633=>"101010100",
  49634=>"110101101",
  49635=>"101000110",
  49636=>"000110000",
  49637=>"101001111",
  49638=>"001000010",
  49639=>"010010000",
  49640=>"110010101",
  49641=>"011000101",
  49642=>"100001011",
  49643=>"011011000",
  49644=>"111100110",
  49645=>"001110000",
  49646=>"000100000",
  49647=>"010010100",
  49648=>"001001111",
  49649=>"111110010",
  49650=>"100000010",
  49651=>"000110010",
  49652=>"111111111",
  49653=>"000111100",
  49654=>"000111010",
  49655=>"000010001",
  49656=>"010100001",
  49657=>"010101010",
  49658=>"001101010",
  49659=>"011110011",
  49660=>"111001111",
  49661=>"001010010",
  49662=>"110011111",
  49663=>"010100101",
  49664=>"110111111",
  49665=>"010101110",
  49666=>"110101110",
  49667=>"100010100",
  49668=>"001000011",
  49669=>"000000000",
  49670=>"011011111",
  49671=>"110101001",
  49672=>"001101001",
  49673=>"011011001",
  49674=>"111101000",
  49675=>"000010000",
  49676=>"101010110",
  49677=>"100110000",
  49678=>"101001000",
  49679=>"001111111",
  49680=>"110010000",
  49681=>"101011101",
  49682=>"011111000",
  49683=>"010110111",
  49684=>"100010010",
  49685=>"000111010",
  49686=>"001111101",
  49687=>"110101011",
  49688=>"100111110",
  49689=>"100000111",
  49690=>"101001001",
  49691=>"001110001",
  49692=>"001011001",
  49693=>"011010011",
  49694=>"111010111",
  49695=>"010011110",
  49696=>"101110011",
  49697=>"010100011",
  49698=>"100010111",
  49699=>"011100111",
  49700=>"111100001",
  49701=>"010101011",
  49702=>"000011011",
  49703=>"010110010",
  49704=>"011010110",
  49705=>"001010011",
  49706=>"110000110",
  49707=>"001111011",
  49708=>"100011010",
  49709=>"000000110",
  49710=>"110110000",
  49711=>"101001101",
  49712=>"111110000",
  49713=>"011101101",
  49714=>"101011111",
  49715=>"110101101",
  49716=>"111110101",
  49717=>"011100011",
  49718=>"001000011",
  49719=>"000001111",
  49720=>"011011110",
  49721=>"011110110",
  49722=>"000111010",
  49723=>"000111111",
  49724=>"010110001",
  49725=>"011010111",
  49726=>"100101110",
  49727=>"111100000",
  49728=>"011001111",
  49729=>"010111101",
  49730=>"001000001",
  49731=>"110110111",
  49732=>"010010111",
  49733=>"010010101",
  49734=>"001110010",
  49735=>"010100001",
  49736=>"110001001",
  49737=>"001001101",
  49738=>"001011101",
  49739=>"111101001",
  49740=>"001110101",
  49741=>"101100111",
  49742=>"111111011",
  49743=>"101000000",
  49744=>"010100101",
  49745=>"111111101",
  49746=>"001101011",
  49747=>"001011100",
  49748=>"000011101",
  49749=>"000011100",
  49750=>"000000000",
  49751=>"100011110",
  49752=>"110010010",
  49753=>"100000000",
  49754=>"001000001",
  49755=>"111000111",
  49756=>"101001101",
  49757=>"100001100",
  49758=>"000110101",
  49759=>"010010010",
  49760=>"100000000",
  49761=>"000101100",
  49762=>"010100101",
  49763=>"010111001",
  49764=>"111101110",
  49765=>"100001101",
  49766=>"100101111",
  49767=>"111001111",
  49768=>"010011110",
  49769=>"010000010",
  49770=>"010100000",
  49771=>"010100111",
  49772=>"001010110",
  49773=>"100011101",
  49774=>"110000010",
  49775=>"101000001",
  49776=>"010111000",
  49777=>"110111111",
  49778=>"000010000",
  49779=>"001011111",
  49780=>"011001111",
  49781=>"110001011",
  49782=>"111100100",
  49783=>"111010000",
  49784=>"101000111",
  49785=>"110101100",
  49786=>"100110011",
  49787=>"011011001",
  49788=>"010001010",
  49789=>"001001110",
  49790=>"100110101",
  49791=>"000110100",
  49792=>"101000100",
  49793=>"000111100",
  49794=>"111100110",
  49795=>"110000000",
  49796=>"000110100",
  49797=>"101110010",
  49798=>"110111010",
  49799=>"010100011",
  49800=>"110100010",
  49801=>"101001101",
  49802=>"100110110",
  49803=>"010101100",
  49804=>"001000011",
  49805=>"000011110",
  49806=>"111101000",
  49807=>"100001100",
  49808=>"010010100",
  49809=>"011110111",
  49810=>"010010110",
  49811=>"010101101",
  49812=>"000010001",
  49813=>"010110101",
  49814=>"011110111",
  49815=>"100101110",
  49816=>"010100101",
  49817=>"111100010",
  49818=>"011100011",
  49819=>"111110011",
  49820=>"001011001",
  49821=>"101110100",
  49822=>"110100000",
  49823=>"101010111",
  49824=>"000000101",
  49825=>"110011000",
  49826=>"000001010",
  49827=>"000011010",
  49828=>"110110000",
  49829=>"000010101",
  49830=>"000010100",
  49831=>"000001111",
  49832=>"010011101",
  49833=>"111110100",
  49834=>"010001101",
  49835=>"001001000",
  49836=>"001110000",
  49837=>"110010111",
  49838=>"101010010",
  49839=>"111111111",
  49840=>"100101000",
  49841=>"010010110",
  49842=>"000101110",
  49843=>"111001001",
  49844=>"011101000",
  49845=>"110111100",
  49846=>"101111010",
  49847=>"101111100",
  49848=>"011100010",
  49849=>"110100100",
  49850=>"111011000",
  49851=>"101010010",
  49852=>"001101000",
  49853=>"101111111",
  49854=>"111000101",
  49855=>"101110110",
  49856=>"111011100",
  49857=>"100100001",
  49858=>"010010100",
  49859=>"001111010",
  49860=>"101011111",
  49861=>"110101100",
  49862=>"101001111",
  49863=>"000101001",
  49864=>"010010000",
  49865=>"000001100",
  49866=>"000100101",
  49867=>"011001000",
  49868=>"011001001",
  49869=>"110000001",
  49870=>"011100101",
  49871=>"000111001",
  49872=>"000000001",
  49873=>"001010111",
  49874=>"010111100",
  49875=>"001011111",
  49876=>"011100100",
  49877=>"000001001",
  49878=>"110111010",
  49879=>"100011000",
  49880=>"101101010",
  49881=>"110100101",
  49882=>"000101100",
  49883=>"101111010",
  49884=>"011011111",
  49885=>"000000000",
  49886=>"001011010",
  49887=>"000110111",
  49888=>"011011001",
  49889=>"101000101",
  49890=>"111111110",
  49891=>"101111010",
  49892=>"001111000",
  49893=>"010010010",
  49894=>"011110001",
  49895=>"111111001",
  49896=>"000101011",
  49897=>"011010001",
  49898=>"010000011",
  49899=>"001110101",
  49900=>"001001001",
  49901=>"100010100",
  49902=>"100111011",
  49903=>"000000000",
  49904=>"011110100",
  49905=>"011110000",
  49906=>"001101101",
  49907=>"010111110",
  49908=>"011100000",
  49909=>"010101110",
  49910=>"010011011",
  49911=>"111011100",
  49912=>"010010110",
  49913=>"110101001",
  49914=>"010001100",
  49915=>"100111001",
  49916=>"010100100",
  49917=>"100010110",
  49918=>"101101010",
  49919=>"110100011",
  49920=>"010001100",
  49921=>"111010011",
  49922=>"010110011",
  49923=>"000011110",
  49924=>"000100011",
  49925=>"010110000",
  49926=>"000100011",
  49927=>"010011110",
  49928=>"101111000",
  49929=>"101110000",
  49930=>"110010110",
  49931=>"100101110",
  49932=>"000110011",
  49933=>"000111100",
  49934=>"001100000",
  49935=>"110110100",
  49936=>"000100111",
  49937=>"110100100",
  49938=>"111000100",
  49939=>"001100100",
  49940=>"000111111",
  49941=>"001110100",
  49942=>"010001111",
  49943=>"100010000",
  49944=>"001001001",
  49945=>"011111001",
  49946=>"111110011",
  49947=>"000001111",
  49948=>"011101110",
  49949=>"000000110",
  49950=>"100100110",
  49951=>"011011010",
  49952=>"100010111",
  49953=>"111001001",
  49954=>"101110111",
  49955=>"001101101",
  49956=>"000111000",
  49957=>"100101001",
  49958=>"001011101",
  49959=>"101011101",
  49960=>"000100011",
  49961=>"010000000",
  49962=>"011011010",
  49963=>"110000100",
  49964=>"000110100",
  49965=>"111010010",
  49966=>"001101101",
  49967=>"110011101",
  49968=>"101011100",
  49969=>"000001001",
  49970=>"110110010",
  49971=>"001001001",
  49972=>"111000111",
  49973=>"010101111",
  49974=>"101001110",
  49975=>"011000010",
  49976=>"001100110",
  49977=>"110011111",
  49978=>"011111100",
  49979=>"100100000",
  49980=>"110001000",
  49981=>"100001011",
  49982=>"001011100",
  49983=>"110110110",
  49984=>"110010111",
  49985=>"011101001",
  49986=>"000010111",
  49987=>"110001111",
  49988=>"101011101",
  49989=>"110000000",
  49990=>"101011000",
  49991=>"111011111",
  49992=>"010101110",
  49993=>"001011011",
  49994=>"101001000",
  49995=>"001000101",
  49996=>"110110100",
  49997=>"000000001",
  49998=>"110000001",
  49999=>"110110000",
  50000=>"100001011",
  50001=>"010111100",
  50002=>"100011101",
  50003=>"110110001",
  50004=>"100110100",
  50005=>"000100110",
  50006=>"111000011",
  50007=>"000010000",
  50008=>"000111111",
  50009=>"101011101",
  50010=>"000010110",
  50011=>"101010101",
  50012=>"100001000",
  50013=>"100001011",
  50014=>"111111101",
  50015=>"110100011",
  50016=>"001111010",
  50017=>"101110011",
  50018=>"001101110",
  50019=>"011001000",
  50020=>"100000110",
  50021=>"011010101",
  50022=>"100100011",
  50023=>"100110100",
  50024=>"000001010",
  50025=>"101001110",
  50026=>"001010011",
  50027=>"000010010",
  50028=>"111100100",
  50029=>"000101000",
  50030=>"001000001",
  50031=>"001111110",
  50032=>"100011011",
  50033=>"110110101",
  50034=>"011010110",
  50035=>"100100001",
  50036=>"101100101",
  50037=>"111100100",
  50038=>"101011001",
  50039=>"010000010",
  50040=>"000000010",
  50041=>"100100000",
  50042=>"011010101",
  50043=>"000010011",
  50044=>"101111110",
  50045=>"111111001",
  50046=>"101100011",
  50047=>"111000111",
  50048=>"010100010",
  50049=>"000111111",
  50050=>"110100100",
  50051=>"010001010",
  50052=>"100100110",
  50053=>"011010111",
  50054=>"100100111",
  50055=>"111100100",
  50056=>"001010111",
  50057=>"100011011",
  50058=>"111111100",
  50059=>"011101011",
  50060=>"111011111",
  50061=>"000001111",
  50062=>"110100010",
  50063=>"001010110",
  50064=>"100100101",
  50065=>"101111111",
  50066=>"100101000",
  50067=>"101000111",
  50068=>"110001001",
  50069=>"010100111",
  50070=>"011101001",
  50071=>"111010000",
  50072=>"101010011",
  50073=>"111011101",
  50074=>"111011111",
  50075=>"100100000",
  50076=>"101100011",
  50077=>"100000111",
  50078=>"001010000",
  50079=>"110010001",
  50080=>"010011111",
  50081=>"111110111",
  50082=>"110010001",
  50083=>"000001010",
  50084=>"001101100",
  50085=>"011001001",
  50086=>"011011100",
  50087=>"010110110",
  50088=>"000010001",
  50089=>"100010010",
  50090=>"011011011",
  50091=>"100001010",
  50092=>"101010101",
  50093=>"111110100",
  50094=>"011111110",
  50095=>"100010111",
  50096=>"010010010",
  50097=>"110111000",
  50098=>"010000011",
  50099=>"001010111",
  50100=>"011000101",
  50101=>"001000011",
  50102=>"011001011",
  50103=>"100100001",
  50104=>"011010101",
  50105=>"010000110",
  50106=>"101011100",
  50107=>"101110010",
  50108=>"001111001",
  50109=>"010000010",
  50110=>"101001111",
  50111=>"000001111",
  50112=>"011011000",
  50113=>"101001110",
  50114=>"101000110",
  50115=>"101101101",
  50116=>"000000101",
  50117=>"000110101",
  50118=>"000010011",
  50119=>"100001100",
  50120=>"110100100",
  50121=>"000000000",
  50122=>"101101110",
  50123=>"100100011",
  50124=>"100110011",
  50125=>"101001011",
  50126=>"010011101",
  50127=>"100111110",
  50128=>"000110110",
  50129=>"100100001",
  50130=>"000010000",
  50131=>"001001000",
  50132=>"011001111",
  50133=>"110001010",
  50134=>"000000010",
  50135=>"010100110",
  50136=>"110010011",
  50137=>"000000100",
  50138=>"100111111",
  50139=>"101011100",
  50140=>"010111100",
  50141=>"000111100",
  50142=>"010011000",
  50143=>"101100001",
  50144=>"111100111",
  50145=>"001011111",
  50146=>"100010111",
  50147=>"001111100",
  50148=>"101101111",
  50149=>"000000000",
  50150=>"011110111",
  50151=>"100000110",
  50152=>"000101111",
  50153=>"101100100",
  50154=>"101100101",
  50155=>"100001010",
  50156=>"101000000",
  50157=>"110011101",
  50158=>"011111010",
  50159=>"110111101",
  50160=>"101101001",
  50161=>"100000001",
  50162=>"101110110",
  50163=>"110001011",
  50164=>"000000011",
  50165=>"010010100",
  50166=>"001010000",
  50167=>"110110110",
  50168=>"000011010",
  50169=>"010111011",
  50170=>"100101011",
  50171=>"011011011",
  50172=>"111101111",
  50173=>"000010010",
  50174=>"000100011",
  50175=>"011000101",
  50176=>"011101011",
  50177=>"000000000",
  50178=>"001010100",
  50179=>"010000101",
  50180=>"100011110",
  50181=>"000001010",
  50182=>"110100000",
  50183=>"101111000",
  50184=>"110110101",
  50185=>"100101000",
  50186=>"101001111",
  50187=>"111010000",
  50188=>"101010110",
  50189=>"101011000",
  50190=>"100101000",
  50191=>"111001111",
  50192=>"111001011",
  50193=>"010111101",
  50194=>"001101101",
  50195=>"011011111",
  50196=>"111000110",
  50197=>"101010010",
  50198=>"111100001",
  50199=>"110010011",
  50200=>"100001100",
  50201=>"010100110",
  50202=>"001011000",
  50203=>"100000000",
  50204=>"101100111",
  50205=>"111011100",
  50206=>"110101011",
  50207=>"110011101",
  50208=>"001010000",
  50209=>"000011110",
  50210=>"010000000",
  50211=>"001011111",
  50212=>"001001100",
  50213=>"100000110",
  50214=>"111000100",
  50215=>"110101001",
  50216=>"001001000",
  50217=>"011111111",
  50218=>"011001001",
  50219=>"110110101",
  50220=>"011000100",
  50221=>"000000110",
  50222=>"101001101",
  50223=>"011111000",
  50224=>"001011110",
  50225=>"111001010",
  50226=>"010011011",
  50227=>"100110011",
  50228=>"000010101",
  50229=>"101110000",
  50230=>"001100100",
  50231=>"001110010",
  50232=>"010001101",
  50233=>"101000100",
  50234=>"101000010",
  50235=>"001110111",
  50236=>"110011110",
  50237=>"000101011",
  50238=>"111101111",
  50239=>"011000011",
  50240=>"110011100",
  50241=>"011101011",
  50242=>"101011111",
  50243=>"010111011",
  50244=>"011111001",
  50245=>"000000111",
  50246=>"000010111",
  50247=>"001000111",
  50248=>"000010111",
  50249=>"111010011",
  50250=>"110010001",
  50251=>"001000010",
  50252=>"101010000",
  50253=>"001010100",
  50254=>"100111111",
  50255=>"101111111",
  50256=>"001010010",
  50257=>"000100011",
  50258=>"111101001",
  50259=>"110001000",
  50260=>"101110110",
  50261=>"110100011",
  50262=>"110011111",
  50263=>"000000011",
  50264=>"000101111",
  50265=>"010111100",
  50266=>"110110101",
  50267=>"011100010",
  50268=>"100001100",
  50269=>"100000110",
  50270=>"111100001",
  50271=>"000111100",
  50272=>"111010010",
  50273=>"100111110",
  50274=>"010100100",
  50275=>"110100111",
  50276=>"110100100",
  50277=>"101101010",
  50278=>"010000101",
  50279=>"110000001",
  50280=>"100000100",
  50281=>"100101111",
  50282=>"101111000",
  50283=>"110001101",
  50284=>"001111110",
  50285=>"001001111",
  50286=>"111100011",
  50287=>"110111001",
  50288=>"110101100",
  50289=>"000010000",
  50290=>"100001110",
  50291=>"001010001",
  50292=>"001110111",
  50293=>"100000111",
  50294=>"001111001",
  50295=>"110010101",
  50296=>"110000010",
  50297=>"000110100",
  50298=>"100001001",
  50299=>"110001110",
  50300=>"000111110",
  50301=>"010010010",
  50302=>"011101100",
  50303=>"100001100",
  50304=>"001001101",
  50305=>"110000000",
  50306=>"101010001",
  50307=>"101011100",
  50308=>"000000111",
  50309=>"101001001",
  50310=>"110111010",
  50311=>"010010101",
  50312=>"000101101",
  50313=>"111101100",
  50314=>"011110000",
  50315=>"011100000",
  50316=>"011110101",
  50317=>"000110001",
  50318=>"010001011",
  50319=>"010011010",
  50320=>"111111100",
  50321=>"111101011",
  50322=>"111100111",
  50323=>"100011100",
  50324=>"000100101",
  50325=>"000100110",
  50326=>"010010011",
  50327=>"010010111",
  50328=>"101111011",
  50329=>"001011111",
  50330=>"101101011",
  50331=>"000011111",
  50332=>"110100011",
  50333=>"010111001",
  50334=>"110111111",
  50335=>"010100110",
  50336=>"100110100",
  50337=>"011010010",
  50338=>"100001000",
  50339=>"000101010",
  50340=>"000110010",
  50341=>"100001000",
  50342=>"010101111",
  50343=>"010001010",
  50344=>"111001001",
  50345=>"010001010",
  50346=>"101010001",
  50347=>"001100000",
  50348=>"110110110",
  50349=>"000101011",
  50350=>"100000100",
  50351=>"100010100",
  50352=>"000111001",
  50353=>"111101110",
  50354=>"000000010",
  50355=>"000101001",
  50356=>"001000101",
  50357=>"110111100",
  50358=>"101111111",
  50359=>"011100111",
  50360=>"011101001",
  50361=>"101100110",
  50362=>"001100101",
  50363=>"000110101",
  50364=>"001010011",
  50365=>"001001000",
  50366=>"111101110",
  50367=>"100011011",
  50368=>"011001110",
  50369=>"100100000",
  50370=>"110100000",
  50371=>"010010101",
  50372=>"101111010",
  50373=>"100011011",
  50374=>"100001101",
  50375=>"001000100",
  50376=>"000111110",
  50377=>"000000111",
  50378=>"000000011",
  50379=>"011000111",
  50380=>"011000000",
  50381=>"101000100",
  50382=>"110100111",
  50383=>"100101010",
  50384=>"001101000",
  50385=>"100011111",
  50386=>"101011100",
  50387=>"111100010",
  50388=>"001011011",
  50389=>"010000110",
  50390=>"101111111",
  50391=>"011011001",
  50392=>"110100001",
  50393=>"100111111",
  50394=>"010110000",
  50395=>"000100010",
  50396=>"101010001",
  50397=>"101001111",
  50398=>"101110011",
  50399=>"100011010",
  50400=>"001001010",
  50401=>"110001100",
  50402=>"010110100",
  50403=>"110111001",
  50404=>"000111100",
  50405=>"000101111",
  50406=>"111000011",
  50407=>"101110101",
  50408=>"000110100",
  50409=>"110111011",
  50410=>"011110111",
  50411=>"111100110",
  50412=>"101000010",
  50413=>"111111110",
  50414=>"110001001",
  50415=>"110101010",
  50416=>"111111111",
  50417=>"000100010",
  50418=>"111100001",
  50419=>"000100111",
  50420=>"001010100",
  50421=>"100101100",
  50422=>"000111000",
  50423=>"110000000",
  50424=>"001110101",
  50425=>"101110111",
  50426=>"010101111",
  50427=>"010000000",
  50428=>"011100101",
  50429=>"110010100",
  50430=>"111110101",
  50431=>"001010010",
  50432=>"000100010",
  50433=>"000110100",
  50434=>"011110101",
  50435=>"000001011",
  50436=>"010101011",
  50437=>"011100010",
  50438=>"111011111",
  50439=>"100011001",
  50440=>"100010100",
  50441=>"010001110",
  50442=>"010100011",
  50443=>"110010110",
  50444=>"011001100",
  50445=>"001101010",
  50446=>"001011101",
  50447=>"101000110",
  50448=>"011000000",
  50449=>"000010001",
  50450=>"100010011",
  50451=>"000110100",
  50452=>"110111000",
  50453=>"001100111",
  50454=>"010101010",
  50455=>"010001101",
  50456=>"101010000",
  50457=>"110011001",
  50458=>"101101010",
  50459=>"011110111",
  50460=>"000010011",
  50461=>"100011000",
  50462=>"101101000",
  50463=>"101011010",
  50464=>"000000010",
  50465=>"011010001",
  50466=>"110101001",
  50467=>"111101111",
  50468=>"000000100",
  50469=>"000100010",
  50470=>"101110010",
  50471=>"011110000",
  50472=>"101100000",
  50473=>"000100101",
  50474=>"000011001",
  50475=>"010100001",
  50476=>"110101101",
  50477=>"110010101",
  50478=>"110101100",
  50479=>"000100110",
  50480=>"010000010",
  50481=>"111111111",
  50482=>"001000010",
  50483=>"011011101",
  50484=>"101011100",
  50485=>"111100010",
  50486=>"111100101",
  50487=>"100001101",
  50488=>"011100001",
  50489=>"011101001",
  50490=>"000000000",
  50491=>"110011010",
  50492=>"111011001",
  50493=>"101110111",
  50494=>"110011101",
  50495=>"001110101",
  50496=>"011100111",
  50497=>"000000000",
  50498=>"000111000",
  50499=>"101000001",
  50500=>"101000111",
  50501=>"010010111",
  50502=>"001110010",
  50503=>"101110111",
  50504=>"110011011",
  50505=>"010110101",
  50506=>"000001010",
  50507=>"000001010",
  50508=>"100001101",
  50509=>"101100011",
  50510=>"110001110",
  50511=>"000110001",
  50512=>"010110101",
  50513=>"110000110",
  50514=>"000110010",
  50515=>"000000001",
  50516=>"010101010",
  50517=>"010010110",
  50518=>"010000101",
  50519=>"110111110",
  50520=>"010111101",
  50521=>"000000100",
  50522=>"010111001",
  50523=>"100010100",
  50524=>"101101111",
  50525=>"110011111",
  50526=>"010010110",
  50527=>"011111011",
  50528=>"011110110",
  50529=>"101110111",
  50530=>"111101111",
  50531=>"101001000",
  50532=>"011011000",
  50533=>"100000010",
  50534=>"110100111",
  50535=>"011001011",
  50536=>"010000111",
  50537=>"110001000",
  50538=>"101100011",
  50539=>"000010111",
  50540=>"100000001",
  50541=>"100100110",
  50542=>"101011010",
  50543=>"100011001",
  50544=>"111110010",
  50545=>"001111101",
  50546=>"011101011",
  50547=>"110000001",
  50548=>"000001010",
  50549=>"011110100",
  50550=>"001011001",
  50551=>"000111001",
  50552=>"100011111",
  50553=>"101000001",
  50554=>"000010001",
  50555=>"100100010",
  50556=>"001100100",
  50557=>"001010001",
  50558=>"110111101",
  50559=>"000101011",
  50560=>"100100100",
  50561=>"110100001",
  50562=>"100110001",
  50563=>"110101101",
  50564=>"000000101",
  50565=>"000110100",
  50566=>"010110001",
  50567=>"000000100",
  50568=>"111111111",
  50569=>"000011110",
  50570=>"111101110",
  50571=>"101000110",
  50572=>"111010001",
  50573=>"011111011",
  50574=>"011011010",
  50575=>"011000010",
  50576=>"010011100",
  50577=>"110011000",
  50578=>"100101100",
  50579=>"101001011",
  50580=>"010011000",
  50581=>"000000000",
  50582=>"110110111",
  50583=>"000001111",
  50584=>"000111001",
  50585=>"111111110",
  50586=>"000110110",
  50587=>"101011001",
  50588=>"101110100",
  50589=>"001111001",
  50590=>"100011100",
  50591=>"110010001",
  50592=>"010001110",
  50593=>"111111010",
  50594=>"100111101",
  50595=>"101100011",
  50596=>"101010011",
  50597=>"011000100",
  50598=>"100000101",
  50599=>"000101001",
  50600=>"110100111",
  50601=>"000010001",
  50602=>"101000100",
  50603=>"010100000",
  50604=>"011101101",
  50605=>"011011000",
  50606=>"010100010",
  50607=>"011001111",
  50608=>"010001000",
  50609=>"111010010",
  50610=>"110000100",
  50611=>"010000010",
  50612=>"111010110",
  50613=>"000100100",
  50614=>"011000001",
  50615=>"111100111",
  50616=>"011000110",
  50617=>"111010111",
  50618=>"111000111",
  50619=>"011000100",
  50620=>"010111100",
  50621=>"010101101",
  50622=>"001100100",
  50623=>"101010000",
  50624=>"111000010",
  50625=>"011110111",
  50626=>"000010110",
  50627=>"000111010",
  50628=>"101000000",
  50629=>"011111100",
  50630=>"101111101",
  50631=>"111111001",
  50632=>"100001001",
  50633=>"101000101",
  50634=>"010001101",
  50635=>"011110101",
  50636=>"011111110",
  50637=>"010001011",
  50638=>"001110100",
  50639=>"110001001",
  50640=>"100000101",
  50641=>"011011101",
  50642=>"001001101",
  50643=>"111010110",
  50644=>"000111000",
  50645=>"001010000",
  50646=>"100011000",
  50647=>"110111011",
  50648=>"001100101",
  50649=>"110000000",
  50650=>"010101001",
  50651=>"110000001",
  50652=>"001000011",
  50653=>"010100111",
  50654=>"111011110",
  50655=>"100111111",
  50656=>"100010100",
  50657=>"100011010",
  50658=>"000001100",
  50659=>"010000000",
  50660=>"101101110",
  50661=>"101100000",
  50662=>"100000001",
  50663=>"110101011",
  50664=>"100011011",
  50665=>"010010011",
  50666=>"000101010",
  50667=>"111100001",
  50668=>"000100000",
  50669=>"100111101",
  50670=>"110111010",
  50671=>"001000000",
  50672=>"110101010",
  50673=>"101111101",
  50674=>"001101100",
  50675=>"011001101",
  50676=>"000100110",
  50677=>"000111111",
  50678=>"111110101",
  50679=>"110001100",
  50680=>"011010110",
  50681=>"101010100",
  50682=>"000110100",
  50683=>"110101001",
  50684=>"111100001",
  50685=>"110100001",
  50686=>"000010100",
  50687=>"101110011",
  50688=>"001010011",
  50689=>"100001111",
  50690=>"100100011",
  50691=>"011101111",
  50692=>"001011101",
  50693=>"001110110",
  50694=>"010100001",
  50695=>"000001010",
  50696=>"001101011",
  50697=>"111110001",
  50698=>"001000010",
  50699=>"001001000",
  50700=>"011111010",
  50701=>"011001111",
  50702=>"110011001",
  50703=>"011001000",
  50704=>"101110110",
  50705=>"011111001",
  50706=>"001010001",
  50707=>"100000110",
  50708=>"101010010",
  50709=>"110001010",
  50710=>"100101100",
  50711=>"111011100",
  50712=>"101101001",
  50713=>"101001011",
  50714=>"001101000",
  50715=>"100001011",
  50716=>"000001101",
  50717=>"110011001",
  50718=>"011110001",
  50719=>"110110111",
  50720=>"101011100",
  50721=>"011010001",
  50722=>"001100010",
  50723=>"001000010",
  50724=>"110101111",
  50725=>"111100111",
  50726=>"011000011",
  50727=>"111100101",
  50728=>"110011001",
  50729=>"111001000",
  50730=>"101011000",
  50731=>"000000011",
  50732=>"000000100",
  50733=>"110101111",
  50734=>"111000100",
  50735=>"111110110",
  50736=>"111000101",
  50737=>"000110101",
  50738=>"010011011",
  50739=>"000000000",
  50740=>"001001000",
  50741=>"100100111",
  50742=>"111000000",
  50743=>"000100000",
  50744=>"101000010",
  50745=>"000111100",
  50746=>"001000110",
  50747=>"101001000",
  50748=>"011110000",
  50749=>"000001111",
  50750=>"001000000",
  50751=>"011000101",
  50752=>"100101001",
  50753=>"001101100",
  50754=>"101000111",
  50755=>"111101000",
  50756=>"001011111",
  50757=>"101101100",
  50758=>"101011010",
  50759=>"110001100",
  50760=>"101010010",
  50761=>"010010000",
  50762=>"101111001",
  50763=>"010110000",
  50764=>"001001000",
  50765=>"111001101",
  50766=>"111011010",
  50767=>"101001101",
  50768=>"110000101",
  50769=>"001010111",
  50770=>"000101101",
  50771=>"001111000",
  50772=>"010100101",
  50773=>"000110110",
  50774=>"101101101",
  50775=>"101111111",
  50776=>"110011011",
  50777=>"000001101",
  50778=>"111111000",
  50779=>"011000110",
  50780=>"100101011",
  50781=>"100000001",
  50782=>"001001110",
  50783=>"110100010",
  50784=>"001010100",
  50785=>"011000100",
  50786=>"110101111",
  50787=>"111100111",
  50788=>"110110011",
  50789=>"110000111",
  50790=>"110101100",
  50791=>"111101100",
  50792=>"100100010",
  50793=>"111110111",
  50794=>"101111001",
  50795=>"101000101",
  50796=>"001001100",
  50797=>"111011100",
  50798=>"011110110",
  50799=>"010011001",
  50800=>"100101010",
  50801=>"011010011",
  50802=>"001110100",
  50803=>"101010110",
  50804=>"001100011",
  50805=>"001110001",
  50806=>"101011001",
  50807=>"011000011",
  50808=>"011011110",
  50809=>"100000010",
  50810=>"011011111",
  50811=>"110101111",
  50812=>"100110011",
  50813=>"010111000",
  50814=>"110010101",
  50815=>"101010110",
  50816=>"010000110",
  50817=>"110000010",
  50818=>"110001101",
  50819=>"000010100",
  50820=>"111101000",
  50821=>"011000100",
  50822=>"000100010",
  50823=>"001110011",
  50824=>"011100001",
  50825=>"101000001",
  50826=>"110010110",
  50827=>"001001011",
  50828=>"101000011",
  50829=>"100001101",
  50830=>"010001001",
  50831=>"111101111",
  50832=>"011011001",
  50833=>"111111101",
  50834=>"001011111",
  50835=>"101011010",
  50836=>"111010101",
  50837=>"111000001",
  50838=>"101111000",
  50839=>"101011010",
  50840=>"000000000",
  50841=>"001001000",
  50842=>"001100100",
  50843=>"011111010",
  50844=>"001010011",
  50845=>"101110110",
  50846=>"101011110",
  50847=>"010100101",
  50848=>"010111001",
  50849=>"110111110",
  50850=>"010101100",
  50851=>"111110010",
  50852=>"100110100",
  50853=>"110101110",
  50854=>"010110000",
  50855=>"000000000",
  50856=>"111101111",
  50857=>"101001010",
  50858=>"111010010",
  50859=>"100010110",
  50860=>"110000000",
  50861=>"010010001",
  50862=>"111101001",
  50863=>"000011000",
  50864=>"001101011",
  50865=>"001010111",
  50866=>"010010000",
  50867=>"010111011",
  50868=>"111101001",
  50869=>"111100100",
  50870=>"011000010",
  50871=>"101100111",
  50872=>"111010001",
  50873=>"100111011",
  50874=>"001010010",
  50875=>"101011001",
  50876=>"000111101",
  50877=>"101011001",
  50878=>"000111101",
  50879=>"111010111",
  50880=>"001000110",
  50881=>"001000000",
  50882=>"101110100",
  50883=>"011011111",
  50884=>"000100011",
  50885=>"110100001",
  50886=>"100111110",
  50887=>"011110101",
  50888=>"010001110",
  50889=>"000011000",
  50890=>"110100110",
  50891=>"011100110",
  50892=>"101000101",
  50893=>"001111011",
  50894=>"011010111",
  50895=>"101010010",
  50896=>"001110110",
  50897=>"111101010",
  50898=>"001101101",
  50899=>"111010011",
  50900=>"000010000",
  50901=>"111111110",
  50902=>"010010101",
  50903=>"100100010",
  50904=>"010011001",
  50905=>"001010110",
  50906=>"110111101",
  50907=>"011111110",
  50908=>"100100110",
  50909=>"000011111",
  50910=>"101100111",
  50911=>"000000101",
  50912=>"110011010",
  50913=>"101001011",
  50914=>"100101010",
  50915=>"100000001",
  50916=>"001000010",
  50917=>"001100000",
  50918=>"110110001",
  50919=>"011000000",
  50920=>"010101000",
  50921=>"100001011",
  50922=>"101001001",
  50923=>"110001010",
  50924=>"000000110",
  50925=>"110010000",
  50926=>"011111010",
  50927=>"101010101",
  50928=>"100110101",
  50929=>"110011010",
  50930=>"011000001",
  50931=>"000010010",
  50932=>"011010000",
  50933=>"001111010",
  50934=>"011001001",
  50935=>"001111010",
  50936=>"110001000",
  50937=>"100111111",
  50938=>"100011000",
  50939=>"110010110",
  50940=>"111110101",
  50941=>"111111100",
  50942=>"111101110",
  50943=>"111001110",
  50944=>"110110101",
  50945=>"000111111",
  50946=>"111110110",
  50947=>"001011100",
  50948=>"010000000",
  50949=>"011000101",
  50950=>"110100110",
  50951=>"111011111",
  50952=>"010000100",
  50953=>"001101100",
  50954=>"011010100",
  50955=>"101000110",
  50956=>"101000000",
  50957=>"110010001",
  50958=>"100110001",
  50959=>"000100111",
  50960=>"111111011",
  50961=>"001000001",
  50962=>"101001111",
  50963=>"010100100",
  50964=>"011001001",
  50965=>"011010100",
  50966=>"010011110",
  50967=>"001001001",
  50968=>"011111000",
  50969=>"100100010",
  50970=>"111011001",
  50971=>"000101111",
  50972=>"001111010",
  50973=>"110110101",
  50974=>"011111100",
  50975=>"100010100",
  50976=>"110001110",
  50977=>"111010011",
  50978=>"011101101",
  50979=>"001100101",
  50980=>"110111111",
  50981=>"010100110",
  50982=>"101000110",
  50983=>"001111110",
  50984=>"101001101",
  50985=>"100011110",
  50986=>"011101111",
  50987=>"011111010",
  50988=>"001001100",
  50989=>"000000000",
  50990=>"110000011",
  50991=>"101101100",
  50992=>"110001000",
  50993=>"010110110",
  50994=>"110010100",
  50995=>"101110010",
  50996=>"101111011",
  50997=>"010110101",
  50998=>"101010111",
  50999=>"101111010",
  51000=>"010101110",
  51001=>"011011111",
  51002=>"010110110",
  51003=>"100101110",
  51004=>"110011111",
  51005=>"011100011",
  51006=>"110011011",
  51007=>"001010010",
  51008=>"100110000",
  51009=>"010101011",
  51010=>"111110011",
  51011=>"101111000",
  51012=>"010111110",
  51013=>"001001010",
  51014=>"000110010",
  51015=>"011100100",
  51016=>"101111101",
  51017=>"001111111",
  51018=>"000000000",
  51019=>"010111000",
  51020=>"101111111",
  51021=>"100000011",
  51022=>"011111010",
  51023=>"101000111",
  51024=>"111011100",
  51025=>"111111000",
  51026=>"100000010",
  51027=>"010011000",
  51028=>"111110101",
  51029=>"010111111",
  51030=>"010100001",
  51031=>"111000100",
  51032=>"011111001",
  51033=>"110000111",
  51034=>"111010011",
  51035=>"010110011",
  51036=>"001110000",
  51037=>"010101110",
  51038=>"010001001",
  51039=>"000100011",
  51040=>"111001000",
  51041=>"011101100",
  51042=>"100000101",
  51043=>"111111011",
  51044=>"001001110",
  51045=>"100101101",
  51046=>"000111010",
  51047=>"110000001",
  51048=>"010110100",
  51049=>"101001011",
  51050=>"100110110",
  51051=>"110000011",
  51052=>"010000110",
  51053=>"100010111",
  51054=>"100011001",
  51055=>"100101110",
  51056=>"010000010",
  51057=>"001001001",
  51058=>"011110011",
  51059=>"110011011",
  51060=>"110101111",
  51061=>"110001010",
  51062=>"110011000",
  51063=>"101101100",
  51064=>"101011000",
  51065=>"111011010",
  51066=>"110100100",
  51067=>"001011111",
  51068=>"001001000",
  51069=>"100101110",
  51070=>"000111010",
  51071=>"010101100",
  51072=>"110000001",
  51073=>"001110011",
  51074=>"101000001",
  51075=>"111010011",
  51076=>"101000001",
  51077=>"000110011",
  51078=>"100000101",
  51079=>"011111100",
  51080=>"100111101",
  51081=>"000101101",
  51082=>"011101010",
  51083=>"111100000",
  51084=>"100010000",
  51085=>"111001111",
  51086=>"000000011",
  51087=>"010111100",
  51088=>"100000000",
  51089=>"000001000",
  51090=>"001110010",
  51091=>"100011111",
  51092=>"110010000",
  51093=>"100011111",
  51094=>"010001111",
  51095=>"100011111",
  51096=>"100100111",
  51097=>"010011000",
  51098=>"011000101",
  51099=>"101110100",
  51100=>"100011111",
  51101=>"010101001",
  51102=>"100101000",
  51103=>"011001010",
  51104=>"000011010",
  51105=>"100011000",
  51106=>"010100000",
  51107=>"000110110",
  51108=>"111011000",
  51109=>"011110110",
  51110=>"111000111",
  51111=>"111001110",
  51112=>"000000110",
  51113=>"111001101",
  51114=>"011111010",
  51115=>"110010101",
  51116=>"000000000",
  51117=>"101101101",
  51118=>"101000000",
  51119=>"111001001",
  51120=>"111001010",
  51121=>"010111111",
  51122=>"000010110",
  51123=>"100001010",
  51124=>"110111111",
  51125=>"111111100",
  51126=>"111101011",
  51127=>"000000010",
  51128=>"000010111",
  51129=>"101001111",
  51130=>"000000011",
  51131=>"000110110",
  51132=>"111100101",
  51133=>"110001010",
  51134=>"110000110",
  51135=>"010011000",
  51136=>"001101001",
  51137=>"011001001",
  51138=>"101101100",
  51139=>"111000000",
  51140=>"000000011",
  51141=>"010000100",
  51142=>"001110101",
  51143=>"001010100",
  51144=>"011111110",
  51145=>"010001110",
  51146=>"011011001",
  51147=>"010101011",
  51148=>"111111101",
  51149=>"101100111",
  51150=>"001101111",
  51151=>"101010010",
  51152=>"001101010",
  51153=>"001000100",
  51154=>"101011111",
  51155=>"001010010",
  51156=>"100111011",
  51157=>"011010011",
  51158=>"010010100",
  51159=>"010100001",
  51160=>"111001011",
  51161=>"001011010",
  51162=>"101011011",
  51163=>"011001110",
  51164=>"101110011",
  51165=>"110011010",
  51166=>"011101010",
  51167=>"110000011",
  51168=>"101001110",
  51169=>"010100110",
  51170=>"000101010",
  51171=>"101111001",
  51172=>"111111000",
  51173=>"010100001",
  51174=>"001000111",
  51175=>"111111000",
  51176=>"110010110",
  51177=>"110100010",
  51178=>"000001011",
  51179=>"110101011",
  51180=>"011001111",
  51181=>"000011001",
  51182=>"101000000",
  51183=>"000000111",
  51184=>"011000010",
  51185=>"000110001",
  51186=>"101011010",
  51187=>"011001001",
  51188=>"001000001",
  51189=>"001010110",
  51190=>"100110110",
  51191=>"011000000",
  51192=>"011001001",
  51193=>"101111100",
  51194=>"110001001",
  51195=>"110111011",
  51196=>"110000111",
  51197=>"011011111",
  51198=>"110101111",
  51199=>"110110110",
  51200=>"000111100",
  51201=>"010000101",
  51202=>"010100011",
  51203=>"011111101",
  51204=>"100011111",
  51205=>"100010110",
  51206=>"000001011",
  51207=>"011000011",
  51208=>"010011101",
  51209=>"001111010",
  51210=>"000101101",
  51211=>"110010100",
  51212=>"100101010",
  51213=>"011011011",
  51214=>"000011000",
  51215=>"101101011",
  51216=>"100100110",
  51217=>"101010111",
  51218=>"000110010",
  51219=>"100100000",
  51220=>"110111110",
  51221=>"101101101",
  51222=>"000101110",
  51223=>"100000001",
  51224=>"101100111",
  51225=>"101010100",
  51226=>"100000101",
  51227=>"110110110",
  51228=>"100001001",
  51229=>"000001101",
  51230=>"101101110",
  51231=>"011100010",
  51232=>"111101000",
  51233=>"100011101",
  51234=>"001100101",
  51235=>"100000100",
  51236=>"100110110",
  51237=>"110001000",
  51238=>"111000110",
  51239=>"000101110",
  51240=>"110010100",
  51241=>"100100010",
  51242=>"110011111",
  51243=>"001001100",
  51244=>"110111000",
  51245=>"000011011",
  51246=>"110011100",
  51247=>"110100001",
  51248=>"100010010",
  51249=>"100111100",
  51250=>"000101100",
  51251=>"000001011",
  51252=>"111111100",
  51253=>"000111000",
  51254=>"001000100",
  51255=>"010101001",
  51256=>"100000001",
  51257=>"110010110",
  51258=>"101011001",
  51259=>"000100110",
  51260=>"001100100",
  51261=>"000000001",
  51262=>"110101100",
  51263=>"101001000",
  51264=>"101100111",
  51265=>"000010000",
  51266=>"001011100",
  51267=>"100100101",
  51268=>"100010110",
  51269=>"101001101",
  51270=>"100101011",
  51271=>"001000101",
  51272=>"101111000",
  51273=>"001010010",
  51274=>"110001001",
  51275=>"100010100",
  51276=>"111101100",
  51277=>"010101111",
  51278=>"010101010",
  51279=>"001110010",
  51280=>"011110100",
  51281=>"111011110",
  51282=>"011100011",
  51283=>"101100100",
  51284=>"010101011",
  51285=>"011110011",
  51286=>"010011010",
  51287=>"110100101",
  51288=>"110101011",
  51289=>"100000111",
  51290=>"110101010",
  51291=>"001101011",
  51292=>"111011011",
  51293=>"101110010",
  51294=>"001110010",
  51295=>"011101110",
  51296=>"001010100",
  51297=>"101010000",
  51298=>"011110111",
  51299=>"000011011",
  51300=>"111100111",
  51301=>"100110100",
  51302=>"010101010",
  51303=>"010111110",
  51304=>"100110101",
  51305=>"011011011",
  51306=>"000000010",
  51307=>"001001111",
  51308=>"111101101",
  51309=>"001011111",
  51310=>"001010110",
  51311=>"110000000",
  51312=>"010010110",
  51313=>"000001010",
  51314=>"001111101",
  51315=>"001010110",
  51316=>"001100010",
  51317=>"011000011",
  51318=>"110111100",
  51319=>"010011011",
  51320=>"000100111",
  51321=>"110101001",
  51322=>"110011001",
  51323=>"000111000",
  51324=>"100000101",
  51325=>"001010100",
  51326=>"100010100",
  51327=>"001111000",
  51328=>"010000100",
  51329=>"001010101",
  51330=>"010000010",
  51331=>"010001001",
  51332=>"110000100",
  51333=>"100001110",
  51334=>"111011001",
  51335=>"010100010",
  51336=>"001011100",
  51337=>"111111101",
  51338=>"101000001",
  51339=>"010101011",
  51340=>"001001011",
  51341=>"101100011",
  51342=>"000110000",
  51343=>"110011001",
  51344=>"000101100",
  51345=>"010010111",
  51346=>"011111100",
  51347=>"101000101",
  51348=>"101100000",
  51349=>"001101110",
  51350=>"010101000",
  51351=>"101011110",
  51352=>"001000100",
  51353=>"100010011",
  51354=>"000110000",
  51355=>"010010101",
  51356=>"100010110",
  51357=>"101010100",
  51358=>"010011101",
  51359=>"010010000",
  51360=>"111110110",
  51361=>"101100110",
  51362=>"110111011",
  51363=>"010101001",
  51364=>"110100001",
  51365=>"101110111",
  51366=>"111101110",
  51367=>"101110010",
  51368=>"101001011",
  51369=>"011011001",
  51370=>"100011101",
  51371=>"110001010",
  51372=>"111101011",
  51373=>"110100010",
  51374=>"100000110",
  51375=>"110110110",
  51376=>"010011000",
  51377=>"001000100",
  51378=>"100011001",
  51379=>"110110011",
  51380=>"110000100",
  51381=>"101001010",
  51382=>"001011000",
  51383=>"001001001",
  51384=>"100011000",
  51385=>"110100001",
  51386=>"011000000",
  51387=>"011111011",
  51388=>"001101100",
  51389=>"011110100",
  51390=>"010110111",
  51391=>"011101001",
  51392=>"111000100",
  51393=>"001000110",
  51394=>"000110101",
  51395=>"011011011",
  51396=>"011111100",
  51397=>"101100101",
  51398=>"011101111",
  51399=>"011000110",
  51400=>"110110011",
  51401=>"010010110",
  51402=>"101111011",
  51403=>"111110101",
  51404=>"000110010",
  51405=>"010101010",
  51406=>"000010000",
  51407=>"101010101",
  51408=>"111011101",
  51409=>"111010001",
  51410=>"100010101",
  51411=>"110111001",
  51412=>"001001001",
  51413=>"011001100",
  51414=>"101110010",
  51415=>"000101111",
  51416=>"010101000",
  51417=>"001101011",
  51418=>"010111110",
  51419=>"001000000",
  51420=>"001001101",
  51421=>"101011101",
  51422=>"000010111",
  51423=>"001100111",
  51424=>"101101000",
  51425=>"000000010",
  51426=>"111000101",
  51427=>"010101011",
  51428=>"001100111",
  51429=>"101101111",
  51430=>"111010001",
  51431=>"011111111",
  51432=>"011100100",
  51433=>"011000111",
  51434=>"000001000",
  51435=>"110111110",
  51436=>"110100101",
  51437=>"010011011",
  51438=>"110110001",
  51439=>"011000111",
  51440=>"111001110",
  51441=>"011011000",
  51442=>"011010101",
  51443=>"011010111",
  51444=>"010010011",
  51445=>"010011001",
  51446=>"010000101",
  51447=>"101110100",
  51448=>"011111101",
  51449=>"101011100",
  51450=>"111111100",
  51451=>"000000101",
  51452=>"010010110",
  51453=>"100100000",
  51454=>"010111000",
  51455=>"000011011",
  51456=>"110001100",
  51457=>"000010110",
  51458=>"010000000",
  51459=>"000001010",
  51460=>"000001101",
  51461=>"110001001",
  51462=>"010001100",
  51463=>"011111000",
  51464=>"011110110",
  51465=>"111011000",
  51466=>"010101001",
  51467=>"001000100",
  51468=>"000111000",
  51469=>"011000110",
  51470=>"110111000",
  51471=>"101100110",
  51472=>"010010101",
  51473=>"100010101",
  51474=>"110000000",
  51475=>"001110010",
  51476=>"000101000",
  51477=>"010001010",
  51478=>"100000001",
  51479=>"101111011",
  51480=>"111000001",
  51481=>"010000101",
  51482=>"110010101",
  51483=>"011011111",
  51484=>"101011111",
  51485=>"100100101",
  51486=>"001100101",
  51487=>"001110001",
  51488=>"010010010",
  51489=>"001101101",
  51490=>"010001111",
  51491=>"101111111",
  51492=>"110101010",
  51493=>"110110001",
  51494=>"110011000",
  51495=>"101011111",
  51496=>"101000100",
  51497=>"000100101",
  51498=>"100101110",
  51499=>"010101011",
  51500=>"111100010",
  51501=>"111100000",
  51502=>"110000000",
  51503=>"010100000",
  51504=>"101110111",
  51505=>"101011000",
  51506=>"010111010",
  51507=>"001010011",
  51508=>"001010010",
  51509=>"001011010",
  51510=>"010000001",
  51511=>"001010101",
  51512=>"001100000",
  51513=>"111111101",
  51514=>"001010111",
  51515=>"100100100",
  51516=>"010001101",
  51517=>"011100101",
  51518=>"101001010",
  51519=>"110010111",
  51520=>"011010101",
  51521=>"001000100",
  51522=>"110110001",
  51523=>"111000100",
  51524=>"001001011",
  51525=>"001001100",
  51526=>"000100010",
  51527=>"000001000",
  51528=>"001000101",
  51529=>"000101000",
  51530=>"011010000",
  51531=>"111100101",
  51532=>"011100101",
  51533=>"101101111",
  51534=>"011110000",
  51535=>"111011111",
  51536=>"001110110",
  51537=>"101011100",
  51538=>"011100001",
  51539=>"111011011",
  51540=>"110101100",
  51541=>"000101011",
  51542=>"011011101",
  51543=>"110110010",
  51544=>"100100001",
  51545=>"100111110",
  51546=>"010011001",
  51547=>"100101010",
  51548=>"100011100",
  51549=>"011101110",
  51550=>"101010000",
  51551=>"110110000",
  51552=>"110100111",
  51553=>"010100001",
  51554=>"001100111",
  51555=>"011001100",
  51556=>"110101111",
  51557=>"001110000",
  51558=>"110111111",
  51559=>"100101110",
  51560=>"101000001",
  51561=>"011111000",
  51562=>"101111110",
  51563=>"111110111",
  51564=>"100111011",
  51565=>"100011110",
  51566=>"101100101",
  51567=>"111111100",
  51568=>"110000010",
  51569=>"111010101",
  51570=>"001011100",
  51571=>"001110111",
  51572=>"001001100",
  51573=>"000111010",
  51574=>"001001000",
  51575=>"100101000",
  51576=>"101011100",
  51577=>"011111000",
  51578=>"001101010",
  51579=>"100000100",
  51580=>"010111001",
  51581=>"011100110",
  51582=>"010010111",
  51583=>"101111101",
  51584=>"100100000",
  51585=>"011000010",
  51586=>"111011010",
  51587=>"011101000",
  51588=>"001000111",
  51589=>"101100110",
  51590=>"011010011",
  51591=>"011010000",
  51592=>"100101001",
  51593=>"011110000",
  51594=>"101111000",
  51595=>"001101010",
  51596=>"000000100",
  51597=>"011000010",
  51598=>"100111010",
  51599=>"101001110",
  51600=>"001110011",
  51601=>"110110001",
  51602=>"101100101",
  51603=>"100001101",
  51604=>"100000110",
  51605=>"110111101",
  51606=>"100110111",
  51607=>"111110010",
  51608=>"110111110",
  51609=>"101000001",
  51610=>"101111101",
  51611=>"101011000",
  51612=>"000111010",
  51613=>"000000011",
  51614=>"100100101",
  51615=>"010100111",
  51616=>"101100110",
  51617=>"001010000",
  51618=>"001001101",
  51619=>"110100100",
  51620=>"101100101",
  51621=>"110100111",
  51622=>"010010101",
  51623=>"010100000",
  51624=>"101101111",
  51625=>"110010101",
  51626=>"110000101",
  51627=>"111000010",
  51628=>"100001111",
  51629=>"001111000",
  51630=>"010101110",
  51631=>"110010001",
  51632=>"000001001",
  51633=>"101011000",
  51634=>"011111110",
  51635=>"101000110",
  51636=>"100001000",
  51637=>"111111000",
  51638=>"011110001",
  51639=>"101111010",
  51640=>"110010101",
  51641=>"010010011",
  51642=>"000010001",
  51643=>"001001100",
  51644=>"101000010",
  51645=>"101111101",
  51646=>"101100111",
  51647=>"000100011",
  51648=>"111001010",
  51649=>"100001100",
  51650=>"000100001",
  51651=>"010101001",
  51652=>"000001010",
  51653=>"111111110",
  51654=>"110001000",
  51655=>"100001110",
  51656=>"110111100",
  51657=>"001001001",
  51658=>"011000111",
  51659=>"111001001",
  51660=>"011100101",
  51661=>"001110100",
  51662=>"101001000",
  51663=>"010110100",
  51664=>"011100110",
  51665=>"010001001",
  51666=>"100001000",
  51667=>"101001010",
  51668=>"111110001",
  51669=>"101100101",
  51670=>"010100000",
  51671=>"101110011",
  51672=>"111010101",
  51673=>"011001010",
  51674=>"101000100",
  51675=>"011101100",
  51676=>"000100110",
  51677=>"010110100",
  51678=>"011001111",
  51679=>"111100010",
  51680=>"101111110",
  51681=>"000010111",
  51682=>"010000100",
  51683=>"010101011",
  51684=>"010111000",
  51685=>"101001001",
  51686=>"100011011",
  51687=>"101010100",
  51688=>"010001001",
  51689=>"110111110",
  51690=>"010100110",
  51691=>"110000110",
  51692=>"011011010",
  51693=>"010001001",
  51694=>"100000010",
  51695=>"111011111",
  51696=>"000110010",
  51697=>"110111110",
  51698=>"100011111",
  51699=>"111010001",
  51700=>"011100110",
  51701=>"100100000",
  51702=>"101110010",
  51703=>"101010001",
  51704=>"001110010",
  51705=>"011110001",
  51706=>"111000000",
  51707=>"101111000",
  51708=>"011111100",
  51709=>"110111101",
  51710=>"100001110",
  51711=>"001000000",
  51712=>"011011000",
  51713=>"010001111",
  51714=>"001101100",
  51715=>"000011010",
  51716=>"000111110",
  51717=>"001010000",
  51718=>"101000011",
  51719=>"011001011",
  51720=>"010101100",
  51721=>"101001101",
  51722=>"110110000",
  51723=>"011100000",
  51724=>"011010000",
  51725=>"001000010",
  51726=>"100111011",
  51727=>"111001001",
  51728=>"111011011",
  51729=>"001011111",
  51730=>"100000000",
  51731=>"101010000",
  51732=>"011010101",
  51733=>"101001111",
  51734=>"010011000",
  51735=>"101110010",
  51736=>"111011000",
  51737=>"001101011",
  51738=>"101000000",
  51739=>"010100011",
  51740=>"010010010",
  51741=>"000100111",
  51742=>"000000000",
  51743=>"010011001",
  51744=>"001111000",
  51745=>"001001110",
  51746=>"010101111",
  51747=>"111100111",
  51748=>"010001110",
  51749=>"001011000",
  51750=>"111100101",
  51751=>"110100001",
  51752=>"000010100",
  51753=>"111100010",
  51754=>"111011110",
  51755=>"111100101",
  51756=>"001010110",
  51757=>"110001011",
  51758=>"100101011",
  51759=>"100010110",
  51760=>"011111100",
  51761=>"101011011",
  51762=>"001011011",
  51763=>"110000111",
  51764=>"011000011",
  51765=>"100100010",
  51766=>"000100000",
  51767=>"110001011",
  51768=>"011000101",
  51769=>"010110011",
  51770=>"001111110",
  51771=>"001010011",
  51772=>"000111101",
  51773=>"000011000",
  51774=>"110101110",
  51775=>"011011000",
  51776=>"011011101",
  51777=>"101101011",
  51778=>"111110011",
  51779=>"000101001",
  51780=>"001110000",
  51781=>"100101001",
  51782=>"000010011",
  51783=>"010100111",
  51784=>"110011010",
  51785=>"110001101",
  51786=>"110010110",
  51787=>"100000111",
  51788=>"011110100",
  51789=>"010100010",
  51790=>"001000011",
  51791=>"101111110",
  51792=>"000011100",
  51793=>"000011001",
  51794=>"110101111",
  51795=>"010011100",
  51796=>"001100101",
  51797=>"000011000",
  51798=>"001011100",
  51799=>"010011011",
  51800=>"000101101",
  51801=>"111100101",
  51802=>"010101001",
  51803=>"100000111",
  51804=>"000100100",
  51805=>"110100000",
  51806=>"101100110",
  51807=>"111100011",
  51808=>"011111000",
  51809=>"100000011",
  51810=>"101100000",
  51811=>"000001100",
  51812=>"111101110",
  51813=>"011100000",
  51814=>"110100101",
  51815=>"010000011",
  51816=>"001011000",
  51817=>"011000100",
  51818=>"000010011",
  51819=>"111110101",
  51820=>"000000011",
  51821=>"011010100",
  51822=>"001100100",
  51823=>"110010101",
  51824=>"101000110",
  51825=>"010001100",
  51826=>"010001111",
  51827=>"101000010",
  51828=>"110110000",
  51829=>"000001001",
  51830=>"011101001",
  51831=>"101010110",
  51832=>"101101110",
  51833=>"100101000",
  51834=>"010101000",
  51835=>"000111010",
  51836=>"101000111",
  51837=>"111001110",
  51838=>"000000001",
  51839=>"000001111",
  51840=>"000100101",
  51841=>"100101111",
  51842=>"000100001",
  51843=>"100101000",
  51844=>"011001100",
  51845=>"101100000",
  51846=>"010010101",
  51847=>"001110011",
  51848=>"000001000",
  51849=>"000010111",
  51850=>"001011111",
  51851=>"001001110",
  51852=>"000000000",
  51853=>"011100000",
  51854=>"000100010",
  51855=>"010000101",
  51856=>"011010001",
  51857=>"110100101",
  51858=>"011010100",
  51859=>"111010101",
  51860=>"100010010",
  51861=>"010011100",
  51862=>"101100010",
  51863=>"111101001",
  51864=>"011000000",
  51865=>"111010111",
  51866=>"010010101",
  51867=>"110111011",
  51868=>"100110001",
  51869=>"010100100",
  51870=>"001000011",
  51871=>"001011011",
  51872=>"101001101",
  51873=>"100011101",
  51874=>"101101011",
  51875=>"011111110",
  51876=>"111011111",
  51877=>"001000011",
  51878=>"100110010",
  51879=>"100100000",
  51880=>"000010011",
  51881=>"001000111",
  51882=>"110111111",
  51883=>"010001100",
  51884=>"000010100",
  51885=>"100100111",
  51886=>"101111001",
  51887=>"110001000",
  51888=>"110010001",
  51889=>"001010011",
  51890=>"111011011",
  51891=>"101010000",
  51892=>"111111111",
  51893=>"100001100",
  51894=>"010000100",
  51895=>"000101111",
  51896=>"100011001",
  51897=>"001101100",
  51898=>"001111001",
  51899=>"100111111",
  51900=>"010000011",
  51901=>"110100010",
  51902=>"110110100",
  51903=>"000010010",
  51904=>"000011011",
  51905=>"101101000",
  51906=>"111000110",
  51907=>"110010011",
  51908=>"011111110",
  51909=>"011110000",
  51910=>"100110100",
  51911=>"110110011",
  51912=>"001000010",
  51913=>"100001010",
  51914=>"011110010",
  51915=>"001101100",
  51916=>"101110100",
  51917=>"010110111",
  51918=>"111101101",
  51919=>"001001010",
  51920=>"110011001",
  51921=>"101101001",
  51922=>"111100010",
  51923=>"000101101",
  51924=>"110100010",
  51925=>"001010010",
  51926=>"000100111",
  51927=>"111001001",
  51928=>"101111001",
  51929=>"000110000",
  51930=>"100011000",
  51931=>"011000101",
  51932=>"101100101",
  51933=>"001111100",
  51934=>"111110010",
  51935=>"111100100",
  51936=>"110000110",
  51937=>"110000000",
  51938=>"111001111",
  51939=>"100101101",
  51940=>"001011110",
  51941=>"011001100",
  51942=>"011000000",
  51943=>"000101111",
  51944=>"100111111",
  51945=>"010000000",
  51946=>"111011100",
  51947=>"001010011",
  51948=>"001000010",
  51949=>"000110011",
  51950=>"011010100",
  51951=>"001101000",
  51952=>"010110011",
  51953=>"001100100",
  51954=>"100101110",
  51955=>"101110110",
  51956=>"011101011",
  51957=>"110010010",
  51958=>"000011110",
  51959=>"111111010",
  51960=>"010111110",
  51961=>"010001101",
  51962=>"010100100",
  51963=>"100101100",
  51964=>"001101011",
  51965=>"111011100",
  51966=>"110101100",
  51967=>"111101100",
  51968=>"000001101",
  51969=>"010100101",
  51970=>"000110000",
  51971=>"100001001",
  51972=>"001111010",
  51973=>"010101010",
  51974=>"011111110",
  51975=>"101011011",
  51976=>"110011101",
  51977=>"001010000",
  51978=>"000011100",
  51979=>"101001100",
  51980=>"101100011",
  51981=>"100000010",
  51982=>"111100111",
  51983=>"010110101",
  51984=>"110100010",
  51985=>"110100011",
  51986=>"111010010",
  51987=>"000101100",
  51988=>"001111111",
  51989=>"001000100",
  51990=>"010011111",
  51991=>"111010000",
  51992=>"011010010",
  51993=>"010100101",
  51994=>"011000000",
  51995=>"000000010",
  51996=>"000000010",
  51997=>"010000101",
  51998=>"000010101",
  51999=>"000011101",
  52000=>"101100011",
  52001=>"001110111",
  52002=>"001001010",
  52003=>"111001100",
  52004=>"001111000",
  52005=>"001110111",
  52006=>"011111001",
  52007=>"000000010",
  52008=>"110111101",
  52009=>"110100100",
  52010=>"100110100",
  52011=>"100111111",
  52012=>"110010101",
  52013=>"111010011",
  52014=>"110000010",
  52015=>"100101000",
  52016=>"101001101",
  52017=>"101110110",
  52018=>"100001001",
  52019=>"100010000",
  52020=>"010101000",
  52021=>"111111011",
  52022=>"100100110",
  52023=>"110010011",
  52024=>"010100001",
  52025=>"111100110",
  52026=>"111101010",
  52027=>"001011000",
  52028=>"111001010",
  52029=>"011010011",
  52030=>"100101110",
  52031=>"100110010",
  52032=>"000111101",
  52033=>"101011010",
  52034=>"111000101",
  52035=>"111101011",
  52036=>"001100010",
  52037=>"010001000",
  52038=>"001111011",
  52039=>"011100100",
  52040=>"111011010",
  52041=>"111111011",
  52042=>"010000100",
  52043=>"110011110",
  52044=>"110110101",
  52045=>"010110010",
  52046=>"111010010",
  52047=>"010100001",
  52048=>"010111011",
  52049=>"001110011",
  52050=>"000011110",
  52051=>"010011111",
  52052=>"011001101",
  52053=>"011110001",
  52054=>"000011100",
  52055=>"011011110",
  52056=>"110011011",
  52057=>"011100000",
  52058=>"101110111",
  52059=>"111101111",
  52060=>"100100000",
  52061=>"101111010",
  52062=>"011000010",
  52063=>"110000110",
  52064=>"101011101",
  52065=>"111110100",
  52066=>"100001010",
  52067=>"010110011",
  52068=>"010101101",
  52069=>"110000111",
  52070=>"111100001",
  52071=>"001010111",
  52072=>"001000001",
  52073=>"101110111",
  52074=>"011100111",
  52075=>"100111001",
  52076=>"110110010",
  52077=>"001001001",
  52078=>"010111001",
  52079=>"011101010",
  52080=>"011111010",
  52081=>"111100000",
  52082=>"100011011",
  52083=>"111101000",
  52084=>"000000100",
  52085=>"000001111",
  52086=>"010010101",
  52087=>"001100111",
  52088=>"011000000",
  52089=>"010101000",
  52090=>"101011000",
  52091=>"000101111",
  52092=>"000000100",
  52093=>"111001111",
  52094=>"011110111",
  52095=>"111111101",
  52096=>"101011111",
  52097=>"101010001",
  52098=>"111110000",
  52099=>"001101101",
  52100=>"010001110",
  52101=>"110100000",
  52102=>"000010000",
  52103=>"001110010",
  52104=>"111001100",
  52105=>"000000111",
  52106=>"101001000",
  52107=>"100000011",
  52108=>"100010110",
  52109=>"100101011",
  52110=>"000110001",
  52111=>"000110111",
  52112=>"101001110",
  52113=>"100000010",
  52114=>"110000010",
  52115=>"110111111",
  52116=>"111101101",
  52117=>"011000110",
  52118=>"000011100",
  52119=>"010110000",
  52120=>"011111100",
  52121=>"000101100",
  52122=>"111011100",
  52123=>"011010011",
  52124=>"000111101",
  52125=>"101011100",
  52126=>"001101011",
  52127=>"000001010",
  52128=>"110100100",
  52129=>"001011001",
  52130=>"111011101",
  52131=>"001001100",
  52132=>"010100000",
  52133=>"010111101",
  52134=>"011000011",
  52135=>"111111001",
  52136=>"010010111",
  52137=>"101110011",
  52138=>"100110011",
  52139=>"111010100",
  52140=>"101110000",
  52141=>"110000111",
  52142=>"101100010",
  52143=>"011001000",
  52144=>"101100101",
  52145=>"101110011",
  52146=>"110001110",
  52147=>"100011111",
  52148=>"010001011",
  52149=>"100100001",
  52150=>"100111100",
  52151=>"011000110",
  52152=>"000101001",
  52153=>"000101010",
  52154=>"011111111",
  52155=>"110011110",
  52156=>"001000000",
  52157=>"000010101",
  52158=>"010010110",
  52159=>"010000101",
  52160=>"001100101",
  52161=>"010110001",
  52162=>"111110100",
  52163=>"001101110",
  52164=>"110110110",
  52165=>"100110010",
  52166=>"100000000",
  52167=>"010001001",
  52168=>"000001110",
  52169=>"101100001",
  52170=>"011110101",
  52171=>"001000110",
  52172=>"111110110",
  52173=>"010111001",
  52174=>"101111110",
  52175=>"010111110",
  52176=>"111110010",
  52177=>"000110100",
  52178=>"001110100",
  52179=>"110100001",
  52180=>"101001111",
  52181=>"000010011",
  52182=>"111001111",
  52183=>"101100011",
  52184=>"100110100",
  52185=>"100101111",
  52186=>"011000000",
  52187=>"001000011",
  52188=>"101000001",
  52189=>"001000111",
  52190=>"111001000",
  52191=>"101000011",
  52192=>"100010111",
  52193=>"100100010",
  52194=>"000011000",
  52195=>"100110111",
  52196=>"000101100",
  52197=>"010010101",
  52198=>"111100001",
  52199=>"101000100",
  52200=>"100000001",
  52201=>"110111011",
  52202=>"111001010",
  52203=>"100110111",
  52204=>"101111100",
  52205=>"001111101",
  52206=>"000101000",
  52207=>"110000011",
  52208=>"000011000",
  52209=>"101000101",
  52210=>"001101111",
  52211=>"011001010",
  52212=>"101011100",
  52213=>"011101111",
  52214=>"010011101",
  52215=>"000101100",
  52216=>"100000100",
  52217=>"111101000",
  52218=>"110001111",
  52219=>"110110010",
  52220=>"001000011",
  52221=>"111011101",
  52222=>"101011010",
  52223=>"011100010",
  52224=>"110111011",
  52225=>"011001001",
  52226=>"010001010",
  52227=>"101101111",
  52228=>"111000000",
  52229=>"001110110",
  52230=>"110101101",
  52231=>"110011111",
  52232=>"100101110",
  52233=>"000100000",
  52234=>"001011111",
  52235=>"000010111",
  52236=>"000101100",
  52237=>"000100000",
  52238=>"111001001",
  52239=>"110011010",
  52240=>"111111000",
  52241=>"100110010",
  52242=>"101000000",
  52243=>"001101000",
  52244=>"111000101",
  52245=>"110001101",
  52246=>"010111111",
  52247=>"010111011",
  52248=>"000000000",
  52249=>"001010000",
  52250=>"011110100",
  52251=>"001000000",
  52252=>"101010101",
  52253=>"011001010",
  52254=>"010000010",
  52255=>"111010111",
  52256=>"000000110",
  52257=>"011100111",
  52258=>"001010011",
  52259=>"010011111",
  52260=>"111011001",
  52261=>"111001100",
  52262=>"001011100",
  52263=>"010000111",
  52264=>"000010100",
  52265=>"001100110",
  52266=>"000101110",
  52267=>"111110011",
  52268=>"001011101",
  52269=>"010101010",
  52270=>"011010010",
  52271=>"111111010",
  52272=>"011000111",
  52273=>"100100111",
  52274=>"000010000",
  52275=>"010011001",
  52276=>"111001111",
  52277=>"111011111",
  52278=>"100000011",
  52279=>"011101011",
  52280=>"001111100",
  52281=>"111101110",
  52282=>"111011000",
  52283=>"000001101",
  52284=>"011100001",
  52285=>"010111111",
  52286=>"100110001",
  52287=>"101011000",
  52288=>"000010100",
  52289=>"010001000",
  52290=>"111010000",
  52291=>"001111111",
  52292=>"011001101",
  52293=>"110011110",
  52294=>"001001000",
  52295=>"110010001",
  52296=>"000100101",
  52297=>"101011111",
  52298=>"111010100",
  52299=>"001110100",
  52300=>"100010001",
  52301=>"101110100",
  52302=>"100000010",
  52303=>"010010000",
  52304=>"111101001",
  52305=>"010011101",
  52306=>"001000100",
  52307=>"010111000",
  52308=>"110000011",
  52309=>"111101110",
  52310=>"001011100",
  52311=>"001100110",
  52312=>"111110010",
  52313=>"001000111",
  52314=>"000111001",
  52315=>"111010110",
  52316=>"011000001",
  52317=>"100010001",
  52318=>"111111111",
  52319=>"100001101",
  52320=>"100011010",
  52321=>"101101001",
  52322=>"010110100",
  52323=>"101000001",
  52324=>"111010001",
  52325=>"011110111",
  52326=>"110001101",
  52327=>"100110001",
  52328=>"001100100",
  52329=>"110111110",
  52330=>"111000110",
  52331=>"100010011",
  52332=>"100110001",
  52333=>"001010100",
  52334=>"110100110",
  52335=>"010000100",
  52336=>"001001001",
  52337=>"110111000",
  52338=>"000111101",
  52339=>"001000110",
  52340=>"111111110",
  52341=>"111000110",
  52342=>"010010101",
  52343=>"001001000",
  52344=>"100001101",
  52345=>"011001001",
  52346=>"101000010",
  52347=>"100010000",
  52348=>"011011000",
  52349=>"100101101",
  52350=>"100000010",
  52351=>"101011011",
  52352=>"011111110",
  52353=>"000111110",
  52354=>"001100001",
  52355=>"110000010",
  52356=>"001001000",
  52357=>"110111111",
  52358=>"101111110",
  52359=>"011011110",
  52360=>"000111111",
  52361=>"000010000",
  52362=>"000001100",
  52363=>"100111111",
  52364=>"100000110",
  52365=>"101011011",
  52366=>"110000010",
  52367=>"011000011",
  52368=>"110101000",
  52369=>"001100101",
  52370=>"010000000",
  52371=>"000110011",
  52372=>"100001111",
  52373=>"011101011",
  52374=>"010100010",
  52375=>"000010001",
  52376=>"110000000",
  52377=>"111110101",
  52378=>"000101100",
  52379=>"101111111",
  52380=>"101010111",
  52381=>"000101110",
  52382=>"100000111",
  52383=>"001101110",
  52384=>"110100110",
  52385=>"101100110",
  52386=>"001100000",
  52387=>"100011101",
  52388=>"111110101",
  52389=>"101000011",
  52390=>"000011000",
  52391=>"010000011",
  52392=>"000101111",
  52393=>"111110111",
  52394=>"000101100",
  52395=>"011010010",
  52396=>"001110100",
  52397=>"110101101",
  52398=>"101111111",
  52399=>"001100101",
  52400=>"101111110",
  52401=>"010000111",
  52402=>"010011101",
  52403=>"010010010",
  52404=>"010001101",
  52405=>"001011000",
  52406=>"011001010",
  52407=>"101100110",
  52408=>"111010111",
  52409=>"111110101",
  52410=>"010001001",
  52411=>"101010110",
  52412=>"010110011",
  52413=>"110011100",
  52414=>"000011000",
  52415=>"100101110",
  52416=>"000111001",
  52417=>"101000001",
  52418=>"000010000",
  52419=>"001010000",
  52420=>"011111010",
  52421=>"001001001",
  52422=>"100101110",
  52423=>"111011000",
  52424=>"110011101",
  52425=>"000010000",
  52426=>"000111101",
  52427=>"010110110",
  52428=>"000111001",
  52429=>"010110100",
  52430=>"111101011",
  52431=>"111101001",
  52432=>"001001101",
  52433=>"101011011",
  52434=>"111100011",
  52435=>"101100101",
  52436=>"000100110",
  52437=>"001011001",
  52438=>"101001101",
  52439=>"100101100",
  52440=>"010001110",
  52441=>"010100011",
  52442=>"001001010",
  52443=>"010100101",
  52444=>"000100100",
  52445=>"010101100",
  52446=>"110110010",
  52447=>"110011001",
  52448=>"100001110",
  52449=>"000110101",
  52450=>"110101011",
  52451=>"101110010",
  52452=>"100111100",
  52453=>"011111011",
  52454=>"000111100",
  52455=>"010000101",
  52456=>"000000001",
  52457=>"111111010",
  52458=>"111011000",
  52459=>"100111001",
  52460=>"011000010",
  52461=>"101010000",
  52462=>"010111111",
  52463=>"011000100",
  52464=>"011000010",
  52465=>"111101111",
  52466=>"100000010",
  52467=>"111010111",
  52468=>"000110000",
  52469=>"101001010",
  52470=>"100111100",
  52471=>"110010110",
  52472=>"110111010",
  52473=>"001111111",
  52474=>"101001100",
  52475=>"001011110",
  52476=>"100110101",
  52477=>"100011001",
  52478=>"111011001",
  52479=>"100011010",
  52480=>"011101011",
  52481=>"011100000",
  52482=>"100001101",
  52483=>"101000001",
  52484=>"110111010",
  52485=>"111010101",
  52486=>"101000101",
  52487=>"101001001",
  52488=>"000000011",
  52489=>"110001101",
  52490=>"111010011",
  52491=>"101010001",
  52492=>"100110110",
  52493=>"011110111",
  52494=>"101111000",
  52495=>"110001111",
  52496=>"111011110",
  52497=>"101101111",
  52498=>"101111001",
  52499=>"001100100",
  52500=>"111010000",
  52501=>"100110111",
  52502=>"010110110",
  52503=>"101101101",
  52504=>"101001101",
  52505=>"111111111",
  52506=>"100001111",
  52507=>"010110011",
  52508=>"111000110",
  52509=>"001111111",
  52510=>"001011000",
  52511=>"111100000",
  52512=>"111101110",
  52513=>"100111101",
  52514=>"011001011",
  52515=>"100100100",
  52516=>"111011101",
  52517=>"011101100",
  52518=>"010011001",
  52519=>"001001110",
  52520=>"000000000",
  52521=>"011010011",
  52522=>"100110101",
  52523=>"010010001",
  52524=>"101100010",
  52525=>"100110101",
  52526=>"111110100",
  52527=>"011010110",
  52528=>"010100110",
  52529=>"001100110",
  52530=>"110011111",
  52531=>"110000010",
  52532=>"100111001",
  52533=>"000111101",
  52534=>"111110100",
  52535=>"110100000",
  52536=>"111101111",
  52537=>"111001110",
  52538=>"001101101",
  52539=>"000111110",
  52540=>"111001010",
  52541=>"011110110",
  52542=>"001111001",
  52543=>"000011001",
  52544=>"100100101",
  52545=>"010011010",
  52546=>"000101011",
  52547=>"110110001",
  52548=>"011010100",
  52549=>"011011110",
  52550=>"010011000",
  52551=>"001011111",
  52552=>"011101100",
  52553=>"011001010",
  52554=>"011100001",
  52555=>"111110100",
  52556=>"010100111",
  52557=>"000101100",
  52558=>"011001100",
  52559=>"001111101",
  52560=>"010101000",
  52561=>"001000000",
  52562=>"100000101",
  52563=>"000111010",
  52564=>"110110000",
  52565=>"011111110",
  52566=>"001010001",
  52567=>"001110101",
  52568=>"010001011",
  52569=>"110101001",
  52570=>"110000110",
  52571=>"111111001",
  52572=>"001100110",
  52573=>"111100110",
  52574=>"101000100",
  52575=>"100000111",
  52576=>"110100000",
  52577=>"010111010",
  52578=>"010111000",
  52579=>"000011111",
  52580=>"100110001",
  52581=>"011101000",
  52582=>"110110101",
  52583=>"111000101",
  52584=>"010100111",
  52585=>"011110110",
  52586=>"100111100",
  52587=>"101001001",
  52588=>"110000001",
  52589=>"010010000",
  52590=>"101001100",
  52591=>"000100011",
  52592=>"011001010",
  52593=>"000111011",
  52594=>"010000001",
  52595=>"110111001",
  52596=>"000101101",
  52597=>"100001111",
  52598=>"011110100",
  52599=>"110111100",
  52600=>"010111111",
  52601=>"100010101",
  52602=>"001001010",
  52603=>"110010111",
  52604=>"000100100",
  52605=>"101101101",
  52606=>"110001010",
  52607=>"100001001",
  52608=>"010010001",
  52609=>"010011010",
  52610=>"101010010",
  52611=>"100100000",
  52612=>"111101101",
  52613=>"010101110",
  52614=>"110110010",
  52615=>"111011101",
  52616=>"110100011",
  52617=>"000010110",
  52618=>"110010001",
  52619=>"101110110",
  52620=>"000000011",
  52621=>"000001001",
  52622=>"000000110",
  52623=>"001011110",
  52624=>"101100010",
  52625=>"000111011",
  52626=>"111110001",
  52627=>"010011011",
  52628=>"111111011",
  52629=>"011000110",
  52630=>"111101110",
  52631=>"000111010",
  52632=>"100101001",
  52633=>"010111101",
  52634=>"010111001",
  52635=>"100001011",
  52636=>"000111000",
  52637=>"101011110",
  52638=>"111011110",
  52639=>"001001011",
  52640=>"000100010",
  52641=>"001010110",
  52642=>"001111111",
  52643=>"011111010",
  52644=>"100100110",
  52645=>"001010111",
  52646=>"110100000",
  52647=>"011101110",
  52648=>"001000100",
  52649=>"101111110",
  52650=>"001000110",
  52651=>"110010111",
  52652=>"000000110",
  52653=>"010100000",
  52654=>"000100101",
  52655=>"011110001",
  52656=>"111110010",
  52657=>"011101011",
  52658=>"001011101",
  52659=>"111001010",
  52660=>"101001110",
  52661=>"101100110",
  52662=>"001000100",
  52663=>"010110000",
  52664=>"100111010",
  52665=>"101010100",
  52666=>"001111101",
  52667=>"011101101",
  52668=>"011100011",
  52669=>"110011010",
  52670=>"010111001",
  52671=>"100010111",
  52672=>"000001000",
  52673=>"111100010",
  52674=>"000011000",
  52675=>"011001001",
  52676=>"100000000",
  52677=>"101101011",
  52678=>"110101100",
  52679=>"110001000",
  52680=>"000000011",
  52681=>"010010110",
  52682=>"001010000",
  52683=>"100101111",
  52684=>"011110010",
  52685=>"001111001",
  52686=>"010100110",
  52687=>"001000101",
  52688=>"011010101",
  52689=>"111111111",
  52690=>"110000101",
  52691=>"110110000",
  52692=>"011010000",
  52693=>"101101101",
  52694=>"011111000",
  52695=>"111000100",
  52696=>"001001110",
  52697=>"010110010",
  52698=>"110011100",
  52699=>"000101010",
  52700=>"000011011",
  52701=>"111111000",
  52702=>"001000010",
  52703=>"100101000",
  52704=>"011011110",
  52705=>"101001111",
  52706=>"001110010",
  52707=>"111011011",
  52708=>"111010111",
  52709=>"111111001",
  52710=>"110000010",
  52711=>"010101000",
  52712=>"010000110",
  52713=>"001010110",
  52714=>"111111100",
  52715=>"101000000",
  52716=>"110100011",
  52717=>"101000010",
  52718=>"110100100",
  52719=>"011100111",
  52720=>"100111011",
  52721=>"111010100",
  52722=>"111010010",
  52723=>"100101110",
  52724=>"100000101",
  52725=>"000110110",
  52726=>"101101101",
  52727=>"001001101",
  52728=>"110110010",
  52729=>"011100101",
  52730=>"000001111",
  52731=>"110110111",
  52732=>"000010011",
  52733=>"011111100",
  52734=>"000111000",
  52735=>"001001111",
  52736=>"111000110",
  52737=>"010000010",
  52738=>"010111101",
  52739=>"010101001",
  52740=>"011101001",
  52741=>"111111111",
  52742=>"000000110",
  52743=>"010000000",
  52744=>"101110000",
  52745=>"101111000",
  52746=>"011001100",
  52747=>"010001100",
  52748=>"001011010",
  52749=>"000010001",
  52750=>"101000111",
  52751=>"111110100",
  52752=>"000110010",
  52753=>"010010000",
  52754=>"110001000",
  52755=>"011100111",
  52756=>"001011100",
  52757=>"010000011",
  52758=>"001111100",
  52759=>"010110010",
  52760=>"000010100",
  52761=>"100011000",
  52762=>"010010011",
  52763=>"111100011",
  52764=>"001100011",
  52765=>"100110010",
  52766=>"000011101",
  52767=>"011110111",
  52768=>"011001001",
  52769=>"100100100",
  52770=>"000001100",
  52771=>"001111011",
  52772=>"011101000",
  52773=>"111100001",
  52774=>"100101010",
  52775=>"111001010",
  52776=>"011010001",
  52777=>"001001011",
  52778=>"011011001",
  52779=>"001100011",
  52780=>"111000101",
  52781=>"110110001",
  52782=>"101010001",
  52783=>"110000010",
  52784=>"111000000",
  52785=>"011010001",
  52786=>"000110001",
  52787=>"010001000",
  52788=>"010111000",
  52789=>"000100000",
  52790=>"100101100",
  52791=>"101010110",
  52792=>"010010011",
  52793=>"101111000",
  52794=>"100001111",
  52795=>"110101100",
  52796=>"110000100",
  52797=>"001100001",
  52798=>"110010000",
  52799=>"001101101",
  52800=>"000111011",
  52801=>"111001111",
  52802=>"001100110",
  52803=>"011011011",
  52804=>"110011011",
  52805=>"000111111",
  52806=>"101010110",
  52807=>"100111100",
  52808=>"111100100",
  52809=>"110011100",
  52810=>"001001111",
  52811=>"001000000",
  52812=>"011011001",
  52813=>"101000000",
  52814=>"001110010",
  52815=>"111011110",
  52816=>"110111011",
  52817=>"010010011",
  52818=>"000010111",
  52819=>"000100010",
  52820=>"110000010",
  52821=>"001010001",
  52822=>"101110101",
  52823=>"001011111",
  52824=>"111111111",
  52825=>"101001110",
  52826=>"011111101",
  52827=>"000100001",
  52828=>"110100010",
  52829=>"110011000",
  52830=>"011010011",
  52831=>"100010011",
  52832=>"111010000",
  52833=>"011100100",
  52834=>"010001111",
  52835=>"100010110",
  52836=>"000111000",
  52837=>"101000001",
  52838=>"110000110",
  52839=>"111111000",
  52840=>"101001110",
  52841=>"001111010",
  52842=>"101000000",
  52843=>"100000101",
  52844=>"111010010",
  52845=>"111100111",
  52846=>"011111010",
  52847=>"110000111",
  52848=>"010000001",
  52849=>"100000110",
  52850=>"100111101",
  52851=>"101100011",
  52852=>"100110111",
  52853=>"000101111",
  52854=>"110100001",
  52855=>"100011101",
  52856=>"101110001",
  52857=>"101100111",
  52858=>"101110100",
  52859=>"011001100",
  52860=>"001100000",
  52861=>"100001000",
  52862=>"110100001",
  52863=>"010111111",
  52864=>"110110011",
  52865=>"101001101",
  52866=>"111101010",
  52867=>"100100101",
  52868=>"011100100",
  52869=>"010111111",
  52870=>"111010001",
  52871=>"100000111",
  52872=>"101001000",
  52873=>"000001010",
  52874=>"101011111",
  52875=>"110111011",
  52876=>"010000000",
  52877=>"000110001",
  52878=>"101100110",
  52879=>"010010100",
  52880=>"010101111",
  52881=>"100101010",
  52882=>"010101100",
  52883=>"001000110",
  52884=>"100100010",
  52885=>"001000101",
  52886=>"001101010",
  52887=>"001110000",
  52888=>"101101110",
  52889=>"000110101",
  52890=>"111101101",
  52891=>"001111011",
  52892=>"110001010",
  52893=>"010100000",
  52894=>"000011101",
  52895=>"011010010",
  52896=>"000001100",
  52897=>"111010101",
  52898=>"000101001",
  52899=>"110011001",
  52900=>"011110010",
  52901=>"101111100",
  52902=>"111010110",
  52903=>"000000011",
  52904=>"100011110",
  52905=>"101100010",
  52906=>"010100000",
  52907=>"000100011",
  52908=>"000001110",
  52909=>"001111111",
  52910=>"011110111",
  52911=>"011110000",
  52912=>"110101100",
  52913=>"110010011",
  52914=>"000100100",
  52915=>"101000011",
  52916=>"101001101",
  52917=>"110111010",
  52918=>"101101111",
  52919=>"001001000",
  52920=>"111110101",
  52921=>"000011111",
  52922=>"111111011",
  52923=>"010011111",
  52924=>"101111011",
  52925=>"111100001",
  52926=>"000011010",
  52927=>"110011100",
  52928=>"101000011",
  52929=>"001000101",
  52930=>"001101000",
  52931=>"000111001",
  52932=>"101111110",
  52933=>"111101110",
  52934=>"100111110",
  52935=>"001011111",
  52936=>"000110011",
  52937=>"011001110",
  52938=>"000100001",
  52939=>"100010110",
  52940=>"000111001",
  52941=>"011111100",
  52942=>"100111000",
  52943=>"111011001",
  52944=>"011110010",
  52945=>"010000000",
  52946=>"001000001",
  52947=>"000001101",
  52948=>"010010011",
  52949=>"101100010",
  52950=>"100001000",
  52951=>"101111110",
  52952=>"101010011",
  52953=>"100110011",
  52954=>"010010001",
  52955=>"111000010",
  52956=>"001110011",
  52957=>"001000010",
  52958=>"101110101",
  52959=>"100111111",
  52960=>"101111000",
  52961=>"101000100",
  52962=>"111000101",
  52963=>"001001111",
  52964=>"101100100",
  52965=>"100010101",
  52966=>"111100100",
  52967=>"100010111",
  52968=>"000010100",
  52969=>"010110010",
  52970=>"111100110",
  52971=>"001001011",
  52972=>"111111001",
  52973=>"110100110",
  52974=>"111101110",
  52975=>"010000001",
  52976=>"010110110",
  52977=>"110110011",
  52978=>"110111001",
  52979=>"010010010",
  52980=>"100110011",
  52981=>"100011011",
  52982=>"100100111",
  52983=>"000101001",
  52984=>"000111001",
  52985=>"100101010",
  52986=>"010001101",
  52987=>"011110011",
  52988=>"001010110",
  52989=>"010001100",
  52990=>"011100110",
  52991=>"100100110",
  52992=>"011111100",
  52993=>"101011111",
  52994=>"001111100",
  52995=>"010001001",
  52996=>"111111010",
  52997=>"111110011",
  52998=>"100011110",
  52999=>"010010011",
  53000=>"001100110",
  53001=>"010010100",
  53002=>"001110010",
  53003=>"001011101",
  53004=>"111000111",
  53005=>"001010100",
  53006=>"010001010",
  53007=>"011010100",
  53008=>"111011101",
  53009=>"110110010",
  53010=>"011100001",
  53011=>"010000001",
  53012=>"100010110",
  53013=>"010010000",
  53014=>"000000010",
  53015=>"011010101",
  53016=>"110100000",
  53017=>"010001000",
  53018=>"110101011",
  53019=>"100111010",
  53020=>"010011100",
  53021=>"011100111",
  53022=>"110111100",
  53023=>"100000110",
  53024=>"100111011",
  53025=>"111100001",
  53026=>"111011011",
  53027=>"001111100",
  53028=>"001000111",
  53029=>"110100010",
  53030=>"101111010",
  53031=>"101011111",
  53032=>"001101010",
  53033=>"101101110",
  53034=>"000101000",
  53035=>"010001110",
  53036=>"000010010",
  53037=>"110001011",
  53038=>"100000001",
  53039=>"010010010",
  53040=>"111111011",
  53041=>"000001000",
  53042=>"011100001",
  53043=>"011001011",
  53044=>"111111111",
  53045=>"100110000",
  53046=>"101110000",
  53047=>"101101111",
  53048=>"100110111",
  53049=>"110011100",
  53050=>"100101111",
  53051=>"100001011",
  53052=>"100100001",
  53053=>"101110010",
  53054=>"111100010",
  53055=>"001110110",
  53056=>"111111110",
  53057=>"111110111",
  53058=>"100000100",
  53059=>"110010111",
  53060=>"000110111",
  53061=>"001101001",
  53062=>"101111001",
  53063=>"111011011",
  53064=>"100100010",
  53065=>"101111010",
  53066=>"111000000",
  53067=>"011000000",
  53068=>"110010000",
  53069=>"111001001",
  53070=>"011111101",
  53071=>"110101010",
  53072=>"111010001",
  53073=>"100001001",
  53074=>"110101100",
  53075=>"110100010",
  53076=>"110010001",
  53077=>"000010010",
  53078=>"011100100",
  53079=>"010011001",
  53080=>"110110100",
  53081=>"100010000",
  53082=>"011001000",
  53083=>"000100010",
  53084=>"010101110",
  53085=>"000010011",
  53086=>"111010100",
  53087=>"100110001",
  53088=>"101001010",
  53089=>"100001101",
  53090=>"001110011",
  53091=>"010111010",
  53092=>"000110110",
  53093=>"111000110",
  53094=>"111111010",
  53095=>"101101111",
  53096=>"001010001",
  53097=>"100100111",
  53098=>"001111001",
  53099=>"000111111",
  53100=>"100010111",
  53101=>"101100010",
  53102=>"000100001",
  53103=>"101101111",
  53104=>"001101010",
  53105=>"000000000",
  53106=>"101100010",
  53107=>"000100000",
  53108=>"010000101",
  53109=>"110110001",
  53110=>"000100100",
  53111=>"011000111",
  53112=>"000001010",
  53113=>"101011100",
  53114=>"010100110",
  53115=>"101110010",
  53116=>"111000110",
  53117=>"001001101",
  53118=>"110010111",
  53119=>"111000010",
  53120=>"001000011",
  53121=>"110111111",
  53122=>"010011110",
  53123=>"011010001",
  53124=>"111110111",
  53125=>"111010001",
  53126=>"000000000",
  53127=>"110100101",
  53128=>"111100010",
  53129=>"100010101",
  53130=>"101101010",
  53131=>"100101010",
  53132=>"101110011",
  53133=>"101000000",
  53134=>"000100000",
  53135=>"101000101",
  53136=>"100010100",
  53137=>"101111111",
  53138=>"010011011",
  53139=>"010010100",
  53140=>"111001101",
  53141=>"111000000",
  53142=>"010101001",
  53143=>"001101000",
  53144=>"100010110",
  53145=>"011100000",
  53146=>"001111000",
  53147=>"000000000",
  53148=>"001000010",
  53149=>"011111111",
  53150=>"111100000",
  53151=>"001111100",
  53152=>"100010000",
  53153=>"001101011",
  53154=>"001010010",
  53155=>"101100111",
  53156=>"100100100",
  53157=>"000100001",
  53158=>"110101000",
  53159=>"010000011",
  53160=>"100000010",
  53161=>"101000111",
  53162=>"000111010",
  53163=>"000110111",
  53164=>"100001011",
  53165=>"000111100",
  53166=>"100000000",
  53167=>"100000100",
  53168=>"001110011",
  53169=>"110011001",
  53170=>"110100011",
  53171=>"000101000",
  53172=>"000001000",
  53173=>"011110001",
  53174=>"110110101",
  53175=>"010001100",
  53176=>"010010111",
  53177=>"111010000",
  53178=>"100001110",
  53179=>"110101001",
  53180=>"000110100",
  53181=>"001001001",
  53182=>"011000111",
  53183=>"111000101",
  53184=>"011000101",
  53185=>"010001101",
  53186=>"010110100",
  53187=>"100100100",
  53188=>"101011110",
  53189=>"010110110",
  53190=>"000010000",
  53191=>"101000001",
  53192=>"111110000",
  53193=>"001001111",
  53194=>"000101000",
  53195=>"110001100",
  53196=>"101111000",
  53197=>"001000010",
  53198=>"101011010",
  53199=>"000101001",
  53200=>"110100000",
  53201=>"010100001",
  53202=>"011000101",
  53203=>"101011110",
  53204=>"100010001",
  53205=>"000011101",
  53206=>"001111101",
  53207=>"011111111",
  53208=>"011100110",
  53209=>"000000010",
  53210=>"110000001",
  53211=>"011101100",
  53212=>"101011110",
  53213=>"100001111",
  53214=>"101100001",
  53215=>"011011111",
  53216=>"111101100",
  53217=>"111101000",
  53218=>"010010111",
  53219=>"101000110",
  53220=>"110101000",
  53221=>"010111010",
  53222=>"010011011",
  53223=>"011001110",
  53224=>"100111011",
  53225=>"011100001",
  53226=>"111110100",
  53227=>"000010110",
  53228=>"101101101",
  53229=>"000000110",
  53230=>"011011101",
  53231=>"000001001",
  53232=>"001011110",
  53233=>"101011101",
  53234=>"111000110",
  53235=>"011110111",
  53236=>"111100101",
  53237=>"000111110",
  53238=>"100010110",
  53239=>"111100011",
  53240=>"000010010",
  53241=>"010011110",
  53242=>"111110110",
  53243=>"010001101",
  53244=>"111010010",
  53245=>"011001000",
  53246=>"001000010",
  53247=>"001110100",
  53248=>"110111110",
  53249=>"111110101",
  53250=>"010110110",
  53251=>"100011010",
  53252=>"101011110",
  53253=>"111010101",
  53254=>"100010110",
  53255=>"001010110",
  53256=>"010001010",
  53257=>"001101001",
  53258=>"101101111",
  53259=>"111110011",
  53260=>"011100101",
  53261=>"101011010",
  53262=>"110111010",
  53263=>"111001001",
  53264=>"110100010",
  53265=>"101100010",
  53266=>"101110100",
  53267=>"111010110",
  53268=>"101011100",
  53269=>"011011101",
  53270=>"000110011",
  53271=>"001001101",
  53272=>"110111001",
  53273=>"000000010",
  53274=>"011001111",
  53275=>"100010000",
  53276=>"000110110",
  53277=>"011001111",
  53278=>"100100101",
  53279=>"101110011",
  53280=>"000110110",
  53281=>"010001101",
  53282=>"101101100",
  53283=>"100011100",
  53284=>"000111100",
  53285=>"001101111",
  53286=>"001100011",
  53287=>"111011001",
  53288=>"011110011",
  53289=>"101110100",
  53290=>"110000111",
  53291=>"010001011",
  53292=>"100001110",
  53293=>"101111101",
  53294=>"100010100",
  53295=>"001010000",
  53296=>"010110101",
  53297=>"010100010",
  53298=>"000000000",
  53299=>"101110000",
  53300=>"000000100",
  53301=>"001010000",
  53302=>"110000111",
  53303=>"100110000",
  53304=>"001101101",
  53305=>"101001010",
  53306=>"000011010",
  53307=>"101100001",
  53308=>"001010001",
  53309=>"001011001",
  53310=>"001100011",
  53311=>"001100100",
  53312=>"110011010",
  53313=>"010001001",
  53314=>"111010010",
  53315=>"001000101",
  53316=>"011101000",
  53317=>"010000000",
  53318=>"001000110",
  53319=>"001011001",
  53320=>"111111011",
  53321=>"000000010",
  53322=>"010001000",
  53323=>"100000001",
  53324=>"011011001",
  53325=>"100110100",
  53326=>"111110000",
  53327=>"001010000",
  53328=>"110111001",
  53329=>"001100110",
  53330=>"100001110",
  53331=>"011111100",
  53332=>"100111001",
  53333=>"101111010",
  53334=>"011110101",
  53335=>"010001010",
  53336=>"101111100",
  53337=>"010110110",
  53338=>"001101010",
  53339=>"011000001",
  53340=>"000110011",
  53341=>"101101100",
  53342=>"000010101",
  53343=>"110000101",
  53344=>"111101000",
  53345=>"011000101",
  53346=>"110001111",
  53347=>"110101111",
  53348=>"001101011",
  53349=>"110001110",
  53350=>"111010111",
  53351=>"010101000",
  53352=>"110101100",
  53353=>"101110100",
  53354=>"011101010",
  53355=>"100101011",
  53356=>"110001100",
  53357=>"111111001",
  53358=>"111000000",
  53359=>"000101110",
  53360=>"000111000",
  53361=>"010011110",
  53362=>"010000001",
  53363=>"001010101",
  53364=>"010110111",
  53365=>"010111001",
  53366=>"001110111",
  53367=>"111100111",
  53368=>"011001111",
  53369=>"001100001",
  53370=>"010100110",
  53371=>"110111010",
  53372=>"000000101",
  53373=>"010110010",
  53374=>"000001111",
  53375=>"001110011",
  53376=>"111001111",
  53377=>"110001011",
  53378=>"110001010",
  53379=>"000100100",
  53380=>"011101011",
  53381=>"110010101",
  53382=>"101111000",
  53383=>"000110111",
  53384=>"001001110",
  53385=>"100000111",
  53386=>"100101000",
  53387=>"110010101",
  53388=>"011000010",
  53389=>"111111000",
  53390=>"100010000",
  53391=>"100011010",
  53392=>"101001100",
  53393=>"001100010",
  53394=>"000001010",
  53395=>"011110011",
  53396=>"011000001",
  53397=>"000000111",
  53398=>"000110011",
  53399=>"101001111",
  53400=>"111000111",
  53401=>"001110001",
  53402=>"011000001",
  53403=>"100101101",
  53404=>"001101101",
  53405=>"100010001",
  53406=>"001100100",
  53407=>"101101000",
  53408=>"111101011",
  53409=>"010111100",
  53410=>"110100010",
  53411=>"011110011",
  53412=>"110001110",
  53413=>"101000010",
  53414=>"100011011",
  53415=>"010110001",
  53416=>"100011101",
  53417=>"111010010",
  53418=>"001001100",
  53419=>"100001111",
  53420=>"000001100",
  53421=>"010100110",
  53422=>"001000100",
  53423=>"010100001",
  53424=>"001001000",
  53425=>"100010001",
  53426=>"010000010",
  53427=>"000100111",
  53428=>"111001011",
  53429=>"001011011",
  53430=>"011001100",
  53431=>"011011111",
  53432=>"011001000",
  53433=>"101101000",
  53434=>"000000011",
  53435=>"000010001",
  53436=>"100001011",
  53437=>"000000001",
  53438=>"010000011",
  53439=>"000100100",
  53440=>"110010011",
  53441=>"100101011",
  53442=>"000000110",
  53443=>"111000110",
  53444=>"101101110",
  53445=>"101111001",
  53446=>"011100110",
  53447=>"000001011",
  53448=>"111011101",
  53449=>"111011111",
  53450=>"100000110",
  53451=>"110011110",
  53452=>"111100000",
  53453=>"101000111",
  53454=>"010100000",
  53455=>"010100010",
  53456=>"101111100",
  53457=>"010101001",
  53458=>"001100000",
  53459=>"000010010",
  53460=>"000110110",
  53461=>"010010111",
  53462=>"111000010",
  53463=>"100000010",
  53464=>"000001111",
  53465=>"010100111",
  53466=>"111011011",
  53467=>"101100001",
  53468=>"011111011",
  53469=>"110000110",
  53470=>"010000101",
  53471=>"011011010",
  53472=>"000001100",
  53473=>"101101111",
  53474=>"010011110",
  53475=>"000011011",
  53476=>"010111010",
  53477=>"001111110",
  53478=>"100001010",
  53479=>"010011000",
  53480=>"111110111",
  53481=>"010100010",
  53482=>"101101101",
  53483=>"000111110",
  53484=>"110100000",
  53485=>"100000011",
  53486=>"111100101",
  53487=>"011010001",
  53488=>"011110010",
  53489=>"010111110",
  53490=>"100110111",
  53491=>"100000001",
  53492=>"100110110",
  53493=>"101010111",
  53494=>"111111000",
  53495=>"011101011",
  53496=>"111011011",
  53497=>"001001011",
  53498=>"101001101",
  53499=>"111011111",
  53500=>"010011001",
  53501=>"001101100",
  53502=>"101010001",
  53503=>"010011101",
  53504=>"110111101",
  53505=>"101110001",
  53506=>"010111001",
  53507=>"110010101",
  53508=>"111000001",
  53509=>"001000011",
  53510=>"010001011",
  53511=>"101000101",
  53512=>"001110111",
  53513=>"000011011",
  53514=>"011111110",
  53515=>"011111100",
  53516=>"111111111",
  53517=>"001101100",
  53518=>"110111011",
  53519=>"100010100",
  53520=>"011111110",
  53521=>"111010111",
  53522=>"011101111",
  53523=>"011101001",
  53524=>"010010010",
  53525=>"000010111",
  53526=>"011110101",
  53527=>"111011110",
  53528=>"010011100",
  53529=>"111000100",
  53530=>"011110000",
  53531=>"101000000",
  53532=>"111000110",
  53533=>"000000010",
  53534=>"100100100",
  53535=>"011110010",
  53536=>"001110011",
  53537=>"010011011",
  53538=>"100011100",
  53539=>"101010010",
  53540=>"000110001",
  53541=>"010100000",
  53542=>"101000101",
  53543=>"011000101",
  53544=>"110001010",
  53545=>"111011110",
  53546=>"111111011",
  53547=>"000101011",
  53548=>"111011110",
  53549=>"101110100",
  53550=>"001000010",
  53551=>"010001000",
  53552=>"000010010",
  53553=>"100101100",
  53554=>"001000111",
  53555=>"010110100",
  53556=>"010000100",
  53557=>"000101000",
  53558=>"100101100",
  53559=>"000101110",
  53560=>"111011011",
  53561=>"000000011",
  53562=>"000011101",
  53563=>"010010110",
  53564=>"100000110",
  53565=>"001010011",
  53566=>"111101010",
  53567=>"011100110",
  53568=>"100100101",
  53569=>"111011011",
  53570=>"111100101",
  53571=>"101011011",
  53572=>"111101111",
  53573=>"010000000",
  53574=>"101110100",
  53575=>"001101111",
  53576=>"110000011",
  53577=>"011001001",
  53578=>"101111110",
  53579=>"001000000",
  53580=>"111001010",
  53581=>"101111010",
  53582=>"010001001",
  53583=>"110101110",
  53584=>"011110001",
  53585=>"000110110",
  53586=>"110001101",
  53587=>"010000011",
  53588=>"000000000",
  53589=>"101111111",
  53590=>"101111001",
  53591=>"000010101",
  53592=>"011010101",
  53593=>"101000111",
  53594=>"011100011",
  53595=>"100000000",
  53596=>"000010100",
  53597=>"110100000",
  53598=>"000000101",
  53599=>"111000100",
  53600=>"001101111",
  53601=>"001110100",
  53602=>"010101110",
  53603=>"100000101",
  53604=>"000101110",
  53605=>"101110111",
  53606=>"000001101",
  53607=>"010110010",
  53608=>"101000100",
  53609=>"011101100",
  53610=>"000010000",
  53611=>"011101101",
  53612=>"010000110",
  53613=>"101110000",
  53614=>"011001111",
  53615=>"000000100",
  53616=>"001101111",
  53617=>"001010101",
  53618=>"110110111",
  53619=>"100000000",
  53620=>"100010011",
  53621=>"110010001",
  53622=>"101010100",
  53623=>"000111001",
  53624=>"001000000",
  53625=>"010110000",
  53626=>"010101111",
  53627=>"011010000",
  53628=>"101100000",
  53629=>"110100010",
  53630=>"111101011",
  53631=>"111100101",
  53632=>"000011111",
  53633=>"010110100",
  53634=>"111101000",
  53635=>"011010001",
  53636=>"101100010",
  53637=>"000001000",
  53638=>"010001101",
  53639=>"001100110",
  53640=>"010001101",
  53641=>"110111000",
  53642=>"000101101",
  53643=>"111010011",
  53644=>"110001001",
  53645=>"001000110",
  53646=>"010010011",
  53647=>"100000000",
  53648=>"000011001",
  53649=>"001001000",
  53650=>"111000010",
  53651=>"001100001",
  53652=>"110110011",
  53653=>"001100110",
  53654=>"111001000",
  53655=>"001000001",
  53656=>"101110101",
  53657=>"100000011",
  53658=>"010001010",
  53659=>"010001101",
  53660=>"010011001",
  53661=>"101110111",
  53662=>"010101000",
  53663=>"100110110",
  53664=>"000011000",
  53665=>"100101011",
  53666=>"100000011",
  53667=>"010010111",
  53668=>"100011010",
  53669=>"110111100",
  53670=>"011110000",
  53671=>"100010110",
  53672=>"110010111",
  53673=>"001000000",
  53674=>"011011000",
  53675=>"100010001",
  53676=>"010010111",
  53677=>"110111000",
  53678=>"101101000",
  53679=>"011011111",
  53680=>"111101001",
  53681=>"001100001",
  53682=>"100011110",
  53683=>"010111010",
  53684=>"010111111",
  53685=>"011101000",
  53686=>"001100001",
  53687=>"111110110",
  53688=>"011111010",
  53689=>"010001000",
  53690=>"110110001",
  53691=>"101100100",
  53692=>"001111110",
  53693=>"101110001",
  53694=>"011001100",
  53695=>"000001110",
  53696=>"110100001",
  53697=>"100011010",
  53698=>"010010011",
  53699=>"111000001",
  53700=>"000000011",
  53701=>"010010101",
  53702=>"001100001",
  53703=>"111101111",
  53704=>"010110000",
  53705=>"110010011",
  53706=>"100010010",
  53707=>"011111011",
  53708=>"001011000",
  53709=>"101111001",
  53710=>"101010000",
  53711=>"111111111",
  53712=>"001101011",
  53713=>"010010110",
  53714=>"011010100",
  53715=>"101000110",
  53716=>"101101101",
  53717=>"000001000",
  53718=>"011001010",
  53719=>"111111110",
  53720=>"100010000",
  53721=>"001101110",
  53722=>"100111101",
  53723=>"100111000",
  53724=>"010111011",
  53725=>"101001010",
  53726=>"110101101",
  53727=>"011110000",
  53728=>"111110010",
  53729=>"110111001",
  53730=>"011101101",
  53731=>"001101110",
  53732=>"110011001",
  53733=>"111111111",
  53734=>"010101110",
  53735=>"101001010",
  53736=>"101010010",
  53737=>"000110110",
  53738=>"000101100",
  53739=>"001100101",
  53740=>"010101010",
  53741=>"011000000",
  53742=>"010001001",
  53743=>"100000100",
  53744=>"010011000",
  53745=>"010110100",
  53746=>"100010100",
  53747=>"001000011",
  53748=>"010101010",
  53749=>"011010101",
  53750=>"110110000",
  53751=>"010010001",
  53752=>"100000111",
  53753=>"101101011",
  53754=>"010100000",
  53755=>"101001100",
  53756=>"001000000",
  53757=>"000101000",
  53758=>"010101111",
  53759=>"010011000",
  53760=>"000100101",
  53761=>"101110001",
  53762=>"111100010",
  53763=>"011001000",
  53764=>"010001100",
  53765=>"101111000",
  53766=>"111101110",
  53767=>"110111010",
  53768=>"000000000",
  53769=>"111101110",
  53770=>"011000101",
  53771=>"011110001",
  53772=>"001100101",
  53773=>"111100000",
  53774=>"011100111",
  53775=>"101010101",
  53776=>"001111110",
  53777=>"011010110",
  53778=>"100111100",
  53779=>"110111010",
  53780=>"000011010",
  53781=>"111000101",
  53782=>"010010101",
  53783=>"011110011",
  53784=>"011000010",
  53785=>"000000011",
  53786=>"001011011",
  53787=>"010010101",
  53788=>"000010001",
  53789=>"111001101",
  53790=>"000110011",
  53791=>"010011001",
  53792=>"110101011",
  53793=>"010101001",
  53794=>"011101001",
  53795=>"001000001",
  53796=>"001110011",
  53797=>"010111011",
  53798=>"010101101",
  53799=>"001100110",
  53800=>"111100100",
  53801=>"111111111",
  53802=>"001100101",
  53803=>"000010010",
  53804=>"100100101",
  53805=>"001000001",
  53806=>"100000110",
  53807=>"110011111",
  53808=>"100110001",
  53809=>"111110100",
  53810=>"001001001",
  53811=>"101100110",
  53812=>"000011001",
  53813=>"001001111",
  53814=>"010011001",
  53815=>"100111111",
  53816=>"110101101",
  53817=>"110010110",
  53818=>"001000111",
  53819=>"100111011",
  53820=>"100101111",
  53821=>"011110011",
  53822=>"000001101",
  53823=>"101000000",
  53824=>"001000011",
  53825=>"000110011",
  53826=>"111000010",
  53827=>"001110001",
  53828=>"101001010",
  53829=>"010100010",
  53830=>"000101001",
  53831=>"011001110",
  53832=>"001100010",
  53833=>"000110011",
  53834=>"010100011",
  53835=>"101011111",
  53836=>"101000101",
  53837=>"111111000",
  53838=>"000001101",
  53839=>"101111101",
  53840=>"110111110",
  53841=>"010001001",
  53842=>"000100110",
  53843=>"000001110",
  53844=>"011100011",
  53845=>"011010100",
  53846=>"001010000",
  53847=>"010100000",
  53848=>"100010001",
  53849=>"101101111",
  53850=>"110000111",
  53851=>"101000011",
  53852=>"011001101",
  53853=>"110011001",
  53854=>"101001010",
  53855=>"011000001",
  53856=>"011101011",
  53857=>"001010001",
  53858=>"000010011",
  53859=>"010011000",
  53860=>"111001001",
  53861=>"110101111",
  53862=>"011100001",
  53863=>"100001011",
  53864=>"110110000",
  53865=>"100101001",
  53866=>"001010010",
  53867=>"011011011",
  53868=>"011110101",
  53869=>"110001000",
  53870=>"001010010",
  53871=>"101000001",
  53872=>"010101001",
  53873=>"100101110",
  53874=>"010010101",
  53875=>"011010010",
  53876=>"010011000",
  53877=>"001101101",
  53878=>"000101001",
  53879=>"110000110",
  53880=>"000000000",
  53881=>"011001010",
  53882=>"100110111",
  53883=>"000010100",
  53884=>"011101100",
  53885=>"110110001",
  53886=>"101001010",
  53887=>"001110010",
  53888=>"001110011",
  53889=>"010000001",
  53890=>"100001000",
  53891=>"001100000",
  53892=>"101110101",
  53893=>"101000011",
  53894=>"011001000",
  53895=>"111110101",
  53896=>"000100101",
  53897=>"011101100",
  53898=>"010000101",
  53899=>"110100100",
  53900=>"111001111",
  53901=>"000011110",
  53902=>"110111100",
  53903=>"100010110",
  53904=>"111010001",
  53905=>"010000011",
  53906=>"001000101",
  53907=>"000111111",
  53908=>"100000111",
  53909=>"001110100",
  53910=>"111001110",
  53911=>"100001010",
  53912=>"010010101",
  53913=>"110011011",
  53914=>"011100010",
  53915=>"111000000",
  53916=>"001101011",
  53917=>"010010100",
  53918=>"100000000",
  53919=>"101011010",
  53920=>"101101110",
  53921=>"000001100",
  53922=>"100101111",
  53923=>"000100011",
  53924=>"010111001",
  53925=>"000010110",
  53926=>"001100100",
  53927=>"100000001",
  53928=>"110110010",
  53929=>"011111000",
  53930=>"001100001",
  53931=>"010011010",
  53932=>"100101001",
  53933=>"001100100",
  53934=>"101010010",
  53935=>"001101010",
  53936=>"000110110",
  53937=>"100001100",
  53938=>"011000100",
  53939=>"000101101",
  53940=>"011011111",
  53941=>"010111010",
  53942=>"000000111",
  53943=>"110000011",
  53944=>"011000001",
  53945=>"110001011",
  53946=>"010000001",
  53947=>"001010000",
  53948=>"000001000",
  53949=>"101111011",
  53950=>"100101001",
  53951=>"011110110",
  53952=>"110111100",
  53953=>"011011000",
  53954=>"110110101",
  53955=>"101111000",
  53956=>"111100101",
  53957=>"001101001",
  53958=>"110110001",
  53959=>"100000010",
  53960=>"000000011",
  53961=>"111100111",
  53962=>"000111001",
  53963=>"001000010",
  53964=>"111111001",
  53965=>"110011110",
  53966=>"011101001",
  53967=>"010110101",
  53968=>"001001111",
  53969=>"000100110",
  53970=>"100010000",
  53971=>"010001101",
  53972=>"010000110",
  53973=>"100100001",
  53974=>"110110000",
  53975=>"111101010",
  53976=>"001101001",
  53977=>"111111101",
  53978=>"100100010",
  53979=>"010001001",
  53980=>"110011001",
  53981=>"101110010",
  53982=>"111001000",
  53983=>"100101101",
  53984=>"010000000",
  53985=>"001101101",
  53986=>"000101101",
  53987=>"100101011",
  53988=>"011100100",
  53989=>"110001100",
  53990=>"010100001",
  53991=>"100110001",
  53992=>"111000111",
  53993=>"110111111",
  53994=>"111110001",
  53995=>"010010010",
  53996=>"010001000",
  53997=>"110100111",
  53998=>"111001010",
  53999=>"000110000",
  54000=>"110001010",
  54001=>"001101110",
  54002=>"001110111",
  54003=>"010000100",
  54004=>"100111111",
  54005=>"001010000",
  54006=>"010100110",
  54007=>"101110011",
  54008=>"001000111",
  54009=>"000010101",
  54010=>"110110000",
  54011=>"111101000",
  54012=>"110000100",
  54013=>"110000000",
  54014=>"111000110",
  54015=>"101011011",
  54016=>"101111001",
  54017=>"000001100",
  54018=>"000000100",
  54019=>"001100000",
  54020=>"000100011",
  54021=>"001000110",
  54022=>"000110011",
  54023=>"100100101",
  54024=>"001000111",
  54025=>"110001011",
  54026=>"100010110",
  54027=>"110100001",
  54028=>"001101001",
  54029=>"110111111",
  54030=>"011110001",
  54031=>"111110001",
  54032=>"110100001",
  54033=>"011001111",
  54034=>"011111100",
  54035=>"011110101",
  54036=>"001101111",
  54037=>"101011010",
  54038=>"101001100",
  54039=>"101000000",
  54040=>"001010111",
  54041=>"000111110",
  54042=>"011100011",
  54043=>"110110010",
  54044=>"000010010",
  54045=>"010111000",
  54046=>"100110101",
  54047=>"000111110",
  54048=>"100011001",
  54049=>"011001111",
  54050=>"111100110",
  54051=>"100001111",
  54052=>"111010010",
  54053=>"100001011",
  54054=>"110000111",
  54055=>"010111110",
  54056=>"000110101",
  54057=>"101100111",
  54058=>"001010000",
  54059=>"100000000",
  54060=>"110111001",
  54061=>"000001101",
  54062=>"001011010",
  54063=>"000010101",
  54064=>"000100001",
  54065=>"101101011",
  54066=>"101011000",
  54067=>"101000010",
  54068=>"010001100",
  54069=>"000100100",
  54070=>"111000110",
  54071=>"101001010",
  54072=>"000001101",
  54073=>"100011110",
  54074=>"001000011",
  54075=>"110101001",
  54076=>"110110101",
  54077=>"000101101",
  54078=>"110000110",
  54079=>"001011001",
  54080=>"111101000",
  54081=>"111011100",
  54082=>"110110101",
  54083=>"000100101",
  54084=>"001001111",
  54085=>"101000000",
  54086=>"000000011",
  54087=>"110001011",
  54088=>"011001000",
  54089=>"110011001",
  54090=>"011010010",
  54091=>"001000111",
  54092=>"100100100",
  54093=>"000010111",
  54094=>"000001001",
  54095=>"101111011",
  54096=>"000011100",
  54097=>"000100011",
  54098=>"000000010",
  54099=>"011010001",
  54100=>"000010011",
  54101=>"000101011",
  54102=>"011011011",
  54103=>"100101111",
  54104=>"100001000",
  54105=>"101110100",
  54106=>"011100010",
  54107=>"101100111",
  54108=>"001001001",
  54109=>"110100110",
  54110=>"111010111",
  54111=>"000111011",
  54112=>"111011111",
  54113=>"011001001",
  54114=>"001101110",
  54115=>"110110111",
  54116=>"101110010",
  54117=>"001000001",
  54118=>"001011111",
  54119=>"001000111",
  54120=>"111001111",
  54121=>"001100001",
  54122=>"010111011",
  54123=>"110101001",
  54124=>"000000000",
  54125=>"010011001",
  54126=>"010000010",
  54127=>"100000111",
  54128=>"010101000",
  54129=>"111001100",
  54130=>"000000100",
  54131=>"011001010",
  54132=>"101011001",
  54133=>"100100110",
  54134=>"000110010",
  54135=>"011011111",
  54136=>"000010010",
  54137=>"111010001",
  54138=>"000100111",
  54139=>"001011011",
  54140=>"000000001",
  54141=>"011000010",
  54142=>"100010000",
  54143=>"110101110",
  54144=>"011011001",
  54145=>"000100110",
  54146=>"110101001",
  54147=>"010001011",
  54148=>"010000010",
  54149=>"110101101",
  54150=>"001110110",
  54151=>"111001101",
  54152=>"010100111",
  54153=>"110011110",
  54154=>"010101110",
  54155=>"100010110",
  54156=>"010000000",
  54157=>"011001011",
  54158=>"001010000",
  54159=>"101010110",
  54160=>"000000100",
  54161=>"010010100",
  54162=>"010011010",
  54163=>"101101001",
  54164=>"000110111",
  54165=>"110010111",
  54166=>"101001101",
  54167=>"000010001",
  54168=>"001000001",
  54169=>"011010111",
  54170=>"111010100",
  54171=>"000010011",
  54172=>"000001010",
  54173=>"010000000",
  54174=>"010000111",
  54175=>"011101001",
  54176=>"011111001",
  54177=>"000000011",
  54178=>"110111010",
  54179=>"000001001",
  54180=>"001101100",
  54181=>"010111111",
  54182=>"110110011",
  54183=>"011100100",
  54184=>"001101101",
  54185=>"001011010",
  54186=>"101101000",
  54187=>"010111101",
  54188=>"011101101",
  54189=>"101100110",
  54190=>"001011100",
  54191=>"010101000",
  54192=>"000010110",
  54193=>"100110011",
  54194=>"101101101",
  54195=>"111101001",
  54196=>"110101111",
  54197=>"111100101",
  54198=>"000110110",
  54199=>"111011100",
  54200=>"011010101",
  54201=>"101011101",
  54202=>"010110011",
  54203=>"101010110",
  54204=>"101101100",
  54205=>"101000010",
  54206=>"011110111",
  54207=>"011110011",
  54208=>"010011011",
  54209=>"101101000",
  54210=>"100101011",
  54211=>"001101111",
  54212=>"000101000",
  54213=>"111000111",
  54214=>"110010100",
  54215=>"101110001",
  54216=>"101000010",
  54217=>"010101111",
  54218=>"010001011",
  54219=>"100011000",
  54220=>"101111010",
  54221=>"101101010",
  54222=>"011001011",
  54223=>"010000000",
  54224=>"100101111",
  54225=>"001000111",
  54226=>"110010011",
  54227=>"110100001",
  54228=>"111101010",
  54229=>"101010100",
  54230=>"010100001",
  54231=>"001001110",
  54232=>"010000000",
  54233=>"001100101",
  54234=>"100010011",
  54235=>"001010101",
  54236=>"100110100",
  54237=>"111101011",
  54238=>"010100010",
  54239=>"000001010",
  54240=>"100000111",
  54241=>"100011110",
  54242=>"011000111",
  54243=>"001011110",
  54244=>"110011001",
  54245=>"010011000",
  54246=>"111011101",
  54247=>"111100010",
  54248=>"010100111",
  54249=>"111011110",
  54250=>"111100001",
  54251=>"100010101",
  54252=>"100000001",
  54253=>"010010100",
  54254=>"110111000",
  54255=>"111011011",
  54256=>"011001111",
  54257=>"100110101",
  54258=>"000101000",
  54259=>"010001000",
  54260=>"011110101",
  54261=>"010001011",
  54262=>"001000111",
  54263=>"011011110",
  54264=>"000000001",
  54265=>"010110111",
  54266=>"000101100",
  54267=>"001011111",
  54268=>"001111000",
  54269=>"000000001",
  54270=>"110101100",
  54271=>"100101100",
  54272=>"101101111",
  54273=>"011001101",
  54274=>"110100001",
  54275=>"101011100",
  54276=>"101011001",
  54277=>"101111111",
  54278=>"111000111",
  54279=>"100100001",
  54280=>"111100011",
  54281=>"000000010",
  54282=>"101010010",
  54283=>"001110100",
  54284=>"100101011",
  54285=>"010101101",
  54286=>"111000100",
  54287=>"001001011",
  54288=>"010100010",
  54289=>"001001111",
  54290=>"010110110",
  54291=>"100101101",
  54292=>"111000001",
  54293=>"100001111",
  54294=>"110011000",
  54295=>"000100000",
  54296=>"111001110",
  54297=>"001101000",
  54298=>"101101001",
  54299=>"010010111",
  54300=>"111111111",
  54301=>"010110001",
  54302=>"111111000",
  54303=>"000111001",
  54304=>"011101010",
  54305=>"011000010",
  54306=>"110000100",
  54307=>"100100000",
  54308=>"111111011",
  54309=>"011111101",
  54310=>"011010101",
  54311=>"010101111",
  54312=>"100110100",
  54313=>"110011010",
  54314=>"111111101",
  54315=>"011110100",
  54316=>"001010000",
  54317=>"011000000",
  54318=>"011010111",
  54319=>"000011010",
  54320=>"000010001",
  54321=>"001000100",
  54322=>"001100011",
  54323=>"011100011",
  54324=>"101100111",
  54325=>"100101100",
  54326=>"101111101",
  54327=>"100010110",
  54328=>"101010110",
  54329=>"101101101",
  54330=>"111110100",
  54331=>"010001011",
  54332=>"111100101",
  54333=>"011110100",
  54334=>"101100000",
  54335=>"000111000",
  54336=>"010000100",
  54337=>"000001100",
  54338=>"010010111",
  54339=>"010111000",
  54340=>"110100111",
  54341=>"111111100",
  54342=>"000110100",
  54343=>"101011001",
  54344=>"000011010",
  54345=>"110011110",
  54346=>"111011111",
  54347=>"001111101",
  54348=>"000000110",
  54349=>"010110011",
  54350=>"011011101",
  54351=>"101110001",
  54352=>"110100011",
  54353=>"000011110",
  54354=>"111010001",
  54355=>"010000000",
  54356=>"000101010",
  54357=>"010111100",
  54358=>"101111011",
  54359=>"000110110",
  54360=>"110101111",
  54361=>"101000011",
  54362=>"111110101",
  54363=>"010000010",
  54364=>"001001111",
  54365=>"111110100",
  54366=>"111011000",
  54367=>"111000000",
  54368=>"001001101",
  54369=>"010000010",
  54370=>"100110101",
  54371=>"100000100",
  54372=>"100110110",
  54373=>"000101010",
  54374=>"110101100",
  54375=>"101000101",
  54376=>"011111101",
  54377=>"011010100",
  54378=>"001010000",
  54379=>"000100110",
  54380=>"111101110",
  54381=>"001011111",
  54382=>"111100100",
  54383=>"110000001",
  54384=>"110101010",
  54385=>"101011011",
  54386=>"001101101",
  54387=>"010100101",
  54388=>"101000011",
  54389=>"001011000",
  54390=>"100001100",
  54391=>"010111101",
  54392=>"101111011",
  54393=>"010011100",
  54394=>"111110111",
  54395=>"000101000",
  54396=>"111101000",
  54397=>"010000010",
  54398=>"111100111",
  54399=>"001111111",
  54400=>"000011110",
  54401=>"000011100",
  54402=>"010000000",
  54403=>"011010000",
  54404=>"000001100",
  54405=>"001000110",
  54406=>"000000001",
  54407=>"110110000",
  54408=>"110010101",
  54409=>"111011101",
  54410=>"100000000",
  54411=>"100100000",
  54412=>"000010101",
  54413=>"011110001",
  54414=>"111110001",
  54415=>"110110000",
  54416=>"110001011",
  54417=>"001110001",
  54418=>"010000100",
  54419=>"110010001",
  54420=>"001101010",
  54421=>"111100110",
  54422=>"001000100",
  54423=>"000101001",
  54424=>"010100000",
  54425=>"100001011",
  54426=>"111111011",
  54427=>"111011110",
  54428=>"111111101",
  54429=>"011110011",
  54430=>"001110101",
  54431=>"010111001",
  54432=>"111111011",
  54433=>"110100011",
  54434=>"110101010",
  54435=>"000100111",
  54436=>"000110110",
  54437=>"110111111",
  54438=>"010011011",
  54439=>"101000101",
  54440=>"011110100",
  54441=>"011101111",
  54442=>"010110101",
  54443=>"101100011",
  54444=>"000001000",
  54445=>"010100000",
  54446=>"001011110",
  54447=>"010100111",
  54448=>"111100101",
  54449=>"001000101",
  54450=>"101000001",
  54451=>"000110101",
  54452=>"111000001",
  54453=>"011011010",
  54454=>"010000100",
  54455=>"011110110",
  54456=>"100000000",
  54457=>"001001000",
  54458=>"001000111",
  54459=>"011000100",
  54460=>"011011110",
  54461=>"111101011",
  54462=>"011100010",
  54463=>"001100011",
  54464=>"001100000",
  54465=>"001111100",
  54466=>"011001000",
  54467=>"111100010",
  54468=>"101100100",
  54469=>"110100000",
  54470=>"010000010",
  54471=>"000110110",
  54472=>"111111101",
  54473=>"010011101",
  54474=>"101011011",
  54475=>"001100001",
  54476=>"110001000",
  54477=>"001011111",
  54478=>"111101000",
  54479=>"100101110",
  54480=>"011101000",
  54481=>"000100010",
  54482=>"000001011",
  54483=>"101000111",
  54484=>"001111111",
  54485=>"111011001",
  54486=>"000010101",
  54487=>"111001111",
  54488=>"001010000",
  54489=>"000011111",
  54490=>"101000000",
  54491=>"000111111",
  54492=>"001110010",
  54493=>"001100001",
  54494=>"100110110",
  54495=>"101000101",
  54496=>"101100101",
  54497=>"011100011",
  54498=>"100110010",
  54499=>"110101000",
  54500=>"101100001",
  54501=>"110101111",
  54502=>"101010001",
  54503=>"001000011",
  54504=>"000001011",
  54505=>"001100000",
  54506=>"101000110",
  54507=>"010101101",
  54508=>"011010011",
  54509=>"001101100",
  54510=>"101100101",
  54511=>"111000110",
  54512=>"001111110",
  54513=>"110100001",
  54514=>"101111010",
  54515=>"010000010",
  54516=>"100100001",
  54517=>"100010001",
  54518=>"101011001",
  54519=>"101010110",
  54520=>"101111111",
  54521=>"111110111",
  54522=>"001101001",
  54523=>"000101010",
  54524=>"110010000",
  54525=>"010100110",
  54526=>"100111010",
  54527=>"100011001",
  54528=>"100101001",
  54529=>"101010101",
  54530=>"111101100",
  54531=>"110111101",
  54532=>"110110000",
  54533=>"010001100",
  54534=>"000110001",
  54535=>"110100001",
  54536=>"111101111",
  54537=>"000110111",
  54538=>"000000001",
  54539=>"000000111",
  54540=>"010000100",
  54541=>"000010110",
  54542=>"010000001",
  54543=>"001101100",
  54544=>"010000010",
  54545=>"111101011",
  54546=>"111111100",
  54547=>"111110100",
  54548=>"110100110",
  54549=>"011101001",
  54550=>"010001010",
  54551=>"111000011",
  54552=>"000100001",
  54553=>"111101101",
  54554=>"110000111",
  54555=>"010000101",
  54556=>"111110101",
  54557=>"001101000",
  54558=>"101011111",
  54559=>"000101101",
  54560=>"110010010",
  54561=>"000000010",
  54562=>"110011111",
  54563=>"001001101",
  54564=>"011110110",
  54565=>"000011001",
  54566=>"011100010",
  54567=>"000001101",
  54568=>"111101101",
  54569=>"001001100",
  54570=>"110011101",
  54571=>"111111001",
  54572=>"100011100",
  54573=>"000111111",
  54574=>"001001111",
  54575=>"010100010",
  54576=>"100010100",
  54577=>"000011101",
  54578=>"100110110",
  54579=>"100101010",
  54580=>"001010111",
  54581=>"110101110",
  54582=>"001000100",
  54583=>"110110000",
  54584=>"100011000",
  54585=>"000001010",
  54586=>"111100111",
  54587=>"001100111",
  54588=>"011111010",
  54589=>"101010100",
  54590=>"101110000",
  54591=>"110000001",
  54592=>"101101100",
  54593=>"101110101",
  54594=>"011100101",
  54595=>"011010110",
  54596=>"101010111",
  54597=>"010100110",
  54598=>"011000000",
  54599=>"101001101",
  54600=>"101100000",
  54601=>"010000000",
  54602=>"111000100",
  54603=>"110111001",
  54604=>"101001111",
  54605=>"100000000",
  54606=>"011010111",
  54607=>"001111111",
  54608=>"011101010",
  54609=>"010000010",
  54610=>"111011111",
  54611=>"111111000",
  54612=>"000000010",
  54613=>"100101000",
  54614=>"000110010",
  54615=>"011110101",
  54616=>"100001010",
  54617=>"000001001",
  54618=>"110000101",
  54619=>"101001111",
  54620=>"110100111",
  54621=>"010010010",
  54622=>"101101101",
  54623=>"100000110",
  54624=>"001001101",
  54625=>"111000110",
  54626=>"101101011",
  54627=>"011101100",
  54628=>"011000011",
  54629=>"111101000",
  54630=>"001011101",
  54631=>"100011110",
  54632=>"010001100",
  54633=>"100111110",
  54634=>"111101100",
  54635=>"101011001",
  54636=>"000110010",
  54637=>"101111000",
  54638=>"100101100",
  54639=>"011001111",
  54640=>"010010001",
  54641=>"110100000",
  54642=>"010000100",
  54643=>"100100101",
  54644=>"000000011",
  54645=>"001101001",
  54646=>"110100110",
  54647=>"011101011",
  54648=>"111001111",
  54649=>"000001011",
  54650=>"101011111",
  54651=>"110100010",
  54652=>"110111001",
  54653=>"111000001",
  54654=>"101100000",
  54655=>"001100111",
  54656=>"000011100",
  54657=>"101101000",
  54658=>"010110011",
  54659=>"000010010",
  54660=>"110111001",
  54661=>"100001011",
  54662=>"100010111",
  54663=>"001000000",
  54664=>"001000001",
  54665=>"111101100",
  54666=>"000000111",
  54667=>"110111000",
  54668=>"111011000",
  54669=>"001001000",
  54670=>"101100111",
  54671=>"001110100",
  54672=>"101001110",
  54673=>"100101101",
  54674=>"011101001",
  54675=>"001110011",
  54676=>"101110010",
  54677=>"010110101",
  54678=>"011001011",
  54679=>"010011111",
  54680=>"111010111",
  54681=>"000001011",
  54682=>"111100001",
  54683=>"000100000",
  54684=>"101100111",
  54685=>"000000010",
  54686=>"001001001",
  54687=>"100000110",
  54688=>"011110010",
  54689=>"000110100",
  54690=>"001000101",
  54691=>"001100110",
  54692=>"010010100",
  54693=>"100010000",
  54694=>"000011111",
  54695=>"010010001",
  54696=>"110110000",
  54697=>"101001111",
  54698=>"010011001",
  54699=>"010001100",
  54700=>"000100110",
  54701=>"001010010",
  54702=>"000010000",
  54703=>"011110011",
  54704=>"100100000",
  54705=>"110000000",
  54706=>"010110000",
  54707=>"010111110",
  54708=>"101101101",
  54709=>"000011111",
  54710=>"000001100",
  54711=>"110110110",
  54712=>"110111111",
  54713=>"100001010",
  54714=>"110000110",
  54715=>"001100111",
  54716=>"110001111",
  54717=>"000011110",
  54718=>"011010110",
  54719=>"100101110",
  54720=>"010001110",
  54721=>"111110100",
  54722=>"100000111",
  54723=>"011101011",
  54724=>"111000111",
  54725=>"001001111",
  54726=>"001110101",
  54727=>"011010101",
  54728=>"001111001",
  54729=>"001000100",
  54730=>"011000001",
  54731=>"100111110",
  54732=>"010011010",
  54733=>"011111001",
  54734=>"101000001",
  54735=>"110101001",
  54736=>"001011110",
  54737=>"011100111",
  54738=>"100110111",
  54739=>"101100111",
  54740=>"000010111",
  54741=>"100001111",
  54742=>"010000001",
  54743=>"110011100",
  54744=>"000000011",
  54745=>"100001000",
  54746=>"110000000",
  54747=>"010011111",
  54748=>"110011111",
  54749=>"000110010",
  54750=>"101100000",
  54751=>"001101010",
  54752=>"110000101",
  54753=>"101000100",
  54754=>"000010011",
  54755=>"010010100",
  54756=>"010011111",
  54757=>"110011010",
  54758=>"010000111",
  54759=>"111011001",
  54760=>"010011001",
  54761=>"100010000",
  54762=>"010011111",
  54763=>"001101101",
  54764=>"101000101",
  54765=>"010001111",
  54766=>"110010000",
  54767=>"001101100",
  54768=>"110110110",
  54769=>"111000010",
  54770=>"110011111",
  54771=>"000001110",
  54772=>"110001101",
  54773=>"100000000",
  54774=>"011101011",
  54775=>"111010010",
  54776=>"011110011",
  54777=>"001101100",
  54778=>"100100000",
  54779=>"111011110",
  54780=>"001011100",
  54781=>"111011010",
  54782=>"111101111",
  54783=>"111111010",
  54784=>"011010010",
  54785=>"111001011",
  54786=>"101010100",
  54787=>"110101111",
  54788=>"011010110",
  54789=>"111111011",
  54790=>"011000001",
  54791=>"000111111",
  54792=>"110100110",
  54793=>"010101001",
  54794=>"101011010",
  54795=>"110101000",
  54796=>"110010000",
  54797=>"011001010",
  54798=>"110100101",
  54799=>"111011011",
  54800=>"100101111",
  54801=>"010000001",
  54802=>"101101100",
  54803=>"110000011",
  54804=>"110100001",
  54805=>"111011011",
  54806=>"110001010",
  54807=>"011011111",
  54808=>"010001111",
  54809=>"111110111",
  54810=>"110000011",
  54811=>"100010111",
  54812=>"110100001",
  54813=>"110010111",
  54814=>"010000010",
  54815=>"111000111",
  54816=>"101111010",
  54817=>"000000001",
  54818=>"001111001",
  54819=>"011011100",
  54820=>"110011100",
  54821=>"011111101",
  54822=>"110100101",
  54823=>"000101001",
  54824=>"101100011",
  54825=>"000000100",
  54826=>"110101111",
  54827=>"000110110",
  54828=>"100100011",
  54829=>"001100011",
  54830=>"111101100",
  54831=>"010000000",
  54832=>"100011000",
  54833=>"101101001",
  54834=>"111100101",
  54835=>"101000111",
  54836=>"100101111",
  54837=>"010011101",
  54838=>"110000010",
  54839=>"001001111",
  54840=>"010000000",
  54841=>"011010101",
  54842=>"100011101",
  54843=>"011000011",
  54844=>"111001110",
  54845=>"100101001",
  54846=>"101011001",
  54847=>"111001001",
  54848=>"110011101",
  54849=>"110000110",
  54850=>"111110000",
  54851=>"100100001",
  54852=>"000111011",
  54853=>"111101010",
  54854=>"000111111",
  54855=>"010110011",
  54856=>"011100100",
  54857=>"010100111",
  54858=>"000000000",
  54859=>"011011110",
  54860=>"101110100",
  54861=>"011100011",
  54862=>"110110110",
  54863=>"001110011",
  54864=>"011011010",
  54865=>"001010000",
  54866=>"000010000",
  54867=>"100101011",
  54868=>"000101000",
  54869=>"111110101",
  54870=>"000000101",
  54871=>"100111110",
  54872=>"111111101",
  54873=>"111110101",
  54874=>"101111101",
  54875=>"011000110",
  54876=>"110101010",
  54877=>"011011000",
  54878=>"011111011",
  54879=>"101000010",
  54880=>"110001010",
  54881=>"100001010",
  54882=>"001101100",
  54883=>"111011100",
  54884=>"100111011",
  54885=>"001100000",
  54886=>"011010000",
  54887=>"010100011",
  54888=>"000101001",
  54889=>"001111101",
  54890=>"111111111",
  54891=>"011001110",
  54892=>"100011110",
  54893=>"100011011",
  54894=>"101000011",
  54895=>"100000001",
  54896=>"101111101",
  54897=>"101010000",
  54898=>"101000000",
  54899=>"111101011",
  54900=>"111010010",
  54901=>"100011000",
  54902=>"000000000",
  54903=>"110101001",
  54904=>"111101000",
  54905=>"111000110",
  54906=>"110011001",
  54907=>"011110000",
  54908=>"011100110",
  54909=>"111001111",
  54910=>"011111000",
  54911=>"011001010",
  54912=>"000101101",
  54913=>"110001010",
  54914=>"111001011",
  54915=>"100011000",
  54916=>"101011111",
  54917=>"010010000",
  54918=>"101000110",
  54919=>"111100001",
  54920=>"011101011",
  54921=>"111010111",
  54922=>"010000001",
  54923=>"011011110",
  54924=>"101001100",
  54925=>"000111100",
  54926=>"101000010",
  54927=>"110101011",
  54928=>"010011001",
  54929=>"100100011",
  54930=>"001110111",
  54931=>"010111100",
  54932=>"010001011",
  54933=>"001001111",
  54934=>"100000100",
  54935=>"010001001",
  54936=>"101111110",
  54937=>"010011000",
  54938=>"111101111",
  54939=>"110110100",
  54940=>"000101011",
  54941=>"001101011",
  54942=>"010011000",
  54943=>"001100100",
  54944=>"110011001",
  54945=>"110010001",
  54946=>"111111010",
  54947=>"011100010",
  54948=>"110010101",
  54949=>"110110000",
  54950=>"010011110",
  54951=>"010000001",
  54952=>"000000111",
  54953=>"001000110",
  54954=>"011111100",
  54955=>"010111101",
  54956=>"011110101",
  54957=>"010101110",
  54958=>"011010101",
  54959=>"000000000",
  54960=>"010111101",
  54961=>"011110001",
  54962=>"010111011",
  54963=>"110101001",
  54964=>"000000111",
  54965=>"000100001",
  54966=>"110110100",
  54967=>"111010110",
  54968=>"110110111",
  54969=>"010110001",
  54970=>"100001011",
  54971=>"000101000",
  54972=>"101101100",
  54973=>"101110100",
  54974=>"101010101",
  54975=>"000100111",
  54976=>"001100100",
  54977=>"110010011",
  54978=>"101110110",
  54979=>"010000101",
  54980=>"111111100",
  54981=>"000001011",
  54982=>"010100100",
  54983=>"111110010",
  54984=>"010011111",
  54985=>"001010001",
  54986=>"101010000",
  54987=>"111010110",
  54988=>"000010011",
  54989=>"100001101",
  54990=>"011001000",
  54991=>"001100111",
  54992=>"111101101",
  54993=>"100011000",
  54994=>"011101111",
  54995=>"100101000",
  54996=>"001011001",
  54997=>"111111101",
  54998=>"010101010",
  54999=>"110000000",
  55000=>"000000011",
  55001=>"111101001",
  55002=>"101011111",
  55003=>"011000110",
  55004=>"100010011",
  55005=>"110101110",
  55006=>"001110111",
  55007=>"110100110",
  55008=>"001000100",
  55009=>"010000111",
  55010=>"111010111",
  55011=>"111000000",
  55012=>"100000100",
  55013=>"000000011",
  55014=>"101000000",
  55015=>"111111010",
  55016=>"110110000",
  55017=>"000010100",
  55018=>"101011101",
  55019=>"101100100",
  55020=>"000100111",
  55021=>"001000101",
  55022=>"100111110",
  55023=>"110010010",
  55024=>"001000010",
  55025=>"111111110",
  55026=>"101100000",
  55027=>"110110001",
  55028=>"011110011",
  55029=>"111111111",
  55030=>"010101101",
  55031=>"001110001",
  55032=>"111001111",
  55033=>"110001110",
  55034=>"000101000",
  55035=>"011100100",
  55036=>"100010000",
  55037=>"011001110",
  55038=>"000100100",
  55039=>"001110101",
  55040=>"000000010",
  55041=>"100111011",
  55042=>"010111010",
  55043=>"010010000",
  55044=>"010101111",
  55045=>"000001010",
  55046=>"100011001",
  55047=>"011010101",
  55048=>"000100001",
  55049=>"111010011",
  55050=>"001111101",
  55051=>"011111000",
  55052=>"111101111",
  55053=>"101001001",
  55054=>"101000111",
  55055=>"100111010",
  55056=>"100111000",
  55057=>"001101000",
  55058=>"011001101",
  55059=>"110101011",
  55060=>"011110000",
  55061=>"010010101",
  55062=>"111101101",
  55063=>"000000010",
  55064=>"001100100",
  55065=>"001111110",
  55066=>"110001100",
  55067=>"000110100",
  55068=>"001111101",
  55069=>"010111100",
  55070=>"101101111",
  55071=>"010110111",
  55072=>"111011101",
  55073=>"110110010",
  55074=>"110111111",
  55075=>"000001010",
  55076=>"100011000",
  55077=>"101100110",
  55078=>"110110011",
  55079=>"000111111",
  55080=>"111110101",
  55081=>"000100111",
  55082=>"110100010",
  55083=>"110000011",
  55084=>"110011101",
  55085=>"101010011",
  55086=>"010000010",
  55087=>"100010010",
  55088=>"101111000",
  55089=>"010011110",
  55090=>"001101110",
  55091=>"000100010",
  55092=>"010000000",
  55093=>"100110111",
  55094=>"010100100",
  55095=>"011110011",
  55096=>"101111101",
  55097=>"010100000",
  55098=>"001110001",
  55099=>"000010001",
  55100=>"000110111",
  55101=>"101100011",
  55102=>"011000110",
  55103=>"111100101",
  55104=>"011101011",
  55105=>"101111100",
  55106=>"111111111",
  55107=>"001000001",
  55108=>"111101111",
  55109=>"001111000",
  55110=>"010000111",
  55111=>"001110110",
  55112=>"110001010",
  55113=>"110100011",
  55114=>"111011111",
  55115=>"001110100",
  55116=>"011001100",
  55117=>"001110110",
  55118=>"011010110",
  55119=>"100010100",
  55120=>"011011011",
  55121=>"111110110",
  55122=>"011010010",
  55123=>"000000110",
  55124=>"100010010",
  55125=>"011110101",
  55126=>"000001111",
  55127=>"011111001",
  55128=>"001000100",
  55129=>"101100111",
  55130=>"101111000",
  55131=>"001111001",
  55132=>"010100011",
  55133=>"010100000",
  55134=>"010001010",
  55135=>"100110101",
  55136=>"010000100",
  55137=>"011010001",
  55138=>"000000110",
  55139=>"110010100",
  55140=>"011010101",
  55141=>"001101110",
  55142=>"011000110",
  55143=>"000010010",
  55144=>"011011010",
  55145=>"000011100",
  55146=>"011000011",
  55147=>"101100011",
  55148=>"011000101",
  55149=>"100111010",
  55150=>"000110110",
  55151=>"000100110",
  55152=>"101111100",
  55153=>"101110110",
  55154=>"101000110",
  55155=>"111100011",
  55156=>"100001010",
  55157=>"011010000",
  55158=>"011000000",
  55159=>"111110110",
  55160=>"010010011",
  55161=>"001011101",
  55162=>"100110101",
  55163=>"011111101",
  55164=>"001101101",
  55165=>"111111111",
  55166=>"010011101",
  55167=>"100001101",
  55168=>"100011001",
  55169=>"110101100",
  55170=>"110110111",
  55171=>"110110110",
  55172=>"100000001",
  55173=>"111111001",
  55174=>"100110100",
  55175=>"000111101",
  55176=>"001001000",
  55177=>"111011100",
  55178=>"101000111",
  55179=>"110100001",
  55180=>"000001110",
  55181=>"111011101",
  55182=>"101111101",
  55183=>"011011000",
  55184=>"001111010",
  55185=>"111110110",
  55186=>"000110001",
  55187=>"011011010",
  55188=>"010101100",
  55189=>"101000110",
  55190=>"100011001",
  55191=>"000110111",
  55192=>"100000001",
  55193=>"010110101",
  55194=>"110010000",
  55195=>"101110011",
  55196=>"111001100",
  55197=>"011011000",
  55198=>"111110000",
  55199=>"110000010",
  55200=>"101000110",
  55201=>"110010101",
  55202=>"010001000",
  55203=>"001100010",
  55204=>"110000011",
  55205=>"110011111",
  55206=>"001111010",
  55207=>"110001101",
  55208=>"110111101",
  55209=>"011000111",
  55210=>"101010000",
  55211=>"011110100",
  55212=>"000100110",
  55213=>"010010010",
  55214=>"010101010",
  55215=>"111101000",
  55216=>"000111100",
  55217=>"111011011",
  55218=>"001110101",
  55219=>"000110100",
  55220=>"010110111",
  55221=>"001011010",
  55222=>"101001110",
  55223=>"111101000",
  55224=>"010001111",
  55225=>"100111000",
  55226=>"001011100",
  55227=>"111011111",
  55228=>"011101111",
  55229=>"011000001",
  55230=>"110011101",
  55231=>"010110110",
  55232=>"001000111",
  55233=>"110111101",
  55234=>"111010110",
  55235=>"100000101",
  55236=>"100110111",
  55237=>"001001000",
  55238=>"010101011",
  55239=>"001001011",
  55240=>"000010000",
  55241=>"101011011",
  55242=>"110101000",
  55243=>"000011101",
  55244=>"001101011",
  55245=>"110110000",
  55246=>"010100100",
  55247=>"110001110",
  55248=>"101011111",
  55249=>"010001011",
  55250=>"010001110",
  55251=>"011100110",
  55252=>"011111101",
  55253=>"111111110",
  55254=>"101111110",
  55255=>"010001011",
  55256=>"010010111",
  55257=>"011000000",
  55258=>"111111100",
  55259=>"101001001",
  55260=>"100111100",
  55261=>"100100010",
  55262=>"010011110",
  55263=>"101001011",
  55264=>"001101100",
  55265=>"011011110",
  55266=>"110101111",
  55267=>"001100111",
  55268=>"010000101",
  55269=>"001011000",
  55270=>"001001100",
  55271=>"010100010",
  55272=>"001001010",
  55273=>"100110011",
  55274=>"111101010",
  55275=>"000101011",
  55276=>"111110110",
  55277=>"001111111",
  55278=>"110000011",
  55279=>"011010010",
  55280=>"111110010",
  55281=>"011101000",
  55282=>"000000110",
  55283=>"011100101",
  55284=>"111110101",
  55285=>"101111101",
  55286=>"000000001",
  55287=>"011000101",
  55288=>"000101111",
  55289=>"001101110",
  55290=>"010100111",
  55291=>"111111000",
  55292=>"100001000",
  55293=>"101001100",
  55294=>"111110000",
  55295=>"111011110",
  55296=>"110000111",
  55297=>"011010100",
  55298=>"000000011",
  55299=>"000000111",
  55300=>"001100010",
  55301=>"010000110",
  55302=>"110011101",
  55303=>"111111111",
  55304=>"100101110",
  55305=>"101100010",
  55306=>"101000010",
  55307=>"010101100",
  55308=>"111100100",
  55309=>"001100010",
  55310=>"110111000",
  55311=>"000100110",
  55312=>"011111101",
  55313=>"101010111",
  55314=>"011001100",
  55315=>"110000110",
  55316=>"000101011",
  55317=>"000110000",
  55318=>"011011011",
  55319=>"101000101",
  55320=>"101111000",
  55321=>"001110001",
  55322=>"010000001",
  55323=>"100000100",
  55324=>"111110011",
  55325=>"011110001",
  55326=>"001110111",
  55327=>"011110100",
  55328=>"101100010",
  55329=>"110011110",
  55330=>"000111101",
  55331=>"011010100",
  55332=>"010001100",
  55333=>"001000001",
  55334=>"001100110",
  55335=>"100010111",
  55336=>"111111110",
  55337=>"100000001",
  55338=>"110111110",
  55339=>"001100100",
  55340=>"011111010",
  55341=>"010111110",
  55342=>"100101100",
  55343=>"010000011",
  55344=>"110100010",
  55345=>"110110101",
  55346=>"110100100",
  55347=>"101001101",
  55348=>"100100111",
  55349=>"000001011",
  55350=>"010000010",
  55351=>"111101010",
  55352=>"111010000",
  55353=>"001010001",
  55354=>"101001111",
  55355=>"001110010",
  55356=>"101001011",
  55357=>"111000001",
  55358=>"101011010",
  55359=>"111101000",
  55360=>"011101110",
  55361=>"011101111",
  55362=>"101001010",
  55363=>"010011010",
  55364=>"101100001",
  55365=>"011101001",
  55366=>"011000000",
  55367=>"000101001",
  55368=>"001001100",
  55369=>"011010011",
  55370=>"100011011",
  55371=>"110100001",
  55372=>"010001101",
  55373=>"110001011",
  55374=>"001010001",
  55375=>"111111101",
  55376=>"111110111",
  55377=>"111111100",
  55378=>"101000110",
  55379=>"010000111",
  55380=>"111111111",
  55381=>"101010000",
  55382=>"000001101",
  55383=>"101101000",
  55384=>"000100000",
  55385=>"111011010",
  55386=>"101110000",
  55387=>"111011000",
  55388=>"111110000",
  55389=>"011011101",
  55390=>"110011111",
  55391=>"000111010",
  55392=>"100101111",
  55393=>"001000011",
  55394=>"101110100",
  55395=>"110100101",
  55396=>"000000101",
  55397=>"010001100",
  55398=>"011011001",
  55399=>"100010000",
  55400=>"110110011",
  55401=>"111101000",
  55402=>"110011110",
  55403=>"001000110",
  55404=>"110011001",
  55405=>"110100010",
  55406=>"110111011",
  55407=>"110110100",
  55408=>"101000001",
  55409=>"111010101",
  55410=>"111011110",
  55411=>"010001010",
  55412=>"100001010",
  55413=>"001011011",
  55414=>"101110011",
  55415=>"000010100",
  55416=>"001111110",
  55417=>"000010101",
  55418=>"011011010",
  55419=>"111110111",
  55420=>"001111101",
  55421=>"000001101",
  55422=>"010000000",
  55423=>"011000000",
  55424=>"000110110",
  55425=>"111001000",
  55426=>"011011010",
  55427=>"100101110",
  55428=>"110001010",
  55429=>"111010101",
  55430=>"111101010",
  55431=>"011100101",
  55432=>"111100010",
  55433=>"010000000",
  55434=>"101010101",
  55435=>"000111000",
  55436=>"101110000",
  55437=>"011010010",
  55438=>"100010011",
  55439=>"010011110",
  55440=>"011101110",
  55441=>"001011100",
  55442=>"011010000",
  55443=>"111001001",
  55444=>"101101111",
  55445=>"010011001",
  55446=>"101101011",
  55447=>"111100101",
  55448=>"110000010",
  55449=>"010111100",
  55450=>"001100111",
  55451=>"111001011",
  55452=>"010000111",
  55453=>"101100001",
  55454=>"101010001",
  55455=>"100110000",
  55456=>"110101011",
  55457=>"101101011",
  55458=>"110111111",
  55459=>"001111101",
  55460=>"011001001",
  55461=>"010010000",
  55462=>"001101101",
  55463=>"001110011",
  55464=>"100001100",
  55465=>"111001110",
  55466=>"100010101",
  55467=>"001101110",
  55468=>"100000000",
  55469=>"000011010",
  55470=>"010111110",
  55471=>"011000100",
  55472=>"001000001",
  55473=>"011001000",
  55474=>"101100101",
  55475=>"100000110",
  55476=>"110100100",
  55477=>"011100001",
  55478=>"011001101",
  55479=>"100000010",
  55480=>"001000000",
  55481=>"000010100",
  55482=>"111110100",
  55483=>"111111010",
  55484=>"001001001",
  55485=>"101011101",
  55486=>"011110011",
  55487=>"101100000",
  55488=>"011101001",
  55489=>"001000100",
  55490=>"111000001",
  55491=>"001001001",
  55492=>"110001100",
  55493=>"101000010",
  55494=>"010101110",
  55495=>"010010101",
  55496=>"011110011",
  55497=>"000000110",
  55498=>"000000001",
  55499=>"010000100",
  55500=>"010100000",
  55501=>"000111111",
  55502=>"010001101",
  55503=>"000100110",
  55504=>"011100110",
  55505=>"001010000",
  55506=>"100111111",
  55507=>"111011011",
  55508=>"010011110",
  55509=>"100011111",
  55510=>"000011010",
  55511=>"110001010",
  55512=>"100001100",
  55513=>"010100110",
  55514=>"110001010",
  55515=>"111011100",
  55516=>"011100111",
  55517=>"010111110",
  55518=>"110110001",
  55519=>"011101011",
  55520=>"111101111",
  55521=>"100000011",
  55522=>"110010010",
  55523=>"010111101",
  55524=>"111111110",
  55525=>"001010001",
  55526=>"101101100",
  55527=>"010000100",
  55528=>"000100100",
  55529=>"110001010",
  55530=>"000001100",
  55531=>"000010000",
  55532=>"101101001",
  55533=>"110110011",
  55534=>"110010100",
  55535=>"101001101",
  55536=>"000001010",
  55537=>"110110101",
  55538=>"001100001",
  55539=>"010010000",
  55540=>"001101111",
  55541=>"011000010",
  55542=>"011100000",
  55543=>"100011001",
  55544=>"101011111",
  55545=>"000110000",
  55546=>"001100001",
  55547=>"100100101",
  55548=>"000100110",
  55549=>"101010110",
  55550=>"111010011",
  55551=>"111111110",
  55552=>"000000110",
  55553=>"101000110",
  55554=>"011110100",
  55555=>"010111000",
  55556=>"111110011",
  55557=>"111100001",
  55558=>"111111001",
  55559=>"000111100",
  55560=>"011101111",
  55561=>"001101100",
  55562=>"011100000",
  55563=>"100100000",
  55564=>"110011000",
  55565=>"111001101",
  55566=>"110010011",
  55567=>"111100010",
  55568=>"110000100",
  55569=>"001000001",
  55570=>"111000000",
  55571=>"100101000",
  55572=>"101001111",
  55573=>"101100001",
  55574=>"001011010",
  55575=>"110111011",
  55576=>"111000000",
  55577=>"000001100",
  55578=>"110110101",
  55579=>"100101010",
  55580=>"000011111",
  55581=>"010100011",
  55582=>"011100010",
  55583=>"010000000",
  55584=>"100111010",
  55585=>"011001110",
  55586=>"001001110",
  55587=>"111100000",
  55588=>"101111111",
  55589=>"111110101",
  55590=>"110110111",
  55591=>"011010001",
  55592=>"100100100",
  55593=>"100010011",
  55594=>"001110111",
  55595=>"110110001",
  55596=>"000100110",
  55597=>"011001101",
  55598=>"111111000",
  55599=>"100010101",
  55600=>"110000000",
  55601=>"000001011",
  55602=>"111111011",
  55603=>"110000000",
  55604=>"111101101",
  55605=>"000000111",
  55606=>"100011100",
  55607=>"011000001",
  55608=>"011001000",
  55609=>"000000110",
  55610=>"101111100",
  55611=>"010100101",
  55612=>"101111101",
  55613=>"110011110",
  55614=>"000000100",
  55615=>"100110011",
  55616=>"100100001",
  55617=>"000100010",
  55618=>"011101101",
  55619=>"000000000",
  55620=>"011111000",
  55621=>"100101100",
  55622=>"101001000",
  55623=>"111111110",
  55624=>"011001100",
  55625=>"010000000",
  55626=>"010001101",
  55627=>"001011101",
  55628=>"111101011",
  55629=>"110000011",
  55630=>"101011010",
  55631=>"110000000",
  55632=>"101101111",
  55633=>"010111111",
  55634=>"011100010",
  55635=>"011101111",
  55636=>"000010011",
  55637=>"011101000",
  55638=>"100011110",
  55639=>"100101100",
  55640=>"010110000",
  55641=>"010101101",
  55642=>"000110101",
  55643=>"000101001",
  55644=>"010111100",
  55645=>"011001000",
  55646=>"011001000",
  55647=>"110110100",
  55648=>"101111010",
  55649=>"110001100",
  55650=>"100101110",
  55651=>"001101110",
  55652=>"001001001",
  55653=>"000010110",
  55654=>"000101111",
  55655=>"011110100",
  55656=>"001000011",
  55657=>"001010110",
  55658=>"000010001",
  55659=>"001000010",
  55660=>"100111101",
  55661=>"111101111",
  55662=>"000101100",
  55663=>"011001001",
  55664=>"111010100",
  55665=>"100001101",
  55666=>"001001010",
  55667=>"000011111",
  55668=>"000011000",
  55669=>"100100111",
  55670=>"001001101",
  55671=>"101010110",
  55672=>"010000101",
  55673=>"000000111",
  55674=>"001100101",
  55675=>"000001010",
  55676=>"101011110",
  55677=>"100111101",
  55678=>"000000001",
  55679=>"011100110",
  55680=>"101100011",
  55681=>"100111111",
  55682=>"110100110",
  55683=>"100111111",
  55684=>"111101111",
  55685=>"001000100",
  55686=>"110010001",
  55687=>"100100000",
  55688=>"010001010",
  55689=>"110000110",
  55690=>"111110000",
  55691=>"010000101",
  55692=>"001001111",
  55693=>"000010110",
  55694=>"010100010",
  55695=>"000010111",
  55696=>"100100010",
  55697=>"101111001",
  55698=>"001100001",
  55699=>"100111010",
  55700=>"001101110",
  55701=>"001010011",
  55702=>"010100000",
  55703=>"000010000",
  55704=>"100010000",
  55705=>"101000011",
  55706=>"011011000",
  55707=>"101000110",
  55708=>"011010111",
  55709=>"011001111",
  55710=>"101100100",
  55711=>"010011100",
  55712=>"101011110",
  55713=>"001110000",
  55714=>"101000010",
  55715=>"000000000",
  55716=>"001111001",
  55717=>"110111101",
  55718=>"100101000",
  55719=>"111001110",
  55720=>"101111111",
  55721=>"110001000",
  55722=>"010110101",
  55723=>"010110100",
  55724=>"101111000",
  55725=>"001111111",
  55726=>"001111100",
  55727=>"001011001",
  55728=>"010011001",
  55729=>"000100010",
  55730=>"111011000",
  55731=>"000001111",
  55732=>"101001110",
  55733=>"001000000",
  55734=>"110111101",
  55735=>"101011111",
  55736=>"111110110",
  55737=>"010111110",
  55738=>"100110010",
  55739=>"001010111",
  55740=>"001000100",
  55741=>"001110001",
  55742=>"011111011",
  55743=>"011111100",
  55744=>"010100111",
  55745=>"010001110",
  55746=>"100100001",
  55747=>"110011111",
  55748=>"111000000",
  55749=>"000110011",
  55750=>"010011001",
  55751=>"000000000",
  55752=>"000000100",
  55753=>"001101111",
  55754=>"110111010",
  55755=>"111011000",
  55756=>"101001010",
  55757=>"111010100",
  55758=>"110001000",
  55759=>"111111011",
  55760=>"111110100",
  55761=>"101101000",
  55762=>"111000000",
  55763=>"011011111",
  55764=>"101111110",
  55765=>"110100101",
  55766=>"100111110",
  55767=>"110001111",
  55768=>"100101010",
  55769=>"001100011",
  55770=>"011101101",
  55771=>"000111100",
  55772=>"111100100",
  55773=>"100100110",
  55774=>"001011110",
  55775=>"100111110",
  55776=>"100000111",
  55777=>"000011011",
  55778=>"100001111",
  55779=>"111101111",
  55780=>"111010101",
  55781=>"001000010",
  55782=>"111100111",
  55783=>"100000010",
  55784=>"001010101",
  55785=>"101001110",
  55786=>"011101011",
  55787=>"111011011",
  55788=>"011110111",
  55789=>"000000001",
  55790=>"100111100",
  55791=>"000011101",
  55792=>"010111000",
  55793=>"000101000",
  55794=>"110010001",
  55795=>"110010001",
  55796=>"010011111",
  55797=>"110011011",
  55798=>"011011001",
  55799=>"110010001",
  55800=>"011000000",
  55801=>"011011100",
  55802=>"101010100",
  55803=>"111111001",
  55804=>"101111111",
  55805=>"011100010",
  55806=>"101101011",
  55807=>"100111110",
  55808=>"001000000",
  55809=>"111100010",
  55810=>"100000111",
  55811=>"000100111",
  55812=>"001010001",
  55813=>"101000010",
  55814=>"101011110",
  55815=>"100111110",
  55816=>"100101100",
  55817=>"111101001",
  55818=>"000111000",
  55819=>"110110001",
  55820=>"000011001",
  55821=>"111000000",
  55822=>"101111011",
  55823=>"100001010",
  55824=>"111011000",
  55825=>"100010010",
  55826=>"110100110",
  55827=>"000100111",
  55828=>"100100000",
  55829=>"101101111",
  55830=>"110011111",
  55831=>"000001001",
  55832=>"101110111",
  55833=>"011000111",
  55834=>"000000011",
  55835=>"000111110",
  55836=>"000110011",
  55837=>"110110101",
  55838=>"110000110",
  55839=>"110111100",
  55840=>"010001011",
  55841=>"111101010",
  55842=>"111000001",
  55843=>"110000000",
  55844=>"010111110",
  55845=>"000100000",
  55846=>"110000101",
  55847=>"101001101",
  55848=>"111001110",
  55849=>"100011000",
  55850=>"101010001",
  55851=>"000000110",
  55852=>"101100001",
  55853=>"011111011",
  55854=>"100001111",
  55855=>"100101101",
  55856=>"110110111",
  55857=>"111101110",
  55858=>"000011110",
  55859=>"011000110",
  55860=>"101100010",
  55861=>"110110100",
  55862=>"011110010",
  55863=>"000001011",
  55864=>"100001101",
  55865=>"101110010",
  55866=>"010101011",
  55867=>"101111001",
  55868=>"001001110",
  55869=>"001111111",
  55870=>"111111001",
  55871=>"011110110",
  55872=>"010100110",
  55873=>"111101010",
  55874=>"111010010",
  55875=>"010001110",
  55876=>"100101111",
  55877=>"101100000",
  55878=>"011010101",
  55879=>"000101101",
  55880=>"000011111",
  55881=>"001100111",
  55882=>"100011100",
  55883=>"111001110",
  55884=>"111100101",
  55885=>"000000010",
  55886=>"110100001",
  55887=>"100111001",
  55888=>"101000111",
  55889=>"101100001",
  55890=>"000110111",
  55891=>"100010001",
  55892=>"100101001",
  55893=>"000111101",
  55894=>"000110000",
  55895=>"100001110",
  55896=>"000101010",
  55897=>"110011010",
  55898=>"110101011",
  55899=>"010010001",
  55900=>"101001000",
  55901=>"110001100",
  55902=>"010011111",
  55903=>"100101001",
  55904=>"110011011",
  55905=>"000111110",
  55906=>"111101111",
  55907=>"000000000",
  55908=>"111110100",
  55909=>"000000011",
  55910=>"100101101",
  55911=>"011101000",
  55912=>"111000000",
  55913=>"110011011",
  55914=>"101010101",
  55915=>"000101100",
  55916=>"100000011",
  55917=>"100010011",
  55918=>"100100110",
  55919=>"101111001",
  55920=>"100011100",
  55921=>"000000011",
  55922=>"110111001",
  55923=>"011111001",
  55924=>"111100100",
  55925=>"100011110",
  55926=>"001101000",
  55927=>"000110011",
  55928=>"001100111",
  55929=>"101011001",
  55930=>"111010101",
  55931=>"101000001",
  55932=>"001010101",
  55933=>"001000000",
  55934=>"101101111",
  55935=>"111111001",
  55936=>"011000100",
  55937=>"001110100",
  55938=>"111001101",
  55939=>"000000100",
  55940=>"000010000",
  55941=>"011000000",
  55942=>"111010100",
  55943=>"000100000",
  55944=>"111110011",
  55945=>"000011001",
  55946=>"000010111",
  55947=>"011000111",
  55948=>"001111111",
  55949=>"110101100",
  55950=>"011100110",
  55951=>"100110111",
  55952=>"111101101",
  55953=>"011001111",
  55954=>"000001100",
  55955=>"100101110",
  55956=>"010110110",
  55957=>"110111101",
  55958=>"110110001",
  55959=>"101100000",
  55960=>"000011101",
  55961=>"000010111",
  55962=>"101111010",
  55963=>"111100101",
  55964=>"101101101",
  55965=>"110100010",
  55966=>"000100010",
  55967=>"111101101",
  55968=>"110011100",
  55969=>"010001111",
  55970=>"100100011",
  55971=>"011001000",
  55972=>"011010100",
  55973=>"000111011",
  55974=>"110101101",
  55975=>"000001010",
  55976=>"100110111",
  55977=>"000000100",
  55978=>"110100110",
  55979=>"101010110",
  55980=>"111001111",
  55981=>"011000101",
  55982=>"001101001",
  55983=>"101110101",
  55984=>"010111100",
  55985=>"101111101",
  55986=>"110000100",
  55987=>"010100010",
  55988=>"000000000",
  55989=>"100111000",
  55990=>"110100010",
  55991=>"010010101",
  55992=>"000000100",
  55993=>"110100000",
  55994=>"101011110",
  55995=>"111011100",
  55996=>"110001001",
  55997=>"001000001",
  55998=>"001100001",
  55999=>"100101100",
  56000=>"000011111",
  56001=>"100100110",
  56002=>"011100000",
  56003=>"100011001",
  56004=>"000100101",
  56005=>"000001000",
  56006=>"011000110",
  56007=>"110000111",
  56008=>"011110100",
  56009=>"111000011",
  56010=>"000000100",
  56011=>"101000010",
  56012=>"111110111",
  56013=>"000100010",
  56014=>"001000110",
  56015=>"000100011",
  56016=>"101011010",
  56017=>"110010110",
  56018=>"011000110",
  56019=>"100111011",
  56020=>"010000000",
  56021=>"001001010",
  56022=>"011100111",
  56023=>"001000011",
  56024=>"000011110",
  56025=>"011001011",
  56026=>"011000001",
  56027=>"101000101",
  56028=>"110100110",
  56029=>"000011001",
  56030=>"001010000",
  56031=>"000010000",
  56032=>"111100101",
  56033=>"101011011",
  56034=>"110010101",
  56035=>"100100100",
  56036=>"100001011",
  56037=>"001100110",
  56038=>"000011111",
  56039=>"110110101",
  56040=>"000011110",
  56041=>"011011111",
  56042=>"000011000",
  56043=>"101010100",
  56044=>"100101000",
  56045=>"000111000",
  56046=>"101011000",
  56047=>"011100000",
  56048=>"110011110",
  56049=>"000001010",
  56050=>"110000111",
  56051=>"011110111",
  56052=>"001000011",
  56053=>"010010010",
  56054=>"011100111",
  56055=>"111011000",
  56056=>"001010100",
  56057=>"000010110",
  56058=>"000011111",
  56059=>"111100100",
  56060=>"010011100",
  56061=>"001001010",
  56062=>"010100000",
  56063=>"111101010",
  56064=>"111110101",
  56065=>"010111001",
  56066=>"010101010",
  56067=>"011100101",
  56068=>"111101111",
  56069=>"001000000",
  56070=>"010001010",
  56071=>"111111101",
  56072=>"010101101",
  56073=>"000101111",
  56074=>"111001110",
  56075=>"000100000",
  56076=>"110011000",
  56077=>"011000011",
  56078=>"100001100",
  56079=>"010100110",
  56080=>"100111100",
  56081=>"111001110",
  56082=>"001000111",
  56083=>"111111111",
  56084=>"000101000",
  56085=>"111100111",
  56086=>"101011110",
  56087=>"000010000",
  56088=>"001011001",
  56089=>"001000001",
  56090=>"110101001",
  56091=>"110110000",
  56092=>"100111001",
  56093=>"101101001",
  56094=>"101100110",
  56095=>"100001010",
  56096=>"100001011",
  56097=>"101011000",
  56098=>"000000100",
  56099=>"010101001",
  56100=>"101111101",
  56101=>"100110000",
  56102=>"001100001",
  56103=>"100010110",
  56104=>"100001011",
  56105=>"111101100",
  56106=>"000111111",
  56107=>"010001101",
  56108=>"011101011",
  56109=>"101000001",
  56110=>"101000010",
  56111=>"101000010",
  56112=>"100110001",
  56113=>"110000100",
  56114=>"001111000",
  56115=>"100100000",
  56116=>"101100111",
  56117=>"000111000",
  56118=>"010101101",
  56119=>"100111101",
  56120=>"111001110",
  56121=>"000110010",
  56122=>"111110011",
  56123=>"110111001",
  56124=>"111101011",
  56125=>"100101011",
  56126=>"001011000",
  56127=>"100100001",
  56128=>"011111111",
  56129=>"001001011",
  56130=>"110011101",
  56131=>"001010100",
  56132=>"101110011",
  56133=>"010101100",
  56134=>"000000101",
  56135=>"111100111",
  56136=>"010010011",
  56137=>"000100011",
  56138=>"010101110",
  56139=>"001011101",
  56140=>"100110100",
  56141=>"011110010",
  56142=>"001010011",
  56143=>"101000011",
  56144=>"110111111",
  56145=>"110000001",
  56146=>"001000101",
  56147=>"100101010",
  56148=>"001111000",
  56149=>"001010011",
  56150=>"111111010",
  56151=>"110010000",
  56152=>"011000011",
  56153=>"011100110",
  56154=>"011111010",
  56155=>"101011110",
  56156=>"101111011",
  56157=>"011111110",
  56158=>"110100100",
  56159=>"001000011",
  56160=>"001110101",
  56161=>"000101100",
  56162=>"000110011",
  56163=>"010001111",
  56164=>"000010101",
  56165=>"101000111",
  56166=>"010000110",
  56167=>"010110110",
  56168=>"000100101",
  56169=>"110010001",
  56170=>"101100001",
  56171=>"001010101",
  56172=>"111111100",
  56173=>"000101011",
  56174=>"010010101",
  56175=>"111111000",
  56176=>"100101111",
  56177=>"011101000",
  56178=>"101001010",
  56179=>"101111111",
  56180=>"101100001",
  56181=>"001010100",
  56182=>"111111101",
  56183=>"101011101",
  56184=>"101101001",
  56185=>"110101101",
  56186=>"100110001",
  56187=>"101000000",
  56188=>"000001001",
  56189=>"100101111",
  56190=>"001110101",
  56191=>"100001100",
  56192=>"000101001",
  56193=>"001101110",
  56194=>"000001010",
  56195=>"100110010",
  56196=>"001100100",
  56197=>"010101001",
  56198=>"000000000",
  56199=>"101011010",
  56200=>"000011100",
  56201=>"100001011",
  56202=>"100111100",
  56203=>"101100111",
  56204=>"111110011",
  56205=>"110100100",
  56206=>"000110001",
  56207=>"101000001",
  56208=>"000110101",
  56209=>"010000011",
  56210=>"000111001",
  56211=>"101111011",
  56212=>"000010010",
  56213=>"001010000",
  56214=>"000001011",
  56215=>"000111100",
  56216=>"110000000",
  56217=>"010011100",
  56218=>"101010101",
  56219=>"011110010",
  56220=>"001000110",
  56221=>"000011000",
  56222=>"010000110",
  56223=>"010100000",
  56224=>"111100100",
  56225=>"100110000",
  56226=>"101111101",
  56227=>"000010011",
  56228=>"001100000",
  56229=>"000111011",
  56230=>"011010000",
  56231=>"101101001",
  56232=>"001100000",
  56233=>"011000000",
  56234=>"110111001",
  56235=>"100111111",
  56236=>"110000110",
  56237=>"000110111",
  56238=>"100001010",
  56239=>"110011110",
  56240=>"000111001",
  56241=>"100100110",
  56242=>"011111100",
  56243=>"111100001",
  56244=>"110010001",
  56245=>"100000100",
  56246=>"000110110",
  56247=>"111011111",
  56248=>"111101000",
  56249=>"111001000",
  56250=>"011101010",
  56251=>"100000001",
  56252=>"101001000",
  56253=>"110100111",
  56254=>"000011100",
  56255=>"101100010",
  56256=>"001001110",
  56257=>"110110000",
  56258=>"100001100",
  56259=>"100000000",
  56260=>"001110110",
  56261=>"010011100",
  56262=>"111011010",
  56263=>"001001010",
  56264=>"100101000",
  56265=>"011010010",
  56266=>"111000111",
  56267=>"101001011",
  56268=>"001101011",
  56269=>"110111111",
  56270=>"011001110",
  56271=>"111011111",
  56272=>"101110111",
  56273=>"111110011",
  56274=>"010000001",
  56275=>"011011110",
  56276=>"001100110",
  56277=>"100111011",
  56278=>"001001100",
  56279=>"100000100",
  56280=>"010010011",
  56281=>"011011110",
  56282=>"011001000",
  56283=>"100000000",
  56284=>"101010010",
  56285=>"011111001",
  56286=>"000001101",
  56287=>"111100010",
  56288=>"100111001",
  56289=>"000000010",
  56290=>"111111111",
  56291=>"101011001",
  56292=>"111000100",
  56293=>"011001111",
  56294=>"001101000",
  56295=>"000000011",
  56296=>"110111101",
  56297=>"001001100",
  56298=>"110011101",
  56299=>"001110000",
  56300=>"000000001",
  56301=>"111110010",
  56302=>"110111000",
  56303=>"100110001",
  56304=>"101101100",
  56305=>"010101110",
  56306=>"101110011",
  56307=>"101110000",
  56308=>"011010010",
  56309=>"101010111",
  56310=>"001101111",
  56311=>"110011101",
  56312=>"110011011",
  56313=>"010010111",
  56314=>"100001001",
  56315=>"010011110",
  56316=>"010011010",
  56317=>"110000011",
  56318=>"100111110",
  56319=>"101010011",
  56320=>"001110111",
  56321=>"011111110",
  56322=>"110110010",
  56323=>"001000111",
  56324=>"111111001",
  56325=>"100010001",
  56326=>"100110111",
  56327=>"111000001",
  56328=>"100010111",
  56329=>"100111111",
  56330=>"000010100",
  56331=>"111101100",
  56332=>"010111001",
  56333=>"100010110",
  56334=>"101000101",
  56335=>"101001100",
  56336=>"111001011",
  56337=>"000001000",
  56338=>"010100001",
  56339=>"110000111",
  56340=>"000001011",
  56341=>"110011011",
  56342=>"100110101",
  56343=>"010011111",
  56344=>"111010111",
  56345=>"100100110",
  56346=>"010001010",
  56347=>"001011101",
  56348=>"011100110",
  56349=>"100111110",
  56350=>"111011111",
  56351=>"111110011",
  56352=>"000100110",
  56353=>"111101000",
  56354=>"000000010",
  56355=>"101011101",
  56356=>"001011110",
  56357=>"101010101",
  56358=>"100011110",
  56359=>"111011001",
  56360=>"000010010",
  56361=>"000110011",
  56362=>"001010000",
  56363=>"010110100",
  56364=>"100111100",
  56365=>"001110101",
  56366=>"000101111",
  56367=>"010001010",
  56368=>"010001000",
  56369=>"001001011",
  56370=>"001011000",
  56371=>"111101010",
  56372=>"011001100",
  56373=>"111010000",
  56374=>"001001001",
  56375=>"111110101",
  56376=>"001010110",
  56377=>"000001010",
  56378=>"000001110",
  56379=>"011111100",
  56380=>"010110111",
  56381=>"110111000",
  56382=>"111011101",
  56383=>"100010011",
  56384=>"010100000",
  56385=>"000001111",
  56386=>"000010011",
  56387=>"101101000",
  56388=>"000010111",
  56389=>"101010011",
  56390=>"101101010",
  56391=>"110100011",
  56392=>"100000010",
  56393=>"100011011",
  56394=>"010010111",
  56395=>"110110001",
  56396=>"101111101",
  56397=>"100010111",
  56398=>"011110000",
  56399=>"010001000",
  56400=>"011101011",
  56401=>"000111010",
  56402=>"111010011",
  56403=>"011010011",
  56404=>"010101100",
  56405=>"111100000",
  56406=>"110001111",
  56407=>"010000001",
  56408=>"001110001",
  56409=>"110100010",
  56410=>"101011101",
  56411=>"000110000",
  56412=>"110000001",
  56413=>"001100010",
  56414=>"100111001",
  56415=>"110100011",
  56416=>"111000000",
  56417=>"011010111",
  56418=>"010000011",
  56419=>"100010001",
  56420=>"001000010",
  56421=>"101010111",
  56422=>"100011100",
  56423=>"000111100",
  56424=>"011100011",
  56425=>"100001111",
  56426=>"000001110",
  56427=>"110111100",
  56428=>"111000100",
  56429=>"011111001",
  56430=>"011000100",
  56431=>"110111011",
  56432=>"000001101",
  56433=>"001111010",
  56434=>"111100011",
  56435=>"111000011",
  56436=>"000001110",
  56437=>"101010110",
  56438=>"001001011",
  56439=>"000001001",
  56440=>"100001111",
  56441=>"100110111",
  56442=>"011001001",
  56443=>"010111010",
  56444=>"101011011",
  56445=>"111110001",
  56446=>"001011010",
  56447=>"001011110",
  56448=>"110101001",
  56449=>"011110111",
  56450=>"111011100",
  56451=>"110011110",
  56452=>"001110110",
  56453=>"110111010",
  56454=>"011111111",
  56455=>"101010110",
  56456=>"000100001",
  56457=>"001111100",
  56458=>"011010010",
  56459=>"111000010",
  56460=>"000001110",
  56461=>"001000010",
  56462=>"100101000",
  56463=>"001110010",
  56464=>"010010001",
  56465=>"100111101",
  56466=>"111110110",
  56467=>"110011011",
  56468=>"110001010",
  56469=>"111110010",
  56470=>"110011011",
  56471=>"010000000",
  56472=>"010010001",
  56473=>"011111110",
  56474=>"110101000",
  56475=>"011000100",
  56476=>"100110111",
  56477=>"010110101",
  56478=>"111110001",
  56479=>"111100100",
  56480=>"111001110",
  56481=>"000111000",
  56482=>"110000000",
  56483=>"001000000",
  56484=>"000010101",
  56485=>"000101100",
  56486=>"000010000",
  56487=>"110010100",
  56488=>"110111001",
  56489=>"000001111",
  56490=>"000011101",
  56491=>"011011000",
  56492=>"011110001",
  56493=>"010100110",
  56494=>"110110111",
  56495=>"000001000",
  56496=>"011110011",
  56497=>"110101001",
  56498=>"001100011",
  56499=>"100001101",
  56500=>"100000000",
  56501=>"100100001",
  56502=>"000110111",
  56503=>"100000100",
  56504=>"011111110",
  56505=>"000100000",
  56506=>"100101100",
  56507=>"111100000",
  56508=>"001000101",
  56509=>"001100000",
  56510=>"001000111",
  56511=>"000000001",
  56512=>"001110001",
  56513=>"110110000",
  56514=>"110000110",
  56515=>"111110111",
  56516=>"110101111",
  56517=>"000101110",
  56518=>"101000011",
  56519=>"011010001",
  56520=>"010011001",
  56521=>"010011111",
  56522=>"101110011",
  56523=>"011100000",
  56524=>"100100000",
  56525=>"100110111",
  56526=>"100010100",
  56527=>"100100000",
  56528=>"111101011",
  56529=>"001110011",
  56530=>"000001001",
  56531=>"110000101",
  56532=>"000110010",
  56533=>"110110001",
  56534=>"110101100",
  56535=>"010101100",
  56536=>"011010000",
  56537=>"101100110",
  56538=>"111111000",
  56539=>"100100010",
  56540=>"001100001",
  56541=>"101110010",
  56542=>"011101100",
  56543=>"110000011",
  56544=>"101001000",
  56545=>"111101011",
  56546=>"000000010",
  56547=>"000111001",
  56548=>"010101111",
  56549=>"000001110",
  56550=>"111010100",
  56551=>"010100110",
  56552=>"100101010",
  56553=>"000011000",
  56554=>"011011101",
  56555=>"100001110",
  56556=>"000100100",
  56557=>"110000101",
  56558=>"000101011",
  56559=>"101001000",
  56560=>"100010110",
  56561=>"111110010",
  56562=>"100101111",
  56563=>"011110011",
  56564=>"011100000",
  56565=>"100101011",
  56566=>"110000111",
  56567=>"110100111",
  56568=>"001110110",
  56569=>"111001001",
  56570=>"000100100",
  56571=>"110100111",
  56572=>"101100101",
  56573=>"101011110",
  56574=>"100101010",
  56575=>"011010100",
  56576=>"101011011",
  56577=>"000001101",
  56578=>"101110011",
  56579=>"100100010",
  56580=>"000111000",
  56581=>"000000111",
  56582=>"000110010",
  56583=>"111001100",
  56584=>"000010101",
  56585=>"110100011",
  56586=>"010110011",
  56587=>"001101101",
  56588=>"101001001",
  56589=>"011001000",
  56590=>"100000111",
  56591=>"111110100",
  56592=>"111000000",
  56593=>"001110001",
  56594=>"001010011",
  56595=>"101110001",
  56596=>"111000101",
  56597=>"100100010",
  56598=>"011000101",
  56599=>"110001000",
  56600=>"100000111",
  56601=>"110100001",
  56602=>"001010000",
  56603=>"111101110",
  56604=>"001111111",
  56605=>"110000110",
  56606=>"101110001",
  56607=>"000000000",
  56608=>"110100001",
  56609=>"011110001",
  56610=>"100011100",
  56611=>"111011100",
  56612=>"000011111",
  56613=>"111100011",
  56614=>"100001100",
  56615=>"001001001",
  56616=>"000101010",
  56617=>"000010001",
  56618=>"010011001",
  56619=>"000111001",
  56620=>"111011011",
  56621=>"101111000",
  56622=>"101111011",
  56623=>"001110110",
  56624=>"001000000",
  56625=>"100001100",
  56626=>"111110011",
  56627=>"000001000",
  56628=>"110101110",
  56629=>"001101011",
  56630=>"011010000",
  56631=>"010000101",
  56632=>"001000000",
  56633=>"101110010",
  56634=>"000010011",
  56635=>"001111101",
  56636=>"101000101",
  56637=>"001100011",
  56638=>"110000111",
  56639=>"100001110",
  56640=>"100110101",
  56641=>"101011111",
  56642=>"110111111",
  56643=>"010010010",
  56644=>"100011100",
  56645=>"110010101",
  56646=>"101100000",
  56647=>"100110010",
  56648=>"110001011",
  56649=>"111010010",
  56650=>"111001001",
  56651=>"000111110",
  56652=>"100010001",
  56653=>"001100101",
  56654=>"101011100",
  56655=>"000111100",
  56656=>"110011011",
  56657=>"001111001",
  56658=>"001100111",
  56659=>"000000110",
  56660=>"000000101",
  56661=>"111001000",
  56662=>"110001010",
  56663=>"011100100",
  56664=>"001111000",
  56665=>"100100011",
  56666=>"110101110",
  56667=>"100000000",
  56668=>"110101101",
  56669=>"100000100",
  56670=>"110010110",
  56671=>"011010111",
  56672=>"000000001",
  56673=>"001111100",
  56674=>"000100000",
  56675=>"000001010",
  56676=>"101111010",
  56677=>"101011111",
  56678=>"000010101",
  56679=>"111101110",
  56680=>"000101001",
  56681=>"000101000",
  56682=>"111000101",
  56683=>"000100100",
  56684=>"111000110",
  56685=>"100000101",
  56686=>"001110101",
  56687=>"001111001",
  56688=>"000111110",
  56689=>"011111101",
  56690=>"001101111",
  56691=>"000111000",
  56692=>"000111011",
  56693=>"101001001",
  56694=>"001001000",
  56695=>"110000111",
  56696=>"000110001",
  56697=>"001111100",
  56698=>"111011000",
  56699=>"110000100",
  56700=>"100111010",
  56701=>"101110110",
  56702=>"111100111",
  56703=>"001001110",
  56704=>"101010101",
  56705=>"011101101",
  56706=>"001001111",
  56707=>"100100111",
  56708=>"111111000",
  56709=>"100111011",
  56710=>"010101001",
  56711=>"010000011",
  56712=>"001000001",
  56713=>"010010100",
  56714=>"010101100",
  56715=>"110011001",
  56716=>"101110101",
  56717=>"000001000",
  56718=>"110111001",
  56719=>"111111001",
  56720=>"001000011",
  56721=>"001011011",
  56722=>"111110000",
  56723=>"000110111",
  56724=>"100110100",
  56725=>"101101111",
  56726=>"011000010",
  56727=>"111011111",
  56728=>"001111010",
  56729=>"101001011",
  56730=>"101111000",
  56731=>"001100110",
  56732=>"100101010",
  56733=>"011001011",
  56734=>"101001100",
  56735=>"011000011",
  56736=>"000010010",
  56737=>"110110011",
  56738=>"011110100",
  56739=>"110001111",
  56740=>"111010001",
  56741=>"000011101",
  56742=>"000000110",
  56743=>"001000101",
  56744=>"011010110",
  56745=>"011000010",
  56746=>"010100010",
  56747=>"101011011",
  56748=>"100010110",
  56749=>"100100101",
  56750=>"000110100",
  56751=>"111110001",
  56752=>"001111011",
  56753=>"000100100",
  56754=>"011000001",
  56755=>"000111110",
  56756=>"110100011",
  56757=>"111011000",
  56758=>"100101101",
  56759=>"100101001",
  56760=>"011110110",
  56761=>"000111101",
  56762=>"100000001",
  56763=>"100001000",
  56764=>"111111100",
  56765=>"101011110",
  56766=>"001010000",
  56767=>"011100000",
  56768=>"111001111",
  56769=>"001001011",
  56770=>"100110101",
  56771=>"011011110",
  56772=>"101010000",
  56773=>"010100010",
  56774=>"000000011",
  56775=>"100001000",
  56776=>"110110011",
  56777=>"011111010",
  56778=>"011110001",
  56779=>"000011010",
  56780=>"000000011",
  56781=>"010110010",
  56782=>"000100100",
  56783=>"111100110",
  56784=>"110111001",
  56785=>"010100011",
  56786=>"111101101",
  56787=>"010110110",
  56788=>"110000111",
  56789=>"000100000",
  56790=>"000100000",
  56791=>"111110111",
  56792=>"011111000",
  56793=>"110010011",
  56794=>"101011001",
  56795=>"100100101",
  56796=>"000011011",
  56797=>"101001010",
  56798=>"100010101",
  56799=>"101111111",
  56800=>"001010101",
  56801=>"000100110",
  56802=>"000001010",
  56803=>"011011100",
  56804=>"010000111",
  56805=>"010011100",
  56806=>"100001000",
  56807=>"100010001",
  56808=>"000100011",
  56809=>"010000001",
  56810=>"000100011",
  56811=>"101001100",
  56812=>"101100100",
  56813=>"010101100",
  56814=>"000010101",
  56815=>"011111000",
  56816=>"101100000",
  56817=>"110001011",
  56818=>"101001010",
  56819=>"001010100",
  56820=>"011111111",
  56821=>"100001011",
  56822=>"100000010",
  56823=>"010110001",
  56824=>"110011111",
  56825=>"000110001",
  56826=>"100100101",
  56827=>"101111000",
  56828=>"111000101",
  56829=>"000001101",
  56830=>"111110101",
  56831=>"000001001",
  56832=>"001010001",
  56833=>"111111111",
  56834=>"101100111",
  56835=>"110111100",
  56836=>"101100110",
  56837=>"101100100",
  56838=>"011110100",
  56839=>"010111001",
  56840=>"111010011",
  56841=>"001101000",
  56842=>"100010110",
  56843=>"010010001",
  56844=>"000111100",
  56845=>"000100011",
  56846=>"100010000",
  56847=>"001011011",
  56848=>"101010001",
  56849=>"100111011",
  56850=>"010111010",
  56851=>"110101000",
  56852=>"010101000",
  56853=>"100011101",
  56854=>"111011010",
  56855=>"110111110",
  56856=>"010011010",
  56857=>"011100001",
  56858=>"000010000",
  56859=>"001111010",
  56860=>"000100000",
  56861=>"100000000",
  56862=>"101100000",
  56863=>"010110001",
  56864=>"011110111",
  56865=>"110001010",
  56866=>"000011011",
  56867=>"110101010",
  56868=>"110101101",
  56869=>"101010101",
  56870=>"111000010",
  56871=>"000111101",
  56872=>"001110100",
  56873=>"101110001",
  56874=>"110001011",
  56875=>"100010010",
  56876=>"001011101",
  56877=>"010101000",
  56878=>"111010000",
  56879=>"111000000",
  56880=>"001100011",
  56881=>"000010101",
  56882=>"001000010",
  56883=>"011010010",
  56884=>"110010010",
  56885=>"010101110",
  56886=>"010001111",
  56887=>"111001101",
  56888=>"001100100",
  56889=>"101011011",
  56890=>"010011100",
  56891=>"011111000",
  56892=>"010101110",
  56893=>"010111101",
  56894=>"111000100",
  56895=>"100110011",
  56896=>"000011111",
  56897=>"011101101",
  56898=>"101010010",
  56899=>"001000000",
  56900=>"101100111",
  56901=>"000001000",
  56902=>"000101001",
  56903=>"000101110",
  56904=>"101111100",
  56905=>"100011001",
  56906=>"001110010",
  56907=>"100101111",
  56908=>"110111110",
  56909=>"110011011",
  56910=>"000010111",
  56911=>"001011000",
  56912=>"101001111",
  56913=>"111001110",
  56914=>"000010100",
  56915=>"110110110",
  56916=>"001101011",
  56917=>"000101110",
  56918=>"011100101",
  56919=>"010001010",
  56920=>"101110111",
  56921=>"011110011",
  56922=>"101101001",
  56923=>"011011001",
  56924=>"000111100",
  56925=>"110000100",
  56926=>"010100001",
  56927=>"010100101",
  56928=>"001001110",
  56929=>"001011001",
  56930=>"010010100",
  56931=>"111111100",
  56932=>"001000000",
  56933=>"001000100",
  56934=>"110011101",
  56935=>"100100111",
  56936=>"001010011",
  56937=>"001101110",
  56938=>"111011110",
  56939=>"001110111",
  56940=>"100111001",
  56941=>"110001010",
  56942=>"110110111",
  56943=>"111001101",
  56944=>"101000011",
  56945=>"011110110",
  56946=>"100111000",
  56947=>"010001000",
  56948=>"010110101",
  56949=>"000101001",
  56950=>"011001000",
  56951=>"101000100",
  56952=>"111100001",
  56953=>"111011000",
  56954=>"111101011",
  56955=>"001001110",
  56956=>"011100110",
  56957=>"100001110",
  56958=>"100111111",
  56959=>"011110111",
  56960=>"111001000",
  56961=>"110110010",
  56962=>"100010111",
  56963=>"001000101",
  56964=>"101101100",
  56965=>"000111011",
  56966=>"010001101",
  56967=>"101001000",
  56968=>"101001000",
  56969=>"100000100",
  56970=>"010011001",
  56971=>"101101101",
  56972=>"000001110",
  56973=>"000000100",
  56974=>"111001001",
  56975=>"011111100",
  56976=>"101100000",
  56977=>"101110001",
  56978=>"101101011",
  56979=>"011100000",
  56980=>"101111111",
  56981=>"001111110",
  56982=>"100111100",
  56983=>"101000100",
  56984=>"111011001",
  56985=>"001011000",
  56986=>"000000001",
  56987=>"001010000",
  56988=>"100101010",
  56989=>"111100111",
  56990=>"011100101",
  56991=>"000000110",
  56992=>"101111110",
  56993=>"101011011",
  56994=>"000000011",
  56995=>"010111101",
  56996=>"100111100",
  56997=>"001010011",
  56998=>"111000100",
  56999=>"010100010",
  57000=>"100101000",
  57001=>"110000000",
  57002=>"011000100",
  57003=>"000110000",
  57004=>"110000000",
  57005=>"101001110",
  57006=>"100010000",
  57007=>"100010111",
  57008=>"000101110",
  57009=>"101100000",
  57010=>"110111010",
  57011=>"100111110",
  57012=>"011100111",
  57013=>"101111110",
  57014=>"111110000",
  57015=>"011000010",
  57016=>"100000001",
  57017=>"100011010",
  57018=>"001101011",
  57019=>"001001001",
  57020=>"010001001",
  57021=>"000110001",
  57022=>"010101011",
  57023=>"000011011",
  57024=>"001111011",
  57025=>"101001001",
  57026=>"000011101",
  57027=>"000101100",
  57028=>"000110111",
  57029=>"001010110",
  57030=>"010100010",
  57031=>"110110101",
  57032=>"111011110",
  57033=>"111101010",
  57034=>"100101111",
  57035=>"011100100",
  57036=>"000111111",
  57037=>"111111101",
  57038=>"100100101",
  57039=>"110000100",
  57040=>"101111010",
  57041=>"011011110",
  57042=>"100000000",
  57043=>"011001011",
  57044=>"101100100",
  57045=>"010110111",
  57046=>"100001110",
  57047=>"110110010",
  57048=>"111100110",
  57049=>"001100100",
  57050=>"100001001",
  57051=>"111000101",
  57052=>"000111011",
  57053=>"110110111",
  57054=>"101110001",
  57055=>"100111111",
  57056=>"000101110",
  57057=>"010100100",
  57058=>"011011100",
  57059=>"010011011",
  57060=>"101010111",
  57061=>"111010101",
  57062=>"011100100",
  57063=>"001000011",
  57064=>"101010101",
  57065=>"111001111",
  57066=>"011110011",
  57067=>"100110010",
  57068=>"000100101",
  57069=>"000111100",
  57070=>"011100011",
  57071=>"001110011",
  57072=>"011111010",
  57073=>"110111101",
  57074=>"100100110",
  57075=>"110101001",
  57076=>"100010111",
  57077=>"010001101",
  57078=>"111111101",
  57079=>"111011111",
  57080=>"110010100",
  57081=>"110110010",
  57082=>"110000000",
  57083=>"000010100",
  57084=>"000000111",
  57085=>"100111000",
  57086=>"111111101",
  57087=>"000100010",
  57088=>"000000100",
  57089=>"100010100",
  57090=>"101010001",
  57091=>"001100000",
  57092=>"101111011",
  57093=>"111000101",
  57094=>"111110000",
  57095=>"011101011",
  57096=>"101001001",
  57097=>"000100111",
  57098=>"011100111",
  57099=>"010011011",
  57100=>"001001100",
  57101=>"011010001",
  57102=>"010110101",
  57103=>"001111110",
  57104=>"100001001",
  57105=>"110101011",
  57106=>"011000001",
  57107=>"111110100",
  57108=>"111101101",
  57109=>"101111101",
  57110=>"101111010",
  57111=>"010011000",
  57112=>"000101111",
  57113=>"001101111",
  57114=>"011001110",
  57115=>"001101001",
  57116=>"111010010",
  57117=>"100101010",
  57118=>"101110001",
  57119=>"001001101",
  57120=>"110011101",
  57121=>"001011011",
  57122=>"101000010",
  57123=>"001101010",
  57124=>"100100110",
  57125=>"000100101",
  57126=>"110010010",
  57127=>"100100101",
  57128=>"011111110",
  57129=>"011010010",
  57130=>"110111101",
  57131=>"101100010",
  57132=>"011001000",
  57133=>"110010001",
  57134=>"010110000",
  57135=>"110111110",
  57136=>"000010100",
  57137=>"101001111",
  57138=>"001110000",
  57139=>"111101011",
  57140=>"011001110",
  57141=>"110000011",
  57142=>"100110010",
  57143=>"001100111",
  57144=>"110001000",
  57145=>"010000000",
  57146=>"000100111",
  57147=>"001110000",
  57148=>"001001010",
  57149=>"000011011",
  57150=>"100101001",
  57151=>"100111111",
  57152=>"100001111",
  57153=>"101001010",
  57154=>"000010111",
  57155=>"111111000",
  57156=>"000011001",
  57157=>"011111101",
  57158=>"000011111",
  57159=>"100110111",
  57160=>"001100000",
  57161=>"011001001",
  57162=>"001111001",
  57163=>"111011110",
  57164=>"000110010",
  57165=>"011001100",
  57166=>"100011001",
  57167=>"011001111",
  57168=>"000010011",
  57169=>"110111111",
  57170=>"111111010",
  57171=>"000100110",
  57172=>"110001100",
  57173=>"000011111",
  57174=>"100100001",
  57175=>"011011000",
  57176=>"110100101",
  57177=>"100000011",
  57178=>"101111001",
  57179=>"011000101",
  57180=>"011100110",
  57181=>"000110111",
  57182=>"011101001",
  57183=>"101001010",
  57184=>"001011001",
  57185=>"010010100",
  57186=>"111111011",
  57187=>"011010011",
  57188=>"100011111",
  57189=>"110000111",
  57190=>"000001111",
  57191=>"110011001",
  57192=>"011110011",
  57193=>"111011011",
  57194=>"001100001",
  57195=>"011111010",
  57196=>"111000110",
  57197=>"010011111",
  57198=>"010111010",
  57199=>"111001010",
  57200=>"101111011",
  57201=>"110010110",
  57202=>"001011010",
  57203=>"011110001",
  57204=>"001100010",
  57205=>"100100111",
  57206=>"001001011",
  57207=>"001110111",
  57208=>"010110101",
  57209=>"010100111",
  57210=>"111111111",
  57211=>"100000011",
  57212=>"001011111",
  57213=>"001110011",
  57214=>"000100101",
  57215=>"010101101",
  57216=>"010010110",
  57217=>"101100000",
  57218=>"000000010",
  57219=>"010110100",
  57220=>"010010010",
  57221=>"011100000",
  57222=>"000101011",
  57223=>"101111101",
  57224=>"000010011",
  57225=>"000110111",
  57226=>"110111000",
  57227=>"001101111",
  57228=>"101011000",
  57229=>"100000011",
  57230=>"100111100",
  57231=>"110100001",
  57232=>"110000110",
  57233=>"110110000",
  57234=>"101001010",
  57235=>"101100011",
  57236=>"001100110",
  57237=>"001100101",
  57238=>"010010000",
  57239=>"011000110",
  57240=>"010100110",
  57241=>"111100011",
  57242=>"000100000",
  57243=>"000110110",
  57244=>"100010110",
  57245=>"111101011",
  57246=>"001110100",
  57247=>"001001101",
  57248=>"110010100",
  57249=>"011100110",
  57250=>"001000001",
  57251=>"111111111",
  57252=>"010001010",
  57253=>"011110001",
  57254=>"001101110",
  57255=>"110011100",
  57256=>"001011001",
  57257=>"001010000",
  57258=>"100001101",
  57259=>"111100111",
  57260=>"011100101",
  57261=>"110011101",
  57262=>"110010000",
  57263=>"011101111",
  57264=>"111010101",
  57265=>"111011100",
  57266=>"101110100",
  57267=>"010001001",
  57268=>"111100110",
  57269=>"000011110",
  57270=>"101011000",
  57271=>"010110101",
  57272=>"010010101",
  57273=>"100111101",
  57274=>"001111110",
  57275=>"100001111",
  57276=>"000110010",
  57277=>"000111110",
  57278=>"000001011",
  57279=>"000011011",
  57280=>"010111011",
  57281=>"101100010",
  57282=>"000011010",
  57283=>"011101000",
  57284=>"100110011",
  57285=>"100011010",
  57286=>"001111000",
  57287=>"110111010",
  57288=>"100001000",
  57289=>"111101111",
  57290=>"010011100",
  57291=>"010111111",
  57292=>"110110110",
  57293=>"001001011",
  57294=>"100001010",
  57295=>"110110111",
  57296=>"000110011",
  57297=>"010011011",
  57298=>"111111011",
  57299=>"000100110",
  57300=>"001111110",
  57301=>"010010001",
  57302=>"011110110",
  57303=>"001111000",
  57304=>"000110110",
  57305=>"101010000",
  57306=>"001110000",
  57307=>"010100001",
  57308=>"101110001",
  57309=>"100011011",
  57310=>"110101100",
  57311=>"001000011",
  57312=>"000001101",
  57313=>"000110100",
  57314=>"100111110",
  57315=>"110110111",
  57316=>"101010010",
  57317=>"110101010",
  57318=>"000010000",
  57319=>"100001000",
  57320=>"010001100",
  57321=>"011110101",
  57322=>"100001101",
  57323=>"110010011",
  57324=>"001011010",
  57325=>"011010111",
  57326=>"011000001",
  57327=>"001000100",
  57328=>"101010001",
  57329=>"011111101",
  57330=>"001010111",
  57331=>"110111110",
  57332=>"010000000",
  57333=>"010001000",
  57334=>"110111010",
  57335=>"101011111",
  57336=>"011001011",
  57337=>"111001010",
  57338=>"001100011",
  57339=>"101000011",
  57340=>"010100111",
  57341=>"111111100",
  57342=>"111110000",
  57343=>"010011010",
  57344=>"111101001",
  57345=>"010010001",
  57346=>"010110110",
  57347=>"100001010",
  57348=>"100101110",
  57349=>"011000101",
  57350=>"101110110",
  57351=>"111110110",
  57352=>"110010011",
  57353=>"101111111",
  57354=>"010000000",
  57355=>"001100011",
  57356=>"010101101",
  57357=>"001100111",
  57358=>"010001111",
  57359=>"111101011",
  57360=>"001110001",
  57361=>"100010110",
  57362=>"011101101",
  57363=>"000100100",
  57364=>"011100011",
  57365=>"000000011",
  57366=>"110110011",
  57367=>"010011010",
  57368=>"011011100",
  57369=>"101100010",
  57370=>"010101000",
  57371=>"000010111",
  57372=>"000000000",
  57373=>"001001001",
  57374=>"000010111",
  57375=>"101101110",
  57376=>"000010011",
  57377=>"001000011",
  57378=>"111101001",
  57379=>"100001010",
  57380=>"000010111",
  57381=>"011010101",
  57382=>"001111111",
  57383=>"011101100",
  57384=>"001011111",
  57385=>"111011111",
  57386=>"001110101",
  57387=>"000001010",
  57388=>"000100100",
  57389=>"011000101",
  57390=>"011110001",
  57391=>"111011011",
  57392=>"100010010",
  57393=>"010101101",
  57394=>"100100100",
  57395=>"100101000",
  57396=>"001110110",
  57397=>"001010100",
  57398=>"101111010",
  57399=>"110001011",
  57400=>"111101100",
  57401=>"000000010",
  57402=>"000011101",
  57403=>"101010010",
  57404=>"111101111",
  57405=>"011001001",
  57406=>"001010100",
  57407=>"101101111",
  57408=>"000000110",
  57409=>"000000000",
  57410=>"100111111",
  57411=>"001001110",
  57412=>"110000110",
  57413=>"001011100",
  57414=>"010000111",
  57415=>"100011011",
  57416=>"011111100",
  57417=>"011110100",
  57418=>"001101101",
  57419=>"001010000",
  57420=>"110001101",
  57421=>"000000001",
  57422=>"111100010",
  57423=>"010111101",
  57424=>"111110100",
  57425=>"000000011",
  57426=>"011001110",
  57427=>"011011111",
  57428=>"001110011",
  57429=>"110000111",
  57430=>"111010110",
  57431=>"011111001",
  57432=>"110101110",
  57433=>"011100000",
  57434=>"111111111",
  57435=>"000101010",
  57436=>"011010110",
  57437=>"110110111",
  57438=>"110000001",
  57439=>"000001011",
  57440=>"000110111",
  57441=>"100110101",
  57442=>"101011000",
  57443=>"000111111",
  57444=>"000000010",
  57445=>"100011100",
  57446=>"111011010",
  57447=>"100111010",
  57448=>"100110100",
  57449=>"110000111",
  57450=>"111111100",
  57451=>"100010110",
  57452=>"010100001",
  57453=>"000100101",
  57454=>"110111110",
  57455=>"000111010",
  57456=>"000100000",
  57457=>"100011101",
  57458=>"000111100",
  57459=>"000100000",
  57460=>"111101100",
  57461=>"111001111",
  57462=>"111101110",
  57463=>"101010110",
  57464=>"001101011",
  57465=>"001100010",
  57466=>"010100110",
  57467=>"101010100",
  57468=>"110001011",
  57469=>"011110110",
  57470=>"010110110",
  57471=>"011101011",
  57472=>"011100010",
  57473=>"011101100",
  57474=>"010011000",
  57475=>"110110000",
  57476=>"100100101",
  57477=>"100000011",
  57478=>"010101111",
  57479=>"000111111",
  57480=>"000100000",
  57481=>"111010110",
  57482=>"001001011",
  57483=>"010001111",
  57484=>"101011110",
  57485=>"100110111",
  57486=>"111001001",
  57487=>"101011010",
  57488=>"101000000",
  57489=>"101011001",
  57490=>"100010100",
  57491=>"000001010",
  57492=>"001111101",
  57493=>"101111101",
  57494=>"011110111",
  57495=>"000110101",
  57496=>"011010100",
  57497=>"100111111",
  57498=>"111001010",
  57499=>"111000001",
  57500=>"110111101",
  57501=>"111010010",
  57502=>"100000110",
  57503=>"010100001",
  57504=>"000010001",
  57505=>"111111110",
  57506=>"111011000",
  57507=>"001001111",
  57508=>"100101010",
  57509=>"000001000",
  57510=>"010111011",
  57511=>"011101001",
  57512=>"000101111",
  57513=>"110000011",
  57514=>"101010001",
  57515=>"110010000",
  57516=>"000010110",
  57517=>"100111000",
  57518=>"111001010",
  57519=>"100001110",
  57520=>"100000010",
  57521=>"110010011",
  57522=>"000101010",
  57523=>"101000000",
  57524=>"010100011",
  57525=>"011100000",
  57526=>"010000011",
  57527=>"111000011",
  57528=>"010111110",
  57529=>"100001010",
  57530=>"111001101",
  57531=>"010111111",
  57532=>"101110010",
  57533=>"101011111",
  57534=>"010111000",
  57535=>"000011111",
  57536=>"011011011",
  57537=>"110110110",
  57538=>"010001000",
  57539=>"000000000",
  57540=>"101000010",
  57541=>"100111010",
  57542=>"000000010",
  57543=>"111110111",
  57544=>"101111101",
  57545=>"111010000",
  57546=>"110000001",
  57547=>"000011110",
  57548=>"110001100",
  57549=>"111000001",
  57550=>"100110001",
  57551=>"010100010",
  57552=>"100001000",
  57553=>"010011001",
  57554=>"101011100",
  57555=>"100001000",
  57556=>"110100001",
  57557=>"101110101",
  57558=>"010011101",
  57559=>"111100010",
  57560=>"011010000",
  57561=>"010010110",
  57562=>"010000100",
  57563=>"000101010",
  57564=>"010001000",
  57565=>"110011100",
  57566=>"100001010",
  57567=>"111001011",
  57568=>"001001100",
  57569=>"111110010",
  57570=>"100011100",
  57571=>"111110001",
  57572=>"111001100",
  57573=>"000100011",
  57574=>"000000001",
  57575=>"011101011",
  57576=>"010101100",
  57577=>"111101001",
  57578=>"000010101",
  57579=>"010010000",
  57580=>"000001001",
  57581=>"100010111",
  57582=>"011001100",
  57583=>"110011101",
  57584=>"010001100",
  57585=>"100010000",
  57586=>"110110001",
  57587=>"110001100",
  57588=>"010011101",
  57589=>"100111011",
  57590=>"010001011",
  57591=>"100000011",
  57592=>"011000001",
  57593=>"010011000",
  57594=>"101100100",
  57595=>"110111000",
  57596=>"101001101",
  57597=>"000001000",
  57598=>"001100111",
  57599=>"100010000",
  57600=>"110011000",
  57601=>"101001011",
  57602=>"001001000",
  57603=>"110000111",
  57604=>"011010110",
  57605=>"100011111",
  57606=>"000110101",
  57607=>"111111100",
  57608=>"100011001",
  57609=>"111100111",
  57610=>"010011111",
  57611=>"001101001",
  57612=>"111111011",
  57613=>"001011010",
  57614=>"010101101",
  57615=>"110011100",
  57616=>"110111010",
  57617=>"100101001",
  57618=>"110000101",
  57619=>"000110100",
  57620=>"110111101",
  57621=>"110101111",
  57622=>"100100100",
  57623=>"001110100",
  57624=>"011000011",
  57625=>"010110101",
  57626=>"101010101",
  57627=>"010001110",
  57628=>"000101110",
  57629=>"011101111",
  57630=>"000010111",
  57631=>"010111111",
  57632=>"111011100",
  57633=>"111001111",
  57634=>"011000110",
  57635=>"011000110",
  57636=>"000101011",
  57637=>"100110110",
  57638=>"111110111",
  57639=>"010001011",
  57640=>"010011100",
  57641=>"110001000",
  57642=>"000100100",
  57643=>"011011100",
  57644=>"011111110",
  57645=>"011111101",
  57646=>"110111111",
  57647=>"110111001",
  57648=>"100010101",
  57649=>"110110111",
  57650=>"101110111",
  57651=>"110010111",
  57652=>"111011001",
  57653=>"100011010",
  57654=>"001011010",
  57655=>"100011000",
  57656=>"100011101",
  57657=>"010111100",
  57658=>"010001001",
  57659=>"011110010",
  57660=>"011110011",
  57661=>"100001001",
  57662=>"110001110",
  57663=>"010111011",
  57664=>"010001001",
  57665=>"111111111",
  57666=>"110000110",
  57667=>"110011010",
  57668=>"111110100",
  57669=>"010011110",
  57670=>"001110111",
  57671=>"101101110",
  57672=>"100100101",
  57673=>"110111010",
  57674=>"100101001",
  57675=>"001001111",
  57676=>"110001101",
  57677=>"010101101",
  57678=>"111110110",
  57679=>"010001011",
  57680=>"011011001",
  57681=>"001110111",
  57682=>"011010001",
  57683=>"001110110",
  57684=>"001001101",
  57685=>"101100000",
  57686=>"111111011",
  57687=>"010110001",
  57688=>"110010010",
  57689=>"101100010",
  57690=>"000011001",
  57691=>"101100100",
  57692=>"001010010",
  57693=>"110110111",
  57694=>"100000111",
  57695=>"010111101",
  57696=>"100011000",
  57697=>"000010010",
  57698=>"000011001",
  57699=>"100101101",
  57700=>"001010110",
  57701=>"101111110",
  57702=>"000000101",
  57703=>"001110100",
  57704=>"111111101",
  57705=>"010101111",
  57706=>"000101100",
  57707=>"111111110",
  57708=>"111010111",
  57709=>"110110011",
  57710=>"100111011",
  57711=>"000100001",
  57712=>"101010010",
  57713=>"101001101",
  57714=>"001000100",
  57715=>"111100001",
  57716=>"110101011",
  57717=>"000010101",
  57718=>"111000010",
  57719=>"001010001",
  57720=>"101110110",
  57721=>"010011100",
  57722=>"000100011",
  57723=>"110011111",
  57724=>"111101000",
  57725=>"100000011",
  57726=>"101011010",
  57727=>"011011001",
  57728=>"000000101",
  57729=>"010100000",
  57730=>"100111110",
  57731=>"111010101",
  57732=>"110100000",
  57733=>"101101111",
  57734=>"110100011",
  57735=>"101100111",
  57736=>"010011011",
  57737=>"011000101",
  57738=>"011011010",
  57739=>"000000010",
  57740=>"011111111",
  57741=>"000000101",
  57742=>"000011011",
  57743=>"101100000",
  57744=>"111100100",
  57745=>"001100000",
  57746=>"111100100",
  57747=>"000101100",
  57748=>"110000011",
  57749=>"100100111",
  57750=>"101010101",
  57751=>"000000100",
  57752=>"010111001",
  57753=>"101010101",
  57754=>"100010100",
  57755=>"011111010",
  57756=>"111101011",
  57757=>"001110001",
  57758=>"110001011",
  57759=>"111111101",
  57760=>"000100100",
  57761=>"110100110",
  57762=>"110100001",
  57763=>"111100001",
  57764=>"110101000",
  57765=>"111110001",
  57766=>"010010010",
  57767=>"010110001",
  57768=>"010001001",
  57769=>"110111110",
  57770=>"111001010",
  57771=>"100100111",
  57772=>"111010000",
  57773=>"101001001",
  57774=>"111111001",
  57775=>"110110011",
  57776=>"111111011",
  57777=>"010101101",
  57778=>"111011100",
  57779=>"100110000",
  57780=>"110011000",
  57781=>"000110010",
  57782=>"010001001",
  57783=>"101011000",
  57784=>"011000001",
  57785=>"111110111",
  57786=>"011010010",
  57787=>"111010001",
  57788=>"000010100",
  57789=>"000010011",
  57790=>"001010111",
  57791=>"010100000",
  57792=>"000101100",
  57793=>"010100001",
  57794=>"001001011",
  57795=>"100110101",
  57796=>"000000100",
  57797=>"111111100",
  57798=>"001010111",
  57799=>"000001100",
  57800=>"011010010",
  57801=>"000011010",
  57802=>"001000111",
  57803=>"011111100",
  57804=>"111110011",
  57805=>"010111100",
  57806=>"101010100",
  57807=>"100101100",
  57808=>"100111011",
  57809=>"001010100",
  57810=>"100110000",
  57811=>"000100110",
  57812=>"111110110",
  57813=>"110111010",
  57814=>"011100010",
  57815=>"110111101",
  57816=>"111010001",
  57817=>"110110110",
  57818=>"110001001",
  57819=>"111111110",
  57820=>"101000110",
  57821=>"111110011",
  57822=>"011111000",
  57823=>"010001101",
  57824=>"000100001",
  57825=>"100000001",
  57826=>"110010100",
  57827=>"011110111",
  57828=>"100101010",
  57829=>"011000100",
  57830=>"100000101",
  57831=>"101111011",
  57832=>"111000111",
  57833=>"101100001",
  57834=>"010110010",
  57835=>"111011111",
  57836=>"011101101",
  57837=>"001100001",
  57838=>"010100101",
  57839=>"000001111",
  57840=>"110010111",
  57841=>"011100011",
  57842=>"100011100",
  57843=>"011011000",
  57844=>"111010011",
  57845=>"100011011",
  57846=>"010011001",
  57847=>"111011011",
  57848=>"111000111",
  57849=>"001000011",
  57850=>"010011010",
  57851=>"011011111",
  57852=>"100111000",
  57853=>"000010110",
  57854=>"011101101",
  57855=>"010111011",
  57856=>"011000111",
  57857=>"001011011",
  57858=>"001101001",
  57859=>"010111110",
  57860=>"100110100",
  57861=>"001110110",
  57862=>"010110011",
  57863=>"101100100",
  57864=>"010111110",
  57865=>"110110110",
  57866=>"101010110",
  57867=>"011010000",
  57868=>"011011100",
  57869=>"010001110",
  57870=>"010010000",
  57871=>"111111010",
  57872=>"111101101",
  57873=>"001101100",
  57874=>"000001010",
  57875=>"010100000",
  57876=>"101111000",
  57877=>"110001011",
  57878=>"101110111",
  57879=>"110011100",
  57880=>"111111010",
  57881=>"111001100",
  57882=>"111001111",
  57883=>"101001010",
  57884=>"000010101",
  57885=>"010100100",
  57886=>"011111111",
  57887=>"001001100",
  57888=>"111000001",
  57889=>"011011010",
  57890=>"111111111",
  57891=>"110101000",
  57892=>"110011001",
  57893=>"101000011",
  57894=>"011101001",
  57895=>"010001100",
  57896=>"110111010",
  57897=>"001100100",
  57898=>"110110110",
  57899=>"000110011",
  57900=>"010010110",
  57901=>"101000110",
  57902=>"101000111",
  57903=>"100100001",
  57904=>"110110000",
  57905=>"100001101",
  57906=>"111101000",
  57907=>"000000000",
  57908=>"001111100",
  57909=>"100110010",
  57910=>"100000101",
  57911=>"000100010",
  57912=>"010000110",
  57913=>"100100011",
  57914=>"011010110",
  57915=>"111110001",
  57916=>"110100100",
  57917=>"100001011",
  57918=>"001000100",
  57919=>"010101010",
  57920=>"100100011",
  57921=>"011111000",
  57922=>"101101111",
  57923=>"110111011",
  57924=>"110110011",
  57925=>"001011010",
  57926=>"100001101",
  57927=>"111100111",
  57928=>"101100111",
  57929=>"100111100",
  57930=>"110001101",
  57931=>"001101110",
  57932=>"111101001",
  57933=>"001011111",
  57934=>"000001100",
  57935=>"100111100",
  57936=>"110010010",
  57937=>"001010101",
  57938=>"001110111",
  57939=>"010000101",
  57940=>"111010110",
  57941=>"100000010",
  57942=>"100011100",
  57943=>"110011011",
  57944=>"011010100",
  57945=>"000111101",
  57946=>"101111000",
  57947=>"011101011",
  57948=>"011000110",
  57949=>"100010110",
  57950=>"111100010",
  57951=>"010101001",
  57952=>"000001101",
  57953=>"001111001",
  57954=>"110110100",
  57955=>"111001111",
  57956=>"111101011",
  57957=>"100010100",
  57958=>"101010101",
  57959=>"110100010",
  57960=>"111000111",
  57961=>"110011110",
  57962=>"011100101",
  57963=>"101001001",
  57964=>"011110101",
  57965=>"110111000",
  57966=>"100001000",
  57967=>"100100000",
  57968=>"100111100",
  57969=>"111001110",
  57970=>"100110010",
  57971=>"001100111",
  57972=>"110101111",
  57973=>"001011001",
  57974=>"111010110",
  57975=>"001000011",
  57976=>"010000110",
  57977=>"111110010",
  57978=>"101110110",
  57979=>"010000011",
  57980=>"111001011",
  57981=>"100101101",
  57982=>"110101100",
  57983=>"101110100",
  57984=>"110001111",
  57985=>"010101010",
  57986=>"001111111",
  57987=>"100001111",
  57988=>"001010000",
  57989=>"010111011",
  57990=>"110110111",
  57991=>"000010110",
  57992=>"101011101",
  57993=>"000100111",
  57994=>"111101100",
  57995=>"000000110",
  57996=>"100001001",
  57997=>"111011011",
  57998=>"100011011",
  57999=>"110011010",
  58000=>"000011110",
  58001=>"001001101",
  58002=>"011001110",
  58003=>"100100000",
  58004=>"101111110",
  58005=>"110010011",
  58006=>"000010010",
  58007=>"111101000",
  58008=>"010111101",
  58009=>"100001111",
  58010=>"110001100",
  58011=>"101111000",
  58012=>"000101011",
  58013=>"000000100",
  58014=>"001110110",
  58015=>"011010111",
  58016=>"000011110",
  58017=>"001001100",
  58018=>"001000010",
  58019=>"011010101",
  58020=>"100101101",
  58021=>"001100110",
  58022=>"110101111",
  58023=>"101010010",
  58024=>"101011010",
  58025=>"001011110",
  58026=>"000001101",
  58027=>"001101000",
  58028=>"001010001",
  58029=>"111000100",
  58030=>"000001101",
  58031=>"111111001",
  58032=>"001000101",
  58033=>"000010111",
  58034=>"001100110",
  58035=>"110001000",
  58036=>"101001010",
  58037=>"101100010",
  58038=>"110100010",
  58039=>"011000011",
  58040=>"100001111",
  58041=>"011000100",
  58042=>"010011000",
  58043=>"001100000",
  58044=>"101101110",
  58045=>"001101101",
  58046=>"100111011",
  58047=>"111111100",
  58048=>"001101010",
  58049=>"100111000",
  58050=>"011101100",
  58051=>"111111101",
  58052=>"101100001",
  58053=>"111011011",
  58054=>"111101000",
  58055=>"000110111",
  58056=>"111010010",
  58057=>"111110000",
  58058=>"011011011",
  58059=>"100000111",
  58060=>"011011100",
  58061=>"011111001",
  58062=>"000101001",
  58063=>"100000011",
  58064=>"010010000",
  58065=>"010011111",
  58066=>"011000111",
  58067=>"100101011",
  58068=>"001010110",
  58069=>"001111100",
  58070=>"110000110",
  58071=>"001000010",
  58072=>"101101111",
  58073=>"100101000",
  58074=>"010100000",
  58075=>"001000000",
  58076=>"110010110",
  58077=>"100110110",
  58078=>"101011101",
  58079=>"011011110",
  58080=>"011000010",
  58081=>"000100101",
  58082=>"011001010",
  58083=>"100011001",
  58084=>"111111111",
  58085=>"001111111",
  58086=>"010111110",
  58087=>"001010110",
  58088=>"101110100",
  58089=>"110111100",
  58090=>"110100110",
  58091=>"111001010",
  58092=>"010101101",
  58093=>"101101010",
  58094=>"001000011",
  58095=>"011100000",
  58096=>"101000000",
  58097=>"101010101",
  58098=>"000100111",
  58099=>"111011100",
  58100=>"001000000",
  58101=>"100001101",
  58102=>"110010000",
  58103=>"111010000",
  58104=>"001111100",
  58105=>"010010110",
  58106=>"100000001",
  58107=>"000111101",
  58108=>"010000000",
  58109=>"101111101",
  58110=>"110111000",
  58111=>"010011110",
  58112=>"111001100",
  58113=>"101010111",
  58114=>"000010110",
  58115=>"000101001",
  58116=>"101111001",
  58117=>"011011110",
  58118=>"100101111",
  58119=>"000000000",
  58120=>"110101010",
  58121=>"010111011",
  58122=>"100010100",
  58123=>"000101110",
  58124=>"111010001",
  58125=>"001100010",
  58126=>"110010000",
  58127=>"000010010",
  58128=>"010111010",
  58129=>"111110100",
  58130=>"000111100",
  58131=>"001001001",
  58132=>"111100100",
  58133=>"100001100",
  58134=>"011001010",
  58135=>"010111110",
  58136=>"001101101",
  58137=>"011101000",
  58138=>"010010010",
  58139=>"001000010",
  58140=>"101011001",
  58141=>"010100111",
  58142=>"011010011",
  58143=>"010010001",
  58144=>"100110000",
  58145=>"001000110",
  58146=>"110010101",
  58147=>"101100001",
  58148=>"000100101",
  58149=>"000100111",
  58150=>"100010111",
  58151=>"011110100",
  58152=>"001100010",
  58153=>"001000011",
  58154=>"111111100",
  58155=>"101101100",
  58156=>"110111101",
  58157=>"100101110",
  58158=>"001111010",
  58159=>"000101111",
  58160=>"011010111",
  58161=>"100011101",
  58162=>"110111011",
  58163=>"010110100",
  58164=>"011111010",
  58165=>"111000011",
  58166=>"111110110",
  58167=>"000010011",
  58168=>"000101011",
  58169=>"111011101",
  58170=>"100111001",
  58171=>"001000111",
  58172=>"100110110",
  58173=>"000101000",
  58174=>"110101111",
  58175=>"101101111",
  58176=>"101110001",
  58177=>"100001110",
  58178=>"001001011",
  58179=>"000110010",
  58180=>"001101110",
  58181=>"101111000",
  58182=>"000000100",
  58183=>"101001000",
  58184=>"001010110",
  58185=>"100110001",
  58186=>"101001110",
  58187=>"100011111",
  58188=>"011011010",
  58189=>"101000100",
  58190=>"111110111",
  58191=>"111010011",
  58192=>"100010110",
  58193=>"010101000",
  58194=>"011000010",
  58195=>"110110110",
  58196=>"101010001",
  58197=>"001001110",
  58198=>"001111100",
  58199=>"011111000",
  58200=>"110010001",
  58201=>"011001101",
  58202=>"010100010",
  58203=>"010001101",
  58204=>"011011110",
  58205=>"110100110",
  58206=>"100000001",
  58207=>"011000111",
  58208=>"101100011",
  58209=>"000101101",
  58210=>"101110111",
  58211=>"010101101",
  58212=>"000100000",
  58213=>"011110001",
  58214=>"100000000",
  58215=>"100100001",
  58216=>"111011111",
  58217=>"010011110",
  58218=>"111111010",
  58219=>"100001001",
  58220=>"000101001",
  58221=>"000110011",
  58222=>"010101011",
  58223=>"111110111",
  58224=>"100000111",
  58225=>"110001111",
  58226=>"111011001",
  58227=>"001111100",
  58228=>"011111110",
  58229=>"110101001",
  58230=>"000111110",
  58231=>"110110111",
  58232=>"111101001",
  58233=>"001100000",
  58234=>"001111110",
  58235=>"111100001",
  58236=>"101000000",
  58237=>"001001000",
  58238=>"110011111",
  58239=>"010010111",
  58240=>"101001110",
  58241=>"000111100",
  58242=>"101001101",
  58243=>"101101100",
  58244=>"001110011",
  58245=>"110000011",
  58246=>"001100010",
  58247=>"001010011",
  58248=>"001000010",
  58249=>"011011011",
  58250=>"101101111",
  58251=>"111111011",
  58252=>"010010010",
  58253=>"001010111",
  58254=>"111101011",
  58255=>"001110100",
  58256=>"111111101",
  58257=>"000101011",
  58258=>"111111010",
  58259=>"100001101",
  58260=>"111010000",
  58261=>"011011111",
  58262=>"101101000",
  58263=>"010011011",
  58264=>"000000100",
  58265=>"101010111",
  58266=>"100100111",
  58267=>"111111010",
  58268=>"111110011",
  58269=>"111001000",
  58270=>"101110000",
  58271=>"010100011",
  58272=>"000000100",
  58273=>"111111101",
  58274=>"000001101",
  58275=>"111111111",
  58276=>"101011110",
  58277=>"000010000",
  58278=>"001110100",
  58279=>"000010000",
  58280=>"111100000",
  58281=>"100000000",
  58282=>"101111110",
  58283=>"010110001",
  58284=>"100101000",
  58285=>"111010101",
  58286=>"010101010",
  58287=>"011010000",
  58288=>"011001010",
  58289=>"000100110",
  58290=>"110000111",
  58291=>"011111100",
  58292=>"111101010",
  58293=>"010110110",
  58294=>"111001001",
  58295=>"010011111",
  58296=>"111110010",
  58297=>"001101101",
  58298=>"101001100",
  58299=>"101111010",
  58300=>"011000010",
  58301=>"001100000",
  58302=>"000111000",
  58303=>"110000010",
  58304=>"000101111",
  58305=>"100101110",
  58306=>"010001000",
  58307=>"111111100",
  58308=>"001010111",
  58309=>"000001110",
  58310=>"101000111",
  58311=>"100101111",
  58312=>"100011000",
  58313=>"001000111",
  58314=>"110100001",
  58315=>"110100000",
  58316=>"000001000",
  58317=>"101000111",
  58318=>"001000111",
  58319=>"110110011",
  58320=>"100110100",
  58321=>"111111111",
  58322=>"000001000",
  58323=>"100001000",
  58324=>"010010000",
  58325=>"100001110",
  58326=>"011100010",
  58327=>"000100011",
  58328=>"000110000",
  58329=>"110000010",
  58330=>"111111110",
  58331=>"011001001",
  58332=>"100000000",
  58333=>"010100000",
  58334=>"110101100",
  58335=>"111101101",
  58336=>"111011010",
  58337=>"111110011",
  58338=>"001010101",
  58339=>"001010001",
  58340=>"101011110",
  58341=>"000101000",
  58342=>"001111011",
  58343=>"111110010",
  58344=>"111011100",
  58345=>"101001000",
  58346=>"001110111",
  58347=>"111010011",
  58348=>"111001111",
  58349=>"010111010",
  58350=>"111111011",
  58351=>"011010111",
  58352=>"000110000",
  58353=>"101101110",
  58354=>"011001110",
  58355=>"010101010",
  58356=>"001010000",
  58357=>"101111110",
  58358=>"110111001",
  58359=>"101011111",
  58360=>"001011011",
  58361=>"110001010",
  58362=>"001111101",
  58363=>"000000000",
  58364=>"011100000",
  58365=>"010010010",
  58366=>"001001000",
  58367=>"000100111",
  58368=>"100000110",
  58369=>"110101111",
  58370=>"110000111",
  58371=>"011111111",
  58372=>"010100101",
  58373=>"010000011",
  58374=>"111110110",
  58375=>"010010100",
  58376=>"001110001",
  58377=>"001000010",
  58378=>"100011010",
  58379=>"001100001",
  58380=>"101110001",
  58381=>"101010111",
  58382=>"000111101",
  58383=>"110100001",
  58384=>"100000010",
  58385=>"011110001",
  58386=>"100111100",
  58387=>"110001010",
  58388=>"011000010",
  58389=>"111001100",
  58390=>"001100010",
  58391=>"111001100",
  58392=>"001011100",
  58393=>"010101010",
  58394=>"110110111",
  58395=>"101101111",
  58396=>"000010100",
  58397=>"000000000",
  58398=>"110011111",
  58399=>"100110001",
  58400=>"010001011",
  58401=>"101111101",
  58402=>"000000100",
  58403=>"110100000",
  58404=>"110111010",
  58405=>"011111110",
  58406=>"010010101",
  58407=>"110110000",
  58408=>"110010110",
  58409=>"011111011",
  58410=>"100011110",
  58411=>"110110101",
  58412=>"101110101",
  58413=>"101110001",
  58414=>"110111010",
  58415=>"000010101",
  58416=>"110101000",
  58417=>"101001110",
  58418=>"011111111",
  58419=>"011000000",
  58420=>"100011001",
  58421=>"111101010",
  58422=>"000111110",
  58423=>"000001111",
  58424=>"101101011",
  58425=>"000001100",
  58426=>"000101100",
  58427=>"101110100",
  58428=>"010010000",
  58429=>"001111001",
  58430=>"101101010",
  58431=>"101000011",
  58432=>"000100010",
  58433=>"011010000",
  58434=>"001010011",
  58435=>"100110110",
  58436=>"000101100",
  58437=>"111011001",
  58438=>"010101110",
  58439=>"100000000",
  58440=>"010010001",
  58441=>"100010101",
  58442=>"100001100",
  58443=>"110110110",
  58444=>"100111010",
  58445=>"011110010",
  58446=>"110001010",
  58447=>"000001100",
  58448=>"001110101",
  58449=>"101111011",
  58450=>"010000011",
  58451=>"101110111",
  58452=>"000111111",
  58453=>"010100001",
  58454=>"111010000",
  58455=>"000001001",
  58456=>"101001001",
  58457=>"000111111",
  58458=>"110000111",
  58459=>"101111000",
  58460=>"111111001",
  58461=>"000100100",
  58462=>"000110110",
  58463=>"100001110",
  58464=>"001000100",
  58465=>"000110110",
  58466=>"011101010",
  58467=>"100010001",
  58468=>"010101100",
  58469=>"000111100",
  58470=>"011110110",
  58471=>"011011001",
  58472=>"000011000",
  58473=>"001001000",
  58474=>"010110000",
  58475=>"101100111",
  58476=>"001111100",
  58477=>"000110110",
  58478=>"000011001",
  58479=>"011011101",
  58480=>"011000010",
  58481=>"101101111",
  58482=>"011001000",
  58483=>"110100010",
  58484=>"100111110",
  58485=>"100011001",
  58486=>"100110000",
  58487=>"010110100",
  58488=>"101010000",
  58489=>"101101011",
  58490=>"110001010",
  58491=>"001001000",
  58492=>"110111001",
  58493=>"010100001",
  58494=>"100011100",
  58495=>"001010000",
  58496=>"010110010",
  58497=>"111011011",
  58498=>"111010110",
  58499=>"001111011",
  58500=>"010001000",
  58501=>"010001111",
  58502=>"000011100",
  58503=>"101001010",
  58504=>"010100111",
  58505=>"000001110",
  58506=>"010101110",
  58507=>"010010001",
  58508=>"000111010",
  58509=>"100111010",
  58510=>"001110100",
  58511=>"111011110",
  58512=>"010111101",
  58513=>"010111000",
  58514=>"011010000",
  58515=>"101111101",
  58516=>"000010001",
  58517=>"101011001",
  58518=>"000010011",
  58519=>"111100101",
  58520=>"011110111",
  58521=>"100000110",
  58522=>"111001001",
  58523=>"101000011",
  58524=>"011101100",
  58525=>"011001000",
  58526=>"100110110",
  58527=>"110110011",
  58528=>"011011000",
  58529=>"011100011",
  58530=>"010010100",
  58531=>"001101111",
  58532=>"101111001",
  58533=>"001000110",
  58534=>"101111101",
  58535=>"100001000",
  58536=>"101000001",
  58537=>"010010111",
  58538=>"111001110",
  58539=>"110011001",
  58540=>"100000011",
  58541=>"111000001",
  58542=>"111100011",
  58543=>"001111010",
  58544=>"000011100",
  58545=>"011110100",
  58546=>"000100001",
  58547=>"011110110",
  58548=>"101110001",
  58549=>"000101100",
  58550=>"001010100",
  58551=>"111000100",
  58552=>"100111011",
  58553=>"111110011",
  58554=>"010111110",
  58555=>"010001111",
  58556=>"111110000",
  58557=>"100111011",
  58558=>"101010110",
  58559=>"100010111",
  58560=>"000000010",
  58561=>"010110001",
  58562=>"010100000",
  58563=>"000000000",
  58564=>"110010010",
  58565=>"100010011",
  58566=>"100001001",
  58567=>"110100000",
  58568=>"101000110",
  58569=>"111000100",
  58570=>"001110011",
  58571=>"000111011",
  58572=>"000000010",
  58573=>"101101101",
  58574=>"001000011",
  58575=>"011000001",
  58576=>"111101000",
  58577=>"001010110",
  58578=>"011011111",
  58579=>"100111011",
  58580=>"010010000",
  58581=>"011110101",
  58582=>"110000110",
  58583=>"001000110",
  58584=>"010000000",
  58585=>"010100011",
  58586=>"110101111",
  58587=>"100000010",
  58588=>"010110111",
  58589=>"101100111",
  58590=>"010101000",
  58591=>"010110110",
  58592=>"101000100",
  58593=>"000111110",
  58594=>"011000110",
  58595=>"000001010",
  58596=>"000011100",
  58597=>"000001110",
  58598=>"101111011",
  58599=>"011101011",
  58600=>"100010000",
  58601=>"010111101",
  58602=>"111101011",
  58603=>"010111011",
  58604=>"111000000",
  58605=>"101000011",
  58606=>"100000010",
  58607=>"011100001",
  58608=>"110100111",
  58609=>"110011101",
  58610=>"010010011",
  58611=>"100011011",
  58612=>"100010100",
  58613=>"111010101",
  58614=>"011011000",
  58615=>"100101010",
  58616=>"111111001",
  58617=>"001000100",
  58618=>"000101000",
  58619=>"101000101",
  58620=>"000110100",
  58621=>"001111110",
  58622=>"101110000",
  58623=>"000011111",
  58624=>"000110110",
  58625=>"111000111",
  58626=>"110000101",
  58627=>"000011000",
  58628=>"100100100",
  58629=>"001111011",
  58630=>"000011110",
  58631=>"000010110",
  58632=>"111111111",
  58633=>"111100101",
  58634=>"011011001",
  58635=>"110010110",
  58636=>"100110000",
  58637=>"001000100",
  58638=>"110000100",
  58639=>"011110101",
  58640=>"101011110",
  58641=>"010000011",
  58642=>"100111110",
  58643=>"100101101",
  58644=>"010100101",
  58645=>"010111010",
  58646=>"000100100",
  58647=>"110000110",
  58648=>"111011010",
  58649=>"111010010",
  58650=>"000101000",
  58651=>"111000101",
  58652=>"001001011",
  58653=>"011000111",
  58654=>"101111000",
  58655=>"011000010",
  58656=>"001001111",
  58657=>"001101111",
  58658=>"001101011",
  58659=>"011101110",
  58660=>"001010111",
  58661=>"110001110",
  58662=>"001011000",
  58663=>"101010111",
  58664=>"000111010",
  58665=>"100100101",
  58666=>"110011010",
  58667=>"110111010",
  58668=>"011000000",
  58669=>"111111110",
  58670=>"101100100",
  58671=>"000010001",
  58672=>"011001111",
  58673=>"110101101",
  58674=>"110111000",
  58675=>"000111110",
  58676=>"011101100",
  58677=>"101110111",
  58678=>"011010100",
  58679=>"010001000",
  58680=>"111000101",
  58681=>"111000000",
  58682=>"101101111",
  58683=>"111011010",
  58684=>"011000110",
  58685=>"001001010",
  58686=>"111101101",
  58687=>"111010111",
  58688=>"110001011",
  58689=>"001001001",
  58690=>"010111111",
  58691=>"101001001",
  58692=>"001011000",
  58693=>"100011111",
  58694=>"100011001",
  58695=>"100111000",
  58696=>"000011100",
  58697=>"111000000",
  58698=>"100000010",
  58699=>"000000100",
  58700=>"110101101",
  58701=>"111101011",
  58702=>"101100011",
  58703=>"011100101",
  58704=>"101000100",
  58705=>"110100000",
  58706=>"100010001",
  58707=>"100100001",
  58708=>"101010001",
  58709=>"011110011",
  58710=>"010011001",
  58711=>"110010010",
  58712=>"011101101",
  58713=>"100110010",
  58714=>"100110111",
  58715=>"011001001",
  58716=>"111010000",
  58717=>"110100001",
  58718=>"011001111",
  58719=>"011001010",
  58720=>"010001000",
  58721=>"101010011",
  58722=>"010001000",
  58723=>"011010111",
  58724=>"111011111",
  58725=>"011100101",
  58726=>"001100010",
  58727=>"111011110",
  58728=>"110010101",
  58729=>"111110000",
  58730=>"100000101",
  58731=>"101110011",
  58732=>"001101010",
  58733=>"101000101",
  58734=>"100100010",
  58735=>"000001011",
  58736=>"011011000",
  58737=>"110111101",
  58738=>"011001011",
  58739=>"111110100",
  58740=>"110110011",
  58741=>"100101011",
  58742=>"010011011",
  58743=>"000110010",
  58744=>"000011001",
  58745=>"111111101",
  58746=>"100110010",
  58747=>"011000111",
  58748=>"101001111",
  58749=>"111110111",
  58750=>"011001110",
  58751=>"001100100",
  58752=>"001101101",
  58753=>"100100000",
  58754=>"011010010",
  58755=>"000011011",
  58756=>"100101101",
  58757=>"111010100",
  58758=>"100001101",
  58759=>"000000011",
  58760=>"000001101",
  58761=>"001101100",
  58762=>"010101100",
  58763=>"110011110",
  58764=>"111111101",
  58765=>"000111110",
  58766=>"110010101",
  58767=>"011100010",
  58768=>"000001010",
  58769=>"000000000",
  58770=>"000000000",
  58771=>"000001110",
  58772=>"111111011",
  58773=>"000101010",
  58774=>"010101110",
  58775=>"111000011",
  58776=>"111100100",
  58777=>"001010110",
  58778=>"000010000",
  58779=>"010011000",
  58780=>"101111001",
  58781=>"110010000",
  58782=>"101010010",
  58783=>"000110001",
  58784=>"101101000",
  58785=>"010011000",
  58786=>"010110101",
  58787=>"011010101",
  58788=>"110111000",
  58789=>"100010000",
  58790=>"001000100",
  58791=>"000100101",
  58792=>"100001110",
  58793=>"011000101",
  58794=>"000001111",
  58795=>"000101100",
  58796=>"101100100",
  58797=>"001011010",
  58798=>"111101111",
  58799=>"111111011",
  58800=>"001010111",
  58801=>"100001001",
  58802=>"101110100",
  58803=>"011000001",
  58804=>"001101000",
  58805=>"000110111",
  58806=>"110111011",
  58807=>"010000010",
  58808=>"001001100",
  58809=>"010000000",
  58810=>"001000101",
  58811=>"010011001",
  58812=>"010111110",
  58813=>"000001001",
  58814=>"110001101",
  58815=>"011011001",
  58816=>"011011010",
  58817=>"010111010",
  58818=>"101111101",
  58819=>"000011100",
  58820=>"110001000",
  58821=>"100100010",
  58822=>"100001000",
  58823=>"000000000",
  58824=>"000010101",
  58825=>"010111011",
  58826=>"000100010",
  58827=>"001101101",
  58828=>"000110101",
  58829=>"111010001",
  58830=>"100000101",
  58831=>"111100100",
  58832=>"011000101",
  58833=>"011000100",
  58834=>"000100111",
  58835=>"101000011",
  58836=>"111100101",
  58837=>"110011011",
  58838=>"010111000",
  58839=>"110001111",
  58840=>"000110011",
  58841=>"101001111",
  58842=>"101010000",
  58843=>"001000001",
  58844=>"110101011",
  58845=>"001001000",
  58846=>"010101000",
  58847=>"011001100",
  58848=>"010011000",
  58849=>"001101111",
  58850=>"001010100",
  58851=>"111101000",
  58852=>"101011100",
  58853=>"010101101",
  58854=>"001000010",
  58855=>"001000001",
  58856=>"111001001",
  58857=>"111001110",
  58858=>"001100111",
  58859=>"001011010",
  58860=>"110010110",
  58861=>"110111100",
  58862=>"010100101",
  58863=>"111011010",
  58864=>"110011111",
  58865=>"011011011",
  58866=>"010001111",
  58867=>"111011010",
  58868=>"000111111",
  58869=>"101000001",
  58870=>"000100001",
  58871=>"111010001",
  58872=>"101111011",
  58873=>"001001011",
  58874=>"000010010",
  58875=>"100001111",
  58876=>"111101001",
  58877=>"101111101",
  58878=>"101111010",
  58879=>"001001011",
  58880=>"110111111",
  58881=>"111001010",
  58882=>"010001010",
  58883=>"101101111",
  58884=>"010100110",
  58885=>"111001000",
  58886=>"001100010",
  58887=>"011001001",
  58888=>"011110111",
  58889=>"101100110",
  58890=>"000110110",
  58891=>"001111110",
  58892=>"101010001",
  58893=>"011101001",
  58894=>"000011111",
  58895=>"000101100",
  58896=>"111000101",
  58897=>"100101000",
  58898=>"000110000",
  58899=>"111111111",
  58900=>"110011001",
  58901=>"000011110",
  58902=>"001101100",
  58903=>"000111001",
  58904=>"000010000",
  58905=>"110100110",
  58906=>"011001001",
  58907=>"001111100",
  58908=>"011101101",
  58909=>"010010110",
  58910=>"100111110",
  58911=>"001110010",
  58912=>"011010000",
  58913=>"100001010",
  58914=>"000000000",
  58915=>"010101101",
  58916=>"010000000",
  58917=>"110110000",
  58918=>"000110110",
  58919=>"111110110",
  58920=>"111011011",
  58921=>"111110001",
  58922=>"000101000",
  58923=>"111011101",
  58924=>"110110000",
  58925=>"011010111",
  58926=>"111111101",
  58927=>"110001110",
  58928=>"111101001",
  58929=>"010000101",
  58930=>"101000110",
  58931=>"000010100",
  58932=>"100010000",
  58933=>"110111001",
  58934=>"011111101",
  58935=>"111100000",
  58936=>"011110100",
  58937=>"000111100",
  58938=>"010010000",
  58939=>"010011010",
  58940=>"101110011",
  58941=>"000010011",
  58942=>"110000000",
  58943=>"111010010",
  58944=>"111100101",
  58945=>"111111010",
  58946=>"000000100",
  58947=>"011101110",
  58948=>"111100010",
  58949=>"111101000",
  58950=>"100101100",
  58951=>"111110001",
  58952=>"110110010",
  58953=>"110010001",
  58954=>"100111101",
  58955=>"111010100",
  58956=>"001011100",
  58957=>"001000011",
  58958=>"010110101",
  58959=>"010111101",
  58960=>"010001001",
  58961=>"001010001",
  58962=>"111111101",
  58963=>"011011101",
  58964=>"111010001",
  58965=>"110001110",
  58966=>"000100101",
  58967=>"000111101",
  58968=>"101110001",
  58969=>"110010110",
  58970=>"111001111",
  58971=>"010010111",
  58972=>"010100110",
  58973=>"111100111",
  58974=>"100000101",
  58975=>"100101100",
  58976=>"011010010",
  58977=>"100011001",
  58978=>"010000101",
  58979=>"011101100",
  58980=>"101001111",
  58981=>"011000111",
  58982=>"000110100",
  58983=>"111111000",
  58984=>"111001011",
  58985=>"101101100",
  58986=>"100110001",
  58987=>"001000010",
  58988=>"000000111",
  58989=>"000101100",
  58990=>"001100011",
  58991=>"010110111",
  58992=>"010000000",
  58993=>"000001010",
  58994=>"110001100",
  58995=>"100010111",
  58996=>"001100000",
  58997=>"100001001",
  58998=>"011111100",
  58999=>"011110111",
  59000=>"011010010",
  59001=>"101001000",
  59002=>"100000000",
  59003=>"011101010",
  59004=>"111010000",
  59005=>"101001110",
  59006=>"100000100",
  59007=>"011111011",
  59008=>"000100001",
  59009=>"010010011",
  59010=>"100111100",
  59011=>"001011011",
  59012=>"110011000",
  59013=>"111000000",
  59014=>"010111011",
  59015=>"101010010",
  59016=>"010101111",
  59017=>"001010000",
  59018=>"010100111",
  59019=>"100110101",
  59020=>"000001111",
  59021=>"001011100",
  59022=>"111110000",
  59023=>"101001110",
  59024=>"101111100",
  59025=>"010111000",
  59026=>"101111000",
  59027=>"000011110",
  59028=>"110000011",
  59029=>"000101011",
  59030=>"111110010",
  59031=>"000001110",
  59032=>"010110100",
  59033=>"110000100",
  59034=>"010010001",
  59035=>"000100110",
  59036=>"011100001",
  59037=>"101100101",
  59038=>"000000101",
  59039=>"101111011",
  59040=>"110100011",
  59041=>"000010111",
  59042=>"001100011",
  59043=>"000011010",
  59044=>"111001100",
  59045=>"100000001",
  59046=>"010010000",
  59047=>"100110000",
  59048=>"111001010",
  59049=>"100010010",
  59050=>"100000010",
  59051=>"011111001",
  59052=>"101000001",
  59053=>"011101100",
  59054=>"110010100",
  59055=>"000001001",
  59056=>"010011100",
  59057=>"111000111",
  59058=>"100100111",
  59059=>"011010000",
  59060=>"011000110",
  59061=>"101000111",
  59062=>"110110010",
  59063=>"100001110",
  59064=>"001110000",
  59065=>"110010101",
  59066=>"011001011",
  59067=>"001110010",
  59068=>"010111111",
  59069=>"111010001",
  59070=>"001001000",
  59071=>"100111000",
  59072=>"110011101",
  59073=>"111010111",
  59074=>"100011110",
  59075=>"110101000",
  59076=>"000111011",
  59077=>"111001101",
  59078=>"011000000",
  59079=>"001111000",
  59080=>"110100001",
  59081=>"011001001",
  59082=>"100111010",
  59083=>"010111000",
  59084=>"000110000",
  59085=>"101110011",
  59086=>"110101010",
  59087=>"010110011",
  59088=>"001100111",
  59089=>"000010010",
  59090=>"100110100",
  59091=>"101001000",
  59092=>"000000100",
  59093=>"010110001",
  59094=>"011101110",
  59095=>"100111110",
  59096=>"110000011",
  59097=>"001010101",
  59098=>"110101000",
  59099=>"000001111",
  59100=>"011000011",
  59101=>"000111000",
  59102=>"010011101",
  59103=>"000001010",
  59104=>"010111111",
  59105=>"110010001",
  59106=>"010100100",
  59107=>"110111000",
  59108=>"101010010",
  59109=>"101110101",
  59110=>"100011110",
  59111=>"110001111",
  59112=>"000001110",
  59113=>"010110110",
  59114=>"001000101",
  59115=>"101000100",
  59116=>"010011111",
  59117=>"000011011",
  59118=>"010000011",
  59119=>"001101111",
  59120=>"110111101",
  59121=>"101011111",
  59122=>"000000011",
  59123=>"011110000",
  59124=>"110000010",
  59125=>"000010100",
  59126=>"010010101",
  59127=>"001011000",
  59128=>"010001010",
  59129=>"000011010",
  59130=>"000011011",
  59131=>"101001111",
  59132=>"010011110",
  59133=>"111000111",
  59134=>"010011010",
  59135=>"101001010",
  59136=>"011011011",
  59137=>"011000100",
  59138=>"110100111",
  59139=>"111101010",
  59140=>"010100001",
  59141=>"100011010",
  59142=>"111100011",
  59143=>"001001101",
  59144=>"010011011",
  59145=>"011000010",
  59146=>"001001111",
  59147=>"001011100",
  59148=>"111011100",
  59149=>"001111001",
  59150=>"010001011",
  59151=>"111000000",
  59152=>"100111111",
  59153=>"011011100",
  59154=>"101101101",
  59155=>"010010100",
  59156=>"001010010",
  59157=>"110110001",
  59158=>"010110101",
  59159=>"000010011",
  59160=>"001001000",
  59161=>"010000110",
  59162=>"000000101",
  59163=>"001001010",
  59164=>"101111111",
  59165=>"100100010",
  59166=>"111100100",
  59167=>"010101000",
  59168=>"000101001",
  59169=>"111100110",
  59170=>"100110100",
  59171=>"111011010",
  59172=>"110101000",
  59173=>"000010000",
  59174=>"000010100",
  59175=>"101101000",
  59176=>"000011001",
  59177=>"111110010",
  59178=>"010101100",
  59179=>"010011100",
  59180=>"110001010",
  59181=>"101111101",
  59182=>"000001001",
  59183=>"111010011",
  59184=>"011001010",
  59185=>"101100101",
  59186=>"111010100",
  59187=>"101101110",
  59188=>"011111111",
  59189=>"100011111",
  59190=>"110100100",
  59191=>"001011101",
  59192=>"011000001",
  59193=>"001011011",
  59194=>"101000010",
  59195=>"111000010",
  59196=>"011000100",
  59197=>"011001100",
  59198=>"000001110",
  59199=>"100000001",
  59200=>"001010011",
  59201=>"110011000",
  59202=>"110000010",
  59203=>"000101110",
  59204=>"010111010",
  59205=>"111010000",
  59206=>"010110101",
  59207=>"000100111",
  59208=>"101011001",
  59209=>"101010001",
  59210=>"110010111",
  59211=>"110101011",
  59212=>"111011010",
  59213=>"010000100",
  59214=>"010110001",
  59215=>"100000111",
  59216=>"001001010",
  59217=>"101000000",
  59218=>"000111001",
  59219=>"111110110",
  59220=>"101100101",
  59221=>"001000100",
  59222=>"000001000",
  59223=>"110111111",
  59224=>"100111001",
  59225=>"011100100",
  59226=>"110000100",
  59227=>"011010000",
  59228=>"010001001",
  59229=>"110011010",
  59230=>"000111000",
  59231=>"101000001",
  59232=>"101101100",
  59233=>"111110001",
  59234=>"110011111",
  59235=>"010010011",
  59236=>"110000000",
  59237=>"111011001",
  59238=>"001011111",
  59239=>"100101100",
  59240=>"011101001",
  59241=>"011111111",
  59242=>"100001001",
  59243=>"010100010",
  59244=>"001101100",
  59245=>"011011010",
  59246=>"100000010",
  59247=>"100100111",
  59248=>"110010101",
  59249=>"101111000",
  59250=>"011110000",
  59251=>"100110010",
  59252=>"000101001",
  59253=>"000011010",
  59254=>"001000111",
  59255=>"111100001",
  59256=>"010111100",
  59257=>"100010011",
  59258=>"000100111",
  59259=>"001001001",
  59260=>"101000000",
  59261=>"010011111",
  59262=>"001101110",
  59263=>"111010010",
  59264=>"001110010",
  59265=>"101010101",
  59266=>"010000010",
  59267=>"010110111",
  59268=>"010001010",
  59269=>"000110011",
  59270=>"110101000",
  59271=>"000100010",
  59272=>"010000101",
  59273=>"110000101",
  59274=>"000100101",
  59275=>"110010000",
  59276=>"100001101",
  59277=>"011110111",
  59278=>"010011101",
  59279=>"101000100",
  59280=>"111000000",
  59281=>"000011011",
  59282=>"101000100",
  59283=>"011100011",
  59284=>"010100001",
  59285=>"000010010",
  59286=>"011001011",
  59287=>"111010000",
  59288=>"001000010",
  59289=>"100010110",
  59290=>"000001111",
  59291=>"110001101",
  59292=>"011010011",
  59293=>"110110111",
  59294=>"000000000",
  59295=>"001001000",
  59296=>"010000000",
  59297=>"101100010",
  59298=>"001111111",
  59299=>"000101100",
  59300=>"000000001",
  59301=>"111010010",
  59302=>"100100000",
  59303=>"101001010",
  59304=>"100101001",
  59305=>"000110100",
  59306=>"111111111",
  59307=>"101010100",
  59308=>"111010101",
  59309=>"000001010",
  59310=>"101111101",
  59311=>"100111000",
  59312=>"101000010",
  59313=>"011110000",
  59314=>"010101110",
  59315=>"110001111",
  59316=>"001001010",
  59317=>"100101011",
  59318=>"110100001",
  59319=>"101110111",
  59320=>"000010111",
  59321=>"111000100",
  59322=>"011111000",
  59323=>"010000010",
  59324=>"101010101",
  59325=>"011000000",
  59326=>"001111111",
  59327=>"000001101",
  59328=>"001111000",
  59329=>"000110011",
  59330=>"001101011",
  59331=>"011111111",
  59332=>"000110100",
  59333=>"111111110",
  59334=>"111101110",
  59335=>"111000111",
  59336=>"110100001",
  59337=>"001111101",
  59338=>"001010011",
  59339=>"010010111",
  59340=>"100110000",
  59341=>"110000101",
  59342=>"001101000",
  59343=>"011100110",
  59344=>"001010001",
  59345=>"101101100",
  59346=>"101000001",
  59347=>"001100000",
  59348=>"000111100",
  59349=>"000100011",
  59350=>"011010000",
  59351=>"000010111",
  59352=>"111100111",
  59353=>"000111101",
  59354=>"100011000",
  59355=>"010101111",
  59356=>"000111000",
  59357=>"001101001",
  59358=>"110010011",
  59359=>"000111010",
  59360=>"011110111",
  59361=>"011100010",
  59362=>"100001000",
  59363=>"011111100",
  59364=>"000001000",
  59365=>"110100101",
  59366=>"000110110",
  59367=>"110110001",
  59368=>"111000010",
  59369=>"111000100",
  59370=>"000011011",
  59371=>"111010010",
  59372=>"110010010",
  59373=>"011110111",
  59374=>"100011100",
  59375=>"110111010",
  59376=>"010101100",
  59377=>"100110110",
  59378=>"110000111",
  59379=>"011111101",
  59380=>"100110101",
  59381=>"101100001",
  59382=>"010001111",
  59383=>"010010010",
  59384=>"011011101",
  59385=>"010001001",
  59386=>"001100101",
  59387=>"011010111",
  59388=>"110100100",
  59389=>"011010011",
  59390=>"010011000",
  59391=>"101110101",
  59392=>"111001111",
  59393=>"010101011",
  59394=>"111011101",
  59395=>"101001000",
  59396=>"110010111",
  59397=>"010010011",
  59398=>"110111111",
  59399=>"010111111",
  59400=>"111011000",
  59401=>"100101000",
  59402=>"000001010",
  59403=>"100111001",
  59404=>"111101010",
  59405=>"011001111",
  59406=>"011111001",
  59407=>"101010110",
  59408=>"100100011",
  59409=>"000000101",
  59410=>"101011001",
  59411=>"001111011",
  59412=>"101100001",
  59413=>"001100111",
  59414=>"110010110",
  59415=>"100000000",
  59416=>"101000000",
  59417=>"111100000",
  59418=>"101111000",
  59419=>"010100010",
  59420=>"111000010",
  59421=>"111001101",
  59422=>"000011101",
  59423=>"100010101",
  59424=>"011000011",
  59425=>"001110000",
  59426=>"110111010",
  59427=>"111111100",
  59428=>"011110111",
  59429=>"110111100",
  59430=>"100001011",
  59431=>"100011101",
  59432=>"000001000",
  59433=>"000111110",
  59434=>"101101000",
  59435=>"111101101",
  59436=>"101100001",
  59437=>"001000010",
  59438=>"111010110",
  59439=>"000001010",
  59440=>"000010000",
  59441=>"110110010",
  59442=>"001000110",
  59443=>"010001110",
  59444=>"101010001",
  59445=>"110110010",
  59446=>"000000010",
  59447=>"000000111",
  59448=>"110101101",
  59449=>"000011000",
  59450=>"011010100",
  59451=>"111111100",
  59452=>"110100110",
  59453=>"111110110",
  59454=>"100010100",
  59455=>"111101011",
  59456=>"111111000",
  59457=>"011100000",
  59458=>"011000000",
  59459=>"100111010",
  59460=>"101011010",
  59461=>"011010101",
  59462=>"111010000",
  59463=>"111010110",
  59464=>"111111001",
  59465=>"011111110",
  59466=>"101000101",
  59467=>"001010011",
  59468=>"101001001",
  59469=>"011011011",
  59470=>"111100100",
  59471=>"011000011",
  59472=>"110101011",
  59473=>"010100010",
  59474=>"100010111",
  59475=>"110110100",
  59476=>"111010000",
  59477=>"000101101",
  59478=>"110010010",
  59479=>"001100010",
  59480=>"111010010",
  59481=>"100010110",
  59482=>"001011101",
  59483=>"011011011",
  59484=>"111111100",
  59485=>"010001100",
  59486=>"101111000",
  59487=>"001011100",
  59488=>"000100110",
  59489=>"101110011",
  59490=>"011100100",
  59491=>"010111001",
  59492=>"000110000",
  59493=>"100011000",
  59494=>"100111010",
  59495=>"111000111",
  59496=>"100010101",
  59497=>"001010111",
  59498=>"010000011",
  59499=>"000000000",
  59500=>"000101011",
  59501=>"110110001",
  59502=>"110011011",
  59503=>"100000111",
  59504=>"010100011",
  59505=>"001110100",
  59506=>"010100100",
  59507=>"111101011",
  59508=>"010111100",
  59509=>"001000101",
  59510=>"000010110",
  59511=>"011011111",
  59512=>"000100001",
  59513=>"100000010",
  59514=>"111110101",
  59515=>"010111011",
  59516=>"100001101",
  59517=>"111100010",
  59518=>"100101101",
  59519=>"100101111",
  59520=>"000011010",
  59521=>"001111000",
  59522=>"101010000",
  59523=>"101110100",
  59524=>"111101000",
  59525=>"100111100",
  59526=>"100000000",
  59527=>"010010010",
  59528=>"101011111",
  59529=>"001000111",
  59530=>"111111111",
  59531=>"100001100",
  59532=>"000100110",
  59533=>"010010000",
  59534=>"000100010",
  59535=>"001011010",
  59536=>"001110100",
  59537=>"111010010",
  59538=>"101010001",
  59539=>"111110100",
  59540=>"011010010",
  59541=>"000100111",
  59542=>"100100001",
  59543=>"110110111",
  59544=>"110101101",
  59545=>"010011000",
  59546=>"010010111",
  59547=>"100010110",
  59548=>"010110011",
  59549=>"100110001",
  59550=>"010001000",
  59551=>"001101000",
  59552=>"000101010",
  59553=>"000001100",
  59554=>"011101010",
  59555=>"100010100",
  59556=>"100011011",
  59557=>"100011100",
  59558=>"100100011",
  59559=>"000101000",
  59560=>"110111010",
  59561=>"011000001",
  59562=>"000011010",
  59563=>"101000011",
  59564=>"111110001",
  59565=>"101111011",
  59566=>"000111011",
  59567=>"100010110",
  59568=>"100011010",
  59569=>"010101110",
  59570=>"010100010",
  59571=>"001001110",
  59572=>"011111001",
  59573=>"110010011",
  59574=>"110101011",
  59575=>"100000110",
  59576=>"101000000",
  59577=>"110001101",
  59578=>"011000100",
  59579=>"000010000",
  59580=>"011101011",
  59581=>"001001111",
  59582=>"100010000",
  59583=>"111011001",
  59584=>"110101100",
  59585=>"001001101",
  59586=>"101000010",
  59587=>"101000110",
  59588=>"011101001",
  59589=>"000101001",
  59590=>"101001100",
  59591=>"101011101",
  59592=>"110011001",
  59593=>"110111111",
  59594=>"110100101",
  59595=>"000011000",
  59596=>"110100101",
  59597=>"001110111",
  59598=>"010111011",
  59599=>"001100110",
  59600=>"011011110",
  59601=>"001100000",
  59602=>"100110101",
  59603=>"011011110",
  59604=>"001000000",
  59605=>"111110001",
  59606=>"110001000",
  59607=>"111110111",
  59608=>"111011101",
  59609=>"010000000",
  59610=>"110000100",
  59611=>"111000000",
  59612=>"111110010",
  59613=>"011110110",
  59614=>"010111000",
  59615=>"011110011",
  59616=>"010010000",
  59617=>"000111100",
  59618=>"101110110",
  59619=>"100000110",
  59620=>"011010001",
  59621=>"001111110",
  59622=>"110000100",
  59623=>"000001001",
  59624=>"000000001",
  59625=>"111000001",
  59626=>"101001011",
  59627=>"010101110",
  59628=>"010011111",
  59629=>"000110010",
  59630=>"000001000",
  59631=>"111101001",
  59632=>"111111111",
  59633=>"000100111",
  59634=>"111011111",
  59635=>"011001111",
  59636=>"110000101",
  59637=>"000100101",
  59638=>"010101110",
  59639=>"011101111",
  59640=>"000010110",
  59641=>"100000100",
  59642=>"000101000",
  59643=>"001000001",
  59644=>"011001110",
  59645=>"001111110",
  59646=>"001101011",
  59647=>"000011100",
  59648=>"101100110",
  59649=>"101011100",
  59650=>"001010001",
  59651=>"000010010",
  59652=>"001100001",
  59653=>"011000100",
  59654=>"010110001",
  59655=>"011100000",
  59656=>"111111001",
  59657=>"110111111",
  59658=>"000011111",
  59659=>"100011101",
  59660=>"011111101",
  59661=>"001001010",
  59662=>"010100110",
  59663=>"111111100",
  59664=>"100011110",
  59665=>"101101000",
  59666=>"111010111",
  59667=>"000010110",
  59668=>"110110111",
  59669=>"011000111",
  59670=>"100110011",
  59671=>"001100110",
  59672=>"111000111",
  59673=>"000111111",
  59674=>"011000101",
  59675=>"011110000",
  59676=>"100000100",
  59677=>"001101100",
  59678=>"000100011",
  59679=>"001111001",
  59680=>"011000010",
  59681=>"011011100",
  59682=>"100100110",
  59683=>"110000010",
  59684=>"000011000",
  59685=>"001100110",
  59686=>"010100100",
  59687=>"000001010",
  59688=>"100001001",
  59689=>"101010000",
  59690=>"101001000",
  59691=>"110110011",
  59692=>"101010110",
  59693=>"101001111",
  59694=>"100011110",
  59695=>"000110100",
  59696=>"100010000",
  59697=>"101110111",
  59698=>"111111101",
  59699=>"001011111",
  59700=>"101111100",
  59701=>"100100111",
  59702=>"010000111",
  59703=>"001001101",
  59704=>"110010011",
  59705=>"010000000",
  59706=>"110100100",
  59707=>"101000010",
  59708=>"010101001",
  59709=>"111001011",
  59710=>"010100000",
  59711=>"010101110",
  59712=>"000001100",
  59713=>"110011001",
  59714=>"111001011",
  59715=>"111101000",
  59716=>"000010010",
  59717=>"111000010",
  59718=>"110111000",
  59719=>"010010001",
  59720=>"101010101",
  59721=>"110010000",
  59722=>"101101101",
  59723=>"011101001",
  59724=>"100101010",
  59725=>"000110101",
  59726=>"001000101",
  59727=>"110000001",
  59728=>"100001010",
  59729=>"100011011",
  59730=>"000011000",
  59731=>"100100100",
  59732=>"010001100",
  59733=>"000011001",
  59734=>"001000110",
  59735=>"001111010",
  59736=>"100111001",
  59737=>"001110100",
  59738=>"000001010",
  59739=>"111110000",
  59740=>"110011101",
  59741=>"100000010",
  59742=>"110111101",
  59743=>"000001111",
  59744=>"100110011",
  59745=>"001000010",
  59746=>"111000110",
  59747=>"000011010",
  59748=>"111110000",
  59749=>"110101010",
  59750=>"101111000",
  59751=>"101100110",
  59752=>"010000000",
  59753=>"000010010",
  59754=>"100111111",
  59755=>"100011010",
  59756=>"000101111",
  59757=>"010111110",
  59758=>"001011010",
  59759=>"000110110",
  59760=>"000111000",
  59761=>"101100100",
  59762=>"010011100",
  59763=>"100001001",
  59764=>"101010010",
  59765=>"011111001",
  59766=>"100010100",
  59767=>"000101101",
  59768=>"110000011",
  59769=>"010111100",
  59770=>"110011101",
  59771=>"000010000",
  59772=>"111111101",
  59773=>"001010100",
  59774=>"010011111",
  59775=>"100011101",
  59776=>"001111001",
  59777=>"111100000",
  59778=>"110011001",
  59779=>"010101001",
  59780=>"011000100",
  59781=>"000100011",
  59782=>"101101111",
  59783=>"001100011",
  59784=>"100110111",
  59785=>"111101110",
  59786=>"011010011",
  59787=>"100111010",
  59788=>"110001100",
  59789=>"110101101",
  59790=>"101100110",
  59791=>"001100011",
  59792=>"111001001",
  59793=>"000010001",
  59794=>"011001000",
  59795=>"100101101",
  59796=>"011101111",
  59797=>"111011010",
  59798=>"010111101",
  59799=>"111111101",
  59800=>"100011000",
  59801=>"100110001",
  59802=>"111000000",
  59803=>"011100011",
  59804=>"110111100",
  59805=>"110101111",
  59806=>"010000010",
  59807=>"000101010",
  59808=>"000101110",
  59809=>"101001011",
  59810=>"011111111",
  59811=>"010000111",
  59812=>"100110101",
  59813=>"001110110",
  59814=>"010000000",
  59815=>"111001101",
  59816=>"011100110",
  59817=>"100011011",
  59818=>"000111100",
  59819=>"011010110",
  59820=>"110101110",
  59821=>"110000100",
  59822=>"100011111",
  59823=>"011001100",
  59824=>"001110100",
  59825=>"010000111",
  59826=>"101001110",
  59827=>"011011111",
  59828=>"110011101",
  59829=>"111100100",
  59830=>"110101000",
  59831=>"100011000",
  59832=>"101100000",
  59833=>"100010010",
  59834=>"011110100",
  59835=>"001110001",
  59836=>"110111110",
  59837=>"011011000",
  59838=>"001000000",
  59839=>"001011000",
  59840=>"100100100",
  59841=>"010100001",
  59842=>"010110110",
  59843=>"000011111",
  59844=>"001000001",
  59845=>"111110110",
  59846=>"000010110",
  59847=>"001000110",
  59848=>"001110000",
  59849=>"100010011",
  59850=>"100111000",
  59851=>"010000010",
  59852=>"001100111",
  59853=>"001110011",
  59854=>"001101110",
  59855=>"011100101",
  59856=>"100010110",
  59857=>"111111100",
  59858=>"001011000",
  59859=>"111111010",
  59860=>"011011100",
  59861=>"101110100",
  59862=>"111110010",
  59863=>"001101100",
  59864=>"001101111",
  59865=>"111100000",
  59866=>"110100110",
  59867=>"011110100",
  59868=>"100011110",
  59869=>"010001101",
  59870=>"111001001",
  59871=>"010010110",
  59872=>"011111110",
  59873=>"011111011",
  59874=>"010101011",
  59875=>"001110000",
  59876=>"111010110",
  59877=>"011001011",
  59878=>"001101001",
  59879=>"000101001",
  59880=>"101111111",
  59881=>"110111010",
  59882=>"010101101",
  59883=>"100000000",
  59884=>"101110110",
  59885=>"011010111",
  59886=>"011000110",
  59887=>"011001101",
  59888=>"110001101",
  59889=>"011000101",
  59890=>"010010011",
  59891=>"100000000",
  59892=>"011111011",
  59893=>"110011111",
  59894=>"000000000",
  59895=>"101010110",
  59896=>"111001001",
  59897=>"111000100",
  59898=>"100001000",
  59899=>"000110101",
  59900=>"011111111",
  59901=>"110011001",
  59902=>"010101001",
  59903=>"011101100",
  59904=>"110111110",
  59905=>"001010111",
  59906=>"001101101",
  59907=>"100000010",
  59908=>"011100001",
  59909=>"101001000",
  59910=>"111100100",
  59911=>"000010000",
  59912=>"011100111",
  59913=>"010011010",
  59914=>"001010111",
  59915=>"110111110",
  59916=>"101111100",
  59917=>"101000111",
  59918=>"100101000",
  59919=>"100011100",
  59920=>"110101001",
  59921=>"100001010",
  59922=>"011111011",
  59923=>"110001100",
  59924=>"110100000",
  59925=>"110100100",
  59926=>"001001100",
  59927=>"010110000",
  59928=>"100000111",
  59929=>"101110100",
  59930=>"111100011",
  59931=>"010011011",
  59932=>"001100111",
  59933=>"111101011",
  59934=>"011001010",
  59935=>"110111011",
  59936=>"101110111",
  59937=>"010000100",
  59938=>"110011001",
  59939=>"110101111",
  59940=>"100100000",
  59941=>"111100101",
  59942=>"010111000",
  59943=>"010110011",
  59944=>"011110000",
  59945=>"111101100",
  59946=>"001001001",
  59947=>"100110010",
  59948=>"010110000",
  59949=>"100001100",
  59950=>"100011100",
  59951=>"011011101",
  59952=>"110010010",
  59953=>"000111001",
  59954=>"110101101",
  59955=>"010001010",
  59956=>"101000100",
  59957=>"000010001",
  59958=>"101100100",
  59959=>"111001010",
  59960=>"000010011",
  59961=>"000100011",
  59962=>"011010111",
  59963=>"100111000",
  59964=>"000010110",
  59965=>"001111010",
  59966=>"010100001",
  59967=>"101110101",
  59968=>"011011111",
  59969=>"100111110",
  59970=>"110001001",
  59971=>"011011101",
  59972=>"101011001",
  59973=>"010011101",
  59974=>"100000001",
  59975=>"010110111",
  59976=>"101001010",
  59977=>"111101100",
  59978=>"110110010",
  59979=>"001101100",
  59980=>"100000000",
  59981=>"001000100",
  59982=>"001000100",
  59983=>"101010111",
  59984=>"101110010",
  59985=>"101001110",
  59986=>"010110011",
  59987=>"001111110",
  59988=>"100010101",
  59989=>"010001011",
  59990=>"111101000",
  59991=>"011001011",
  59992=>"101101011",
  59993=>"100110001",
  59994=>"011111001",
  59995=>"111111010",
  59996=>"101101001",
  59997=>"000011101",
  59998=>"010000101",
  59999=>"000000111",
  60000=>"111010011",
  60001=>"010111000",
  60002=>"010111101",
  60003=>"001011010",
  60004=>"001100000",
  60005=>"100001001",
  60006=>"000000110",
  60007=>"000100001",
  60008=>"001100100",
  60009=>"110100100",
  60010=>"001010000",
  60011=>"111000000",
  60012=>"001111001",
  60013=>"101100101",
  60014=>"111000111",
  60015=>"101111000",
  60016=>"011001000",
  60017=>"011110011",
  60018=>"101011010",
  60019=>"101010011",
  60020=>"010010111",
  60021=>"000101001",
  60022=>"010100111",
  60023=>"011111001",
  60024=>"010100011",
  60025=>"010111010",
  60026=>"100001001",
  60027=>"101011101",
  60028=>"010111101",
  60029=>"111001010",
  60030=>"010111000",
  60031=>"011110110",
  60032=>"111111000",
  60033=>"010011111",
  60034=>"111111101",
  60035=>"110011111",
  60036=>"100000011",
  60037=>"101110000",
  60038=>"111011111",
  60039=>"000100001",
  60040=>"100100000",
  60041=>"001000010",
  60042=>"101010111",
  60043=>"100010001",
  60044=>"001010101",
  60045=>"000011000",
  60046=>"110010001",
  60047=>"111111101",
  60048=>"101011101",
  60049=>"110010001",
  60050=>"000100110",
  60051=>"100011000",
  60052=>"000011011",
  60053=>"011000101",
  60054=>"110110111",
  60055=>"000000100",
  60056=>"111111100",
  60057=>"010100101",
  60058=>"011011101",
  60059=>"100010110",
  60060=>"100111010",
  60061=>"001110010",
  60062=>"000001000",
  60063=>"010011100",
  60064=>"110010110",
  60065=>"001001101",
  60066=>"001101110",
  60067=>"111101100",
  60068=>"111000100",
  60069=>"100110000",
  60070=>"101011011",
  60071=>"001101101",
  60072=>"100001110",
  60073=>"111110100",
  60074=>"001101101",
  60075=>"010110111",
  60076=>"100011111",
  60077=>"001001100",
  60078=>"101010001",
  60079=>"110000000",
  60080=>"010110101",
  60081=>"000010101",
  60082=>"111011000",
  60083=>"110011011",
  60084=>"001000001",
  60085=>"100011000",
  60086=>"000001101",
  60087=>"110000011",
  60088=>"000011011",
  60089=>"101000011",
  60090=>"000011000",
  60091=>"011111010",
  60092=>"001111101",
  60093=>"010111100",
  60094=>"101100110",
  60095=>"011100011",
  60096=>"111011100",
  60097=>"101010101",
  60098=>"010000000",
  60099=>"010001000",
  60100=>"111011111",
  60101=>"001111011",
  60102=>"001100101",
  60103=>"111111110",
  60104=>"111010111",
  60105=>"111001010",
  60106=>"111001000",
  60107=>"111001011",
  60108=>"000000111",
  60109=>"111110101",
  60110=>"001001110",
  60111=>"011110010",
  60112=>"111101101",
  60113=>"110100100",
  60114=>"011111010",
  60115=>"100000111",
  60116=>"101001010",
  60117=>"001000000",
  60118=>"110001101",
  60119=>"001111101",
  60120=>"000100010",
  60121=>"100101011",
  60122=>"101001101",
  60123=>"110100011",
  60124=>"101110110",
  60125=>"111000011",
  60126=>"100111100",
  60127=>"100100011",
  60128=>"110100100",
  60129=>"010001010",
  60130=>"100001001",
  60131=>"001000111",
  60132=>"110011000",
  60133=>"000101000",
  60134=>"000111101",
  60135=>"011111000",
  60136=>"100011001",
  60137=>"110110010",
  60138=>"101100100",
  60139=>"000101001",
  60140=>"000100101",
  60141=>"011101000",
  60142=>"010111111",
  60143=>"111000111",
  60144=>"010000111",
  60145=>"111101011",
  60146=>"110100000",
  60147=>"100100100",
  60148=>"111111101",
  60149=>"011110001",
  60150=>"111101001",
  60151=>"010011000",
  60152=>"111101011",
  60153=>"001111110",
  60154=>"010011011",
  60155=>"001110101",
  60156=>"101011111",
  60157=>"100111010",
  60158=>"000100100",
  60159=>"011100101",
  60160=>"001011011",
  60161=>"000010001",
  60162=>"001101001",
  60163=>"110000100",
  60164=>"100001100",
  60165=>"001010001",
  60166=>"001100011",
  60167=>"001100011",
  60168=>"101011000",
  60169=>"001110111",
  60170=>"010101101",
  60171=>"101001001",
  60172=>"010101111",
  60173=>"001011100",
  60174=>"010011100",
  60175=>"101101101",
  60176=>"101110011",
  60177=>"101101010",
  60178=>"000011011",
  60179=>"100100011",
  60180=>"000100111",
  60181=>"000010110",
  60182=>"101100010",
  60183=>"010000010",
  60184=>"101101110",
  60185=>"000000000",
  60186=>"001111101",
  60187=>"111111001",
  60188=>"110001001",
  60189=>"010001001",
  60190=>"011101000",
  60191=>"001000101",
  60192=>"000000010",
  60193=>"010100111",
  60194=>"000101011",
  60195=>"101010110",
  60196=>"100110010",
  60197=>"001011110",
  60198=>"111100110",
  60199=>"101000001",
  60200=>"010001001",
  60201=>"000010011",
  60202=>"000110111",
  60203=>"110101111",
  60204=>"001100011",
  60205=>"000100000",
  60206=>"110010110",
  60207=>"111011010",
  60208=>"011000101",
  60209=>"101010000",
  60210=>"001111000",
  60211=>"000010111",
  60212=>"000001100",
  60213=>"011001111",
  60214=>"000100001",
  60215=>"101110011",
  60216=>"010111100",
  60217=>"101010110",
  60218=>"111100000",
  60219=>"101000000",
  60220=>"010011010",
  60221=>"001100111",
  60222=>"001010001",
  60223=>"100010111",
  60224=>"010001001",
  60225=>"111011101",
  60226=>"001100001",
  60227=>"011100111",
  60228=>"101110000",
  60229=>"001101101",
  60230=>"100101001",
  60231=>"110011101",
  60232=>"001000100",
  60233=>"110111100",
  60234=>"110100011",
  60235=>"100111100",
  60236=>"101000110",
  60237=>"111110101",
  60238=>"111000001",
  60239=>"100001101",
  60240=>"000010000",
  60241=>"001100011",
  60242=>"010010011",
  60243=>"101010000",
  60244=>"001110000",
  60245=>"001011010",
  60246=>"000110100",
  60247=>"010000110",
  60248=>"111001011",
  60249=>"110111111",
  60250=>"001100100",
  60251=>"011001100",
  60252=>"100001110",
  60253=>"111100110",
  60254=>"111011010",
  60255=>"100001001",
  60256=>"101010110",
  60257=>"001000001",
  60258=>"010010110",
  60259=>"001000100",
  60260=>"001100111",
  60261=>"110111101",
  60262=>"111101111",
  60263=>"100000001",
  60264=>"010010000",
  60265=>"010000100",
  60266=>"011011010",
  60267=>"110000101",
  60268=>"111101000",
  60269=>"010000111",
  60270=>"110000110",
  60271=>"100000010",
  60272=>"111000001",
  60273=>"100000000",
  60274=>"010100010",
  60275=>"110110010",
  60276=>"101110110",
  60277=>"010110111",
  60278=>"010101010",
  60279=>"100101011",
  60280=>"011111101",
  60281=>"000100100",
  60282=>"000010011",
  60283=>"000110000",
  60284=>"000011101",
  60285=>"111000101",
  60286=>"011101001",
  60287=>"111010101",
  60288=>"011011000",
  60289=>"010000101",
  60290=>"001010000",
  60291=>"100110110",
  60292=>"010000100",
  60293=>"110111011",
  60294=>"000100000",
  60295=>"011001101",
  60296=>"110011100",
  60297=>"001001011",
  60298=>"111110110",
  60299=>"110000011",
  60300=>"111100100",
  60301=>"110000101",
  60302=>"100011011",
  60303=>"100011001",
  60304=>"100011001",
  60305=>"010010110",
  60306=>"000011110",
  60307=>"011010110",
  60308=>"001110000",
  60309=>"011001010",
  60310=>"100000111",
  60311=>"001001100",
  60312=>"100110110",
  60313=>"100010011",
  60314=>"010011100",
  60315=>"010101000",
  60316=>"000110010",
  60317=>"000111011",
  60318=>"101000011",
  60319=>"010000101",
  60320=>"100101100",
  60321=>"101000000",
  60322=>"110010011",
  60323=>"000011110",
  60324=>"000010111",
  60325=>"111001000",
  60326=>"010110100",
  60327=>"010010010",
  60328=>"110000000",
  60329=>"011000101",
  60330=>"110011101",
  60331=>"110011000",
  60332=>"000010000",
  60333=>"010111011",
  60334=>"100101100",
  60335=>"100111000",
  60336=>"011100110",
  60337=>"111110100",
  60338=>"100010111",
  60339=>"100011001",
  60340=>"010110010",
  60341=>"011001011",
  60342=>"011101010",
  60343=>"100000010",
  60344=>"111000110",
  60345=>"110101001",
  60346=>"100100000",
  60347=>"111101001",
  60348=>"001011000",
  60349=>"000000000",
  60350=>"101111111",
  60351=>"010000000",
  60352=>"011011010",
  60353=>"000100100",
  60354=>"011001000",
  60355=>"111110110",
  60356=>"110100001",
  60357=>"101111111",
  60358=>"110001111",
  60359=>"010010010",
  60360=>"111000001",
  60361=>"001111011",
  60362=>"111010010",
  60363=>"101011001",
  60364=>"010010100",
  60365=>"010001111",
  60366=>"001001000",
  60367=>"101110111",
  60368=>"100011111",
  60369=>"000011100",
  60370=>"000101010",
  60371=>"101000101",
  60372=>"010100000",
  60373=>"100101101",
  60374=>"010001011",
  60375=>"100110010",
  60376=>"001011100",
  60377=>"000000101",
  60378=>"011011000",
  60379=>"111101111",
  60380=>"001100011",
  60381=>"111011011",
  60382=>"010100110",
  60383=>"001010011",
  60384=>"000100001",
  60385=>"111111101",
  60386=>"011000001",
  60387=>"011010111",
  60388=>"100011010",
  60389=>"010110101",
  60390=>"001010010",
  60391=>"110100101",
  60392=>"101101001",
  60393=>"011100100",
  60394=>"000100111",
  60395=>"101111010",
  60396=>"001101100",
  60397=>"010111011",
  60398=>"000111011",
  60399=>"000000011",
  60400=>"111111011",
  60401=>"110010110",
  60402=>"001110010",
  60403=>"010011001",
  60404=>"111000110",
  60405=>"101000100",
  60406=>"000010111",
  60407=>"110111011",
  60408=>"000001001",
  60409=>"000101100",
  60410=>"000101000",
  60411=>"100111011",
  60412=>"101111101",
  60413=>"000000000",
  60414=>"000101011",
  60415=>"111000010",
  60416=>"011011100",
  60417=>"110001010",
  60418=>"100010000",
  60419=>"111010010",
  60420=>"100001101",
  60421=>"011101111",
  60422=>"001000100",
  60423=>"111100010",
  60424=>"100111111",
  60425=>"011000010",
  60426=>"000010010",
  60427=>"110110000",
  60428=>"000110110",
  60429=>"111101001",
  60430=>"010100101",
  60431=>"000001010",
  60432=>"100111011",
  60433=>"011110010",
  60434=>"000001110",
  60435=>"111110101",
  60436=>"000000100",
  60437=>"101110001",
  60438=>"001110001",
  60439=>"010000111",
  60440=>"010011001",
  60441=>"101000111",
  60442=>"100100101",
  60443=>"011000000",
  60444=>"110001001",
  60445=>"111011000",
  60446=>"100000100",
  60447=>"111111111",
  60448=>"100110101",
  60449=>"010100011",
  60450=>"010101001",
  60451=>"111101110",
  60452=>"011001001",
  60453=>"101111100",
  60454=>"011001011",
  60455=>"110011100",
  60456=>"000001110",
  60457=>"110011100",
  60458=>"101101011",
  60459=>"001010100",
  60460=>"110011011",
  60461=>"010000001",
  60462=>"000111001",
  60463=>"101011010",
  60464=>"000001111",
  60465=>"001000001",
  60466=>"010100101",
  60467=>"110011000",
  60468=>"010010011",
  60469=>"001000010",
  60470=>"001000010",
  60471=>"000001001",
  60472=>"111010101",
  60473=>"011111110",
  60474=>"111110010",
  60475=>"011000000",
  60476=>"001010110",
  60477=>"100100111",
  60478=>"100000010",
  60479=>"010101100",
  60480=>"111100110",
  60481=>"000000111",
  60482=>"110001100",
  60483=>"000111100",
  60484=>"001010000",
  60485=>"110011111",
  60486=>"010000100",
  60487=>"101100101",
  60488=>"111001011",
  60489=>"010101110",
  60490=>"100110010",
  60491=>"001000111",
  60492=>"011010100",
  60493=>"011010110",
  60494=>"100011100",
  60495=>"001100010",
  60496=>"101001011",
  60497=>"000100111",
  60498=>"101100100",
  60499=>"010001101",
  60500=>"001110100",
  60501=>"111100000",
  60502=>"111010001",
  60503=>"100111000",
  60504=>"001100101",
  60505=>"110001111",
  60506=>"010110000",
  60507=>"111000111",
  60508=>"001011000",
  60509=>"001001101",
  60510=>"010000010",
  60511=>"111001011",
  60512=>"110000001",
  60513=>"100001110",
  60514=>"111001011",
  60515=>"000100101",
  60516=>"001100100",
  60517=>"101111111",
  60518=>"000100000",
  60519=>"000100111",
  60520=>"110101111",
  60521=>"010110010",
  60522=>"010000111",
  60523=>"100010100",
  60524=>"110001001",
  60525=>"000100010",
  60526=>"010100011",
  60527=>"000010100",
  60528=>"101001010",
  60529=>"110001100",
  60530=>"001011001",
  60531=>"001101001",
  60532=>"011011000",
  60533=>"000001101",
  60534=>"110011011",
  60535=>"111101001",
  60536=>"111101000",
  60537=>"001110100",
  60538=>"101001011",
  60539=>"110010110",
  60540=>"100001111",
  60541=>"010000000",
  60542=>"101101011",
  60543=>"000000111",
  60544=>"100100110",
  60545=>"011110011",
  60546=>"011100001",
  60547=>"100001100",
  60548=>"111001111",
  60549=>"011101111",
  60550=>"000110000",
  60551=>"101110100",
  60552=>"100000100",
  60553=>"001100000",
  60554=>"000100100",
  60555=>"010000111",
  60556=>"100010010",
  60557=>"001001001",
  60558=>"110011111",
  60559=>"010000000",
  60560=>"001101010",
  60561=>"001000010",
  60562=>"001010100",
  60563=>"011100001",
  60564=>"000110101",
  60565=>"100100110",
  60566=>"110111101",
  60567=>"011001000",
  60568=>"110011000",
  60569=>"100111100",
  60570=>"111001010",
  60571=>"110010000",
  60572=>"110100100",
  60573=>"110000111",
  60574=>"111110010",
  60575=>"110111011",
  60576=>"101011110",
  60577=>"001001101",
  60578=>"100001001",
  60579=>"100100101",
  60580=>"001000000",
  60581=>"010111011",
  60582=>"100101111",
  60583=>"000110100",
  60584=>"011110100",
  60585=>"001100110",
  60586=>"001000001",
  60587=>"110001100",
  60588=>"010011001",
  60589=>"010011010",
  60590=>"001011110",
  60591=>"010010111",
  60592=>"011101001",
  60593=>"000111101",
  60594=>"011110001",
  60595=>"000010011",
  60596=>"100001001",
  60597=>"101111001",
  60598=>"011011100",
  60599=>"000000110",
  60600=>"000010010",
  60601=>"011111011",
  60602=>"110000001",
  60603=>"111101111",
  60604=>"010011100",
  60605=>"000000001",
  60606=>"011100001",
  60607=>"011100100",
  60608=>"010110000",
  60609=>"111011001",
  60610=>"110010101",
  60611=>"001010111",
  60612=>"011110110",
  60613=>"001010100",
  60614=>"101011110",
  60615=>"011011111",
  60616=>"010110001",
  60617=>"000100011",
  60618=>"011110100",
  60619=>"001100101",
  60620=>"001010000",
  60621=>"100101111",
  60622=>"111001111",
  60623=>"011101001",
  60624=>"110100000",
  60625=>"110110110",
  60626=>"110100110",
  60627=>"001010011",
  60628=>"111100000",
  60629=>"011100100",
  60630=>"010001001",
  60631=>"110001101",
  60632=>"000010000",
  60633=>"110110000",
  60634=>"100110110",
  60635=>"110001101",
  60636=>"010001010",
  60637=>"010000101",
  60638=>"101100001",
  60639=>"100000011",
  60640=>"111011000",
  60641=>"110110000",
  60642=>"101001000",
  60643=>"011111110",
  60644=>"000110100",
  60645=>"001001001",
  60646=>"010000000",
  60647=>"110000111",
  60648=>"011010111",
  60649=>"011000101",
  60650=>"011001000",
  60651=>"010011000",
  60652=>"000110110",
  60653=>"001110100",
  60654=>"101001100",
  60655=>"100100100",
  60656=>"001001100",
  60657=>"000111010",
  60658=>"100000111",
  60659=>"010011000",
  60660=>"100100100",
  60661=>"011010100",
  60662=>"000010100",
  60663=>"110001101",
  60664=>"011111110",
  60665=>"100111001",
  60666=>"011000111",
  60667=>"000011101",
  60668=>"000000110",
  60669=>"111000101",
  60670=>"001010100",
  60671=>"111111100",
  60672=>"011101011",
  60673=>"110111000",
  60674=>"101110001",
  60675=>"010100111",
  60676=>"110011101",
  60677=>"000110001",
  60678=>"110101111",
  60679=>"011111100",
  60680=>"111111000",
  60681=>"111011011",
  60682=>"010111101",
  60683=>"010010111",
  60684=>"011111100",
  60685=>"001000001",
  60686=>"100000011",
  60687=>"100011011",
  60688=>"101000011",
  60689=>"100011011",
  60690=>"010001110",
  60691=>"111110010",
  60692=>"111100001",
  60693=>"110010101",
  60694=>"111110101",
  60695=>"101101110",
  60696=>"111000011",
  60697=>"001010000",
  60698=>"110100000",
  60699=>"110001100",
  60700=>"100011000",
  60701=>"110111100",
  60702=>"011111010",
  60703=>"000111101",
  60704=>"000110111",
  60705=>"110011111",
  60706=>"000001000",
  60707=>"101000001",
  60708=>"011010010",
  60709=>"010000000",
  60710=>"010110010",
  60711=>"111101000",
  60712=>"111101100",
  60713=>"111011010",
  60714=>"000110100",
  60715=>"011001011",
  60716=>"100101000",
  60717=>"000110010",
  60718=>"000011000",
  60719=>"101000000",
  60720=>"001100000",
  60721=>"110000011",
  60722=>"000101010",
  60723=>"110010001",
  60724=>"111000001",
  60725=>"000000000",
  60726=>"110011010",
  60727=>"010011110",
  60728=>"000001111",
  60729=>"101000111",
  60730=>"110001010",
  60731=>"010001011",
  60732=>"000000110",
  60733=>"000011100",
  60734=>"001000000",
  60735=>"001100000",
  60736=>"100111111",
  60737=>"111010011",
  60738=>"000100101",
  60739=>"010100000",
  60740=>"101101001",
  60741=>"100010011",
  60742=>"100001000",
  60743=>"101101111",
  60744=>"000000000",
  60745=>"110001111",
  60746=>"101110000",
  60747=>"000001111",
  60748=>"010001111",
  60749=>"110010010",
  60750=>"111101000",
  60751=>"011111101",
  60752=>"101001110",
  60753=>"111101001",
  60754=>"001001000",
  60755=>"111001101",
  60756=>"001000001",
  60757=>"011010000",
  60758=>"100001110",
  60759=>"100001110",
  60760=>"010100000",
  60761=>"000101111",
  60762=>"100000111",
  60763=>"100100000",
  60764=>"111110110",
  60765=>"010011100",
  60766=>"011100001",
  60767=>"001101111",
  60768=>"001011111",
  60769=>"001110011",
  60770=>"111100110",
  60771=>"101100010",
  60772=>"011100111",
  60773=>"010000001",
  60774=>"101111100",
  60775=>"000001001",
  60776=>"111000100",
  60777=>"111111011",
  60778=>"000110101",
  60779=>"100100010",
  60780=>"101000010",
  60781=>"101011110",
  60782=>"010110001",
  60783=>"011001010",
  60784=>"011110100",
  60785=>"001001000",
  60786=>"111110011",
  60787=>"000010000",
  60788=>"001101100",
  60789=>"000101000",
  60790=>"000110111",
  60791=>"010000100",
  60792=>"101100001",
  60793=>"001010001",
  60794=>"101101010",
  60795=>"011001100",
  60796=>"011010001",
  60797=>"010010011",
  60798=>"110000101",
  60799=>"100001011",
  60800=>"100010101",
  60801=>"000100000",
  60802=>"100000101",
  60803=>"010001111",
  60804=>"000000101",
  60805=>"000010100",
  60806=>"011101011",
  60807=>"010001010",
  60808=>"111011111",
  60809=>"010111110",
  60810=>"011101001",
  60811=>"010111010",
  60812=>"000110100",
  60813=>"111011110",
  60814=>"010111100",
  60815=>"111011010",
  60816=>"100000010",
  60817=>"001001001",
  60818=>"010011010",
  60819=>"110111000",
  60820=>"101101100",
  60821=>"110000011",
  60822=>"110000100",
  60823=>"000011011",
  60824=>"000111001",
  60825=>"000000011",
  60826=>"111100111",
  60827=>"100011101",
  60828=>"011110101",
  60829=>"000100110",
  60830=>"110100001",
  60831=>"100001011",
  60832=>"110100111",
  60833=>"000100100",
  60834=>"000100011",
  60835=>"110000000",
  60836=>"110001110",
  60837=>"010010011",
  60838=>"111010110",
  60839=>"000011101",
  60840=>"111001111",
  60841=>"101010100",
  60842=>"010101010",
  60843=>"011011011",
  60844=>"100001111",
  60845=>"111001101",
  60846=>"001010111",
  60847=>"110111000",
  60848=>"110011100",
  60849=>"111100001",
  60850=>"000001110",
  60851=>"001111101",
  60852=>"001010000",
  60853=>"011111101",
  60854=>"011101001",
  60855=>"101000001",
  60856=>"100001101",
  60857=>"001010101",
  60858=>"000111100",
  60859=>"100100000",
  60860=>"111100011",
  60861=>"100011010",
  60862=>"000001101",
  60863=>"000101010",
  60864=>"001111110",
  60865=>"111110001",
  60866=>"001000010",
  60867=>"000001100",
  60868=>"000111111",
  60869=>"101101101",
  60870=>"001100100",
  60871=>"000010110",
  60872=>"011011100",
  60873=>"010001011",
  60874=>"010110001",
  60875=>"010111101",
  60876=>"110111011",
  60877=>"101000100",
  60878=>"000101001",
  60879=>"101111111",
  60880=>"010000101",
  60881=>"010000000",
  60882=>"000001001",
  60883=>"101111010",
  60884=>"110010101",
  60885=>"001011101",
  60886=>"100111000",
  60887=>"000111001",
  60888=>"101100000",
  60889=>"000010111",
  60890=>"000000100",
  60891=>"101000001",
  60892=>"011010011",
  60893=>"101111100",
  60894=>"011110001",
  60895=>"001111101",
  60896=>"110100100",
  60897=>"000110001",
  60898=>"011010001",
  60899=>"010101100",
  60900=>"011001100",
  60901=>"000111111",
  60902=>"000000010",
  60903=>"010000011",
  60904=>"101001000",
  60905=>"110110011",
  60906=>"101100111",
  60907=>"100110001",
  60908=>"000010110",
  60909=>"011110010",
  60910=>"100000000",
  60911=>"110001010",
  60912=>"110010100",
  60913=>"101010100",
  60914=>"111101010",
  60915=>"101001101",
  60916=>"101000000",
  60917=>"010011001",
  60918=>"110111101",
  60919=>"011111110",
  60920=>"110110000",
  60921=>"101110010",
  60922=>"110110101",
  60923=>"000010100",
  60924=>"010000100",
  60925=>"000100000",
  60926=>"011100011",
  60927=>"011110111",
  60928=>"111001000",
  60929=>"101000000",
  60930=>"001010001",
  60931=>"011111101",
  60932=>"101100110",
  60933=>"111101001",
  60934=>"111101001",
  60935=>"001100111",
  60936=>"000011101",
  60937=>"110011000",
  60938=>"010111111",
  60939=>"111010101",
  60940=>"000000011",
  60941=>"010001001",
  60942=>"010010000",
  60943=>"000111111",
  60944=>"100100100",
  60945=>"000010001",
  60946=>"100101010",
  60947=>"110110001",
  60948=>"001010110",
  60949=>"001001011",
  60950=>"111011000",
  60951=>"001111101",
  60952=>"001101001",
  60953=>"111100010",
  60954=>"000001000",
  60955=>"101101000",
  60956=>"011010111",
  60957=>"001000111",
  60958=>"111001100",
  60959=>"101111111",
  60960=>"101111111",
  60961=>"000000000",
  60962=>"000000111",
  60963=>"001011010",
  60964=>"111110011",
  60965=>"001001100",
  60966=>"011001111",
  60967=>"111100100",
  60968=>"011110011",
  60969=>"111001111",
  60970=>"101001110",
  60971=>"011000110",
  60972=>"010111100",
  60973=>"101100100",
  60974=>"110101111",
  60975=>"000100100",
  60976=>"101101000",
  60977=>"000010100",
  60978=>"111000000",
  60979=>"100000111",
  60980=>"100110011",
  60981=>"000010000",
  60982=>"101000001",
  60983=>"000111111",
  60984=>"010101000",
  60985=>"111010100",
  60986=>"101100101",
  60987=>"111111111",
  60988=>"001111011",
  60989=>"001101111",
  60990=>"111101000",
  60991=>"110011000",
  60992=>"001100001",
  60993=>"000000010",
  60994=>"101010100",
  60995=>"010001110",
  60996=>"111110110",
  60997=>"110111100",
  60998=>"011001101",
  60999=>"001010100",
  61000=>"101001001",
  61001=>"001101110",
  61002=>"001100111",
  61003=>"000001011",
  61004=>"111101011",
  61005=>"000000100",
  61006=>"010111000",
  61007=>"000110100",
  61008=>"010000001",
  61009=>"110001101",
  61010=>"001011001",
  61011=>"000011010",
  61012=>"101101110",
  61013=>"101000001",
  61014=>"101101111",
  61015=>"111011100",
  61016=>"110101010",
  61017=>"110101001",
  61018=>"100000001",
  61019=>"000010111",
  61020=>"100011110",
  61021=>"010110001",
  61022=>"100000111",
  61023=>"101011011",
  61024=>"000110010",
  61025=>"010101111",
  61026=>"000101110",
  61027=>"000011110",
  61028=>"000001000",
  61029=>"110111011",
  61030=>"111010001",
  61031=>"011111101",
  61032=>"001101101",
  61033=>"001010110",
  61034=>"100100000",
  61035=>"110100111",
  61036=>"111100001",
  61037=>"000111110",
  61038=>"010011010",
  61039=>"000101111",
  61040=>"110110000",
  61041=>"011011000",
  61042=>"110100101",
  61043=>"000010000",
  61044=>"001001110",
  61045=>"111111100",
  61046=>"001111000",
  61047=>"011010111",
  61048=>"010111011",
  61049=>"000010111",
  61050=>"100011111",
  61051=>"000111011",
  61052=>"110011101",
  61053=>"101111110",
  61054=>"101010000",
  61055=>"101001100",
  61056=>"011011011",
  61057=>"110001101",
  61058=>"011001111",
  61059=>"001101001",
  61060=>"111100001",
  61061=>"000101110",
  61062=>"111100001",
  61063=>"111010011",
  61064=>"100110011",
  61065=>"000010011",
  61066=>"111011000",
  61067=>"000101100",
  61068=>"001011101",
  61069=>"100010100",
  61070=>"000001011",
  61071=>"000000011",
  61072=>"100010100",
  61073=>"011011010",
  61074=>"000101010",
  61075=>"001011001",
  61076=>"111111101",
  61077=>"001000100",
  61078=>"101111001",
  61079=>"101001110",
  61080=>"010001010",
  61081=>"111100010",
  61082=>"010111110",
  61083=>"110001101",
  61084=>"000110110",
  61085=>"111010001",
  61086=>"111110010",
  61087=>"000010001",
  61088=>"100110001",
  61089=>"100011000",
  61090=>"010011000",
  61091=>"011001001",
  61092=>"001000100",
  61093=>"110011001",
  61094=>"011010010",
  61095=>"000010000",
  61096=>"111110111",
  61097=>"100001010",
  61098=>"111001101",
  61099=>"101111000",
  61100=>"100000100",
  61101=>"000110010",
  61102=>"000011111",
  61103=>"000010001",
  61104=>"011100111",
  61105=>"001111111",
  61106=>"111001111",
  61107=>"111111000",
  61108=>"101100110",
  61109=>"011011101",
  61110=>"011100011",
  61111=>"110101111",
  61112=>"101111110",
  61113=>"001000111",
  61114=>"111011000",
  61115=>"101100011",
  61116=>"100000101",
  61117=>"101001101",
  61118=>"001100010",
  61119=>"100010000",
  61120=>"111111010",
  61121=>"111110000",
  61122=>"100010001",
  61123=>"001000100",
  61124=>"100101010",
  61125=>"011110111",
  61126=>"101110100",
  61127=>"010000001",
  61128=>"010000010",
  61129=>"111101001",
  61130=>"011001111",
  61131=>"100000001",
  61132=>"010110001",
  61133=>"011010110",
  61134=>"101001110",
  61135=>"110110111",
  61136=>"000101001",
  61137=>"101101111",
  61138=>"101000110",
  61139=>"010010111",
  61140=>"011000100",
  61141=>"001000000",
  61142=>"110101111",
  61143=>"010101100",
  61144=>"101110110",
  61145=>"100011011",
  61146=>"011110100",
  61147=>"111101100",
  61148=>"010110110",
  61149=>"111111010",
  61150=>"011101010",
  61151=>"100000000",
  61152=>"001001000",
  61153=>"101010000",
  61154=>"000010111",
  61155=>"101111011",
  61156=>"001000010",
  61157=>"100001111",
  61158=>"110100111",
  61159=>"011001001",
  61160=>"000001000",
  61161=>"000011110",
  61162=>"011111001",
  61163=>"000011101",
  61164=>"001000010",
  61165=>"010111111",
  61166=>"001101010",
  61167=>"101100011",
  61168=>"111100100",
  61169=>"101101000",
  61170=>"001111110",
  61171=>"001100110",
  61172=>"100100100",
  61173=>"000111101",
  61174=>"110111001",
  61175=>"011100100",
  61176=>"110000110",
  61177=>"111110100",
  61178=>"111010111",
  61179=>"001001101",
  61180=>"011000101",
  61181=>"010111011",
  61182=>"011010000",
  61183=>"101101111",
  61184=>"111011000",
  61185=>"000011110",
  61186=>"111010001",
  61187=>"110001101",
  61188=>"111100111",
  61189=>"101011011",
  61190=>"000011111",
  61191=>"110100100",
  61192=>"100011000",
  61193=>"000100101",
  61194=>"111100111",
  61195=>"101010101",
  61196=>"011110111",
  61197=>"000110100",
  61198=>"110101111",
  61199=>"100001010",
  61200=>"111110001",
  61201=>"101011000",
  61202=>"001011000",
  61203=>"100111011",
  61204=>"100010000",
  61205=>"111111010",
  61206=>"001100110",
  61207=>"011000010",
  61208=>"110101101",
  61209=>"001101101",
  61210=>"101101101",
  61211=>"010010000",
  61212=>"111011011",
  61213=>"101111111",
  61214=>"010110111",
  61215=>"101101011",
  61216=>"110101010",
  61217=>"010001101",
  61218=>"100100000",
  61219=>"001001111",
  61220=>"011111101",
  61221=>"011010001",
  61222=>"111010000",
  61223=>"100101110",
  61224=>"011000100",
  61225=>"010110111",
  61226=>"010100110",
  61227=>"100001110",
  61228=>"001000110",
  61229=>"000010100",
  61230=>"100101101",
  61231=>"100001110",
  61232=>"011000101",
  61233=>"010011100",
  61234=>"101110001",
  61235=>"111100111",
  61236=>"011011001",
  61237=>"111110010",
  61238=>"110111110",
  61239=>"111111010",
  61240=>"110110111",
  61241=>"000100110",
  61242=>"100111001",
  61243=>"111111111",
  61244=>"000000111",
  61245=>"010110011",
  61246=>"100111001",
  61247=>"001100011",
  61248=>"000010000",
  61249=>"110010101",
  61250=>"000001100",
  61251=>"100100000",
  61252=>"111100111",
  61253=>"110011011",
  61254=>"010001100",
  61255=>"100111010",
  61256=>"110101111",
  61257=>"010010000",
  61258=>"111111101",
  61259=>"111110000",
  61260=>"110001100",
  61261=>"101000111",
  61262=>"110110011",
  61263=>"100100100",
  61264=>"000111010",
  61265=>"111001010",
  61266=>"001011001",
  61267=>"010000110",
  61268=>"111101101",
  61269=>"111111111",
  61270=>"010010000",
  61271=>"101011010",
  61272=>"000110111",
  61273=>"111011011",
  61274=>"001011001",
  61275=>"001001011",
  61276=>"000010111",
  61277=>"011000011",
  61278=>"001100000",
  61279=>"000101010",
  61280=>"010010010",
  61281=>"011011110",
  61282=>"001100000",
  61283=>"010001111",
  61284=>"110101101",
  61285=>"100101010",
  61286=>"100000000",
  61287=>"001111111",
  61288=>"001001100",
  61289=>"010000000",
  61290=>"101011101",
  61291=>"011001000",
  61292=>"011000001",
  61293=>"010000000",
  61294=>"110110111",
  61295=>"010011010",
  61296=>"100010000",
  61297=>"110001111",
  61298=>"011110101",
  61299=>"111100010",
  61300=>"010110101",
  61301=>"010110111",
  61302=>"110111110",
  61303=>"011011011",
  61304=>"001110000",
  61305=>"001000111",
  61306=>"011100110",
  61307=>"001010011",
  61308=>"110010000",
  61309=>"010001110",
  61310=>"011010101",
  61311=>"100110101",
  61312=>"100111011",
  61313=>"011010101",
  61314=>"011110101",
  61315=>"110100010",
  61316=>"110111111",
  61317=>"111101010",
  61318=>"000010010",
  61319=>"010010000",
  61320=>"010101110",
  61321=>"101111101",
  61322=>"000010110",
  61323=>"001101111",
  61324=>"111101111",
  61325=>"011111010",
  61326=>"110000010",
  61327=>"110001011",
  61328=>"101010001",
  61329=>"111001001",
  61330=>"001000001",
  61331=>"011011100",
  61332=>"100100101",
  61333=>"000111000",
  61334=>"100001101",
  61335=>"100001000",
  61336=>"011010000",
  61337=>"000000011",
  61338=>"010100000",
  61339=>"100010111",
  61340=>"101110000",
  61341=>"111100100",
  61342=>"001100101",
  61343=>"001011111",
  61344=>"001011000",
  61345=>"101111000",
  61346=>"001111111",
  61347=>"000101111",
  61348=>"100000100",
  61349=>"110000111",
  61350=>"110100001",
  61351=>"011011111",
  61352=>"110011010",
  61353=>"111101001",
  61354=>"011111011",
  61355=>"101010100",
  61356=>"111100111",
  61357=>"010011010",
  61358=>"110000000",
  61359=>"111111110",
  61360=>"101001111",
  61361=>"111000001",
  61362=>"101011010",
  61363=>"101011000",
  61364=>"011110011",
  61365=>"001110110",
  61366=>"011111001",
  61367=>"011101111",
  61368=>"111001001",
  61369=>"111100111",
  61370=>"011100110",
  61371=>"000010100",
  61372=>"111111000",
  61373=>"110001100",
  61374=>"000011110",
  61375=>"101000100",
  61376=>"011111110",
  61377=>"011110010",
  61378=>"101010001",
  61379=>"001111100",
  61380=>"001001001",
  61381=>"110111101",
  61382=>"111000000",
  61383=>"111001110",
  61384=>"111101101",
  61385=>"001010000",
  61386=>"110110110",
  61387=>"111101010",
  61388=>"100100111",
  61389=>"101011001",
  61390=>"101110110",
  61391=>"010011111",
  61392=>"011111010",
  61393=>"101111010",
  61394=>"101111111",
  61395=>"000110110",
  61396=>"011110110",
  61397=>"111111100",
  61398=>"000001101",
  61399=>"011001010",
  61400=>"010001010",
  61401=>"101111100",
  61402=>"110010001",
  61403=>"100101011",
  61404=>"111010001",
  61405=>"010000110",
  61406=>"010010011",
  61407=>"010010001",
  61408=>"100000110",
  61409=>"100110010",
  61410=>"001101111",
  61411=>"000000010",
  61412=>"010111011",
  61413=>"110010001",
  61414=>"101100110",
  61415=>"001011010",
  61416=>"001101111",
  61417=>"011010101",
  61418=>"110111101",
  61419=>"100100100",
  61420=>"011100001",
  61421=>"110011111",
  61422=>"011101100",
  61423=>"100010110",
  61424=>"010000000",
  61425=>"001000101",
  61426=>"101001110",
  61427=>"100000100",
  61428=>"000001010",
  61429=>"110111111",
  61430=>"001011010",
  61431=>"000110001",
  61432=>"100110011",
  61433=>"101011101",
  61434=>"101110110",
  61435=>"111001001",
  61436=>"000001000",
  61437=>"101111000",
  61438=>"110011110",
  61439=>"000011011",
  61440=>"000110111",
  61441=>"100000001",
  61442=>"111100010",
  61443=>"011010001",
  61444=>"001011101",
  61445=>"100001001",
  61446=>"010010010",
  61447=>"000001111",
  61448=>"111100110",
  61449=>"111010101",
  61450=>"101101010",
  61451=>"010010100",
  61452=>"001111001",
  61453=>"011010011",
  61454=>"101100100",
  61455=>"100010000",
  61456=>"110100000",
  61457=>"111100001",
  61458=>"110110000",
  61459=>"100100110",
  61460=>"011001011",
  61461=>"001000010",
  61462=>"101010100",
  61463=>"100001011",
  61464=>"011001101",
  61465=>"011100001",
  61466=>"000100101",
  61467=>"111000101",
  61468=>"111101111",
  61469=>"110101101",
  61470=>"100111001",
  61471=>"100010010",
  61472=>"111001000",
  61473=>"010111100",
  61474=>"010000100",
  61475=>"110001010",
  61476=>"000001100",
  61477=>"001010101",
  61478=>"010011000",
  61479=>"001000111",
  61480=>"001000011",
  61481=>"011110010",
  61482=>"000000101",
  61483=>"010100101",
  61484=>"111000001",
  61485=>"101101010",
  61486=>"100010001",
  61487=>"100011110",
  61488=>"010111111",
  61489=>"110111101",
  61490=>"010101111",
  61491=>"111101000",
  61492=>"100111011",
  61493=>"001100101",
  61494=>"110011010",
  61495=>"111011000",
  61496=>"001010100",
  61497=>"000110000",
  61498=>"101101000",
  61499=>"111000001",
  61500=>"010001000",
  61501=>"100101111",
  61502=>"000110010",
  61503=>"010010001",
  61504=>"111100100",
  61505=>"010010101",
  61506=>"111111011",
  61507=>"001011010",
  61508=>"010101100",
  61509=>"111110100",
  61510=>"110010010",
  61511=>"111100010",
  61512=>"101001001",
  61513=>"000011110",
  61514=>"001110010",
  61515=>"110011010",
  61516=>"011101110",
  61517=>"001111111",
  61518=>"011011010",
  61519=>"000001010",
  61520=>"000111101",
  61521=>"111000001",
  61522=>"111101011",
  61523=>"111111101",
  61524=>"011001011",
  61525=>"110001101",
  61526=>"100100101",
  61527=>"011111111",
  61528=>"010000001",
  61529=>"001000101",
  61530=>"011111110",
  61531=>"000010110",
  61532=>"101000000",
  61533=>"100010100",
  61534=>"000110111",
  61535=>"110011101",
  61536=>"111101110",
  61537=>"100100001",
  61538=>"001001100",
  61539=>"000010101",
  61540=>"011001111",
  61541=>"101111110",
  61542=>"011010101",
  61543=>"011001100",
  61544=>"100001110",
  61545=>"100001111",
  61546=>"100001010",
  61547=>"011001001",
  61548=>"001100101",
  61549=>"111110110",
  61550=>"101100001",
  61551=>"010000010",
  61552=>"011011110",
  61553=>"101010001",
  61554=>"010000000",
  61555=>"010110011",
  61556=>"010010010",
  61557=>"011011110",
  61558=>"000100101",
  61559=>"011010110",
  61560=>"011001000",
  61561=>"110111111",
  61562=>"110011110",
  61563=>"000000000",
  61564=>"111010000",
  61565=>"111010111",
  61566=>"010101101",
  61567=>"110011110",
  61568=>"111101010",
  61569=>"111011111",
  61570=>"100101111",
  61571=>"000100000",
  61572=>"110101110",
  61573=>"011110100",
  61574=>"100010101",
  61575=>"101001101",
  61576=>"010100010",
  61577=>"011110101",
  61578=>"011110101",
  61579=>"010011100",
  61580=>"101011111",
  61581=>"101100100",
  61582=>"011110011",
  61583=>"000011000",
  61584=>"111111010",
  61585=>"100000101",
  61586=>"110000000",
  61587=>"110010111",
  61588=>"100111010",
  61589=>"100000000",
  61590=>"100110101",
  61591=>"011011101",
  61592=>"000001011",
  61593=>"000010110",
  61594=>"011111110",
  61595=>"011110000",
  61596=>"001000110",
  61597=>"011011010",
  61598=>"100110011",
  61599=>"100100111",
  61600=>"010010010",
  61601=>"111001000",
  61602=>"110110111",
  61603=>"001100000",
  61604=>"100100101",
  61605=>"010101010",
  61606=>"011100001",
  61607=>"110101011",
  61608=>"001011010",
  61609=>"000011010",
  61610=>"000011001",
  61611=>"111100101",
  61612=>"010010100",
  61613=>"110100100",
  61614=>"011010001",
  61615=>"011101111",
  61616=>"000111100",
  61617=>"111101111",
  61618=>"011100101",
  61619=>"100001001",
  61620=>"000001011",
  61621=>"110000100",
  61622=>"010011110",
  61623=>"111011001",
  61624=>"100100100",
  61625=>"100010111",
  61626=>"001110111",
  61627=>"001010100",
  61628=>"011011001",
  61629=>"010001011",
  61630=>"010000010",
  61631=>"001111010",
  61632=>"010010101",
  61633=>"101110110",
  61634=>"100001011",
  61635=>"000101011",
  61636=>"011000100",
  61637=>"110000111",
  61638=>"000101010",
  61639=>"110101111",
  61640=>"100100100",
  61641=>"011010100",
  61642=>"111101100",
  61643=>"110000001",
  61644=>"001001011",
  61645=>"010001100",
  61646=>"010101110",
  61647=>"101101101",
  61648=>"001110101",
  61649=>"001111101",
  61650=>"001111101",
  61651=>"001000001",
  61652=>"001010100",
  61653=>"011011100",
  61654=>"101001010",
  61655=>"110000001",
  61656=>"000100011",
  61657=>"011101110",
  61658=>"000010100",
  61659=>"011101010",
  61660=>"000110100",
  61661=>"000110110",
  61662=>"100001000",
  61663=>"011110111",
  61664=>"000000011",
  61665=>"111100011",
  61666=>"000001001",
  61667=>"001011100",
  61668=>"100001100",
  61669=>"000110111",
  61670=>"100000010",
  61671=>"110101111",
  61672=>"101010101",
  61673=>"111011010",
  61674=>"001111100",
  61675=>"001000011",
  61676=>"010001101",
  61677=>"010010011",
  61678=>"010001111",
  61679=>"011000010",
  61680=>"000100110",
  61681=>"000101011",
  61682=>"111111111",
  61683=>"001000100",
  61684=>"110110011",
  61685=>"110111000",
  61686=>"101001010",
  61687=>"000111011",
  61688=>"000010011",
  61689=>"000100010",
  61690=>"011000100",
  61691=>"101011011",
  61692=>"111100011",
  61693=>"000110000",
  61694=>"110101110",
  61695=>"111001001",
  61696=>"001101011",
  61697=>"010100001",
  61698=>"110101110",
  61699=>"010100101",
  61700=>"111010101",
  61701=>"001000010",
  61702=>"110111001",
  61703=>"100010101",
  61704=>"010111111",
  61705=>"000110110",
  61706=>"101110101",
  61707=>"000101001",
  61708=>"101001001",
  61709=>"011001000",
  61710=>"111011110",
  61711=>"111110011",
  61712=>"001111100",
  61713=>"000110101",
  61714=>"111101110",
  61715=>"011011010",
  61716=>"101111111",
  61717=>"001111100",
  61718=>"001011111",
  61719=>"111010111",
  61720=>"010010011",
  61721=>"101110110",
  61722=>"110001110",
  61723=>"110101101",
  61724=>"001100101",
  61725=>"110000010",
  61726=>"110001011",
  61727=>"110110011",
  61728=>"001101000",
  61729=>"101000001",
  61730=>"111110101",
  61731=>"000111111",
  61732=>"000101100",
  61733=>"101100010",
  61734=>"100111101",
  61735=>"111000010",
  61736=>"000011001",
  61737=>"101010101",
  61738=>"001110110",
  61739=>"110110010",
  61740=>"011101101",
  61741=>"011001000",
  61742=>"000111110",
  61743=>"000000001",
  61744=>"011001000",
  61745=>"011101011",
  61746=>"111011101",
  61747=>"100001010",
  61748=>"100000110",
  61749=>"110010101",
  61750=>"110100111",
  61751=>"111111111",
  61752=>"011011110",
  61753=>"111100100",
  61754=>"010101110",
  61755=>"010010101",
  61756=>"101011110",
  61757=>"000011010",
  61758=>"010101100",
  61759=>"001111101",
  61760=>"010001100",
  61761=>"110110000",
  61762=>"100001011",
  61763=>"100100011",
  61764=>"110101101",
  61765=>"101100001",
  61766=>"110000111",
  61767=>"101110101",
  61768=>"110001001",
  61769=>"100000101",
  61770=>"111111001",
  61771=>"100000101",
  61772=>"111000010",
  61773=>"000101101",
  61774=>"110011101",
  61775=>"100110000",
  61776=>"110111100",
  61777=>"101001100",
  61778=>"000100110",
  61779=>"000001110",
  61780=>"111000110",
  61781=>"001100000",
  61782=>"111100011",
  61783=>"100000010",
  61784=>"000010001",
  61785=>"010001011",
  61786=>"010101010",
  61787=>"001100110",
  61788=>"001101010",
  61789=>"100000101",
  61790=>"111001110",
  61791=>"010100001",
  61792=>"100000101",
  61793=>"110111011",
  61794=>"011001011",
  61795=>"101000101",
  61796=>"011101101",
  61797=>"110111001",
  61798=>"111001011",
  61799=>"011111000",
  61800=>"110000001",
  61801=>"111100011",
  61802=>"011100110",
  61803=>"100100000",
  61804=>"001101000",
  61805=>"110111011",
  61806=>"111111110",
  61807=>"000110111",
  61808=>"101101111",
  61809=>"000001001",
  61810=>"000011010",
  61811=>"101111101",
  61812=>"011100010",
  61813=>"111101101",
  61814=>"001101101",
  61815=>"110101100",
  61816=>"101001111",
  61817=>"110101000",
  61818=>"000110110",
  61819=>"101011000",
  61820=>"111101110",
  61821=>"110101011",
  61822=>"011010011",
  61823=>"111111101",
  61824=>"111101111",
  61825=>"111011000",
  61826=>"010001101",
  61827=>"010001001",
  61828=>"111100110",
  61829=>"011110001",
  61830=>"110110111",
  61831=>"001001010",
  61832=>"000001011",
  61833=>"111111100",
  61834=>"101000000",
  61835=>"001001111",
  61836=>"111011110",
  61837=>"001001010",
  61838=>"111011001",
  61839=>"101111010",
  61840=>"101110000",
  61841=>"011001011",
  61842=>"110110000",
  61843=>"110001001",
  61844=>"011111101",
  61845=>"000000100",
  61846=>"101000100",
  61847=>"001010000",
  61848=>"101010101",
  61849=>"100011101",
  61850=>"011100001",
  61851=>"100110100",
  61852=>"101100101",
  61853=>"110011001",
  61854=>"010000100",
  61855=>"110010000",
  61856=>"000010010",
  61857=>"011000001",
  61858=>"011010111",
  61859=>"010101000",
  61860=>"100000100",
  61861=>"000011101",
  61862=>"001111001",
  61863=>"111111110",
  61864=>"110001001",
  61865=>"010010111",
  61866=>"000000111",
  61867=>"100100010",
  61868=>"100111100",
  61869=>"001011111",
  61870=>"111000101",
  61871=>"000001110",
  61872=>"000011110",
  61873=>"000110101",
  61874=>"001100000",
  61875=>"101000011",
  61876=>"110011000",
  61877=>"101111101",
  61878=>"110110101",
  61879=>"001001101",
  61880=>"001110001",
  61881=>"100110111",
  61882=>"001110010",
  61883=>"001111111",
  61884=>"110110010",
  61885=>"001000011",
  61886=>"111110111",
  61887=>"101000110",
  61888=>"000011101",
  61889=>"001110110",
  61890=>"111001110",
  61891=>"010010101",
  61892=>"100001001",
  61893=>"010100110",
  61894=>"000011101",
  61895=>"101110110",
  61896=>"100111110",
  61897=>"000111100",
  61898=>"101101000",
  61899=>"110100010",
  61900=>"011111000",
  61901=>"001111011",
  61902=>"100000011",
  61903=>"101100010",
  61904=>"100011001",
  61905=>"000000100",
  61906=>"011101111",
  61907=>"101100011",
  61908=>"101000110",
  61909=>"001100001",
  61910=>"110101101",
  61911=>"101101011",
  61912=>"000111000",
  61913=>"010110100",
  61914=>"010011101",
  61915=>"010111000",
  61916=>"111010111",
  61917=>"000101011",
  61918=>"100100101",
  61919=>"110011111",
  61920=>"000011010",
  61921=>"010111001",
  61922=>"100110111",
  61923=>"111101000",
  61924=>"100001000",
  61925=>"110100010",
  61926=>"000101010",
  61927=>"010001110",
  61928=>"000010000",
  61929=>"101110111",
  61930=>"110010111",
  61931=>"010000111",
  61932=>"101000000",
  61933=>"101011001",
  61934=>"000010110",
  61935=>"001000010",
  61936=>"010010010",
  61937=>"000111110",
  61938=>"100001110",
  61939=>"001001000",
  61940=>"110010110",
  61941=>"111100110",
  61942=>"100110111",
  61943=>"000101011",
  61944=>"000011010",
  61945=>"011110101",
  61946=>"000111110",
  61947=>"011000010",
  61948=>"010001010",
  61949=>"110011111",
  61950=>"111101001",
  61951=>"010100010",
  61952=>"000111011",
  61953=>"011001111",
  61954=>"010110000",
  61955=>"110111100",
  61956=>"110010100",
  61957=>"110100001",
  61958=>"011111010",
  61959=>"101111100",
  61960=>"000100001",
  61961=>"111011010",
  61962=>"011110110",
  61963=>"101010111",
  61964=>"111000001",
  61965=>"110110101",
  61966=>"010010111",
  61967=>"011100000",
  61968=>"101010001",
  61969=>"001100011",
  61970=>"001000101",
  61971=>"111011110",
  61972=>"110100101",
  61973=>"000001110",
  61974=>"100000001",
  61975=>"001101111",
  61976=>"011110111",
  61977=>"000100010",
  61978=>"111100010",
  61979=>"110111000",
  61980=>"000011110",
  61981=>"001111011",
  61982=>"010010110",
  61983=>"110000010",
  61984=>"011010000",
  61985=>"101011101",
  61986=>"000010110",
  61987=>"100101111",
  61988=>"100001110",
  61989=>"111011111",
  61990=>"000100001",
  61991=>"110011110",
  61992=>"111000010",
  61993=>"101000101",
  61994=>"001111011",
  61995=>"010110011",
  61996=>"100111100",
  61997=>"001100001",
  61998=>"010110000",
  61999=>"111000101",
  62000=>"110011110",
  62001=>"001100000",
  62002=>"110101100",
  62003=>"100100000",
  62004=>"101101000",
  62005=>"111011100",
  62006=>"110100000",
  62007=>"011101001",
  62008=>"000011000",
  62009=>"011110101",
  62010=>"001110100",
  62011=>"111110111",
  62012=>"001101110",
  62013=>"011110100",
  62014=>"100111000",
  62015=>"010011111",
  62016=>"101001000",
  62017=>"011011001",
  62018=>"011110100",
  62019=>"000010101",
  62020=>"101011100",
  62021=>"111010100",
  62022=>"000110101",
  62023=>"100100100",
  62024=>"010001100",
  62025=>"100100110",
  62026=>"100110110",
  62027=>"101101111",
  62028=>"110000100",
  62029=>"010010010",
  62030=>"111000101",
  62031=>"000001010",
  62032=>"110010100",
  62033=>"111011001",
  62034=>"010001000",
  62035=>"011000010",
  62036=>"100100001",
  62037=>"011111010",
  62038=>"100000101",
  62039=>"010001101",
  62040=>"010101111",
  62041=>"100110111",
  62042=>"010101010",
  62043=>"011001011",
  62044=>"111011001",
  62045=>"000000001",
  62046=>"011111111",
  62047=>"000110011",
  62048=>"000111010",
  62049=>"100000010",
  62050=>"100000100",
  62051=>"110100001",
  62052=>"101101010",
  62053=>"000010101",
  62054=>"100110010",
  62055=>"010011011",
  62056=>"011001011",
  62057=>"001001101",
  62058=>"001101110",
  62059=>"111011000",
  62060=>"101010000",
  62061=>"111111000",
  62062=>"011010010",
  62063=>"010011011",
  62064=>"001111011",
  62065=>"001100010",
  62066=>"111110111",
  62067=>"011101111",
  62068=>"101001000",
  62069=>"011100001",
  62070=>"110000010",
  62071=>"010110001",
  62072=>"000011000",
  62073=>"010000100",
  62074=>"010011111",
  62075=>"001101001",
  62076=>"110010110",
  62077=>"100000011",
  62078=>"011110101",
  62079=>"111000111",
  62080=>"001000101",
  62081=>"001010101",
  62082=>"000111010",
  62083=>"111100010",
  62084=>"100011110",
  62085=>"100001100",
  62086=>"110110101",
  62087=>"110101110",
  62088=>"100111010",
  62089=>"101011010",
  62090=>"111101011",
  62091=>"111001110",
  62092=>"001000000",
  62093=>"110010101",
  62094=>"000000101",
  62095=>"000111111",
  62096=>"111111010",
  62097=>"111001100",
  62098=>"000101010",
  62099=>"100000000",
  62100=>"001100010",
  62101=>"011001100",
  62102=>"011010101",
  62103=>"101011101",
  62104=>"011110101",
  62105=>"011000000",
  62106=>"111011110",
  62107=>"110000011",
  62108=>"111001001",
  62109=>"110110011",
  62110=>"111001111",
  62111=>"101110100",
  62112=>"001001110",
  62113=>"110111010",
  62114=>"011101000",
  62115=>"110101101",
  62116=>"111111001",
  62117=>"101101010",
  62118=>"000110010",
  62119=>"000110010",
  62120=>"111100111",
  62121=>"100010110",
  62122=>"011111000",
  62123=>"100001000",
  62124=>"000101101",
  62125=>"000011100",
  62126=>"000101101",
  62127=>"000110001",
  62128=>"010111010",
  62129=>"011011111",
  62130=>"111000101",
  62131=>"101111000",
  62132=>"110011101",
  62133=>"000101110",
  62134=>"000101110",
  62135=>"010110111",
  62136=>"010001000",
  62137=>"010111010",
  62138=>"101011100",
  62139=>"110100000",
  62140=>"110101011",
  62141=>"000111000",
  62142=>"110000010",
  62143=>"001011011",
  62144=>"101010100",
  62145=>"100001101",
  62146=>"111001011",
  62147=>"111111101",
  62148=>"111101101",
  62149=>"000010000",
  62150=>"100001011",
  62151=>"111000101",
  62152=>"101100111",
  62153=>"101000010",
  62154=>"111110111",
  62155=>"111010101",
  62156=>"000010001",
  62157=>"010011000",
  62158=>"000000001",
  62159=>"111001001",
  62160=>"100000010",
  62161=>"010011000",
  62162=>"101010011",
  62163=>"000000011",
  62164=>"111111110",
  62165=>"100101010",
  62166=>"010101110",
  62167=>"011110110",
  62168=>"010000001",
  62169=>"110010100",
  62170=>"101100101",
  62171=>"011101111",
  62172=>"010111111",
  62173=>"111101000",
  62174=>"100100110",
  62175=>"101000101",
  62176=>"010100111",
  62177=>"001100000",
  62178=>"101010100",
  62179=>"100110011",
  62180=>"101110010",
  62181=>"001111111",
  62182=>"111110010",
  62183=>"101000000",
  62184=>"100010101",
  62185=>"100011100",
  62186=>"010010000",
  62187=>"110000001",
  62188=>"010110011",
  62189=>"010011000",
  62190=>"111001001",
  62191=>"110001011",
  62192=>"010000011",
  62193=>"010111000",
  62194=>"000011011",
  62195=>"110101100",
  62196=>"011001010",
  62197=>"000011111",
  62198=>"100010100",
  62199=>"001000100",
  62200=>"000111010",
  62201=>"110010100",
  62202=>"000010000",
  62203=>"001110111",
  62204=>"111111001",
  62205=>"111111011",
  62206=>"101011000",
  62207=>"101011010",
  62208=>"111010110",
  62209=>"010101010",
  62210=>"010101001",
  62211=>"011001100",
  62212=>"010001100",
  62213=>"010000111",
  62214=>"100001010",
  62215=>"111011011",
  62216=>"010101101",
  62217=>"001100111",
  62218=>"101110001",
  62219=>"000100110",
  62220=>"111110011",
  62221=>"000010110",
  62222=>"110111111",
  62223=>"011101111",
  62224=>"100000110",
  62225=>"001001001",
  62226=>"011110101",
  62227=>"001111000",
  62228=>"101100111",
  62229=>"111011000",
  62230=>"011001111",
  62231=>"100110100",
  62232=>"000111110",
  62233=>"111000010",
  62234=>"010100101",
  62235=>"010010111",
  62236=>"001111000",
  62237=>"011000000",
  62238=>"101001100",
  62239=>"010000110",
  62240=>"100101110",
  62241=>"011101011",
  62242=>"000000000",
  62243=>"010000101",
  62244=>"010001011",
  62245=>"111100111",
  62246=>"110001001",
  62247=>"011001011",
  62248=>"111001110",
  62249=>"101001101",
  62250=>"101011111",
  62251=>"001001100",
  62252=>"100111101",
  62253=>"000110100",
  62254=>"111111000",
  62255=>"000011110",
  62256=>"100100101",
  62257=>"011100000",
  62258=>"000001110",
  62259=>"111110010",
  62260=>"011001011",
  62261=>"000100111",
  62262=>"000100100",
  62263=>"100001001",
  62264=>"011000001",
  62265=>"111011101",
  62266=>"000101100",
  62267=>"110111010",
  62268=>"110000111",
  62269=>"010111011",
  62270=>"001001101",
  62271=>"010000011",
  62272=>"100100100",
  62273=>"011000001",
  62274=>"111011101",
  62275=>"100000111",
  62276=>"111001100",
  62277=>"001010000",
  62278=>"110110100",
  62279=>"000000000",
  62280=>"110100011",
  62281=>"111111111",
  62282=>"010000100",
  62283=>"101101001",
  62284=>"110000101",
  62285=>"011110101",
  62286=>"001100001",
  62287=>"100111001",
  62288=>"111111010",
  62289=>"010001011",
  62290=>"100110110",
  62291=>"110000010",
  62292=>"110000110",
  62293=>"110100100",
  62294=>"011001010",
  62295=>"100001101",
  62296=>"001111100",
  62297=>"000000001",
  62298=>"010010010",
  62299=>"001000000",
  62300=>"101011010",
  62301=>"001000011",
  62302=>"011111001",
  62303=>"000000010",
  62304=>"000010110",
  62305=>"011001111",
  62306=>"110001010",
  62307=>"100111110",
  62308=>"000111010",
  62309=>"001111111",
  62310=>"001110010",
  62311=>"110010001",
  62312=>"011011000",
  62313=>"100110110",
  62314=>"110011011",
  62315=>"001001110",
  62316=>"011110011",
  62317=>"100010010",
  62318=>"111000010",
  62319=>"101011000",
  62320=>"010110000",
  62321=>"011001010",
  62322=>"111111100",
  62323=>"100110011",
  62324=>"001111100",
  62325=>"000110000",
  62326=>"011001110",
  62327=>"000010111",
  62328=>"100110011",
  62329=>"111000101",
  62330=>"000000000",
  62331=>"101100110",
  62332=>"001011101",
  62333=>"111110111",
  62334=>"000010000",
  62335=>"000000000",
  62336=>"100010011",
  62337=>"001110101",
  62338=>"000111000",
  62339=>"000110000",
  62340=>"100010010",
  62341=>"010011110",
  62342=>"010000100",
  62343=>"001111110",
  62344=>"001000010",
  62345=>"100010101",
  62346=>"011101010",
  62347=>"010100001",
  62348=>"110001011",
  62349=>"001000101",
  62350=>"001101111",
  62351=>"001111010",
  62352=>"001010011",
  62353=>"011111011",
  62354=>"101001100",
  62355=>"000110100",
  62356=>"111110000",
  62357=>"110100001",
  62358=>"001111110",
  62359=>"000000010",
  62360=>"100000011",
  62361=>"110000100",
  62362=>"100001111",
  62363=>"011010100",
  62364=>"010101110",
  62365=>"010111111",
  62366=>"111010100",
  62367=>"010011100",
  62368=>"001101000",
  62369=>"000101110",
  62370=>"111111011",
  62371=>"100000001",
  62372=>"000110110",
  62373=>"000000000",
  62374=>"001000101",
  62375=>"001101000",
  62376=>"001110110",
  62377=>"000010000",
  62378=>"110101001",
  62379=>"101101110",
  62380=>"100001010",
  62381=>"111000111",
  62382=>"100110011",
  62383=>"010011010",
  62384=>"011011110",
  62385=>"010100000",
  62386=>"101111010",
  62387=>"101011100",
  62388=>"110101110",
  62389=>"000001010",
  62390=>"111110110",
  62391=>"110101000",
  62392=>"000000101",
  62393=>"010000001",
  62394=>"100111110",
  62395=>"100100100",
  62396=>"011101001",
  62397=>"010100010",
  62398=>"101100010",
  62399=>"001111001",
  62400=>"101100111",
  62401=>"000000000",
  62402=>"000111000",
  62403=>"100001000",
  62404=>"101001010",
  62405=>"101000001",
  62406=>"100001110",
  62407=>"001111110",
  62408=>"110010111",
  62409=>"010101100",
  62410=>"101001111",
  62411=>"100000011",
  62412=>"000110111",
  62413=>"000100001",
  62414=>"000001000",
  62415=>"111101011",
  62416=>"011011001",
  62417=>"110000000",
  62418=>"111010000",
  62419=>"110001011",
  62420=>"111001111",
  62421=>"111011111",
  62422=>"100010110",
  62423=>"001111100",
  62424=>"010100100",
  62425=>"100010000",
  62426=>"010110100",
  62427=>"110101111",
  62428=>"010010110",
  62429=>"110000000",
  62430=>"101111111",
  62431=>"000000110",
  62432=>"010000111",
  62433=>"011001111",
  62434=>"010101010",
  62435=>"001000011",
  62436=>"110010011",
  62437=>"111100100",
  62438=>"101110111",
  62439=>"100111101",
  62440=>"100000111",
  62441=>"110101100",
  62442=>"110010100",
  62443=>"100000110",
  62444=>"100111110",
  62445=>"010000111",
  62446=>"010111101",
  62447=>"010110111",
  62448=>"100000001",
  62449=>"101101111",
  62450=>"110000111",
  62451=>"010110010",
  62452=>"010100011",
  62453=>"011001000",
  62454=>"001100010",
  62455=>"100000001",
  62456=>"111010001",
  62457=>"101001100",
  62458=>"110110100",
  62459=>"111111000",
  62460=>"100001101",
  62461=>"110011010",
  62462=>"111101111",
  62463=>"011100000",
  62464=>"101101000",
  62465=>"000011010",
  62466=>"001110110",
  62467=>"110011011",
  62468=>"110001100",
  62469=>"111110010",
  62470=>"101011010",
  62471=>"010010000",
  62472=>"111001001",
  62473=>"000001000",
  62474=>"110000101",
  62475=>"010011010",
  62476=>"110101111",
  62477=>"101001001",
  62478=>"000001110",
  62479=>"000100011",
  62480=>"110100110",
  62481=>"011100011",
  62482=>"111111110",
  62483=>"011110001",
  62484=>"111110111",
  62485=>"011110000",
  62486=>"001011010",
  62487=>"100101001",
  62488=>"011001110",
  62489=>"101000111",
  62490=>"010011101",
  62491=>"001011011",
  62492=>"111101100",
  62493=>"101011110",
  62494=>"011011100",
  62495=>"100111010",
  62496=>"000100010",
  62497=>"000110000",
  62498=>"010100100",
  62499=>"101110101",
  62500=>"101100101",
  62501=>"000001010",
  62502=>"010100000",
  62503=>"101011100",
  62504=>"110110101",
  62505=>"111010101",
  62506=>"011100011",
  62507=>"001101111",
  62508=>"001001100",
  62509=>"001110101",
  62510=>"110101111",
  62511=>"000010110",
  62512=>"101010111",
  62513=>"001001101",
  62514=>"010101000",
  62515=>"100111110",
  62516=>"110000001",
  62517=>"111111111",
  62518=>"100011000",
  62519=>"100011011",
  62520=>"100101110",
  62521=>"010100011",
  62522=>"110110110",
  62523=>"101010110",
  62524=>"001100101",
  62525=>"010101011",
  62526=>"111111011",
  62527=>"100110111",
  62528=>"100000101",
  62529=>"000010100",
  62530=>"000100011",
  62531=>"000000011",
  62532=>"111000101",
  62533=>"010011001",
  62534=>"011100000",
  62535=>"100000011",
  62536=>"111110100",
  62537=>"001000110",
  62538=>"111111011",
  62539=>"101000011",
  62540=>"010110100",
  62541=>"011111100",
  62542=>"011100001",
  62543=>"000011011",
  62544=>"101101000",
  62545=>"001001000",
  62546=>"010101000",
  62547=>"000001010",
  62548=>"111111010",
  62549=>"010001101",
  62550=>"100000001",
  62551=>"101000100",
  62552=>"010001101",
  62553=>"110110111",
  62554=>"001100001",
  62555=>"010100111",
  62556=>"101111100",
  62557=>"000010111",
  62558=>"111110111",
  62559=>"000101100",
  62560=>"000000011",
  62561=>"110001100",
  62562=>"100001100",
  62563=>"011101000",
  62564=>"111011011",
  62565=>"111000010",
  62566=>"101011101",
  62567=>"010100100",
  62568=>"101001000",
  62569=>"101000101",
  62570=>"100001111",
  62571=>"000000010",
  62572=>"101111110",
  62573=>"111100110",
  62574=>"110111111",
  62575=>"011001111",
  62576=>"100000011",
  62577=>"011100000",
  62578=>"111101011",
  62579=>"111000111",
  62580=>"111000111",
  62581=>"001011011",
  62582=>"011111110",
  62583=>"111001111",
  62584=>"100100010",
  62585=>"000100111",
  62586=>"100100110",
  62587=>"001100101",
  62588=>"010000111",
  62589=>"111010100",
  62590=>"100001001",
  62591=>"010011000",
  62592=>"100110101",
  62593=>"110100011",
  62594=>"111101100",
  62595=>"010111010",
  62596=>"010000001",
  62597=>"010100111",
  62598=>"011000000",
  62599=>"010110001",
  62600=>"111010110",
  62601=>"100001000",
  62602=>"101110010",
  62603=>"100110010",
  62604=>"000011111",
  62605=>"101111100",
  62606=>"111100011",
  62607=>"111110001",
  62608=>"011101000",
  62609=>"011000000",
  62610=>"110001111",
  62611=>"011001100",
  62612=>"100000111",
  62613=>"000111101",
  62614=>"011000101",
  62615=>"011100011",
  62616=>"010000001",
  62617=>"001011111",
  62618=>"011101011",
  62619=>"010001100",
  62620=>"101100011",
  62621=>"001000010",
  62622=>"000101110",
  62623=>"100101100",
  62624=>"111010101",
  62625=>"011011000",
  62626=>"000011011",
  62627=>"001111101",
  62628=>"101101111",
  62629=>"011100101",
  62630=>"011001011",
  62631=>"111010000",
  62632=>"011001001",
  62633=>"000000110",
  62634=>"100011001",
  62635=>"001111110",
  62636=>"010000001",
  62637=>"011111100",
  62638=>"100001110",
  62639=>"100110000",
  62640=>"011000001",
  62641=>"010101001",
  62642=>"101001110",
  62643=>"111101001",
  62644=>"100101110",
  62645=>"111110100",
  62646=>"011001100",
  62647=>"011001100",
  62648=>"100010101",
  62649=>"110111110",
  62650=>"111100110",
  62651=>"000101100",
  62652=>"100100111",
  62653=>"110011111",
  62654=>"111111000",
  62655=>"101111011",
  62656=>"011011010",
  62657=>"110101010",
  62658=>"011111101",
  62659=>"111100001",
  62660=>"111000001",
  62661=>"000010000",
  62662=>"111111001",
  62663=>"101100011",
  62664=>"111111110",
  62665=>"100101111",
  62666=>"101100111",
  62667=>"100111100",
  62668=>"100110010",
  62669=>"110111111",
  62670=>"101101110",
  62671=>"101000001",
  62672=>"100000110",
  62673=>"001101001",
  62674=>"101010110",
  62675=>"001100010",
  62676=>"000111011",
  62677=>"000010100",
  62678=>"100001000",
  62679=>"011011110",
  62680=>"010010110",
  62681=>"010010111",
  62682=>"011010000",
  62683=>"101011000",
  62684=>"100100001",
  62685=>"101001011",
  62686=>"011000110",
  62687=>"101011111",
  62688=>"110110011",
  62689=>"110111000",
  62690=>"101111001",
  62691=>"001110001",
  62692=>"110010000",
  62693=>"000100011",
  62694=>"000100000",
  62695=>"110101101",
  62696=>"011010010",
  62697=>"000000101",
  62698=>"111110011",
  62699=>"101010010",
  62700=>"000010000",
  62701=>"101100000",
  62702=>"001011100",
  62703=>"000110110",
  62704=>"100011111",
  62705=>"111110111",
  62706=>"000010001",
  62707=>"111101000",
  62708=>"100100000",
  62709=>"010011000",
  62710=>"001000101",
  62711=>"101010100",
  62712=>"100100010",
  62713=>"010111001",
  62714=>"001010011",
  62715=>"000001100",
  62716=>"001110100",
  62717=>"100110000",
  62718=>"100111010",
  62719=>"111110101",
  62720=>"101111001",
  62721=>"110111010",
  62722=>"111001101",
  62723=>"100100001",
  62724=>"100100101",
  62725=>"000001000",
  62726=>"100101110",
  62727=>"100111110",
  62728=>"000101010",
  62729=>"000001111",
  62730=>"111111001",
  62731=>"000001110",
  62732=>"000001011",
  62733=>"111100101",
  62734=>"010010100",
  62735=>"010001011",
  62736=>"111000001",
  62737=>"010001001",
  62738=>"010100000",
  62739=>"101111100",
  62740=>"100100100",
  62741=>"011101100",
  62742=>"110100101",
  62743=>"001000101",
  62744=>"010011000",
  62745=>"110101000",
  62746=>"000101110",
  62747=>"110010001",
  62748=>"001100001",
  62749=>"010110100",
  62750=>"110101011",
  62751=>"001000001",
  62752=>"100111100",
  62753=>"001111000",
  62754=>"110100001",
  62755=>"110101110",
  62756=>"111111000",
  62757=>"000101110",
  62758=>"101110101",
  62759=>"110111111",
  62760=>"101100000",
  62761=>"110011111",
  62762=>"011101000",
  62763=>"001110011",
  62764=>"111111010",
  62765=>"110001001",
  62766=>"100001001",
  62767=>"010100100",
  62768=>"010101110",
  62769=>"000001000",
  62770=>"001100001",
  62771=>"100111011",
  62772=>"011010101",
  62773=>"001111000",
  62774=>"010001001",
  62775=>"111110010",
  62776=>"100100101",
  62777=>"000011110",
  62778=>"101101010",
  62779=>"111000101",
  62780=>"011011000",
  62781=>"011111100",
  62782=>"010011100",
  62783=>"010101000",
  62784=>"010100111",
  62785=>"110111110",
  62786=>"111111101",
  62787=>"010010000",
  62788=>"100011010",
  62789=>"101001110",
  62790=>"100110111",
  62791=>"111001011",
  62792=>"010011111",
  62793=>"110001010",
  62794=>"111011010",
  62795=>"001100001",
  62796=>"111111010",
  62797=>"010101000",
  62798=>"010010010",
  62799=>"011011010",
  62800=>"110001011",
  62801=>"100000011",
  62802=>"010100010",
  62803=>"111011111",
  62804=>"010110001",
  62805=>"000011110",
  62806=>"010010101",
  62807=>"011011011",
  62808=>"101000110",
  62809=>"101101111",
  62810=>"101100010",
  62811=>"001101010",
  62812=>"101101100",
  62813=>"111001100",
  62814=>"001001011",
  62815=>"101010110",
  62816=>"100011110",
  62817=>"111111100",
  62818=>"101101001",
  62819=>"010101001",
  62820=>"101110110",
  62821=>"010100000",
  62822=>"010000111",
  62823=>"111011001",
  62824=>"001010101",
  62825=>"000001100",
  62826=>"001011101",
  62827=>"100010100",
  62828=>"011110100",
  62829=>"111111111",
  62830=>"011000000",
  62831=>"101101001",
  62832=>"000100111",
  62833=>"110010110",
  62834=>"100010001",
  62835=>"111111101",
  62836=>"111001100",
  62837=>"110011001",
  62838=>"010001110",
  62839=>"101100111",
  62840=>"011000000",
  62841=>"111000001",
  62842=>"010011001",
  62843=>"110010111",
  62844=>"010110000",
  62845=>"111011100",
  62846=>"000011011",
  62847=>"001000001",
  62848=>"111100000",
  62849=>"110000001",
  62850=>"000011110",
  62851=>"001010010",
  62852=>"101101101",
  62853=>"000011101",
  62854=>"111100001",
  62855=>"101111011",
  62856=>"001100000",
  62857=>"000111111",
  62858=>"110100000",
  62859=>"011010011",
  62860=>"000000001",
  62861=>"111110101",
  62862=>"110001111",
  62863=>"011101110",
  62864=>"000010100",
  62865=>"011001011",
  62866=>"010001111",
  62867=>"111111001",
  62868=>"001101101",
  62869=>"011110010",
  62870=>"010111011",
  62871=>"010010100",
  62872=>"111000100",
  62873=>"000000001",
  62874=>"010001001",
  62875=>"000110000",
  62876=>"110011001",
  62877=>"100000010",
  62878=>"010101011",
  62879=>"011001101",
  62880=>"010010001",
  62881=>"011111010",
  62882=>"100011010",
  62883=>"001100100",
  62884=>"010100100",
  62885=>"001100011",
  62886=>"101100011",
  62887=>"111101111",
  62888=>"011001000",
  62889=>"001000000",
  62890=>"000010110",
  62891=>"101010111",
  62892=>"111100111",
  62893=>"111010010",
  62894=>"000111000",
  62895=>"000110010",
  62896=>"010100011",
  62897=>"000111011",
  62898=>"101101101",
  62899=>"111110111",
  62900=>"110100110",
  62901=>"011111110",
  62902=>"010010110",
  62903=>"101101110",
  62904=>"001001010",
  62905=>"011011000",
  62906=>"110010101",
  62907=>"101010000",
  62908=>"010111001",
  62909=>"001100100",
  62910=>"010101010",
  62911=>"100001011",
  62912=>"000100010",
  62913=>"110010111",
  62914=>"101111111",
  62915=>"000001011",
  62916=>"001100100",
  62917=>"111010101",
  62918=>"111001101",
  62919=>"011001001",
  62920=>"000000000",
  62921=>"001100101",
  62922=>"110101000",
  62923=>"000001000",
  62924=>"001110100",
  62925=>"010100000",
  62926=>"001001111",
  62927=>"000010011",
  62928=>"000100001",
  62929=>"001000101",
  62930=>"111101111",
  62931=>"011010010",
  62932=>"010001101",
  62933=>"100111000",
  62934=>"001000011",
  62935=>"010100001",
  62936=>"011111001",
  62937=>"110010011",
  62938=>"110111110",
  62939=>"000100011",
  62940=>"000110110",
  62941=>"010100110",
  62942=>"001101100",
  62943=>"101111111",
  62944=>"001000000",
  62945=>"111000001",
  62946=>"011010001",
  62947=>"000001010",
  62948=>"001100101",
  62949=>"001010010",
  62950=>"101101100",
  62951=>"101010110",
  62952=>"010101000",
  62953=>"000010000",
  62954=>"101000100",
  62955=>"100001001",
  62956=>"000101011",
  62957=>"010011111",
  62958=>"000001000",
  62959=>"001000001",
  62960=>"001010010",
  62961=>"011011100",
  62962=>"001001111",
  62963=>"000000110",
  62964=>"101001100",
  62965=>"010001000",
  62966=>"101001110",
  62967=>"001000100",
  62968=>"001010101",
  62969=>"000010000",
  62970=>"001000000",
  62971=>"001100001",
  62972=>"110101111",
  62973=>"001000010",
  62974=>"011000011",
  62975=>"001010001",
  62976=>"101001010",
  62977=>"101100111",
  62978=>"110010110",
  62979=>"001000111",
  62980=>"111101000",
  62981=>"101011100",
  62982=>"101010010",
  62983=>"010001000",
  62984=>"001000000",
  62985=>"100100100",
  62986=>"001111011",
  62987=>"000100111",
  62988=>"100100000",
  62989=>"000100010",
  62990=>"001011010",
  62991=>"001000010",
  62992=>"001111100",
  62993=>"011010010",
  62994=>"101010111",
  62995=>"111011100",
  62996=>"110010011",
  62997=>"101010101",
  62998=>"011111010",
  62999=>"110001011",
  63000=>"000001111",
  63001=>"011111010",
  63002=>"011010110",
  63003=>"000011111",
  63004=>"100111000",
  63005=>"111101101",
  63006=>"111011110",
  63007=>"010000111",
  63008=>"000100100",
  63009=>"111110110",
  63010=>"001000111",
  63011=>"000001100",
  63012=>"010011110",
  63013=>"010001100",
  63014=>"001011010",
  63015=>"011011010",
  63016=>"010010111",
  63017=>"011000011",
  63018=>"001110001",
  63019=>"101011011",
  63020=>"111010111",
  63021=>"101100011",
  63022=>"000000000",
  63023=>"010001100",
  63024=>"000000111",
  63025=>"000110100",
  63026=>"111110110",
  63027=>"011110111",
  63028=>"110000001",
  63029=>"111000110",
  63030=>"100111000",
  63031=>"110010010",
  63032=>"111100010",
  63033=>"100100011",
  63034=>"101111100",
  63035=>"100101110",
  63036=>"001011110",
  63037=>"110110110",
  63038=>"011000000",
  63039=>"111111101",
  63040=>"001110111",
  63041=>"000101001",
  63042=>"000101101",
  63043=>"110000110",
  63044=>"111101001",
  63045=>"110111100",
  63046=>"000000010",
  63047=>"100111000",
  63048=>"000100111",
  63049=>"011111110",
  63050=>"100111110",
  63051=>"100101011",
  63052=>"010000111",
  63053=>"100101101",
  63054=>"100010111",
  63055=>"101000110",
  63056=>"011100011",
  63057=>"111011111",
  63058=>"111010101",
  63059=>"010011010",
  63060=>"010001100",
  63061=>"001000110",
  63062=>"001000010",
  63063=>"001110111",
  63064=>"000001101",
  63065=>"001100011",
  63066=>"101101101",
  63067=>"010101010",
  63068=>"101101010",
  63069=>"111001000",
  63070=>"010100011",
  63071=>"110000010",
  63072=>"100000011",
  63073=>"000001000",
  63074=>"111000010",
  63075=>"010110001",
  63076=>"000100111",
  63077=>"110110100",
  63078=>"101011001",
  63079=>"100001100",
  63080=>"100010110",
  63081=>"110000101",
  63082=>"110000111",
  63083=>"110100110",
  63084=>"000011110",
  63085=>"011001010",
  63086=>"100111101",
  63087=>"001101100",
  63088=>"101011100",
  63089=>"110101101",
  63090=>"000001001",
  63091=>"000011010",
  63092=>"111101110",
  63093=>"010000011",
  63094=>"000100000",
  63095=>"011111011",
  63096=>"001010101",
  63097=>"011001000",
  63098=>"001010000",
  63099=>"110110010",
  63100=>"111111011",
  63101=>"001001000",
  63102=>"100100001",
  63103=>"001100100",
  63104=>"001011000",
  63105=>"100101110",
  63106=>"100011001",
  63107=>"101111010",
  63108=>"010111001",
  63109=>"111011000",
  63110=>"101101110",
  63111=>"001011000",
  63112=>"000011110",
  63113=>"110101101",
  63114=>"111101101",
  63115=>"111000101",
  63116=>"000110111",
  63117=>"110101111",
  63118=>"100100100",
  63119=>"011000110",
  63120=>"110111001",
  63121=>"011001101",
  63122=>"100000010",
  63123=>"100111100",
  63124=>"000101111",
  63125=>"101101100",
  63126=>"111011001",
  63127=>"001001010",
  63128=>"111100100",
  63129=>"101110110",
  63130=>"001001110",
  63131=>"111111001",
  63132=>"010100000",
  63133=>"111001100",
  63134=>"000110111",
  63135=>"001011001",
  63136=>"000001000",
  63137=>"000111111",
  63138=>"010100101",
  63139=>"001010000",
  63140=>"011001000",
  63141=>"001001000",
  63142=>"100000000",
  63143=>"001111011",
  63144=>"000010011",
  63145=>"010000011",
  63146=>"110011111",
  63147=>"001110110",
  63148=>"001000000",
  63149=>"100011011",
  63150=>"000111001",
  63151=>"101001111",
  63152=>"111010010",
  63153=>"010001110",
  63154=>"100110001",
  63155=>"010110100",
  63156=>"010000000",
  63157=>"010100110",
  63158=>"010110010",
  63159=>"011010000",
  63160=>"111100011",
  63161=>"110010110",
  63162=>"001111011",
  63163=>"000111011",
  63164=>"111000010",
  63165=>"100110101",
  63166=>"000001000",
  63167=>"000101101",
  63168=>"010101110",
  63169=>"000011110",
  63170=>"000000100",
  63171=>"100001111",
  63172=>"010001001",
  63173=>"100101001",
  63174=>"000110100",
  63175=>"000110000",
  63176=>"101011110",
  63177=>"101111100",
  63178=>"101010111",
  63179=>"011111001",
  63180=>"001110001",
  63181=>"010111000",
  63182=>"001011000",
  63183=>"010100110",
  63184=>"100100110",
  63185=>"100111010",
  63186=>"111010111",
  63187=>"000001010",
  63188=>"011100111",
  63189=>"101100010",
  63190=>"100001101",
  63191=>"100110100",
  63192=>"100000000",
  63193=>"011111101",
  63194=>"011110000",
  63195=>"001111101",
  63196=>"100110000",
  63197=>"110000011",
  63198=>"100000110",
  63199=>"110001100",
  63200=>"001001011",
  63201=>"101011110",
  63202=>"110100010",
  63203=>"100001001",
  63204=>"111100100",
  63205=>"000111001",
  63206=>"010111011",
  63207=>"101101011",
  63208=>"100000000",
  63209=>"101000111",
  63210=>"111111110",
  63211=>"010111011",
  63212=>"111010100",
  63213=>"010111101",
  63214=>"000001100",
  63215=>"010011010",
  63216=>"011011010",
  63217=>"000011000",
  63218=>"010000000",
  63219=>"001100111",
  63220=>"000010011",
  63221=>"111011100",
  63222=>"010001100",
  63223=>"111111110",
  63224=>"100111011",
  63225=>"010110110",
  63226=>"000100110",
  63227=>"000110101",
  63228=>"011000001",
  63229=>"100011101",
  63230=>"010000010",
  63231=>"001011001",
  63232=>"010011110",
  63233=>"001111000",
  63234=>"000001101",
  63235=>"000000101",
  63236=>"101100100",
  63237=>"100110110",
  63238=>"110000010",
  63239=>"111011110",
  63240=>"010100010",
  63241=>"001011100",
  63242=>"111110010",
  63243=>"011001010",
  63244=>"111110100",
  63245=>"110101001",
  63246=>"111110000",
  63247=>"010001001",
  63248=>"000001110",
  63249=>"110011101",
  63250=>"110111000",
  63251=>"001000010",
  63252=>"011001110",
  63253=>"100001001",
  63254=>"011011010",
  63255=>"000001011",
  63256=>"000110000",
  63257=>"001001010",
  63258=>"010111110",
  63259=>"100011000",
  63260=>"011110001",
  63261=>"111110001",
  63262=>"101010011",
  63263=>"011100011",
  63264=>"100001001",
  63265=>"100100111",
  63266=>"111101011",
  63267=>"001100010",
  63268=>"100000111",
  63269=>"000110000",
  63270=>"000111011",
  63271=>"000001100",
  63272=>"011100111",
  63273=>"101000001",
  63274=>"000111111",
  63275=>"111111110",
  63276=>"110010010",
  63277=>"100001000",
  63278=>"110111100",
  63279=>"101111101",
  63280=>"010001111",
  63281=>"111111010",
  63282=>"001010011",
  63283=>"000111000",
  63284=>"111111111",
  63285=>"010110100",
  63286=>"000110000",
  63287=>"010000001",
  63288=>"010101001",
  63289=>"101000011",
  63290=>"100101010",
  63291=>"110001000",
  63292=>"010010000",
  63293=>"100100011",
  63294=>"000010110",
  63295=>"101111111",
  63296=>"011011111",
  63297=>"111110111",
  63298=>"011000000",
  63299=>"101111100",
  63300=>"011010000",
  63301=>"000000010",
  63302=>"001010011",
  63303=>"011001011",
  63304=>"101011100",
  63305=>"101011111",
  63306=>"110100111",
  63307=>"010101000",
  63308=>"001001001",
  63309=>"100000110",
  63310=>"011001000",
  63311=>"111010000",
  63312=>"111101111",
  63313=>"000010001",
  63314=>"100000010",
  63315=>"011000101",
  63316=>"000101011",
  63317=>"011110110",
  63318=>"111110001",
  63319=>"110100101",
  63320=>"110001001",
  63321=>"110000001",
  63322=>"011011000",
  63323=>"000011001",
  63324=>"000111011",
  63325=>"001000001",
  63326=>"110000001",
  63327=>"001010011",
  63328=>"110111100",
  63329=>"000000001",
  63330=>"001010011",
  63331=>"000001111",
  63332=>"111110000",
  63333=>"100010100",
  63334=>"000110001",
  63335=>"001110110",
  63336=>"100111001",
  63337=>"100001101",
  63338=>"001001101",
  63339=>"010011110",
  63340=>"111111100",
  63341=>"011001100",
  63342=>"100100011",
  63343=>"101001110",
  63344=>"110000101",
  63345=>"101100110",
  63346=>"011000110",
  63347=>"000101111",
  63348=>"000100110",
  63349=>"111111110",
  63350=>"111010001",
  63351=>"101010000",
  63352=>"100011010",
  63353=>"100101101",
  63354=>"000001110",
  63355=>"000010000",
  63356=>"001010111",
  63357=>"110111101",
  63358=>"000101000",
  63359=>"010111100",
  63360=>"000111001",
  63361=>"101111000",
  63362=>"100010110",
  63363=>"010111101",
  63364=>"100100010",
  63365=>"000011100",
  63366=>"101110001",
  63367=>"100110100",
  63368=>"111111001",
  63369=>"101111001",
  63370=>"000011011",
  63371=>"000111000",
  63372=>"011100001",
  63373=>"101110011",
  63374=>"011100101",
  63375=>"000010000",
  63376=>"100011000",
  63377=>"110011010",
  63378=>"000000010",
  63379=>"101111010",
  63380=>"101110100",
  63381=>"101011010",
  63382=>"001110111",
  63383=>"111111111",
  63384=>"111111111",
  63385=>"111101100",
  63386=>"110000101",
  63387=>"110001100",
  63388=>"001110011",
  63389=>"101001110",
  63390=>"100011100",
  63391=>"111111011",
  63392=>"010011100",
  63393=>"110101101",
  63394=>"111110100",
  63395=>"010000001",
  63396=>"001010100",
  63397=>"110100101",
  63398=>"010100100",
  63399=>"100110100",
  63400=>"001010111",
  63401=>"101101111",
  63402=>"101100000",
  63403=>"100111101",
  63404=>"100000000",
  63405=>"011100101",
  63406=>"001001110",
  63407=>"000100111",
  63408=>"001010111",
  63409=>"111001001",
  63410=>"000101000",
  63411=>"001000010",
  63412=>"100010100",
  63413=>"010010111",
  63414=>"110100011",
  63415=>"110001010",
  63416=>"101011000",
  63417=>"100010110",
  63418=>"101011101",
  63419=>"001101111",
  63420=>"100010001",
  63421=>"111101110",
  63422=>"000001100",
  63423=>"101001010",
  63424=>"001010011",
  63425=>"110000001",
  63426=>"000010000",
  63427=>"011100011",
  63428=>"111001101",
  63429=>"010000010",
  63430=>"101000111",
  63431=>"001111101",
  63432=>"010100101",
  63433=>"010110011",
  63434=>"110111110",
  63435=>"011011011",
  63436=>"100111011",
  63437=>"001111000",
  63438=>"100010111",
  63439=>"010001000",
  63440=>"010110111",
  63441=>"010111010",
  63442=>"011001000",
  63443=>"000111111",
  63444=>"110010101",
  63445=>"101111111",
  63446=>"000101110",
  63447=>"100011111",
  63448=>"101101111",
  63449=>"110000110",
  63450=>"001001011",
  63451=>"110011111",
  63452=>"100010000",
  63453=>"100101110",
  63454=>"100010111",
  63455=>"010001111",
  63456=>"000111111",
  63457=>"111010000",
  63458=>"010011100",
  63459=>"100100110",
  63460=>"001001100",
  63461=>"000011001",
  63462=>"111000010",
  63463=>"111101001",
  63464=>"000000100",
  63465=>"111010011",
  63466=>"000111110",
  63467=>"000011111",
  63468=>"110001110",
  63469=>"000111110",
  63470=>"101100000",
  63471=>"110111011",
  63472=>"010110010",
  63473=>"000101100",
  63474=>"101001100",
  63475=>"000001100",
  63476=>"111010110",
  63477=>"100111110",
  63478=>"000001010",
  63479=>"011110110",
  63480=>"111010111",
  63481=>"011011000",
  63482=>"010010100",
  63483=>"101110111",
  63484=>"101100011",
  63485=>"111110100",
  63486=>"001111011",
  63487=>"011011100",
  63488=>"001101100",
  63489=>"001111101",
  63490=>"100011101",
  63491=>"111110110",
  63492=>"000111100",
  63493=>"100011101",
  63494=>"101011111",
  63495=>"111110011",
  63496=>"000011101",
  63497=>"111000101",
  63498=>"101010110",
  63499=>"101110010",
  63500=>"001100001",
  63501=>"000111001",
  63502=>"100001110",
  63503=>"000100110",
  63504=>"001010001",
  63505=>"010110010",
  63506=>"000000001",
  63507=>"000101011",
  63508=>"000011001",
  63509=>"100011100",
  63510=>"111001110",
  63511=>"000011000",
  63512=>"000101111",
  63513=>"101001101",
  63514=>"100110000",
  63515=>"010011100",
  63516=>"101000100",
  63517=>"010001111",
  63518=>"101010010",
  63519=>"011110110",
  63520=>"000000110",
  63521=>"100000001",
  63522=>"101111000",
  63523=>"011010101",
  63524=>"110001011",
  63525=>"101110110",
  63526=>"000001011",
  63527=>"110001111",
  63528=>"000110110",
  63529=>"010011101",
  63530=>"110101110",
  63531=>"000100100",
  63532=>"111110100",
  63533=>"100000110",
  63534=>"001001100",
  63535=>"000000001",
  63536=>"111110011",
  63537=>"001110011",
  63538=>"110100111",
  63539=>"111101100",
  63540=>"001101010",
  63541=>"100110110",
  63542=>"001001110",
  63543=>"110110001",
  63544=>"001100001",
  63545=>"010110010",
  63546=>"110000111",
  63547=>"100111100",
  63548=>"111111100",
  63549=>"001100011",
  63550=>"010111110",
  63551=>"001110011",
  63552=>"101100011",
  63553=>"110110110",
  63554=>"111001111",
  63555=>"010110100",
  63556=>"000010000",
  63557=>"101100100",
  63558=>"001001100",
  63559=>"101111111",
  63560=>"000011101",
  63561=>"111101111",
  63562=>"000000011",
  63563=>"010010011",
  63564=>"000100010",
  63565=>"010110101",
  63566=>"000110101",
  63567=>"011100000",
  63568=>"000101000",
  63569=>"100110000",
  63570=>"000001110",
  63571=>"010101100",
  63572=>"111111100",
  63573=>"001010111",
  63574=>"101111010",
  63575=>"110110001",
  63576=>"000100001",
  63577=>"110001001",
  63578=>"101001010",
  63579=>"000000011",
  63580=>"101110000",
  63581=>"000111001",
  63582=>"110101100",
  63583=>"010110101",
  63584=>"111011100",
  63585=>"101011101",
  63586=>"100110011",
  63587=>"011011010",
  63588=>"100011001",
  63589=>"100011010",
  63590=>"111000000",
  63591=>"000011111",
  63592=>"101010010",
  63593=>"100010010",
  63594=>"001110001",
  63595=>"001101100",
  63596=>"010010010",
  63597=>"010100001",
  63598=>"000010100",
  63599=>"111010011",
  63600=>"111101010",
  63601=>"010001000",
  63602=>"101010111",
  63603=>"001000001",
  63604=>"100100000",
  63605=>"011101111",
  63606=>"000011101",
  63607=>"001111010",
  63608=>"011110000",
  63609=>"111000100",
  63610=>"000000111",
  63611=>"101011101",
  63612=>"111100111",
  63613=>"101100100",
  63614=>"000000100",
  63615=>"010110100",
  63616=>"011011110",
  63617=>"011010010",
  63618=>"111011111",
  63619=>"110000001",
  63620=>"001101001",
  63621=>"010110110",
  63622=>"111101111",
  63623=>"010100111",
  63624=>"011111101",
  63625=>"010011000",
  63626=>"101101101",
  63627=>"000111101",
  63628=>"010110001",
  63629=>"100001000",
  63630=>"111101110",
  63631=>"111110100",
  63632=>"100001011",
  63633=>"011001111",
  63634=>"111001110",
  63635=>"001010100",
  63636=>"111101111",
  63637=>"011000100",
  63638=>"100101011",
  63639=>"010110100",
  63640=>"010101000",
  63641=>"101100111",
  63642=>"110011000",
  63643=>"011001010",
  63644=>"000000011",
  63645=>"010100101",
  63646=>"100010011",
  63647=>"100001010",
  63648=>"000001101",
  63649=>"100100101",
  63650=>"001100011",
  63651=>"011010011",
  63652=>"000001011",
  63653=>"000010010",
  63654=>"111101000",
  63655=>"110011010",
  63656=>"100011101",
  63657=>"110000010",
  63658=>"100010000",
  63659=>"100110101",
  63660=>"001010000",
  63661=>"100011100",
  63662=>"011011111",
  63663=>"100000000",
  63664=>"010000010",
  63665=>"111101111",
  63666=>"000001011",
  63667=>"100111010",
  63668=>"011110001",
  63669=>"000111111",
  63670=>"100111110",
  63671=>"111101111",
  63672=>"000100011",
  63673=>"110101101",
  63674=>"010101101",
  63675=>"101001100",
  63676=>"100001110",
  63677=>"000100101",
  63678=>"111010001",
  63679=>"001010000",
  63680=>"011011110",
  63681=>"110001110",
  63682=>"010011100",
  63683=>"001110011",
  63684=>"100011011",
  63685=>"111100100",
  63686=>"100011100",
  63687=>"111101001",
  63688=>"011100001",
  63689=>"101100101",
  63690=>"001110000",
  63691=>"110011110",
  63692=>"000101111",
  63693=>"010100100",
  63694=>"001101100",
  63695=>"100001101",
  63696=>"001000001",
  63697=>"111100100",
  63698=>"011110010",
  63699=>"011111001",
  63700=>"111001000",
  63701=>"100000001",
  63702=>"011110010",
  63703=>"001001000",
  63704=>"010000011",
  63705=>"010001110",
  63706=>"000110111",
  63707=>"011001101",
  63708=>"000100010",
  63709=>"110011110",
  63710=>"100111111",
  63711=>"010010111",
  63712=>"110001011",
  63713=>"001000001",
  63714=>"011010010",
  63715=>"000001111",
  63716=>"100100000",
  63717=>"000011101",
  63718=>"000100100",
  63719=>"000110100",
  63720=>"011010001",
  63721=>"101000110",
  63722=>"101011010",
  63723=>"001100100",
  63724=>"000000001",
  63725=>"011100110",
  63726=>"101010010",
  63727=>"100101001",
  63728=>"100101010",
  63729=>"110100111",
  63730=>"011001111",
  63731=>"000011111",
  63732=>"010110101",
  63733=>"101100101",
  63734=>"111111001",
  63735=>"000000011",
  63736=>"110110000",
  63737=>"011101001",
  63738=>"101110110",
  63739=>"000111011",
  63740=>"100001100",
  63741=>"011001101",
  63742=>"111010000",
  63743=>"110110011",
  63744=>"001001100",
  63745=>"010011111",
  63746=>"001111110",
  63747=>"111010100",
  63748=>"001010001",
  63749=>"010000111",
  63750=>"111111100",
  63751=>"111001111",
  63752=>"111101111",
  63753=>"001001010",
  63754=>"101101101",
  63755=>"000100010",
  63756=>"010101111",
  63757=>"000001001",
  63758=>"110000111",
  63759=>"000100100",
  63760=>"011100010",
  63761=>"111100001",
  63762=>"110001100",
  63763=>"100000101",
  63764=>"100001000",
  63765=>"100110100",
  63766=>"111111010",
  63767=>"110010001",
  63768=>"101001001",
  63769=>"001001101",
  63770=>"111100111",
  63771=>"011111010",
  63772=>"000101100",
  63773=>"100011100",
  63774=>"101101011",
  63775=>"000000101",
  63776=>"101111001",
  63777=>"000000011",
  63778=>"010100001",
  63779=>"110110010",
  63780=>"010110000",
  63781=>"111011001",
  63782=>"010101111",
  63783=>"011010110",
  63784=>"110001000",
  63785=>"000100111",
  63786=>"110100111",
  63787=>"001001111",
  63788=>"111110111",
  63789=>"111110101",
  63790=>"100101001",
  63791=>"111101000",
  63792=>"000101000",
  63793=>"101011100",
  63794=>"111010100",
  63795=>"100011001",
  63796=>"011111101",
  63797=>"100111010",
  63798=>"000111110",
  63799=>"001000100",
  63800=>"101011000",
  63801=>"000100001",
  63802=>"111101000",
  63803=>"100000100",
  63804=>"101010101",
  63805=>"101111001",
  63806=>"010000000",
  63807=>"010100011",
  63808=>"011011110",
  63809=>"001100001",
  63810=>"110001000",
  63811=>"111111010",
  63812=>"110010010",
  63813=>"110010100",
  63814=>"101000110",
  63815=>"011110100",
  63816=>"010000111",
  63817=>"011100000",
  63818=>"000010110",
  63819=>"011010100",
  63820=>"100001000",
  63821=>"111010110",
  63822=>"010001111",
  63823=>"100000010",
  63824=>"011010011",
  63825=>"011111111",
  63826=>"000000010",
  63827=>"101001110",
  63828=>"010111101",
  63829=>"110001011",
  63830=>"100111101",
  63831=>"101100001",
  63832=>"110000010",
  63833=>"000010100",
  63834=>"000000101",
  63835=>"101101000",
  63836=>"010100100",
  63837=>"010111010",
  63838=>"110100000",
  63839=>"111111101",
  63840=>"000001111",
  63841=>"011010101",
  63842=>"010000011",
  63843=>"110100010",
  63844=>"100100110",
  63845=>"011111001",
  63846=>"000000010",
  63847=>"110011010",
  63848=>"000110101",
  63849=>"001110000",
  63850=>"010100101",
  63851=>"100100010",
  63852=>"011010110",
  63853=>"110000000",
  63854=>"001010110",
  63855=>"101010010",
  63856=>"110111010",
  63857=>"000101110",
  63858=>"001100010",
  63859=>"010110101",
  63860=>"000101010",
  63861=>"101111111",
  63862=>"000000111",
  63863=>"100111101",
  63864=>"000010010",
  63865=>"001001100",
  63866=>"011010010",
  63867=>"011001001",
  63868=>"101111000",
  63869=>"010001011",
  63870=>"011100110",
  63871=>"010001000",
  63872=>"110110001",
  63873=>"100110110",
  63874=>"011101001",
  63875=>"110111000",
  63876=>"111010001",
  63877=>"010100010",
  63878=>"011100001",
  63879=>"110001000",
  63880=>"000010110",
  63881=>"100000100",
  63882=>"011010011",
  63883=>"001100110",
  63884=>"110010111",
  63885=>"000000111",
  63886=>"001111001",
  63887=>"011111100",
  63888=>"111100101",
  63889=>"111101010",
  63890=>"110010001",
  63891=>"111111011",
  63892=>"101111010",
  63893=>"001100110",
  63894=>"110101110",
  63895=>"000110100",
  63896=>"101101100",
  63897=>"001011101",
  63898=>"011101111",
  63899=>"011010001",
  63900=>"101110111",
  63901=>"111000000",
  63902=>"111111100",
  63903=>"100001010",
  63904=>"011000000",
  63905=>"111100110",
  63906=>"000010100",
  63907=>"010010000",
  63908=>"111110000",
  63909=>"101101111",
  63910=>"000111001",
  63911=>"011000000",
  63912=>"111000100",
  63913=>"100100100",
  63914=>"000010111",
  63915=>"110001000",
  63916=>"001111110",
  63917=>"011000111",
  63918=>"100111101",
  63919=>"100000110",
  63920=>"111010111",
  63921=>"001000001",
  63922=>"110100111",
  63923=>"001000001",
  63924=>"101100101",
  63925=>"111101100",
  63926=>"000000001",
  63927=>"001010011",
  63928=>"111111101",
  63929=>"101101100",
  63930=>"000011001",
  63931=>"001000000",
  63932=>"001011110",
  63933=>"110000100",
  63934=>"100110011",
  63935=>"000010010",
  63936=>"111101101",
  63937=>"000100110",
  63938=>"011100100",
  63939=>"001100011",
  63940=>"110101111",
  63941=>"010010011",
  63942=>"010010000",
  63943=>"000000101",
  63944=>"100101111",
  63945=>"010010000",
  63946=>"101110001",
  63947=>"011100110",
  63948=>"111101100",
  63949=>"000011110",
  63950=>"010100000",
  63951=>"100111100",
  63952=>"001101110",
  63953=>"000101001",
  63954=>"010101101",
  63955=>"100101111",
  63956=>"010100111",
  63957=>"111101011",
  63958=>"000010000",
  63959=>"110001101",
  63960=>"101001011",
  63961=>"100110100",
  63962=>"101101111",
  63963=>"111001001",
  63964=>"001100011",
  63965=>"101101111",
  63966=>"001010001",
  63967=>"011010110",
  63968=>"000000101",
  63969=>"010001101",
  63970=>"111111110",
  63971=>"111011111",
  63972=>"000100000",
  63973=>"111111111",
  63974=>"100001101",
  63975=>"000100111",
  63976=>"011001011",
  63977=>"100111111",
  63978=>"111111110",
  63979=>"000100001",
  63980=>"000100001",
  63981=>"101110000",
  63982=>"101110000",
  63983=>"010100011",
  63984=>"100110001",
  63985=>"010000001",
  63986=>"111101111",
  63987=>"001001011",
  63988=>"011001011",
  63989=>"111000010",
  63990=>"110100101",
  63991=>"110010001",
  63992=>"011101001",
  63993=>"001001001",
  63994=>"110111001",
  63995=>"100000000",
  63996=>"101010001",
  63997=>"111111011",
  63998=>"010001000",
  63999=>"111000101",
  64000=>"010111111",
  64001=>"110001100",
  64002=>"101100100",
  64003=>"101000000",
  64004=>"011001011",
  64005=>"010000000",
  64006=>"010100011",
  64007=>"111101000",
  64008=>"011101010",
  64009=>"010100110",
  64010=>"111101100",
  64011=>"011110000",
  64012=>"111011001",
  64013=>"010111100",
  64014=>"010001111",
  64015=>"111000001",
  64016=>"100001010",
  64017=>"001111111",
  64018=>"111000110",
  64019=>"111111110",
  64020=>"101100101",
  64021=>"111010111",
  64022=>"111011111",
  64023=>"100111010",
  64024=>"110111011",
  64025=>"000001110",
  64026=>"011101001",
  64027=>"010000000",
  64028=>"000101110",
  64029=>"110110011",
  64030=>"001101000",
  64031=>"110111100",
  64032=>"111110101",
  64033=>"110110010",
  64034=>"001110001",
  64035=>"011101100",
  64036=>"111110000",
  64037=>"111001011",
  64038=>"011111101",
  64039=>"000101000",
  64040=>"110000100",
  64041=>"100010110",
  64042=>"101100100",
  64043=>"010011011",
  64044=>"000000000",
  64045=>"101111001",
  64046=>"011101111",
  64047=>"111011111",
  64048=>"001000001",
  64049=>"100100010",
  64050=>"111010010",
  64051=>"000011001",
  64052=>"000001010",
  64053=>"100100101",
  64054=>"001010101",
  64055=>"101100011",
  64056=>"101101001",
  64057=>"000100000",
  64058=>"000001110",
  64059=>"001111110",
  64060=>"010011011",
  64061=>"010100111",
  64062=>"000011010",
  64063=>"001001100",
  64064=>"010011010",
  64065=>"111000111",
  64066=>"100100001",
  64067=>"101010010",
  64068=>"001010110",
  64069=>"111111111",
  64070=>"000111111",
  64071=>"010011100",
  64072=>"000001011",
  64073=>"111111011",
  64074=>"000111111",
  64075=>"011111101",
  64076=>"100101101",
  64077=>"100011110",
  64078=>"101011111",
  64079=>"011100010",
  64080=>"111101101",
  64081=>"000101111",
  64082=>"000011000",
  64083=>"011100011",
  64084=>"011100011",
  64085=>"011110011",
  64086=>"000001010",
  64087=>"011100111",
  64088=>"000001101",
  64089=>"111111100",
  64090=>"001101101",
  64091=>"001101000",
  64092=>"011110100",
  64093=>"000000001",
  64094=>"010010011",
  64095=>"001101000",
  64096=>"101001000",
  64097=>"100000111",
  64098=>"111011100",
  64099=>"010000111",
  64100=>"100101011",
  64101=>"010011010",
  64102=>"101000111",
  64103=>"010101001",
  64104=>"100000001",
  64105=>"100011010",
  64106=>"000000001",
  64107=>"001100100",
  64108=>"110101010",
  64109=>"110101100",
  64110=>"011111101",
  64111=>"000100100",
  64112=>"101000001",
  64113=>"011011111",
  64114=>"101010000",
  64115=>"001001000",
  64116=>"110011001",
  64117=>"110001011",
  64118=>"000111111",
  64119=>"111101111",
  64120=>"111111010",
  64121=>"010101100",
  64122=>"010100100",
  64123=>"000001110",
  64124=>"100100100",
  64125=>"011001100",
  64126=>"101011010",
  64127=>"110010101",
  64128=>"101011000",
  64129=>"110001110",
  64130=>"110011011",
  64131=>"111000001",
  64132=>"011011110",
  64133=>"001000001",
  64134=>"001101101",
  64135=>"110111000",
  64136=>"011110001",
  64137=>"111010000",
  64138=>"101111100",
  64139=>"110001001",
  64140=>"001110100",
  64141=>"101110000",
  64142=>"101100101",
  64143=>"100111000",
  64144=>"110111000",
  64145=>"101010110",
  64146=>"010000010",
  64147=>"100010011",
  64148=>"101000000",
  64149=>"001011111",
  64150=>"011000100",
  64151=>"011110101",
  64152=>"100110101",
  64153=>"001000011",
  64154=>"001111000",
  64155=>"011100100",
  64156=>"011001100",
  64157=>"001010101",
  64158=>"111110011",
  64159=>"101111001",
  64160=>"010001011",
  64161=>"100011100",
  64162=>"010011111",
  64163=>"110100011",
  64164=>"110101101",
  64165=>"100011010",
  64166=>"111111010",
  64167=>"000000101",
  64168=>"111011011",
  64169=>"100000001",
  64170=>"010101010",
  64171=>"110001101",
  64172=>"100001011",
  64173=>"000000100",
  64174=>"000001110",
  64175=>"110001100",
  64176=>"111101110",
  64177=>"001100111",
  64178=>"110110010",
  64179=>"011000110",
  64180=>"101100110",
  64181=>"111111111",
  64182=>"101000100",
  64183=>"110011000",
  64184=>"000110000",
  64185=>"101111010",
  64186=>"110100001",
  64187=>"000100000",
  64188=>"001001011",
  64189=>"001010001",
  64190=>"110101000",
  64191=>"001111100",
  64192=>"111010001",
  64193=>"111011101",
  64194=>"100010000",
  64195=>"001010010",
  64196=>"100110011",
  64197=>"110110110",
  64198=>"001011001",
  64199=>"010101001",
  64200=>"000010110",
  64201=>"100001101",
  64202=>"101011100",
  64203=>"000010100",
  64204=>"011111010",
  64205=>"101001000",
  64206=>"011000001",
  64207=>"111101010",
  64208=>"011110000",
  64209=>"000110010",
  64210=>"011001101",
  64211=>"001111101",
  64212=>"111110111",
  64213=>"110010010",
  64214=>"110101000",
  64215=>"011101000",
  64216=>"011111011",
  64217=>"010011101",
  64218=>"100010001",
  64219=>"110011011",
  64220=>"010111000",
  64221=>"111111000",
  64222=>"001010100",
  64223=>"001111111",
  64224=>"010101011",
  64225=>"111001001",
  64226=>"011000011",
  64227=>"011001011",
  64228=>"100001100",
  64229=>"100110000",
  64230=>"110011001",
  64231=>"001001001",
  64232=>"000001111",
  64233=>"101011101",
  64234=>"011111101",
  64235=>"100111111",
  64236=>"110000011",
  64237=>"110000100",
  64238=>"110001110",
  64239=>"101000011",
  64240=>"100111100",
  64241=>"110101011",
  64242=>"111100111",
  64243=>"001110100",
  64244=>"110100101",
  64245=>"010001000",
  64246=>"001100000",
  64247=>"110000001",
  64248=>"011000111",
  64249=>"000010110",
  64250=>"101110000",
  64251=>"001111101",
  64252=>"110100111",
  64253=>"111101111",
  64254=>"100101110",
  64255=>"000000110",
  64256=>"111110100",
  64257=>"010100000",
  64258=>"010001100",
  64259=>"110001000",
  64260=>"000001010",
  64261=>"001111011",
  64262=>"011011110",
  64263=>"010000101",
  64264=>"111001101",
  64265=>"111110101",
  64266=>"111110101",
  64267=>"000000100",
  64268=>"101000100",
  64269=>"100111001",
  64270=>"100111111",
  64271=>"111001010",
  64272=>"011101100",
  64273=>"001000111",
  64274=>"011110111",
  64275=>"011100000",
  64276=>"000100110",
  64277=>"100110001",
  64278=>"010000100",
  64279=>"011010010",
  64280=>"001110101",
  64281=>"111011101",
  64282=>"100100110",
  64283=>"010000010",
  64284=>"000101111",
  64285=>"010000001",
  64286=>"101000000",
  64287=>"001010111",
  64288=>"100110111",
  64289=>"001101100",
  64290=>"111000110",
  64291=>"011110000",
  64292=>"000100010",
  64293=>"111111110",
  64294=>"101111001",
  64295=>"011010010",
  64296=>"101010000",
  64297=>"110001110",
  64298=>"100111111",
  64299=>"110100011",
  64300=>"000101001",
  64301=>"101110011",
  64302=>"001110001",
  64303=>"000010110",
  64304=>"000010011",
  64305=>"110010011",
  64306=>"011100100",
  64307=>"000010100",
  64308=>"001110100",
  64309=>"001111101",
  64310=>"000100010",
  64311=>"110101000",
  64312=>"101001110",
  64313=>"011111011",
  64314=>"011100001",
  64315=>"101001000",
  64316=>"111111100",
  64317=>"101100000",
  64318=>"100001011",
  64319=>"001011111",
  64320=>"110111100",
  64321=>"100100111",
  64322=>"110101000",
  64323=>"100111001",
  64324=>"110100000",
  64325=>"100001001",
  64326=>"010000101",
  64327=>"001011110",
  64328=>"101011001",
  64329=>"010011010",
  64330=>"110010010",
  64331=>"100110110",
  64332=>"100101001",
  64333=>"000010111",
  64334=>"110010010",
  64335=>"100000111",
  64336=>"110111100",
  64337=>"010111011",
  64338=>"110001001",
  64339=>"011010010",
  64340=>"100101100",
  64341=>"000010111",
  64342=>"011001100",
  64343=>"010101111",
  64344=>"110000011",
  64345=>"010100101",
  64346=>"101000111",
  64347=>"001010001",
  64348=>"101011000",
  64349=>"111011000",
  64350=>"111010110",
  64351=>"000111110",
  64352=>"100000010",
  64353=>"100111111",
  64354=>"111011010",
  64355=>"100001110",
  64356=>"101001101",
  64357=>"111010101",
  64358=>"000100001",
  64359=>"101001111",
  64360=>"101111001",
  64361=>"001010011",
  64362=>"110010010",
  64363=>"111011001",
  64364=>"100110101",
  64365=>"111100110",
  64366=>"010100010",
  64367=>"010111111",
  64368=>"101100111",
  64369=>"001011100",
  64370=>"011011001",
  64371=>"100111001",
  64372=>"110110001",
  64373=>"100111111",
  64374=>"100110001",
  64375=>"111001111",
  64376=>"101101110",
  64377=>"111010001",
  64378=>"100011001",
  64379=>"001011001",
  64380=>"101011100",
  64381=>"111101111",
  64382=>"101101010",
  64383=>"011010110",
  64384=>"100001100",
  64385=>"000110001",
  64386=>"110110111",
  64387=>"010101000",
  64388=>"011011011",
  64389=>"110011100",
  64390=>"100001111",
  64391=>"000100010",
  64392=>"001001000",
  64393=>"110000010",
  64394=>"011011010",
  64395=>"111000000",
  64396=>"100000100",
  64397=>"110110110",
  64398=>"001101101",
  64399=>"101001100",
  64400=>"001000011",
  64401=>"110000001",
  64402=>"111010010",
  64403=>"011010110",
  64404=>"000101100",
  64405=>"000100100",
  64406=>"010011010",
  64407=>"010001111",
  64408=>"011010110",
  64409=>"001000111",
  64410=>"001100001",
  64411=>"111110000",
  64412=>"101100011",
  64413=>"001011110",
  64414=>"010010000",
  64415=>"011001000",
  64416=>"110001100",
  64417=>"101011000",
  64418=>"001011100",
  64419=>"101100110",
  64420=>"001100111",
  64421=>"010110101",
  64422=>"100110111",
  64423=>"111000010",
  64424=>"000101001",
  64425=>"000010010",
  64426=>"100101011",
  64427=>"111111010",
  64428=>"111101011",
  64429=>"110100101",
  64430=>"100111100",
  64431=>"000100000",
  64432=>"001010000",
  64433=>"010101100",
  64434=>"011110110",
  64435=>"001001011",
  64436=>"110111010",
  64437=>"000011101",
  64438=>"001001111",
  64439=>"111000101",
  64440=>"010111001",
  64441=>"101101010",
  64442=>"101100001",
  64443=>"100111001",
  64444=>"000100100",
  64445=>"000001001",
  64446=>"010011100",
  64447=>"101010001",
  64448=>"001010000",
  64449=>"111100011",
  64450=>"101010111",
  64451=>"001110110",
  64452=>"100010110",
  64453=>"010010011",
  64454=>"001011100",
  64455=>"000110000",
  64456=>"000101000",
  64457=>"001010100",
  64458=>"101001011",
  64459=>"111000001",
  64460=>"100001001",
  64461=>"100110011",
  64462=>"100111010",
  64463=>"110010111",
  64464=>"101010101",
  64465=>"111101010",
  64466=>"100111010",
  64467=>"011101000",
  64468=>"101010011",
  64469=>"010110011",
  64470=>"111111001",
  64471=>"000011000",
  64472=>"000110111",
  64473=>"010110011",
  64474=>"010010100",
  64475=>"100111001",
  64476=>"000100000",
  64477=>"001000110",
  64478=>"111111111",
  64479=>"110110111",
  64480=>"001110111",
  64481=>"010010010",
  64482=>"101100110",
  64483=>"110110011",
  64484=>"010000011",
  64485=>"111111101",
  64486=>"111010001",
  64487=>"111000101",
  64488=>"100111010",
  64489=>"111110011",
  64490=>"000011100",
  64491=>"010010000",
  64492=>"111011100",
  64493=>"100111011",
  64494=>"011001001",
  64495=>"111010011",
  64496=>"101101100",
  64497=>"110101110",
  64498=>"100111100",
  64499=>"001100101",
  64500=>"010011100",
  64501=>"011000100",
  64502=>"100101101",
  64503=>"010100100",
  64504=>"010010001",
  64505=>"011100100",
  64506=>"011110011",
  64507=>"111101011",
  64508=>"001011000",
  64509=>"010100011",
  64510=>"101010111",
  64511=>"010010110",
  64512=>"111100011",
  64513=>"010010110",
  64514=>"001111110",
  64515=>"011111111",
  64516=>"101011010",
  64517=>"111111101",
  64518=>"001011000",
  64519=>"111110010",
  64520=>"111100011",
  64521=>"000010110",
  64522=>"100001110",
  64523=>"001011010",
  64524=>"000111000",
  64525=>"010110010",
  64526=>"011111101",
  64527=>"001110110",
  64528=>"110000001",
  64529=>"010110100",
  64530=>"010001000",
  64531=>"111010010",
  64532=>"101001110",
  64533=>"100110000",
  64534=>"101111001",
  64535=>"111001000",
  64536=>"110110001",
  64537=>"000101101",
  64538=>"011100100",
  64539=>"111101000",
  64540=>"101011100",
  64541=>"110001000",
  64542=>"110100101",
  64543=>"000010100",
  64544=>"111110001",
  64545=>"101111011",
  64546=>"100010101",
  64547=>"010010110",
  64548=>"010010110",
  64549=>"011000011",
  64550=>"111001011",
  64551=>"010000001",
  64552=>"100101110",
  64553=>"000001010",
  64554=>"010110011",
  64555=>"000100011",
  64556=>"011001000",
  64557=>"011110111",
  64558=>"011100100",
  64559=>"000101110",
  64560=>"000100000",
  64561=>"001001101",
  64562=>"000010001",
  64563=>"010000011",
  64564=>"011101000",
  64565=>"011011010",
  64566=>"010101110",
  64567=>"000110101",
  64568=>"110111000",
  64569=>"101101101",
  64570=>"101001001",
  64571=>"111111111",
  64572=>"011101100",
  64573=>"101111101",
  64574=>"101001000",
  64575=>"010100000",
  64576=>"011000101",
  64577=>"001010000",
  64578=>"110111011",
  64579=>"101101111",
  64580=>"011101111",
  64581=>"010111110",
  64582=>"100110011",
  64583=>"000110111",
  64584=>"100000000",
  64585=>"001110101",
  64586=>"011101000",
  64587=>"011000111",
  64588=>"101001010",
  64589=>"010010110",
  64590=>"010100010",
  64591=>"110100100",
  64592=>"000110010",
  64593=>"011000111",
  64594=>"100010011",
  64595=>"000111100",
  64596=>"000110011",
  64597=>"000001000",
  64598=>"010111100",
  64599=>"001001001",
  64600=>"101010100",
  64601=>"100000101",
  64602=>"001011000",
  64603=>"111101110",
  64604=>"101101100",
  64605=>"111001011",
  64606=>"101010111",
  64607=>"000101011",
  64608=>"100001100",
  64609=>"100100111",
  64610=>"001101110",
  64611=>"011000010",
  64612=>"010001100",
  64613=>"101101001",
  64614=>"001001000",
  64615=>"000111010",
  64616=>"110001111",
  64617=>"001001010",
  64618=>"111100110",
  64619=>"110111011",
  64620=>"101011001",
  64621=>"100010110",
  64622=>"111100110",
  64623=>"011101111",
  64624=>"010010110",
  64625=>"000111010",
  64626=>"100000001",
  64627=>"010011101",
  64628=>"110101111",
  64629=>"000010011",
  64630=>"100011001",
  64631=>"011011001",
  64632=>"010101010",
  64633=>"000001001",
  64634=>"111001101",
  64635=>"100000110",
  64636=>"011100000",
  64637=>"110100000",
  64638=>"101011111",
  64639=>"011101000",
  64640=>"100010111",
  64641=>"111010111",
  64642=>"101111101",
  64643=>"010010110",
  64644=>"001000000",
  64645=>"110101010",
  64646=>"110010101",
  64647=>"001100111",
  64648=>"101111111",
  64649=>"001010100",
  64650=>"101111001",
  64651=>"000100001",
  64652=>"100111111",
  64653=>"010000100",
  64654=>"111111001",
  64655=>"010000001",
  64656=>"111110001",
  64657=>"101101000",
  64658=>"100111110",
  64659=>"111010110",
  64660=>"011101101",
  64661=>"001010101",
  64662=>"000011111",
  64663=>"101001100",
  64664=>"010000110",
  64665=>"001111010",
  64666=>"100101111",
  64667=>"000101100",
  64668=>"001100001",
  64669=>"100011000",
  64670=>"110100101",
  64671=>"101101010",
  64672=>"101011101",
  64673=>"111110111",
  64674=>"001001110",
  64675=>"100010100",
  64676=>"110100001",
  64677=>"100111111",
  64678=>"001100000",
  64679=>"000000110",
  64680=>"101011110",
  64681=>"000010010",
  64682=>"011100011",
  64683=>"000100010",
  64684=>"001110110",
  64685=>"010100000",
  64686=>"000000000",
  64687=>"000010001",
  64688=>"111001001",
  64689=>"001100100",
  64690=>"011111111",
  64691=>"001011111",
  64692=>"001011001",
  64693=>"101101101",
  64694=>"001101111",
  64695=>"011101110",
  64696=>"001010011",
  64697=>"111000111",
  64698=>"100101000",
  64699=>"001111100",
  64700=>"001111100",
  64701=>"100010111",
  64702=>"010100000",
  64703=>"100001010",
  64704=>"000000010",
  64705=>"101111100",
  64706=>"011111011",
  64707=>"001010110",
  64708=>"000001000",
  64709=>"011000001",
  64710=>"101000111",
  64711=>"001010101",
  64712=>"111011011",
  64713=>"110100110",
  64714=>"111110011",
  64715=>"011110100",
  64716=>"010111010",
  64717=>"001101010",
  64718=>"111000100",
  64719=>"010100100",
  64720=>"001000010",
  64721=>"100110011",
  64722=>"001111111",
  64723=>"000010101",
  64724=>"100001010",
  64725=>"100001011",
  64726=>"110111111",
  64727=>"011110000",
  64728=>"010111100",
  64729=>"001000110",
  64730=>"110010110",
  64731=>"100000111",
  64732=>"011011000",
  64733=>"000001111",
  64734=>"001001111",
  64735=>"001011000",
  64736=>"010011001",
  64737=>"000100101",
  64738=>"010000000",
  64739=>"101001110",
  64740=>"110010110",
  64741=>"001000100",
  64742=>"000001010",
  64743=>"000100000",
  64744=>"111000100",
  64745=>"001001111",
  64746=>"101110010",
  64747=>"110100111",
  64748=>"110010001",
  64749=>"111101001",
  64750=>"000001101",
  64751=>"010010100",
  64752=>"100100011",
  64753=>"001101111",
  64754=>"101011100",
  64755=>"100111011",
  64756=>"011100111",
  64757=>"010000011",
  64758=>"100000000",
  64759=>"001001110",
  64760=>"101011100",
  64761=>"101100000",
  64762=>"111001000",
  64763=>"001000010",
  64764=>"100101001",
  64765=>"100000000",
  64766=>"101001001",
  64767=>"000000111",
  64768=>"000001111",
  64769=>"010110001",
  64770=>"100101111",
  64771=>"011100011",
  64772=>"001110000",
  64773=>"000001010",
  64774=>"110001011",
  64775=>"100001100",
  64776=>"101111011",
  64777=>"101011001",
  64778=>"111111000",
  64779=>"101111100",
  64780=>"001001001",
  64781=>"000100100",
  64782=>"110100001",
  64783=>"110101111",
  64784=>"111110010",
  64785=>"101100000",
  64786=>"111001101",
  64787=>"000101111",
  64788=>"100011011",
  64789=>"010001010",
  64790=>"101001100",
  64791=>"100100110",
  64792=>"010000000",
  64793=>"000101010",
  64794=>"010010001",
  64795=>"110101000",
  64796=>"011101101",
  64797=>"001111111",
  64798=>"000110010",
  64799=>"111100001",
  64800=>"111100111",
  64801=>"010110010",
  64802=>"011011110",
  64803=>"010110111",
  64804=>"100011100",
  64805=>"000111011",
  64806=>"101011011",
  64807=>"110000110",
  64808=>"000110100",
  64809=>"001110111",
  64810=>"110011100",
  64811=>"011000100",
  64812=>"110101010",
  64813=>"111001111",
  64814=>"001000011",
  64815=>"101111110",
  64816=>"101010101",
  64817=>"110101011",
  64818=>"100111000",
  64819=>"110010010",
  64820=>"010100010",
  64821=>"101101010",
  64822=>"001100000",
  64823=>"101110000",
  64824=>"011111111",
  64825=>"011000000",
  64826=>"101011011",
  64827=>"011101010",
  64828=>"001010000",
  64829=>"111110011",
  64830=>"110000000",
  64831=>"101011100",
  64832=>"011101110",
  64833=>"101110001",
  64834=>"101001000",
  64835=>"111100111",
  64836=>"011101001",
  64837=>"000100100",
  64838=>"001111011",
  64839=>"111010101",
  64840=>"111111110",
  64841=>"110001011",
  64842=>"111000010",
  64843=>"010010100",
  64844=>"111111101",
  64845=>"101111010",
  64846=>"011001100",
  64847=>"101111100",
  64848=>"100000110",
  64849=>"011000001",
  64850=>"010010000",
  64851=>"101111001",
  64852=>"011111101",
  64853=>"001000111",
  64854=>"001111011",
  64855=>"001001001",
  64856=>"011100101",
  64857=>"111101011",
  64858=>"001001000",
  64859=>"110110111",
  64860=>"111111000",
  64861=>"011100110",
  64862=>"010110001",
  64863=>"101001011",
  64864=>"010010011",
  64865=>"010001111",
  64866=>"001010110",
  64867=>"101100010",
  64868=>"101100111",
  64869=>"100010000",
  64870=>"011110001",
  64871=>"101011100",
  64872=>"001001001",
  64873=>"100010111",
  64874=>"011100111",
  64875=>"111111011",
  64876=>"010001001",
  64877=>"110001100",
  64878=>"000101000",
  64879=>"110111000",
  64880=>"101111010",
  64881=>"010000000",
  64882=>"000101001",
  64883=>"101100100",
  64884=>"000000010",
  64885=>"100111000",
  64886=>"011110100",
  64887=>"111001010",
  64888=>"000010010",
  64889=>"000000000",
  64890=>"011110011",
  64891=>"101011011",
  64892=>"100100111",
  64893=>"111111100",
  64894=>"000100111",
  64895=>"101111011",
  64896=>"100011011",
  64897=>"000101100",
  64898=>"001101000",
  64899=>"111111000",
  64900=>"010110101",
  64901=>"101101011",
  64902=>"000100111",
  64903=>"111110100",
  64904=>"000010110",
  64905=>"010010000",
  64906=>"000011110",
  64907=>"010001101",
  64908=>"110011111",
  64909=>"100010001",
  64910=>"010100010",
  64911=>"110010000",
  64912=>"011110010",
  64913=>"100110000",
  64914=>"011001101",
  64915=>"111100101",
  64916=>"001110111",
  64917=>"010110000",
  64918=>"001101001",
  64919=>"100101010",
  64920=>"111010100",
  64921=>"011011011",
  64922=>"110100101",
  64923=>"000001100",
  64924=>"001110100",
  64925=>"011011000",
  64926=>"000101101",
  64927=>"100001010",
  64928=>"101000011",
  64929=>"110000111",
  64930=>"010001110",
  64931=>"001100011",
  64932=>"110110111",
  64933=>"110100111",
  64934=>"000111010",
  64935=>"100011100",
  64936=>"000110000",
  64937=>"011100101",
  64938=>"101111011",
  64939=>"111011001",
  64940=>"111101110",
  64941=>"110110010",
  64942=>"001001100",
  64943=>"100010010",
  64944=>"111100101",
  64945=>"111100100",
  64946=>"001101011",
  64947=>"010100011",
  64948=>"111001010",
  64949=>"001111010",
  64950=>"000111010",
  64951=>"011100110",
  64952=>"110111000",
  64953=>"000100001",
  64954=>"001110111",
  64955=>"000111110",
  64956=>"110111110",
  64957=>"000100000",
  64958=>"100101010",
  64959=>"110011011",
  64960=>"000010011",
  64961=>"110110010",
  64962=>"010111111",
  64963=>"100000101",
  64964=>"101101110",
  64965=>"100001001",
  64966=>"110001111",
  64967=>"100001010",
  64968=>"011110110",
  64969=>"101010111",
  64970=>"101001110",
  64971=>"000100100",
  64972=>"100010110",
  64973=>"100101001",
  64974=>"111100110",
  64975=>"100000001",
  64976=>"100101011",
  64977=>"010011111",
  64978=>"011000110",
  64979=>"111001101",
  64980=>"110110010",
  64981=>"011010101",
  64982=>"110000111",
  64983=>"001010110",
  64984=>"111111110",
  64985=>"111100101",
  64986=>"000110110",
  64987=>"110111101",
  64988=>"000101110",
  64989=>"111011110",
  64990=>"000100111",
  64991=>"111000000",
  64992=>"010000110",
  64993=>"111110010",
  64994=>"000011110",
  64995=>"100011111",
  64996=>"110110101",
  64997=>"100110110",
  64998=>"110100110",
  64999=>"000001010",
  65000=>"011000100",
  65001=>"101111010",
  65002=>"101110000",
  65003=>"110011000",
  65004=>"000010110",
  65005=>"011010111",
  65006=>"001100010",
  65007=>"011000011",
  65008=>"100100001",
  65009=>"110011011",
  65010=>"110010111",
  65011=>"100001111",
  65012=>"000010100",
  65013=>"010000101",
  65014=>"001010010",
  65015=>"010110001",
  65016=>"101100100",
  65017=>"101101000",
  65018=>"110001000",
  65019=>"100001110",
  65020=>"100001011",
  65021=>"100000001",
  65022=>"100000110",
  65023=>"110000100",
  65024=>"110111111",
  65025=>"001100111",
  65026=>"100111100",
  65027=>"001111100",
  65028=>"000111001",
  65029=>"111111111",
  65030=>"001010000",
  65031=>"101011100",
  65032=>"111101100",
  65033=>"000100101",
  65034=>"100101011",
  65035=>"000011011",
  65036=>"111000101",
  65037=>"001010111",
  65038=>"000001011",
  65039=>"110100110",
  65040=>"110110111",
  65041=>"001101011",
  65042=>"011110011",
  65043=>"001100111",
  65044=>"011111001",
  65045=>"010010110",
  65046=>"011111011",
  65047=>"011010111",
  65048=>"000010011",
  65049=>"110110010",
  65050=>"000010111",
  65051=>"011101001",
  65052=>"000000110",
  65053=>"100010101",
  65054=>"101101001",
  65055=>"001111011",
  65056=>"100001010",
  65057=>"101111101",
  65058=>"011110111",
  65059=>"110000110",
  65060=>"000110010",
  65061=>"101000010",
  65062=>"101011100",
  65063=>"111000011",
  65064=>"100110001",
  65065=>"110100010",
  65066=>"110010011",
  65067=>"001011111",
  65068=>"001100011",
  65069=>"000100001",
  65070=>"000001101",
  65071=>"010101011",
  65072=>"010101011",
  65073=>"010100101",
  65074=>"010101100",
  65075=>"111111011",
  65076=>"001000001",
  65077=>"010001000",
  65078=>"010010000",
  65079=>"111110111",
  65080=>"100111110",
  65081=>"100001001",
  65082=>"110101101",
  65083=>"111111100",
  65084=>"100111101",
  65085=>"110001100",
  65086=>"010010101",
  65087=>"000110010",
  65088=>"110001101",
  65089=>"011101011",
  65090=>"000000000",
  65091=>"110101001",
  65092=>"110100111",
  65093=>"001110111",
  65094=>"000011111",
  65095=>"000100110",
  65096=>"100110011",
  65097=>"101001011",
  65098=>"010011010",
  65099=>"101100111",
  65100=>"000110011",
  65101=>"101001000",
  65102=>"011001101",
  65103=>"111010111",
  65104=>"001011000",
  65105=>"101001000",
  65106=>"000011001",
  65107=>"011110000",
  65108=>"110110111",
  65109=>"110101110",
  65110=>"101000000",
  65111=>"011101000",
  65112=>"110000111",
  65113=>"010001010",
  65114=>"101001000",
  65115=>"110011110",
  65116=>"100011000",
  65117=>"000110111",
  65118=>"101101101",
  65119=>"111010001",
  65120=>"011000001",
  65121=>"101111111",
  65122=>"100100000",
  65123=>"110110110",
  65124=>"100110100",
  65125=>"111001110",
  65126=>"100101000",
  65127=>"001011111",
  65128=>"000010000",
  65129=>"010000001",
  65130=>"001011001",
  65131=>"001101111",
  65132=>"101000000",
  65133=>"011110100",
  65134=>"101101000",
  65135=>"000110001",
  65136=>"011011110",
  65137=>"111100000",
  65138=>"011001010",
  65139=>"100000010",
  65140=>"111001101",
  65141=>"010100000",
  65142=>"011001001",
  65143=>"001000001",
  65144=>"111100001",
  65145=>"001001010",
  65146=>"001101110",
  65147=>"001100011",
  65148=>"011010101",
  65149=>"101101000",
  65150=>"000000000",
  65151=>"110000000",
  65152=>"110000000",
  65153=>"000011000",
  65154=>"111110110",
  65155=>"110000100",
  65156=>"011010110",
  65157=>"011010100",
  65158=>"111001011",
  65159=>"001010100",
  65160=>"011011110",
  65161=>"011010010",
  65162=>"000011110",
  65163=>"001100110",
  65164=>"000101111",
  65165=>"100000010",
  65166=>"001110000",
  65167=>"100111000",
  65168=>"100101101",
  65169=>"111101101",
  65170=>"110111110",
  65171=>"011011000",
  65172=>"101110000",
  65173=>"010111001",
  65174=>"010100011",
  65175=>"001011111",
  65176=>"111101101",
  65177=>"101111101",
  65178=>"010100100",
  65179=>"100011010",
  65180=>"010111100",
  65181=>"000000110",
  65182=>"001110111",
  65183=>"100100001",
  65184=>"111001101",
  65185=>"111111111",
  65186=>"001001100",
  65187=>"100001000",
  65188=>"101110010",
  65189=>"011111111",
  65190=>"111100111",
  65191=>"000111000",
  65192=>"010111010",
  65193=>"110001111",
  65194=>"111000011",
  65195=>"110001011",
  65196=>"001110011",
  65197=>"111110010",
  65198=>"000000100",
  65199=>"100001000",
  65200=>"101100011",
  65201=>"101110110",
  65202=>"000001101",
  65203=>"000110010",
  65204=>"100110010",
  65205=>"111110110",
  65206=>"111101101",
  65207=>"100101110",
  65208=>"001010000",
  65209=>"000110000",
  65210=>"010111101",
  65211=>"001001111",
  65212=>"010000110",
  65213=>"001101100",
  65214=>"110110001",
  65215=>"010100100",
  65216=>"000111011",
  65217=>"110100010",
  65218=>"010000000",
  65219=>"110000010",
  65220=>"001000110",
  65221=>"001111100",
  65222=>"110000100",
  65223=>"000101101",
  65224=>"111111101",
  65225=>"101101001",
  65226=>"000111001",
  65227=>"110000010",
  65228=>"000100100",
  65229=>"000010110",
  65230=>"010110101",
  65231=>"001000100",
  65232=>"001100110",
  65233=>"001001110",
  65234=>"111001010",
  65235=>"011001010",
  65236=>"011011001",
  65237=>"001110101",
  65238=>"100000100",
  65239=>"000011001",
  65240=>"010010100",
  65241=>"000111001",
  65242=>"010111101",
  65243=>"110101011",
  65244=>"000010010",
  65245=>"010001101",
  65246=>"000010011",
  65247=>"111110100",
  65248=>"111001000",
  65249=>"110110110",
  65250=>"001101110",
  65251=>"000000000",
  65252=>"011111000",
  65253=>"000000100",
  65254=>"000101010",
  65255=>"101000101",
  65256=>"001110000",
  65257=>"111011001",
  65258=>"000011100",
  65259=>"010101110",
  65260=>"010000101",
  65261=>"010010110",
  65262=>"011111011",
  65263=>"101111011",
  65264=>"000110011",
  65265=>"011001110",
  65266=>"010100100",
  65267=>"001001000",
  65268=>"000011011",
  65269=>"101001001",
  65270=>"111110110",
  65271=>"001111110",
  65272=>"100110001",
  65273=>"100000001",
  65274=>"001110001",
  65275=>"111011001",
  65276=>"101110100",
  65277=>"111001010",
  65278=>"000010010",
  65279=>"101111001",
  65280=>"100011110",
  65281=>"001101011",
  65282=>"011111111",
  65283=>"010110100",
  65284=>"110100100",
  65285=>"101010011",
  65286=>"001110100",
  65287=>"000000101",
  65288=>"110011011",
  65289=>"000001010",
  65290=>"111110101",
  65291=>"011100101",
  65292=>"001111111",
  65293=>"011111011",
  65294=>"101000000",
  65295=>"111110111",
  65296=>"001011100",
  65297=>"011101011",
  65298=>"000100110",
  65299=>"010110000",
  65300=>"101011100",
  65301=>"011001001",
  65302=>"111100111",
  65303=>"011011111",
  65304=>"111101001",
  65305=>"111100111",
  65306=>"000100010",
  65307=>"011100000",
  65308=>"010110000",
  65309=>"000100001",
  65310=>"001010000",
  65311=>"000111001",
  65312=>"110111110",
  65313=>"010101101",
  65314=>"010010111",
  65315=>"100000100",
  65316=>"011011011",
  65317=>"000101101",
  65318=>"010111101",
  65319=>"111011011",
  65320=>"000101011",
  65321=>"011111000",
  65322=>"101000001",
  65323=>"000100001",
  65324=>"010111001",
  65325=>"110000010",
  65326=>"101000101",
  65327=>"011111010",
  65328=>"000001110",
  65329=>"101011010",
  65330=>"000111111",
  65331=>"011001110",
  65332=>"101101101",
  65333=>"000001101",
  65334=>"110000001",
  65335=>"100000110",
  65336=>"101010001",
  65337=>"001111101",
  65338=>"000101101",
  65339=>"001010111",
  65340=>"111101111",
  65341=>"001010111",
  65342=>"001000111",
  65343=>"100000000",
  65344=>"010001011",
  65345=>"000011110",
  65346=>"011101010",
  65347=>"100000111",
  65348=>"010101100",
  65349=>"100101110",
  65350=>"001111000",
  65351=>"011110000",
  65352=>"111101011",
  65353=>"111101111",
  65354=>"110101101",
  65355=>"101010100",
  65356=>"111011011",
  65357=>"000110000",
  65358=>"010110101",
  65359=>"010100111",
  65360=>"101101011",
  65361=>"001001101",
  65362=>"111001010",
  65363=>"010010110",
  65364=>"010100000",
  65365=>"010110000",
  65366=>"110011011",
  65367=>"000000110",
  65368=>"100000000",
  65369=>"101100000",
  65370=>"110101000",
  65371=>"100110101",
  65372=>"011100101",
  65373=>"001000111",
  65374=>"011100100",
  65375=>"010111010",
  65376=>"000100111",
  65377=>"000101101",
  65378=>"111111111",
  65379=>"100100100",
  65380=>"011010111",
  65381=>"011111111",
  65382=>"110000101",
  65383=>"000100100",
  65384=>"100000000",
  65385=>"101010110",
  65386=>"101111111",
  65387=>"100001111",
  65388=>"011111011",
  65389=>"010110001",
  65390=>"010011111",
  65391=>"011111110",
  65392=>"010100001",
  65393=>"001011101",
  65394=>"001010010",
  65395=>"010101110",
  65396=>"010001011",
  65397=>"101000010",
  65398=>"110001111",
  65399=>"000010011",
  65400=>"110010101",
  65401=>"001011000",
  65402=>"110101000",
  65403=>"110011101",
  65404=>"101111011",
  65405=>"001001011",
  65406=>"010001110",
  65407=>"100001110",
  65408=>"000110000",
  65409=>"010110101",
  65410=>"001010111",
  65411=>"100011001",
  65412=>"111111000",
  65413=>"000010010",
  65414=>"001100001",
  65415=>"010101101",
  65416=>"001110101",
  65417=>"001001000",
  65418=>"110010010",
  65419=>"000111111",
  65420=>"110110001",
  65421=>"010101000",
  65422=>"011111100",
  65423=>"111111110",
  65424=>"001011001",
  65425=>"101011101",
  65426=>"000101010",
  65427=>"011010011",
  65428=>"110111110",
  65429=>"011101001",
  65430=>"010100001",
  65431=>"101010110",
  65432=>"000011111",
  65433=>"000100011",
  65434=>"000010100",
  65435=>"011100101",
  65436=>"000011010",
  65437=>"001100111",
  65438=>"000001011",
  65439=>"011001001",
  65440=>"010010011",
  65441=>"010000001",
  65442=>"001010111",
  65443=>"101001111",
  65444=>"010110010",
  65445=>"001110111",
  65446=>"100011001",
  65447=>"111110010",
  65448=>"010111011",
  65449=>"010100010",
  65450=>"010001101",
  65451=>"010010000",
  65452=>"110111110",
  65453=>"011001000",
  65454=>"111110000",
  65455=>"011000101",
  65456=>"010000010",
  65457=>"100101100",
  65458=>"110101011",
  65459=>"001010111",
  65460=>"100000101",
  65461=>"100010111",
  65462=>"010111000",
  65463=>"110110100",
  65464=>"000001101",
  65465=>"100011000",
  65466=>"111011001",
  65467=>"001111000",
  65468=>"011010011",
  65469=>"000100001",
  65470=>"010111011",
  65471=>"011101110",
  65472=>"000000010",
  65473=>"111010100",
  65474=>"001101000",
  65475=>"011100111",
  65476=>"100011100",
  65477=>"010001011",
  65478=>"111010101",
  65479=>"011010111",
  65480=>"011000101",
  65481=>"100000101",
  65482=>"001100111",
  65483=>"001011101",
  65484=>"000001101",
  65485=>"101000100",
  65486=>"100011011",
  65487=>"010101101",
  65488=>"010000010",
  65489=>"001111000",
  65490=>"100011101",
  65491=>"010001100",
  65492=>"101010000",
  65493=>"011000100",
  65494=>"111101111",
  65495=>"100010111",
  65496=>"111110101",
  65497=>"001000011",
  65498=>"110001000",
  65499=>"100110000",
  65500=>"001101011",
  65501=>"101110001",
  65502=>"110010100",
  65503=>"001001110",
  65504=>"111101101",
  65505=>"100110101",
  65506=>"011010000",
  65507=>"100101100",
  65508=>"111111100",
  65509=>"111011111",
  65510=>"001010010",
  65511=>"000101011",
  65512=>"111000001",
  65513=>"101001011",
  65514=>"010001100",
  65515=>"000000111",
  65516=>"010101000",
  65517=>"111011100",
  65518=>"110001000",
  65519=>"111001100",
  65520=>"100101011",
  65521=>"010010111",
  65522=>"010101111",
  65523=>"000011110",
  65524=>"111111110",
  65525=>"011110101",
  65526=>"000010000",
  65527=>"010000011",
  65528=>"111110011",
  65529=>"110111101",
  65530=>"010111111",
  65531=>"001001010",
  65532=>"001101110",
  65533=>"010101010",
  65534=>"110001001",
  65535=>"001111100");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;