LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L7_8_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(7) - 1 DOWNTO 0));
END L7_8_WROM;

ARCHITECTURE RTL OF L7_8_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"011111111",
  1=>"110110110",
  2=>"111001111",
  3=>"000000000",
  4=>"111111011",
  5=>"000000001",
  6=>"000110110",
  7=>"111111111",
  8=>"111111100",
  9=>"111111100",
  10=>"111111111",
  11=>"000000000",
  12=>"000110110",
  13=>"000001010",
  14=>"100111101",
  15=>"000010000",
  16=>"111000000",
  17=>"111101001",
  18=>"000011000",
  19=>"111111111",
  20=>"101000101",
  21=>"000000000",
  22=>"000000000",
  23=>"000001001",
  24=>"101111111",
  25=>"000001111",
  26=>"001000000",
  27=>"001001000",
  28=>"111100000",
  29=>"011111111",
  30=>"000000100",
  31=>"111111101",
  32=>"100000100",
  33=>"011111111",
  34=>"000000000",
  35=>"010111100",
  36=>"000100111",
  37=>"000000000",
  38=>"000000101",
  39=>"111111111",
  40=>"000001011",
  41=>"111000000",
  42=>"000000000",
  43=>"111111111",
  44=>"111000000",
  45=>"111111011",
  46=>"000010010",
  47=>"000000000",
  48=>"000000100",
  49=>"000000000",
  50=>"010111111",
  51=>"000000000",
  52=>"000111011",
  53=>"111111011",
  54=>"000000000",
  55=>"010000111",
  56=>"111111111",
  57=>"111111110",
  58=>"000000011",
  59=>"011011011",
  60=>"111100101",
  61=>"111111100",
  62=>"000100111",
  63=>"000000100",
  64=>"100100111",
  65=>"000000000",
  66=>"011111111",
  67=>"000110100",
  68=>"110010111",
  69=>"010111110",
  70=>"000010010",
  71=>"111110010",
  72=>"100111111",
  73=>"000000111",
  74=>"111111110",
  75=>"111111110",
  76=>"000000111",
  77=>"111101000",
  78=>"111000100",
  79=>"111111111",
  80=>"111111110",
  81=>"111111110",
  82=>"001000001",
  83=>"001111010",
  84=>"100000000",
  85=>"111111111",
  86=>"000000101",
  87=>"000000000",
  88=>"000000000",
  89=>"101001111",
  90=>"111111111",
  91=>"111111100",
  92=>"101101111",
  93=>"100000111",
  94=>"101111111",
  95=>"110000000",
  96=>"000111011",
  97=>"101000111",
  98=>"000000000",
  99=>"100000000",
  100=>"111011000",
  101=>"001000000",
  102=>"111000000",
  103=>"111110110",
  104=>"110111111",
  105=>"111001000",
  106=>"111110000",
  107=>"000000111",
  108=>"001011111",
  109=>"111111111",
  110=>"100110110",
  111=>"111000111",
  112=>"111111111",
  113=>"111111111",
  114=>"000000000",
  115=>"110000000",
  116=>"010110111",
  117=>"011111000",
  118=>"000000100",
  119=>"000010111",
  120=>"000100000",
  121=>"100111111",
  122=>"011001001",
  123=>"000001111",
  124=>"111111111",
  125=>"000000111",
  126=>"000000000",
  127=>"000000000",
  128=>"000000000",
  129=>"010010011",
  130=>"000000000",
  131=>"000000001",
  132=>"110000000",
  133=>"000001001",
  134=>"110110111",
  135=>"001011000",
  136=>"000000000",
  137=>"000000000",
  138=>"101110000",
  139=>"000111000",
  140=>"111111011",
  141=>"001000000",
  142=>"111111111",
  143=>"000000000",
  144=>"000000100",
  145=>"000000100",
  146=>"100000100",
  147=>"001001010",
  148=>"100111111",
  149=>"110111000",
  150=>"111000010",
  151=>"111000111",
  152=>"000000000",
  153=>"001001011",
  154=>"000000001",
  155=>"000000000",
  156=>"010000111",
  157=>"000000111",
  158=>"111111100",
  159=>"010010111",
  160=>"111111011",
  161=>"011011011",
  162=>"111000000",
  163=>"000000000",
  164=>"111111000",
  165=>"101001111",
  166=>"111000000",
  167=>"000111111",
  168=>"111000000",
  169=>"100011011",
  170=>"000100111",
  171=>"111111011",
  172=>"111111111",
  173=>"000110110",
  174=>"000000000",
  175=>"000010000",
  176=>"111111011",
  177=>"000100000",
  178=>"111111010",
  179=>"111000100",
  180=>"000000011",
  181=>"011000110",
  182=>"000000111",
  183=>"000000000",
  184=>"111000111",
  185=>"000000000",
  186=>"001000101",
  187=>"111111111",
  188=>"000000111",
  189=>"111111000",
  190=>"000000111",
  191=>"111111111",
  192=>"000111111",
  193=>"111111111",
  194=>"111111111",
  195=>"000000000",
  196=>"011000000",
  197=>"000001000",
  198=>"110111111",
  199=>"000000000",
  200=>"000011111",
  201=>"010011001",
  202=>"111010111",
  203=>"000000000",
  204=>"100001011",
  205=>"110111001",
  206=>"010110000",
  207=>"011011011",
  208=>"111111000",
  209=>"111010111",
  210=>"111100100",
  211=>"000111111",
  212=>"000000110",
  213=>"000000111",
  214=>"111000000",
  215=>"101110000",
  216=>"000000000",
  217=>"111111111",
  218=>"001000000",
  219=>"000000000",
  220=>"111111111",
  221=>"110110111",
  222=>"111010000",
  223=>"000000001",
  224=>"001001111",
  225=>"100000000",
  226=>"111111111",
  227=>"111001001",
  228=>"000000001",
  229=>"110110010",
  230=>"000011011",
  231=>"111111111",
  232=>"111110000",
  233=>"111111011",
  234=>"011011001",
  235=>"011110110",
  236=>"100110000",
  237=>"000000111",
  238=>"111110111",
  239=>"101111101",
  240=>"100011011",
  241=>"111111000",
  242=>"000001011",
  243=>"011000000",
  244=>"000000111",
  245=>"111001011",
  246=>"111000000",
  247=>"111111111",
  248=>"010111110",
  249=>"000000000",
  250=>"101001111",
  251=>"111000111",
  252=>"000011011",
  253=>"001100001",
  254=>"111111111",
  255=>"000111111",
  256=>"011111111",
  257=>"010110100",
  258=>"111111011",
  259=>"111000111",
  260=>"000000000",
  261=>"010011001",
  262=>"111110000",
  263=>"101111110",
  264=>"111000000",
  265=>"001000000",
  266=>"010111110",
  267=>"100000000",
  268=>"000000011",
  269=>"001011111",
  270=>"101001001",
  271=>"000000010",
  272=>"111111111",
  273=>"000000000",
  274=>"101001001",
  275=>"110110111",
  276=>"000000111",
  277=>"001010111",
  278=>"001001001",
  279=>"000000000",
  280=>"001111100",
  281=>"111111100",
  282=>"001000101",
  283=>"100000000",
  284=>"111111110",
  285=>"111111000",
  286=>"000000010",
  287=>"111011000",
  288=>"000011001",
  289=>"100100000",
  290=>"110111111",
  291=>"000011001",
  292=>"000001000",
  293=>"000111111",
  294=>"110100100",
  295=>"111111111",
  296=>"000100110",
  297=>"000000110",
  298=>"011000010",
  299=>"000000000",
  300=>"011111001",
  301=>"001111111",
  302=>"000000000",
  303=>"000000000",
  304=>"011111111",
  305=>"000000000",
  306=>"001001111",
  307=>"011111111",
  308=>"100110011",
  309=>"111111101",
  310=>"111111111",
  311=>"001011011",
  312=>"000111000",
  313=>"111000101",
  314=>"111100111",
  315=>"111111111",
  316=>"000100110",
  317=>"000011000",
  318=>"000000100",
  319=>"000101101",
  320=>"110111000",
  321=>"111110010",
  322=>"000000111",
  323=>"001111111",
  324=>"000001000",
  325=>"111111111",
  326=>"000000110",
  327=>"100100111",
  328=>"111000111",
  329=>"100000010",
  330=>"000000100",
  331=>"101000000",
  332=>"000000000",
  333=>"000000000",
  334=>"000001111",
  335=>"111011011",
  336=>"110111111",
  337=>"000000101",
  338=>"001111111",
  339=>"111110110",
  340=>"100000000",
  341=>"010011011",
  342=>"000000001",
  343=>"100000001",
  344=>"000000000",
  345=>"111000000",
  346=>"000000100",
  347=>"001101111",
  348=>"000000000",
  349=>"111111111",
  350=>"000000000",
  351=>"111111111",
  352=>"111011000",
  353=>"011000111",
  354=>"110000011",
  355=>"000000000",
  356=>"000110111",
  357=>"111100110",
  358=>"111111000",
  359=>"000000000",
  360=>"000000110",
  361=>"001000010",
  362=>"000110000",
  363=>"111000110",
  364=>"000000000",
  365=>"001000111",
  366=>"110111110",
  367=>"101000000",
  368=>"001001100",
  369=>"000000000",
  370=>"110000000",
  371=>"111011011",
  372=>"110110111",
  373=>"000000001",
  374=>"100000111",
  375=>"011011001",
  376=>"000000110",
  377=>"111111011",
  378=>"111100111",
  379=>"001010000",
  380=>"111000000",
  381=>"001000111",
  382=>"110100100",
  383=>"010110000",
  384=>"111100111",
  385=>"000000000",
  386=>"111111111",
  387=>"001001111",
  388=>"111111111",
  389=>"001011011",
  390=>"000000000",
  391=>"100011011",
  392=>"101011000",
  393=>"001111111",
  394=>"000000000",
  395=>"010110000",
  396=>"000100111",
  397=>"001001001",
  398=>"111111010",
  399=>"000000000",
  400=>"100000000",
  401=>"000111111",
  402=>"111111001",
  403=>"001000001",
  404=>"111100100",
  405=>"000000000",
  406=>"000000000",
  407=>"111011000",
  408=>"000011000",
  409=>"011011000",
  410=>"011101111",
  411=>"100000001",
  412=>"110000110",
  413=>"000010000",
  414=>"111111111",
  415=>"000111000",
  416=>"000111111",
  417=>"110001000",
  418=>"011000001",
  419=>"111000000",
  420=>"001011111",
  421=>"111111110",
  422=>"000000000",
  423=>"001011000",
  424=>"000010000",
  425=>"101000000",
  426=>"000000000",
  427=>"111000000",
  428=>"000000000",
  429=>"100000110",
  430=>"110100111",
  431=>"101000000",
  432=>"111011000",
  433=>"100111111",
  434=>"111111111",
  435=>"000111111",
  436=>"011000000",
  437=>"010110110",
  438=>"111111111",
  439=>"000001000",
  440=>"000000011",
  441=>"111111110",
  442=>"000000000",
  443=>"000000110",
  444=>"000010000",
  445=>"010111111",
  446=>"111111001",
  447=>"110001000",
  448=>"000000000",
  449=>"000110110",
  450=>"111111011",
  451=>"000111000",
  452=>"111111111",
  453=>"011011100",
  454=>"001000000",
  455=>"101001101",
  456=>"111111111",
  457=>"111111100",
  458=>"000000001",
  459=>"001011011",
  460=>"010010000",
  461=>"001000111",
  462=>"000001011",
  463=>"100000101",
  464=>"000011001",
  465=>"000000011",
  466=>"111110010",
  467=>"000000110",
  468=>"000110000",
  469=>"111000101",
  470=>"111111001",
  471=>"001111111",
  472=>"001000000",
  473=>"000001001",
  474=>"000000110",
  475=>"111111101",
  476=>"011011001",
  477=>"011011000",
  478=>"000000000",
  479=>"111100000",
  480=>"111111000",
  481=>"111111111",
  482=>"000111111",
  483=>"011100100",
  484=>"111111111",
  485=>"000000000",
  486=>"111111111",
  487=>"100100111",
  488=>"100010111",
  489=>"111111111",
  490=>"011111100",
  491=>"111011001",
  492=>"000010110",
  493=>"000011011",
  494=>"000000001",
  495=>"111011000",
  496=>"000000000",
  497=>"000000000",
  498=>"000001100",
  499=>"001111011",
  500=>"011111110",
  501=>"001000001",
  502=>"111111000",
  503=>"101111111",
  504=>"000000000",
  505=>"000011011",
  506=>"011000000",
  507=>"000111111",
  508=>"111111000",
  509=>"000000100",
  510=>"100110110",
  511=>"000000100",
  512=>"000000000",
  513=>"000000000",
  514=>"111000110",
  515=>"000000000",
  516=>"111111110",
  517=>"001000000",
  518=>"000000001",
  519=>"111000110",
  520=>"111111111",
  521=>"100100000",
  522=>"001111001",
  523=>"001001111",
  524=>"000111000",
  525=>"110100000",
  526=>"111111111",
  527=>"111111111",
  528=>"110000000",
  529=>"111000000",
  530=>"000000000",
  531=>"111111111",
  532=>"000111000",
  533=>"111111111",
  534=>"111111111",
  535=>"000111111",
  536=>"000000110",
  537=>"101001100",
  538=>"100000000",
  539=>"101111110",
  540=>"000000000",
  541=>"111101101",
  542=>"011110110",
  543=>"100100100",
  544=>"111110111",
  545=>"000000010",
  546=>"110111111",
  547=>"001001001",
  548=>"111111001",
  549=>"000000000",
  550=>"111000101",
  551=>"000110100",
  552=>"111000000",
  553=>"111000000",
  554=>"110111000",
  555=>"111111111",
  556=>"111000000",
  557=>"110111111",
  558=>"111011011",
  559=>"000000011",
  560=>"111111100",
  561=>"000000000",
  562=>"000001001",
  563=>"000000000",
  564=>"111111011",
  565=>"111001000",
  566=>"001111111",
  567=>"000000000",
  568=>"111111010",
  569=>"111111000",
  570=>"111101111",
  571=>"011000000",
  572=>"111111000",
  573=>"111000000",
  574=>"110110010",
  575=>"111000111",
  576=>"000110111",
  577=>"101111111",
  578=>"000111111",
  579=>"111111000",
  580=>"000000000",
  581=>"110111111",
  582=>"110111111",
  583=>"111111111",
  584=>"011011000",
  585=>"001111111",
  586=>"111111111",
  587=>"111100100",
  588=>"111100111",
  589=>"000000101",
  590=>"011000010",
  591=>"000000000",
  592=>"111111111",
  593=>"001110110",
  594=>"111111111",
  595=>"000111111",
  596=>"111111111",
  597=>"000000110",
  598=>"110000000",
  599=>"000000011",
  600=>"111011000",
  601=>"111111111",
  602=>"111110111",
  603=>"111001001",
  604=>"001001110",
  605=>"111111111",
  606=>"010110110",
  607=>"100000000",
  608=>"000000100",
  609=>"000010000",
  610=>"010010000",
  611=>"000000000",
  612=>"001111111",
  613=>"111100000",
  614=>"100000110",
  615=>"011111000",
  616=>"011111111",
  617=>"010000111",
  618=>"000000101",
  619=>"000000000",
  620=>"001000000",
  621=>"111011110",
  622=>"111000000",
  623=>"111111111",
  624=>"111111110",
  625=>"000000000",
  626=>"111010010",
  627=>"000100100",
  628=>"000110010",
  629=>"000000000",
  630=>"111111011",
  631=>"000110111",
  632=>"000000111",
  633=>"000000001",
  634=>"000000011",
  635=>"000000000",
  636=>"001000111",
  637=>"111001011",
  638=>"110111100",
  639=>"000000001",
  640=>"000000011",
  641=>"111111010",
  642=>"111110100",
  643=>"100000000",
  644=>"111011111",
  645=>"100100000",
  646=>"111111111",
  647=>"111111010",
  648=>"111000000",
  649=>"000000000",
  650=>"000101101",
  651=>"111111111",
  652=>"111000100",
  653=>"111111010",
  654=>"100000000",
  655=>"111111110",
  656=>"000111110",
  657=>"001000111",
  658=>"111111111",
  659=>"100000000",
  660=>"110000000",
  661=>"001000000",
  662=>"000111111",
  663=>"110100000",
  664=>"100100100",
  665=>"111111111",
  666=>"111101110",
  667=>"000000000",
  668=>"101110111",
  669=>"111000000",
  670=>"001111111",
  671=>"000010111",
  672=>"011000001",
  673=>"001111111",
  674=>"000000000",
  675=>"000110111",
  676=>"001000000",
  677=>"100000000",
  678=>"000111110",
  679=>"110110110",
  680=>"101111111",
  681=>"000000000",
  682=>"111111000",
  683=>"111000010",
  684=>"000110111",
  685=>"001111110",
  686=>"111111011",
  687=>"110100100",
  688=>"000000111",
  689=>"000000000",
  690=>"110111110",
  691=>"101100101",
  692=>"000111111",
  693=>"000000111",
  694=>"000000000",
  695=>"111000000",
  696=>"111111111",
  697=>"111011000",
  698=>"111000010",
  699=>"100000000",
  700=>"111011011",
  701=>"101001111",
  702=>"100000000",
  703=>"111111111",
  704=>"110000000",
  705=>"111111111",
  706=>"000000010",
  707=>"000111111",
  708=>"111111010",
  709=>"000111111",
  710=>"000000001",
  711=>"111111111",
  712=>"111000000",
  713=>"001011111",
  714=>"111011011",
  715=>"111000000",
  716=>"000000010",
  717=>"111111100",
  718=>"110100000",
  719=>"011010001",
  720=>"111111111",
  721=>"000000110",
  722=>"001000000",
  723=>"011000000",
  724=>"111101001",
  725=>"111111110",
  726=>"010111111",
  727=>"110100111",
  728=>"101001000",
  729=>"111100111",
  730=>"111100000",
  731=>"111000110",
  732=>"000100111",
  733=>"111111111",
  734=>"111111111",
  735=>"111111111",
  736=>"001101111",
  737=>"111111011",
  738=>"000000101",
  739=>"111000000",
  740=>"000111111",
  741=>"110100100",
  742=>"000100100",
  743=>"111000100",
  744=>"111011000",
  745=>"000000000",
  746=>"101000000",
  747=>"000000000",
  748=>"111111111",
  749=>"000000000",
  750=>"011111111",
  751=>"000000000",
  752=>"000001111",
  753=>"111111100",
  754=>"100100000",
  755=>"111110100",
  756=>"100000000",
  757=>"100100111",
  758=>"110000000",
  759=>"000111111",
  760=>"000111000",
  761=>"111000000",
  762=>"000000000",
  763=>"001001100",
  764=>"011011010",
  765=>"111110000",
  766=>"000000000",
  767=>"111111111",
  768=>"000000101",
  769=>"000111101",
  770=>"111111000",
  771=>"000000100",
  772=>"111111111",
  773=>"100101111",
  774=>"110111111",
  775=>"111111000",
  776=>"000000000",
  777=>"000000000",
  778=>"001111111",
  779=>"111111111",
  780=>"000000000",
  781=>"000001111",
  782=>"111111100",
  783=>"001000111",
  784=>"010111110",
  785=>"011000000",
  786=>"000000111",
  787=>"000000111",
  788=>"000111111",
  789=>"111111000",
  790=>"111111100",
  791=>"101000001",
  792=>"111101011",
  793=>"000000110",
  794=>"000000000",
  795=>"100000000",
  796=>"001000000",
  797=>"000001110",
  798=>"000000000",
  799=>"111111000",
  800=>"000111111",
  801=>"010000101",
  802=>"000111111",
  803=>"000101111",
  804=>"101000000",
  805=>"000100111",
  806=>"000111111",
  807=>"101101000",
  808=>"111000000",
  809=>"111111010",
  810=>"010001001",
  811=>"011000000",
  812=>"111000000",
  813=>"111000000",
  814=>"101111011",
  815=>"000100001",
  816=>"011000110",
  817=>"000000000",
  818=>"010111111",
  819=>"000100110",
  820=>"011101000",
  821=>"001000101",
  822=>"011001111",
  823=>"111000100",
  824=>"111111000",
  825=>"111011111",
  826=>"111001000",
  827=>"000111111",
  828=>"000100100",
  829=>"100000000",
  830=>"011111111",
  831=>"000000000",
  832=>"000000000",
  833=>"000111111",
  834=>"101000000",
  835=>"000000111",
  836=>"000000111",
  837=>"000100101",
  838=>"000000000",
  839=>"011000000",
  840=>"000000000",
  841=>"111111000",
  842=>"000000111",
  843=>"010110110",
  844=>"000100110",
  845=>"000000000",
  846=>"100111111",
  847=>"000111111",
  848=>"000000100",
  849=>"110001111",
  850=>"000111111",
  851=>"111111111",
  852=>"111001000",
  853=>"000000001",
  854=>"000000111",
  855=>"000000100",
  856=>"000000101",
  857=>"000000000",
  858=>"110101000",
  859=>"000111111",
  860=>"000000000",
  861=>"111111001",
  862=>"100100001",
  863=>"000000111",
  864=>"000000000",
  865=>"111011011",
  866=>"000000111",
  867=>"111000000",
  868=>"011011000",
  869=>"110000000",
  870=>"101111111",
  871=>"001000111",
  872=>"100000000",
  873=>"111111110",
  874=>"000000000",
  875=>"111100000",
  876=>"111110110",
  877=>"111000011",
  878=>"011111011",
  879=>"110100000",
  880=>"111000000",
  881=>"011011111",
  882=>"111111111",
  883=>"110110111",
  884=>"111111111",
  885=>"111111111",
  886=>"111111111",
  887=>"000111111",
  888=>"000000000",
  889=>"111100000",
  890=>"111000000",
  891=>"110100000",
  892=>"101111101",
  893=>"111111111",
  894=>"000000000",
  895=>"111111011",
  896=>"001111111",
  897=>"101000011",
  898=>"111111111",
  899=>"111011000",
  900=>"011000000",
  901=>"100111111",
  902=>"110110000",
  903=>"011111110",
  904=>"000000000",
  905=>"000100000",
  906=>"111000001",
  907=>"100111111",
  908=>"111111111",
  909=>"000110111",
  910=>"100001000",
  911=>"000100111",
  912=>"111000000",
  913=>"111111110",
  914=>"110111111",
  915=>"011011011",
  916=>"110111111",
  917=>"000000000",
  918=>"000000000",
  919=>"111011110",
  920=>"000000111",
  921=>"100000000",
  922=>"001011111",
  923=>"000000111",
  924=>"000001000",
  925=>"111101000",
  926=>"001000111",
  927=>"000000000",
  928=>"011011111",
  929=>"001110111",
  930=>"011011011",
  931=>"010111111",
  932=>"000010111",
  933=>"111111010",
  934=>"000000000",
  935=>"011000000",
  936=>"000011111",
  937=>"100110110",
  938=>"101101110",
  939=>"001000000",
  940=>"000110111",
  941=>"000000101",
  942=>"111111111",
  943=>"001000000",
  944=>"111111111",
  945=>"011000000",
  946=>"111000000",
  947=>"110110110",
  948=>"000000101",
  949=>"101100011",
  950=>"001111111",
  951=>"000000100",
  952=>"101100111",
  953=>"000000000",
  954=>"000000100",
  955=>"100000000",
  956=>"110000111",
  957=>"111111111",
  958=>"110111111",
  959=>"101001111",
  960=>"111011000",
  961=>"011000000",
  962=>"010011111",
  963=>"101111111",
  964=>"000000000",
  965=>"110000000",
  966=>"000000001",
  967=>"000001111",
  968=>"000000101",
  969=>"100000000",
  970=>"000110110",
  971=>"110110111",
  972=>"100111000",
  973=>"000000001",
  974=>"100000000",
  975=>"000110111",
  976=>"100111111",
  977=>"000111111",
  978=>"000000111",
  979=>"111100000",
  980=>"000000000",
  981=>"000011111",
  982=>"111011011",
  983=>"111111000",
  984=>"000000000",
  985=>"110010111",
  986=>"111111000",
  987=>"011000000",
  988=>"000011111",
  989=>"100000111",
  990=>"111001001",
  991=>"000100000",
  992=>"110100110",
  993=>"011000001",
  994=>"000000000",
  995=>"000100011",
  996=>"010110000",
  997=>"011111111",
  998=>"111100000",
  999=>"000110110",
  1000=>"111000000",
  1001=>"101101111",
  1002=>"000000111",
  1003=>"100000010",
  1004=>"000111111",
  1005=>"100000001",
  1006=>"000000001",
  1007=>"001000000",
  1008=>"101000000",
  1009=>"011000000",
  1010=>"111111111",
  1011=>"111011111",
  1012=>"111000000",
  1013=>"110000000",
  1014=>"111110100",
  1015=>"111110111",
  1016=>"111111001",
  1017=>"000100111",
  1018=>"000000000",
  1019=>"111111111",
  1020=>"000000010",
  1021=>"111110111",
  1022=>"110111111",
  1023=>"000111111",
  1024=>"100110111",
  1025=>"101111110",
  1026=>"101100100",
  1027=>"000100111",
  1028=>"111110110",
  1029=>"000000000",
  1030=>"010010010",
  1031=>"101001111",
  1032=>"000000111",
  1033=>"000000100",
  1034=>"001001001",
  1035=>"011111000",
  1036=>"110110110",
  1037=>"000010110",
  1038=>"110100100",
  1039=>"111000000",
  1040=>"000100110",
  1041=>"111111111",
  1042=>"000000000",
  1043=>"000000010",
  1044=>"000000000",
  1045=>"000000000",
  1046=>"101101101",
  1047=>"000100101",
  1048=>"000000100",
  1049=>"110101111",
  1050=>"111100111",
  1051=>"100110111",
  1052=>"111111111",
  1053=>"110011000",
  1054=>"100000100",
  1055=>"111111000",
  1056=>"100101101",
  1057=>"101000111",
  1058=>"110110111",
  1059=>"111111111",
  1060=>"011000000",
  1061=>"111111101",
  1062=>"001000110",
  1063=>"000000000",
  1064=>"111111111",
  1065=>"100000100",
  1066=>"001001111",
  1067=>"100100001",
  1068=>"100110110",
  1069=>"000000000",
  1070=>"000000101",
  1071=>"000010000",
  1072=>"001001000",
  1073=>"010110010",
  1074=>"111111110",
  1075=>"111111001",
  1076=>"110010001",
  1077=>"110110111",
  1078=>"110001011",
  1079=>"000000101",
  1080=>"111110000",
  1081=>"111100111",
  1082=>"001010111",
  1083=>"011001111",
  1084=>"001001111",
  1085=>"111000000",
  1086=>"011001000",
  1087=>"111111111",
  1088=>"000110111",
  1089=>"111111111",
  1090=>"111110100",
  1091=>"111000000",
  1092=>"110110110",
  1093=>"011001101",
  1094=>"111111001",
  1095=>"111111111",
  1096=>"000001000",
  1097=>"001000000",
  1098=>"110111111",
  1099=>"101000010",
  1100=>"100000010",
  1101=>"000110111",
  1102=>"010110110",
  1103=>"000000000",
  1104=>"001000000",
  1105=>"001111101",
  1106=>"000001111",
  1107=>"110100000",
  1108=>"010111110",
  1109=>"001001000",
  1110=>"001000011",
  1111=>"101101101",
  1112=>"010110000",
  1113=>"101000000",
  1114=>"001001111",
  1115=>"000000100",
  1116=>"000000000",
  1117=>"111101111",
  1118=>"111111110",
  1119=>"000011011",
  1120=>"001111111",
  1121=>"000111111",
  1122=>"111111010",
  1123=>"111010000",
  1124=>"111000000",
  1125=>"111001100",
  1126=>"110111110",
  1127=>"000000000",
  1128=>"001001000",
  1129=>"000000000",
  1130=>"011001011",
  1131=>"111111010",
  1132=>"110110110",
  1133=>"111111010",
  1134=>"000000000",
  1135=>"111111101",
  1136=>"000000000",
  1137=>"001101001",
  1138=>"000000000",
  1139=>"111100111",
  1140=>"000000000",
  1141=>"000000110",
  1142=>"000111111",
  1143=>"111101100",
  1144=>"101000000",
  1145=>"110111110",
  1146=>"100000000",
  1147=>"100111111",
  1148=>"000001001",
  1149=>"000000000",
  1150=>"010111110",
  1151=>"000100000",
  1152=>"101000000",
  1153=>"000010000",
  1154=>"111111110",
  1155=>"111011001",
  1156=>"111111111",
  1157=>"000000111",
  1158=>"100000110",
  1159=>"111011000",
  1160=>"111010000",
  1161=>"001001111",
  1162=>"111110000",
  1163=>"001001001",
  1164=>"001001000",
  1165=>"000001101",
  1166=>"011101101",
  1167=>"111111010",
  1168=>"101101101",
  1169=>"000110000",
  1170=>"000111111",
  1171=>"111111110",
  1172=>"000000011",
  1173=>"000000110",
  1174=>"000000001",
  1175=>"101000001",
  1176=>"001001101",
  1177=>"000000000",
  1178=>"111111110",
  1179=>"000100100",
  1180=>"111111111",
  1181=>"000000001",
  1182=>"111110000",
  1183=>"111111111",
  1184=>"111111111",
  1185=>"100000000",
  1186=>"111111110",
  1187=>"000000111",
  1188=>"110110110",
  1189=>"111111110",
  1190=>"000000000",
  1191=>"101001111",
  1192=>"101000111",
  1193=>"001111111",
  1194=>"000000000",
  1195=>"100100000",
  1196=>"111111111",
  1197=>"100100100",
  1198=>"010111111",
  1199=>"110111111",
  1200=>"011111111",
  1201=>"111110110",
  1202=>"010111010",
  1203=>"111101000",
  1204=>"100010111",
  1205=>"010000000",
  1206=>"000000000",
  1207=>"101111110",
  1208=>"111111111",
  1209=>"011111101",
  1210=>"111001000",
  1211=>"001001000",
  1212=>"001011011",
  1213=>"000000111",
  1214=>"001000000",
  1215=>"000000000",
  1216=>"011000010",
  1217=>"001001000",
  1218=>"000100110",
  1219=>"101000000",
  1220=>"001111110",
  1221=>"000000000",
  1222=>"110000111",
  1223=>"000000001",
  1224=>"001111000",
  1225=>"111101111",
  1226=>"000000100",
  1227=>"001111111",
  1228=>"111110100",
  1229=>"000111111",
  1230=>"111111111",
  1231=>"000000001",
  1232=>"000111111",
  1233=>"000101101",
  1234=>"000000001",
  1235=>"000000000",
  1236=>"111101100",
  1237=>"110110000",
  1238=>"111111011",
  1239=>"000101000",
  1240=>"000000000",
  1241=>"000000101",
  1242=>"110110111",
  1243=>"000001111",
  1244=>"000000000",
  1245=>"101011011",
  1246=>"110110000",
  1247=>"111101111",
  1248=>"111111111",
  1249=>"000000111",
  1250=>"000000000",
  1251=>"111110111",
  1252=>"000000000",
  1253=>"001001011",
  1254=>"000000000",
  1255=>"000000101",
  1256=>"000000110",
  1257=>"011011000",
  1258=>"011110110",
  1259=>"000100100",
  1260=>"111101101",
  1261=>"101111000",
  1262=>"111110111",
  1263=>"111100000",
  1264=>"000001111",
  1265=>"110000100",
  1266=>"000000000",
  1267=>"111110110",
  1268=>"111111111",
  1269=>"001111111",
  1270=>"110110111",
  1271=>"111100111",
  1272=>"111011000",
  1273=>"000001101",
  1274=>"111000001",
  1275=>"111111111",
  1276=>"001011001",
  1277=>"001001001",
  1278=>"000000111",
  1279=>"000000010",
  1280=>"000000000",
  1281=>"100000101",
  1282=>"000011111",
  1283=>"000101111",
  1284=>"111111000",
  1285=>"001111111",
  1286=>"001000000",
  1287=>"011011011",
  1288=>"111111110",
  1289=>"000000001",
  1290=>"111111101",
  1291=>"111111011",
  1292=>"101000000",
  1293=>"000110111",
  1294=>"000110110",
  1295=>"000011111",
  1296=>"100100110",
  1297=>"000111110",
  1298=>"000101111",
  1299=>"111111110",
  1300=>"010110110",
  1301=>"000001011",
  1302=>"111111111",
  1303=>"000000101",
  1304=>"111111001",
  1305=>"111010000",
  1306=>"000000111",
  1307=>"000111111",
  1308=>"000000001",
  1309=>"001001001",
  1310=>"000000000",
  1311=>"111111111",
  1312=>"010000000",
  1313=>"001001101",
  1314=>"000000101",
  1315=>"011111111",
  1316=>"110100100",
  1317=>"010111000",
  1318=>"001000000",
  1319=>"010000000",
  1320=>"100100110",
  1321=>"111111011",
  1322=>"010110000",
  1323=>"000011000",
  1324=>"111111110",
  1325=>"100110110",
  1326=>"000000000",
  1327=>"001001010",
  1328=>"000000000",
  1329=>"000000001",
  1330=>"011000000",
  1331=>"100000010",
  1332=>"000000111",
  1333=>"000011111",
  1334=>"100000101",
  1335=>"000010000",
  1336=>"010000010",
  1337=>"111111111",
  1338=>"101000101",
  1339=>"000000111",
  1340=>"111000000",
  1341=>"111101001",
  1342=>"111110000",
  1343=>"111000000",
  1344=>"101101100",
  1345=>"001001000",
  1346=>"111000000",
  1347=>"001001101",
  1348=>"001111111",
  1349=>"111100111",
  1350=>"111000000",
  1351=>"001001010",
  1352=>"100000100",
  1353=>"000000000",
  1354=>"000110100",
  1355=>"111100000",
  1356=>"000000000",
  1357=>"000000111",
  1358=>"111001001",
  1359=>"111111011",
  1360=>"001001011",
  1361=>"001001000",
  1362=>"111111000",
  1363=>"000000110",
  1364=>"000000000",
  1365=>"011011000",
  1366=>"111111111",
  1367=>"001100000",
  1368=>"111111111",
  1369=>"000000000",
  1370=>"111111111",
  1371=>"000111110",
  1372=>"000000101",
  1373=>"000000000",
  1374=>"000000000",
  1375=>"000000111",
  1376=>"000111111",
  1377=>"001000000",
  1378=>"011001001",
  1379=>"000000011",
  1380=>"110110100",
  1381=>"111111111",
  1382=>"000001111",
  1383=>"001001001",
  1384=>"101000000",
  1385=>"001001000",
  1386=>"000000000",
  1387=>"111111111",
  1388=>"110110100",
  1389=>"111101000",
  1390=>"000000001",
  1391=>"101001101",
  1392=>"111101101",
  1393=>"100100111",
  1394=>"011110111",
  1395=>"011011011",
  1396=>"011000111",
  1397=>"000000101",
  1398=>"100111111",
  1399=>"000000001",
  1400=>"001001001",
  1401=>"111111111",
  1402=>"101000100",
  1403=>"110110110",
  1404=>"010000000",
  1405=>"000111111",
  1406=>"111110111",
  1407=>"101001111",
  1408=>"111011000",
  1409=>"000001000",
  1410=>"100000000",
  1411=>"000000000",
  1412=>"000000000",
  1413=>"100001101",
  1414=>"000100111",
  1415=>"110110000",
  1416=>"101000000",
  1417=>"000010110",
  1418=>"111110000",
  1419=>"000000000",
  1420=>"101111111",
  1421=>"100100111",
  1422=>"100110010",
  1423=>"010010000",
  1424=>"100000000",
  1425=>"110111101",
  1426=>"000001101",
  1427=>"111001011",
  1428=>"000000000",
  1429=>"000000000",
  1430=>"111010010",
  1431=>"110110111",
  1432=>"000000000",
  1433=>"001111111",
  1434=>"111111011",
  1435=>"111111000",
  1436=>"001001001",
  1437=>"111111000",
  1438=>"101001001",
  1439=>"111111111",
  1440=>"000100000",
  1441=>"001001000",
  1442=>"101000001",
  1443=>"100000011",
  1444=>"111111101",
  1445=>"000000000",
  1446=>"101111111",
  1447=>"000000100",
  1448=>"001001001",
  1449=>"101111111",
  1450=>"110111110",
  1451=>"001111100",
  1452=>"000000000",
  1453=>"000100001",
  1454=>"000000111",
  1455=>"111111101",
  1456=>"001110110",
  1457=>"110110000",
  1458=>"010010010",
  1459=>"000000100",
  1460=>"001001101",
  1461=>"001000001",
  1462=>"111110000",
  1463=>"000000100",
  1464=>"001001101",
  1465=>"000000110",
  1466=>"111011001",
  1467=>"001011111",
  1468=>"000011011",
  1469=>"111011011",
  1470=>"010010000",
  1471=>"000000100",
  1472=>"011011001",
  1473=>"111111111",
  1474=>"001000000",
  1475=>"000000000",
  1476=>"111110000",
  1477=>"011001011",
  1478=>"000000101",
  1479=>"000000000",
  1480=>"001001011",
  1481=>"111000010",
  1482=>"001001101",
  1483=>"111111001",
  1484=>"011011001",
  1485=>"000000010",
  1486=>"000000000",
  1487=>"110111110",
  1488=>"001000100",
  1489=>"101100000",
  1490=>"100000000",
  1491=>"000000001",
  1492=>"000011111",
  1493=>"111001000",
  1494=>"111111111",
  1495=>"011011011",
  1496=>"001111110",
  1497=>"000000000",
  1498=>"100000000",
  1499=>"111010011",
  1500=>"000000101",
  1501=>"000000001",
  1502=>"100000000",
  1503=>"100100110",
  1504=>"001000001",
  1505=>"111011000",
  1506=>"010111111",
  1507=>"001011111",
  1508=>"111111000",
  1509=>"010010000",
  1510=>"000001111",
  1511=>"000000000",
  1512=>"001000001",
  1513=>"100110000",
  1514=>"000000101",
  1515=>"101100101",
  1516=>"001000000",
  1517=>"111111111",
  1518=>"101101111",
  1519=>"001000000",
  1520=>"111111010",
  1521=>"000000000",
  1522=>"000001000",
  1523=>"000000000",
  1524=>"000000000",
  1525=>"000000000",
  1526=>"000000000",
  1527=>"000100100",
  1528=>"010000011",
  1529=>"011101111",
  1530=>"110110110",
  1531=>"000000000",
  1532=>"000000111",
  1533=>"000000101",
  1534=>"111000100",
  1535=>"000000000",
  1536=>"001011111",
  1537=>"111111111",
  1538=>"000111111",
  1539=>"000000000",
  1540=>"000000000",
  1541=>"011011001",
  1542=>"100111010",
  1543=>"111101111",
  1544=>"111100000",
  1545=>"011011011",
  1546=>"001000101",
  1547=>"111111111",
  1548=>"011011011",
  1549=>"111111111",
  1550=>"000011011",
  1551=>"111111000",
  1552=>"110110111",
  1553=>"000110111",
  1554=>"000000001",
  1555=>"000000000",
  1556=>"111001000",
  1557=>"111111111",
  1558=>"000100110",
  1559=>"111111111",
  1560=>"011011011",
  1561=>"111001000",
  1562=>"010111111",
  1563=>"111111111",
  1564=>"000000000",
  1565=>"011000111",
  1566=>"011001001",
  1567=>"000000100",
  1568=>"111001001",
  1569=>"000111111",
  1570=>"000000100",
  1571=>"000000110",
  1572=>"000000000",
  1573=>"001100110",
  1574=>"000001001",
  1575=>"111001001",
  1576=>"011111111",
  1577=>"111111111",
  1578=>"111011001",
  1579=>"110111111",
  1580=>"111111111",
  1581=>"111000000",
  1582=>"100101110",
  1583=>"000001011",
  1584=>"100000100",
  1585=>"100000000",
  1586=>"111000000",
  1587=>"011111111",
  1588=>"000000000",
  1589=>"011011101",
  1590=>"001101001",
  1591=>"111111111",
  1592=>"111111100",
  1593=>"000001111",
  1594=>"011111111",
  1595=>"001000000",
  1596=>"111111111",
  1597=>"000000010",
  1598=>"111110110",
  1599=>"111111111",
  1600=>"010000000",
  1601=>"011011011",
  1602=>"000000111",
  1603=>"111111111",
  1604=>"000000100",
  1605=>"111111110",
  1606=>"000000101",
  1607=>"111111111",
  1608=>"111111011",
  1609=>"111001111",
  1610=>"010111111",
  1611=>"000110000",
  1612=>"111011110",
  1613=>"100100100",
  1614=>"001001001",
  1615=>"111000000",
  1616=>"100000000",
  1617=>"111111111",
  1618=>"001111000",
  1619=>"010111010",
  1620=>"110110111",
  1621=>"000110110",
  1622=>"001101101",
  1623=>"111111111",
  1624=>"000001011",
  1625=>"000000000",
  1626=>"000100000",
  1627=>"100000001",
  1628=>"000000011",
  1629=>"000111111",
  1630=>"111111101",
  1631=>"000111100",
  1632=>"000000000",
  1633=>"000000000",
  1634=>"000000000",
  1635=>"000000000",
  1636=>"111111111",
  1637=>"000100100",
  1638=>"000100111",
  1639=>"000000000",
  1640=>"001000111",
  1641=>"000000000",
  1642=>"011011110",
  1643=>"100100110",
  1644=>"111111111",
  1645=>"000000000",
  1646=>"001000111",
  1647=>"111111101",
  1648=>"000010110",
  1649=>"111111111",
  1650=>"111100100",
  1651=>"000000000",
  1652=>"100111111",
  1653=>"000111110",
  1654=>"010110000",
  1655=>"000000000",
  1656=>"111111111",
  1657=>"000010000",
  1658=>"000000000",
  1659=>"000000000",
  1660=>"011011000",
  1661=>"000010111",
  1662=>"000000000",
  1663=>"110010000",
  1664=>"001001011",
  1665=>"111010000",
  1666=>"111111111",
  1667=>"111101001",
  1668=>"000000000",
  1669=>"001001000",
  1670=>"111110000",
  1671=>"000000000",
  1672=>"101111011",
  1673=>"000000000",
  1674=>"011000000",
  1675=>"011011001",
  1676=>"000000011",
  1677=>"111111000",
  1678=>"111111111",
  1679=>"000000000",
  1680=>"010010000",
  1681=>"110100100",
  1682=>"000010000",
  1683=>"000000000",
  1684=>"001001111",
  1685=>"001001001",
  1686=>"110110000",
  1687=>"011111111",
  1688=>"101000000",
  1689=>"000000000",
  1690=>"000000000",
  1691=>"010010111",
  1692=>"111111111",
  1693=>"110110101",
  1694=>"111111111",
  1695=>"111111000",
  1696=>"111100000",
  1697=>"101001111",
  1698=>"000111111",
  1699=>"000000000",
  1700=>"000001001",
  1701=>"001001111",
  1702=>"111111111",
  1703=>"111100100",
  1704=>"100000011",
  1705=>"000000000",
  1706=>"000000000",
  1707=>"000000000",
  1708=>"101000000",
  1709=>"010000000",
  1710=>"111111111",
  1711=>"101000000",
  1712=>"000000111",
  1713=>"001010110",
  1714=>"000000000",
  1715=>"000000000",
  1716=>"100000000",
  1717=>"110110110",
  1718=>"000000001",
  1719=>"111111111",
  1720=>"111100111",
  1721=>"111111000",
  1722=>"000110111",
  1723=>"000000100",
  1724=>"000000100",
  1725=>"011111111",
  1726=>"000000100",
  1727=>"000000000",
  1728=>"111111111",
  1729=>"000000111",
  1730=>"100010110",
  1731=>"001000000",
  1732=>"100100000",
  1733=>"011111111",
  1734=>"001000111",
  1735=>"000000000",
  1736=>"100100000",
  1737=>"111101101",
  1738=>"010000000",
  1739=>"111111111",
  1740=>"111100101",
  1741=>"111111111",
  1742=>"000000010",
  1743=>"100000000",
  1744=>"000000001",
  1745=>"000000111",
  1746=>"110111100",
  1747=>"001000101",
  1748=>"001001001",
  1749=>"001001001",
  1750=>"000111111",
  1751=>"010000101",
  1752=>"000000000",
  1753=>"111001001",
  1754=>"111111111",
  1755=>"111111111",
  1756=>"000000000",
  1757=>"001011111",
  1758=>"000011000",
  1759=>"001001001",
  1760=>"111111111",
  1761=>"000000100",
  1762=>"000100100",
  1763=>"111111111",
  1764=>"101111111",
  1765=>"011100100",
  1766=>"111111111",
  1767=>"111111111",
  1768=>"111111111",
  1769=>"000000011",
  1770=>"111111111",
  1771=>"111111111",
  1772=>"000000011",
  1773=>"111111001",
  1774=>"000000000",
  1775=>"000000100",
  1776=>"111111001",
  1777=>"000000111",
  1778=>"000000100",
  1779=>"100000000",
  1780=>"111111111",
  1781=>"000000000",
  1782=>"111111110",
  1783=>"000100110",
  1784=>"111111111",
  1785=>"101101000",
  1786=>"110111111",
  1787=>"000100101",
  1788=>"111111111",
  1789=>"010110110",
  1790=>"100111111",
  1791=>"100111111",
  1792=>"111111111",
  1793=>"111001100",
  1794=>"011111111",
  1795=>"000000000",
  1796=>"100001101",
  1797=>"001011111",
  1798=>"111111011",
  1799=>"001000001",
  1800=>"000000000",
  1801=>"000000000",
  1802=>"100100001",
  1803=>"111101101",
  1804=>"110110100",
  1805=>"110111111",
  1806=>"101101101",
  1807=>"111100000",
  1808=>"111011001",
  1809=>"111111111",
  1810=>"111111111",
  1811=>"000000001",
  1812=>"111110100",
  1813=>"111111111",
  1814=>"000110000",
  1815=>"110111111",
  1816=>"000100000",
  1817=>"111111110",
  1818=>"111111111",
  1819=>"111111111",
  1820=>"001001001",
  1821=>"111111111",
  1822=>"000000011",
  1823=>"111110111",
  1824=>"011001001",
  1825=>"100111111",
  1826=>"100000101",
  1827=>"100101011",
  1828=>"001001111",
  1829=>"000000001",
  1830=>"101111101",
  1831=>"001001011",
  1832=>"001011100",
  1833=>"011000000",
  1834=>"000000001",
  1835=>"110011000",
  1836=>"011001000",
  1837=>"111110110",
  1838=>"000100000",
  1839=>"010000000",
  1840=>"001001101",
  1841=>"000000000",
  1842=>"000000010",
  1843=>"111111110",
  1844=>"000000000",
  1845=>"111111111",
  1846=>"000100111",
  1847=>"111111111",
  1848=>"000000000",
  1849=>"110110111",
  1850=>"000000000",
  1851=>"000011011",
  1852=>"000000000",
  1853=>"001110111",
  1854=>"111110110",
  1855=>"111111111",
  1856=>"000000000",
  1857=>"111111111",
  1858=>"000000100",
  1859=>"000000000",
  1860=>"001011011",
  1861=>"101001111",
  1862=>"110111000",
  1863=>"111111111",
  1864=>"100000000",
  1865=>"111111111",
  1866=>"111101001",
  1867=>"100000000",
  1868=>"111111000",
  1869=>"111101000",
  1870=>"001101000",
  1871=>"111111111",
  1872=>"111111010",
  1873=>"111111111",
  1874=>"111111111",
  1875=>"111111111",
  1876=>"111111111",
  1877=>"111100001",
  1878=>"000000000",
  1879=>"111111111",
  1880=>"111101101",
  1881=>"111101101",
  1882=>"011001000",
  1883=>"000000000",
  1884=>"111111111",
  1885=>"000000000",
  1886=>"111111111",
  1887=>"111001000",
  1888=>"001111111",
  1889=>"100100100",
  1890=>"000000000",
  1891=>"000000011",
  1892=>"110100100",
  1893=>"111111111",
  1894=>"111111111",
  1895=>"101101000",
  1896=>"111011001",
  1897=>"110110000",
  1898=>"000000111",
  1899=>"000100100",
  1900=>"111001001",
  1901=>"110111000",
  1902=>"111111111",
  1903=>"000011111",
  1904=>"000000101",
  1905=>"000000000",
  1906=>"111011001",
  1907=>"000000000",
  1908=>"111111101",
  1909=>"111111111",
  1910=>"000000000",
  1911=>"000000100",
  1912=>"101000111",
  1913=>"111111111",
  1914=>"111111111",
  1915=>"001000000",
  1916=>"001001111",
  1917=>"000000111",
  1918=>"111000000",
  1919=>"000000000",
  1920=>"011011011",
  1921=>"000100100",
  1922=>"111111111",
  1923=>"110011001",
  1924=>"110100000",
  1925=>"110100000",
  1926=>"000100100",
  1927=>"011011011",
  1928=>"000000001",
  1929=>"011111010",
  1930=>"111111101",
  1931=>"000000111",
  1932=>"000110111",
  1933=>"000000010",
  1934=>"101111111",
  1935=>"001111111",
  1936=>"111111111",
  1937=>"000000000",
  1938=>"101111111",
  1939=>"000000000",
  1940=>"000000101",
  1941=>"111011001",
  1942=>"100100111",
  1943=>"100100000",
  1944=>"111111111",
  1945=>"000000000",
  1946=>"000110000",
  1947=>"111111111",
  1948=>"000000000",
  1949=>"110111010",
  1950=>"100100100",
  1951=>"000000000",
  1952=>"000000000",
  1953=>"011101101",
  1954=>"100000111",
  1955=>"110111111",
  1956=>"111111111",
  1957=>"001000000",
  1958=>"111111111",
  1959=>"000010111",
  1960=>"001001101",
  1961=>"011001111",
  1962=>"000000000",
  1963=>"110100100",
  1964=>"000000000",
  1965=>"111111111",
  1966=>"111101001",
  1967=>"011001001",
  1968=>"100111111",
  1969=>"111110100",
  1970=>"000000101",
  1971=>"110111111",
  1972=>"000000000",
  1973=>"000000001",
  1974=>"111011111",
  1975=>"111111111",
  1976=>"011111011",
  1977=>"110000111",
  1978=>"001001001",
  1979=>"000000010",
  1980=>"111111111",
  1981=>"111001000",
  1982=>"000011111",
  1983=>"000001000",
  1984=>"000001000",
  1985=>"111011000",
  1986=>"000000000",
  1987=>"000000000",
  1988=>"111100000",
  1989=>"111111000",
  1990=>"010010000",
  1991=>"000111111",
  1992=>"111111111",
  1993=>"111111111",
  1994=>"111111111",
  1995=>"111111111",
  1996=>"000000000",
  1997=>"111111111",
  1998=>"111111110",
  1999=>"100000000",
  2000=>"110111101",
  2001=>"000100100",
  2002=>"000000000",
  2003=>"000000000",
  2004=>"110110111",
  2005=>"111111111",
  2006=>"000000100",
  2007=>"110110111",
  2008=>"111111101",
  2009=>"100000001",
  2010=>"111110110",
  2011=>"111111111",
  2012=>"100000100",
  2013=>"000001011",
  2014=>"111100111",
  2015=>"001011111",
  2016=>"111111111",
  2017=>"000000000",
  2018=>"111111111",
  2019=>"000001111",
  2020=>"100111110",
  2021=>"111111111",
  2022=>"001000001",
  2023=>"111111111",
  2024=>"110110110",
  2025=>"000000111",
  2026=>"100000011",
  2027=>"111111111",
  2028=>"100001111",
  2029=>"111000000",
  2030=>"000000111",
  2031=>"000011111",
  2032=>"000000000",
  2033=>"000000001",
  2034=>"111111111",
  2035=>"100000000",
  2036=>"000000000",
  2037=>"000000000",
  2038=>"111111111",
  2039=>"010011011",
  2040=>"111101111",
  2041=>"110010010",
  2042=>"110111111",
  2043=>"000010010",
  2044=>"111111111",
  2045=>"000000000",
  2046=>"111111111",
  2047=>"111111111",
  2048=>"111111111",
  2049=>"010010111",
  2050=>"111111111",
  2051=>"000000011",
  2052=>"111001111",
  2053=>"111111001",
  2054=>"000001111",
  2055=>"111001000",
  2056=>"011111111",
  2057=>"000000000",
  2058=>"011001011",
  2059=>"000000111",
  2060=>"100100000",
  2061=>"000100111",
  2062=>"111010000",
  2063=>"000111111",
  2064=>"110000000",
  2065=>"000000000",
  2066=>"100110111",
  2067=>"111111111",
  2068=>"101111111",
  2069=>"111111111",
  2070=>"111111111",
  2071=>"100100100",
  2072=>"110011001",
  2073=>"100010010",
  2074=>"100000110",
  2075=>"010111111",
  2076=>"001000011",
  2077=>"001101111",
  2078=>"000110100",
  2079=>"111111110",
  2080=>"000000000",
  2081=>"000000000",
  2082=>"111111111",
  2083=>"011111100",
  2084=>"111111111",
  2085=>"100110000",
  2086=>"111111101",
  2087=>"100000000",
  2088=>"001000000",
  2089=>"111111111",
  2090=>"111111011",
  2091=>"100111000",
  2092=>"000000000",
  2093=>"000000111",
  2094=>"000100111",
  2095=>"001000000",
  2096=>"110010100",
  2097=>"111111111",
  2098=>"100100100",
  2099=>"000000000",
  2100=>"000011011",
  2101=>"000000000",
  2102=>"011011000",
  2103=>"100100000",
  2104=>"111111111",
  2105=>"111000110",
  2106=>"011111111",
  2107=>"000111111",
  2108=>"000000000",
  2109=>"000100100",
  2110=>"010000100",
  2111=>"111111111",
  2112=>"110000000",
  2113=>"111010100",
  2114=>"111111000",
  2115=>"111100000",
  2116=>"111111111",
  2117=>"000000110",
  2118=>"111111111",
  2119=>"010000000",
  2120=>"000000000",
  2121=>"111010010",
  2122=>"111111111",
  2123=>"000000000",
  2124=>"001001110",
  2125=>"111111111",
  2126=>"000000000",
  2127=>"000000000",
  2128=>"000000000",
  2129=>"000000100",
  2130=>"000000000",
  2131=>"101000000",
  2132=>"111110000",
  2133=>"000000110",
  2134=>"110100100",
  2135=>"110000000",
  2136=>"000000000",
  2137=>"111111111",
  2138=>"011001111",
  2139=>"000100000",
  2140=>"111111111",
  2141=>"000000000",
  2142=>"000000000",
  2143=>"001000111",
  2144=>"010111010",
  2145=>"111110100",
  2146=>"100111100",
  2147=>"001000100",
  2148=>"000000011",
  2149=>"110111111",
  2150=>"100100000",
  2151=>"000110111",
  2152=>"111111111",
  2153=>"000000000",
  2154=>"111000000",
  2155=>"111111111",
  2156=>"000000000",
  2157=>"000000101",
  2158=>"100100111",
  2159=>"111111111",
  2160=>"100100000",
  2161=>"111101110",
  2162=>"000000000",
  2163=>"000000000",
  2164=>"000000100",
  2165=>"000001001",
  2166=>"000010110",
  2167=>"000000000",
  2168=>"100100111",
  2169=>"110110100",
  2170=>"000100100",
  2171=>"100000000",
  2172=>"100110101",
  2173=>"111111111",
  2174=>"000000110",
  2175=>"000001000",
  2176=>"110110000",
  2177=>"000000100",
  2178=>"000000010",
  2179=>"000000000",
  2180=>"000111111",
  2181=>"000000101",
  2182=>"111111111",
  2183=>"000000110",
  2184=>"111111111",
  2185=>"000000000",
  2186=>"001111111",
  2187=>"111111111",
  2188=>"111111111",
  2189=>"000000000",
  2190=>"100100100",
  2191=>"111111111",
  2192=>"000000000",
  2193=>"000000000",
  2194=>"100111111",
  2195=>"100000111",
  2196=>"111110110",
  2197=>"000000000",
  2198=>"101001000",
  2199=>"000000000",
  2200=>"110110110",
  2201=>"111111110",
  2202=>"001000000",
  2203=>"000000000",
  2204=>"110100101",
  2205=>"110010011",
  2206=>"111101111",
  2207=>"000000000",
  2208=>"100100111",
  2209=>"111110111",
  2210=>"011001100",
  2211=>"000001111",
  2212=>"000000000",
  2213=>"110000000",
  2214=>"111001110",
  2215=>"000010110",
  2216=>"100111111",
  2217=>"111111111",
  2218=>"001000000",
  2219=>"111101000",
  2220=>"001000000",
  2221=>"011001011",
  2222=>"000000001",
  2223=>"100100001",
  2224=>"111011111",
  2225=>"000100110",
  2226=>"111111110",
  2227=>"100000000",
  2228=>"110111111",
  2229=>"100000000",
  2230=>"000000000",
  2231=>"000000100",
  2232=>"000000000",
  2233=>"111001001",
  2234=>"000000000",
  2235=>"000000100",
  2236=>"111011010",
  2237=>"000000000",
  2238=>"000110111",
  2239=>"000010110",
  2240=>"000000111",
  2241=>"011001111",
  2242=>"111111111",
  2243=>"111111111",
  2244=>"000001000",
  2245=>"000000000",
  2246=>"000000000",
  2247=>"100000000",
  2248=>"000011011",
  2249=>"101101101",
  2250=>"100000000",
  2251=>"001011011",
  2252=>"111111111",
  2253=>"010110100",
  2254=>"100000000",
  2255=>"000000000",
  2256=>"000000111",
  2257=>"100101101",
  2258=>"000000101",
  2259=>"000010111",
  2260=>"001000000",
  2261=>"110111111",
  2262=>"011000100",
  2263=>"000000001",
  2264=>"001101000",
  2265=>"000100110",
  2266=>"000000000",
  2267=>"000000000",
  2268=>"000000000",
  2269=>"111111111",
  2270=>"111111111",
  2271=>"100100001",
  2272=>"111111111",
  2273=>"001000111",
  2274=>"010110111",
  2275=>"000000000",
  2276=>"111111110",
  2277=>"011010101",
  2278=>"000000000",
  2279=>"011111111",
  2280=>"100101111",
  2281=>"000000000",
  2282=>"000101111",
  2283=>"111111111",
  2284=>"111111111",
  2285=>"111111111",
  2286=>"101111110",
  2287=>"011000000",
  2288=>"111000000",
  2289=>"000000110",
  2290=>"111111111",
  2291=>"100100001",
  2292=>"111111111",
  2293=>"111000110",
  2294=>"000110100",
  2295=>"010110001",
  2296=>"111000000",
  2297=>"000000000",
  2298=>"111111111",
  2299=>"000000111",
  2300=>"000000001",
  2301=>"001001000",
  2302=>"111000000",
  2303=>"111111111",
  2304=>"101101111",
  2305=>"011011011",
  2306=>"100110100",
  2307=>"111111111",
  2308=>"000000100",
  2309=>"000000011",
  2310=>"000010111",
  2311=>"101101001",
  2312=>"111111011",
  2313=>"000000000",
  2314=>"111111111",
  2315=>"001001111",
  2316=>"111100100",
  2317=>"111111111",
  2318=>"000000000",
  2319=>"010111000",
  2320=>"000011111",
  2321=>"000000000",
  2322=>"000000000",
  2323=>"010110111",
  2324=>"111111111",
  2325=>"000000000",
  2326=>"110110111",
  2327=>"000010011",
  2328=>"000000001",
  2329=>"000000000",
  2330=>"110100111",
  2331=>"000000110",
  2332=>"011011011",
  2333=>"111010111",
  2334=>"000000001",
  2335=>"110110111",
  2336=>"111111111",
  2337=>"000001011",
  2338=>"110111111",
  2339=>"101000110",
  2340=>"100110100",
  2341=>"110001101",
  2342=>"000001011",
  2343=>"001111101",
  2344=>"110110000",
  2345=>"010000000",
  2346=>"111111111",
  2347=>"111111111",
  2348=>"001011000",
  2349=>"111111101",
  2350=>"111000111",
  2351=>"000000000",
  2352=>"100000000",
  2353=>"010010111",
  2354=>"000000001",
  2355=>"000010011",
  2356=>"111111111",
  2357=>"000100110",
  2358=>"111111111",
  2359=>"000000000",
  2360=>"000000001",
  2361=>"000000000",
  2362=>"010010000",
  2363=>"111111011",
  2364=>"001000001",
  2365=>"100100000",
  2366=>"111111001",
  2367=>"111111001",
  2368=>"000000000",
  2369=>"000000000",
  2370=>"100100001",
  2371=>"000111111",
  2372=>"000110111",
  2373=>"000001000",
  2374=>"100111111",
  2375=>"100000001",
  2376=>"000000000",
  2377=>"000000001",
  2378=>"000000011",
  2379=>"111110000",
  2380=>"000101101",
  2381=>"000100100",
  2382=>"111100101",
  2383=>"000010000",
  2384=>"000000000",
  2385=>"111110110",
  2386=>"011110000",
  2387=>"110110000",
  2388=>"111111111",
  2389=>"011011011",
  2390=>"000000000",
  2391=>"000000111",
  2392=>"101111111",
  2393=>"001111111",
  2394=>"000000000",
  2395=>"110000000",
  2396=>"000000000",
  2397=>"100100111",
  2398=>"000000000",
  2399=>"001111111",
  2400=>"100000000",
  2401=>"000000000",
  2402=>"000110100",
  2403=>"111111111",
  2404=>"000000000",
  2405=>"000000000",
  2406=>"000011111",
  2407=>"000000000",
  2408=>"011011000",
  2409=>"111111111",
  2410=>"111111000",
  2411=>"111111011",
  2412=>"111001011",
  2413=>"111000000",
  2414=>"011111000",
  2415=>"000000000",
  2416=>"000000111",
  2417=>"111111111",
  2418=>"110110111",
  2419=>"010000100",
  2420=>"000000000",
  2421=>"011010110",
  2422=>"111111110",
  2423=>"011111111",
  2424=>"000000000",
  2425=>"111111111",
  2426=>"100111111",
  2427=>"111111000",
  2428=>"000000000",
  2429=>"000000000",
  2430=>"000000000",
  2431=>"001001111",
  2432=>"000100000",
  2433=>"110100000",
  2434=>"110100001",
  2435=>"000000000",
  2436=>"000000000",
  2437=>"111111111",
  2438=>"000000000",
  2439=>"100111111",
  2440=>"000000000",
  2441=>"000000000",
  2442=>"111111101",
  2443=>"000000000",
  2444=>"000000000",
  2445=>"010011111",
  2446=>"100100110",
  2447=>"010010000",
  2448=>"111111111",
  2449=>"111000000",
  2450=>"000000000",
  2451=>"110100100",
  2452=>"111111111",
  2453=>"010000000",
  2454=>"001000000",
  2455=>"101111011",
  2456=>"100100000",
  2457=>"000000111",
  2458=>"101101101",
  2459=>"101000010",
  2460=>"111111000",
  2461=>"000000000",
  2462=>"000000000",
  2463=>"000000110",
  2464=>"000110100",
  2465=>"110011000",
  2466=>"010010000",
  2467=>"101111111",
  2468=>"111111111",
  2469=>"010011010",
  2470=>"111111000",
  2471=>"000000101",
  2472=>"000000011",
  2473=>"000000111",
  2474=>"111111111",
  2475=>"111111111",
  2476=>"000000000",
  2477=>"110111111",
  2478=>"110000000",
  2479=>"000000000",
  2480=>"111111111",
  2481=>"000000000",
  2482=>"101111111",
  2483=>"111101101",
  2484=>"100000000",
  2485=>"101111111",
  2486=>"111111111",
  2487=>"001111111",
  2488=>"000100101",
  2489=>"111111101",
  2490=>"000000110",
  2491=>"111111111",
  2492=>"011001000",
  2493=>"000000000",
  2494=>"111111111",
  2495=>"101001000",
  2496=>"110111111",
  2497=>"000000111",
  2498=>"111111111",
  2499=>"111111110",
  2500=>"111111111",
  2501=>"110110000",
  2502=>"000000000",
  2503=>"001000000",
  2504=>"000000000",
  2505=>"111111000",
  2506=>"110000100",
  2507=>"111100000",
  2508=>"100000000",
  2509=>"111111011",
  2510=>"100100100",
  2511=>"000100000",
  2512=>"100111111",
  2513=>"011011001",
  2514=>"111111111",
  2515=>"000010110",
  2516=>"111111110",
  2517=>"000000000",
  2518=>"000101101",
  2519=>"000100100",
  2520=>"100000100",
  2521=>"101101000",
  2522=>"000000000",
  2523=>"000000000",
  2524=>"000000000",
  2525=>"110110111",
  2526=>"001100110",
  2527=>"011011011",
  2528=>"111100111",
  2529=>"000000000",
  2530=>"111111111",
  2531=>"111111111",
  2532=>"111101001",
  2533=>"111111000",
  2534=>"000110111",
  2535=>"111111111",
  2536=>"100111111",
  2537=>"100100100",
  2538=>"111111111",
  2539=>"000000000",
  2540=>"000011111",
  2541=>"111010110",
  2542=>"000000000",
  2543=>"111111110",
  2544=>"000000000",
  2545=>"000000000",
  2546=>"111111111",
  2547=>"000010000",
  2548=>"111111111",
  2549=>"111011111",
  2550=>"000000000",
  2551=>"000000000",
  2552=>"000000100",
  2553=>"100100100",
  2554=>"111111111",
  2555=>"000000001",
  2556=>"001000000",
  2557=>"110111111",
  2558=>"111100000",
  2559=>"000000000",
  2560=>"000000000",
  2561=>"000000000",
  2562=>"000000111",
  2563=>"000011111",
  2564=>"101001000",
  2565=>"111001000",
  2566=>"000000000",
  2567=>"000000110",
  2568=>"111000000",
  2569=>"001111011",
  2570=>"110110000",
  2571=>"111110000",
  2572=>"000100100",
  2573=>"000000000",
  2574=>"111111011",
  2575=>"000000000",
  2576=>"111011011",
  2577=>"110111111",
  2578=>"111111011",
  2579=>"000000110",
  2580=>"000000000",
  2581=>"110111111",
  2582=>"010000000",
  2583=>"111111000",
  2584=>"100100000",
  2585=>"110111100",
  2586=>"000000000",
  2587=>"000000111",
  2588=>"010111111",
  2589=>"111111111",
  2590=>"111111111",
  2591=>"000000000",
  2592=>"000000000",
  2593=>"111111110",
  2594=>"000000000",
  2595=>"111011000",
  2596=>"000000000",
  2597=>"001000000",
  2598=>"111111111",
  2599=>"111111110",
  2600=>"111111101",
  2601=>"000000000",
  2602=>"000000000",
  2603=>"111110000",
  2604=>"111111000",
  2605=>"111111011",
  2606=>"000000000",
  2607=>"000100110",
  2608=>"000111110",
  2609=>"000000000",
  2610=>"000000000",
  2611=>"000000101",
  2612=>"000001000",
  2613=>"010000000",
  2614=>"100111111",
  2615=>"011000111",
  2616=>"000000011",
  2617=>"001000000",
  2618=>"111111100",
  2619=>"111111000",
  2620=>"100100001",
  2621=>"111111111",
  2622=>"101000000",
  2623=>"000000000",
  2624=>"000000000",
  2625=>"000000000",
  2626=>"111111011",
  2627=>"111111111",
  2628=>"000100000",
  2629=>"000000001",
  2630=>"001000000",
  2631=>"000000000",
  2632=>"000001001",
  2633=>"100001111",
  2634=>"011111110",
  2635=>"100100000",
  2636=>"000001000",
  2637=>"111111011",
  2638=>"111111111",
  2639=>"001110100",
  2640=>"001000000",
  2641=>"111001001",
  2642=>"000000110",
  2643=>"100001101",
  2644=>"000000000",
  2645=>"000000101",
  2646=>"111111111",
  2647=>"000000000",
  2648=>"111111111",
  2649=>"111111111",
  2650=>"111111000",
  2651=>"111111011",
  2652=>"000100100",
  2653=>"111111111",
  2654=>"111111000",
  2655=>"000000000",
  2656=>"111111111",
  2657=>"111000001",
  2658=>"101000000",
  2659=>"000000001",
  2660=>"111101111",
  2661=>"000000000",
  2662=>"110100111",
  2663=>"000100100",
  2664=>"111111111",
  2665=>"111111111",
  2666=>"000000000",
  2667=>"111000000",
  2668=>"111001001",
  2669=>"000000000",
  2670=>"111001000",
  2671=>"001101001",
  2672=>"000000000",
  2673=>"111111111",
  2674=>"111111011",
  2675=>"100000000",
  2676=>"000000000",
  2677=>"000000000",
  2678=>"111001001",
  2679=>"000000000",
  2680=>"000000000",
  2681=>"000000000",
  2682=>"000000000",
  2683=>"000000011",
  2684=>"100100101",
  2685=>"000000000",
  2686=>"000000000",
  2687=>"011011011",
  2688=>"000001111",
  2689=>"101001000",
  2690=>"111111100",
  2691=>"000111111",
  2692=>"001111111",
  2693=>"111000000",
  2694=>"111111111",
  2695=>"111111000",
  2696=>"000000000",
  2697=>"001001000",
  2698=>"111111000",
  2699=>"010111111",
  2700=>"111111100",
  2701=>"111000111",
  2702=>"111110110",
  2703=>"100100000",
  2704=>"000000000",
  2705=>"111111010",
  2706=>"000010110",
  2707=>"110111111",
  2708=>"000000000",
  2709=>"011000000",
  2710=>"111111111",
  2711=>"000000000",
  2712=>"101001101",
  2713=>"000000000",
  2714=>"010111111",
  2715=>"000000010",
  2716=>"011000010",
  2717=>"000000000",
  2718=>"110000000",
  2719=>"000100111",
  2720=>"000000000",
  2721=>"000000000",
  2722=>"000000000",
  2723=>"111111010",
  2724=>"000001001",
  2725=>"001000000",
  2726=>"000000000",
  2727=>"000000000",
  2728=>"000000000",
  2729=>"000000000",
  2730=>"000111111",
  2731=>"001000000",
  2732=>"000000000",
  2733=>"100100111",
  2734=>"000000000",
  2735=>"000000000",
  2736=>"000000101",
  2737=>"110110100",
  2738=>"000110110",
  2739=>"111000000",
  2740=>"001001111",
  2741=>"001001111",
  2742=>"001000000",
  2743=>"000000000",
  2744=>"100000101",
  2745=>"000101111",
  2746=>"000000000",
  2747=>"111011000",
  2748=>"111111110",
  2749=>"111111111",
  2750=>"000000000",
  2751=>"111011001",
  2752=>"111111010",
  2753=>"110110011",
  2754=>"111111101",
  2755=>"111001001",
  2756=>"011000000",
  2757=>"000000000",
  2758=>"111011000",
  2759=>"001000000",
  2760=>"111111111",
  2761=>"000000101",
  2762=>"111111100",
  2763=>"011000000",
  2764=>"100100110",
  2765=>"001010110",
  2766=>"111111110",
  2767=>"000101111",
  2768=>"111110111",
  2769=>"111111111",
  2770=>"001111110",
  2771=>"000100111",
  2772=>"111111111",
  2773=>"000000010",
  2774=>"000000111",
  2775=>"111101101",
  2776=>"111000001",
  2777=>"111111101",
  2778=>"100000000",
  2779=>"000110111",
  2780=>"111111100",
  2781=>"100100111",
  2782=>"111110000",
  2783=>"011000111",
  2784=>"111111111",
  2785=>"000000000",
  2786=>"111010000",
  2787=>"011000000",
  2788=>"010000000",
  2789=>"111110110",
  2790=>"111111000",
  2791=>"000000000",
  2792=>"100111111",
  2793=>"000001111",
  2794=>"000000000",
  2795=>"000000000",
  2796=>"000011000",
  2797=>"100000111",
  2798=>"101111111",
  2799=>"010000000",
  2800=>"001111001",
  2801=>"111111111",
  2802=>"111100000",
  2803=>"001001001",
  2804=>"011011111",
  2805=>"000000000",
  2806=>"011010000",
  2807=>"110100100",
  2808=>"111000100",
  2809=>"111111010",
  2810=>"111111101",
  2811=>"111111111",
  2812=>"000000000",
  2813=>"110111011",
  2814=>"000000000",
  2815=>"000000000",
  2816=>"000000000",
  2817=>"011011011",
  2818=>"000000111",
  2819=>"110110000",
  2820=>"000001001",
  2821=>"000000000",
  2822=>"000000000",
  2823=>"001111111",
  2824=>"110110011",
  2825=>"111111111",
  2826=>"110111110",
  2827=>"111111111",
  2828=>"111110000",
  2829=>"111111111",
  2830=>"001001000",
  2831=>"111000000",
  2832=>"000000000",
  2833=>"101111111",
  2834=>"111001111",
  2835=>"101111111",
  2836=>"000000000",
  2837=>"011110110",
  2838=>"110101110",
  2839=>"111111111",
  2840=>"000000001",
  2841=>"000000111",
  2842=>"111101111",
  2843=>"011010111",
  2844=>"000100000",
  2845=>"111111111",
  2846=>"001010000",
  2847=>"001000000",
  2848=>"111110111",
  2849=>"000000000",
  2850=>"110110111",
  2851=>"011111111",
  2852=>"111101111",
  2853=>"000000000",
  2854=>"000000001",
  2855=>"001000000",
  2856=>"000000000",
  2857=>"000010010",
  2858=>"111100000",
  2859=>"011011001",
  2860=>"111001001",
  2861=>"110100000",
  2862=>"111111111",
  2863=>"100000101",
  2864=>"001000001",
  2865=>"111111111",
  2866=>"000000001",
  2867=>"110000010",
  2868=>"000111111",
  2869=>"111000000",
  2870=>"111111111",
  2871=>"011110101",
  2872=>"111111111",
  2873=>"111000011",
  2874=>"111111111",
  2875=>"111111111",
  2876=>"111110100",
  2877=>"000000000",
  2878=>"001111111",
  2879=>"001000000",
  2880=>"000000000",
  2881=>"100011000",
  2882=>"000000011",
  2883=>"111111111",
  2884=>"111111000",
  2885=>"111111100",
  2886=>"000000111",
  2887=>"001000000",
  2888=>"100100100",
  2889=>"111111110",
  2890=>"110000100",
  2891=>"111110011",
  2892=>"111111111",
  2893=>"101000111",
  2894=>"111101111",
  2895=>"111111111",
  2896=>"011001001",
  2897=>"000000111",
  2898=>"111111000",
  2899=>"000011111",
  2900=>"000000000",
  2901=>"000010011",
  2902=>"111111000",
  2903=>"110000111",
  2904=>"000000000",
  2905=>"111111111",
  2906=>"111111000",
  2907=>"000000001",
  2908=>"000010011",
  2909=>"000100100",
  2910=>"101000111",
  2911=>"000000000",
  2912=>"111111111",
  2913=>"111000000",
  2914=>"011001001",
  2915=>"111111111",
  2916=>"110100100",
  2917=>"011000000",
  2918=>"111000000",
  2919=>"111111111",
  2920=>"111111111",
  2921=>"110100000",
  2922=>"000000000",
  2923=>"111111111",
  2924=>"110111011",
  2925=>"000000000",
  2926=>"000000000",
  2927=>"111111000",
  2928=>"011000000",
  2929=>"000111111",
  2930=>"000011111",
  2931=>"000110111",
  2932=>"111111111",
  2933=>"111111111",
  2934=>"000000000",
  2935=>"111111001",
  2936=>"111111111",
  2937=>"000000000",
  2938=>"000111111",
  2939=>"000000000",
  2940=>"111100111",
  2941=>"000000110",
  2942=>"111111111",
  2943=>"111111111",
  2944=>"110110111",
  2945=>"000000100",
  2946=>"011110110",
  2947=>"111011000",
  2948=>"000001111",
  2949=>"000011110",
  2950=>"011100000",
  2951=>"110111111",
  2952=>"001110110",
  2953=>"100000000",
  2954=>"110000000",
  2955=>"111110110",
  2956=>"111111111",
  2957=>"001000111",
  2958=>"000000000",
  2959=>"110111111",
  2960=>"001100000",
  2961=>"111111000",
  2962=>"111111111",
  2963=>"111111001",
  2964=>"000000000",
  2965=>"011011010",
  2966=>"011000000",
  2967=>"110110000",
  2968=>"101001011",
  2969=>"000000100",
  2970=>"111111111",
  2971=>"100110111",
  2972=>"000100100",
  2973=>"000010111",
  2974=>"000000000",
  2975=>"000000000",
  2976=>"111101001",
  2977=>"001001000",
  2978=>"000000000",
  2979=>"111101001",
  2980=>"100111111",
  2981=>"111111111",
  2982=>"000000000",
  2983=>"111100100",
  2984=>"000000100",
  2985=>"111110011",
  2986=>"000001111",
  2987=>"011111000",
  2988=>"000000000",
  2989=>"000000000",
  2990=>"000000000",
  2991=>"111111111",
  2992=>"000000000",
  2993=>"000100000",
  2994=>"111000000",
  2995=>"000000110",
  2996=>"011111111",
  2997=>"111111011",
  2998=>"100101101",
  2999=>"000000000",
  3000=>"001000110",
  3001=>"010000000",
  3002=>"000000100",
  3003=>"010000000",
  3004=>"000000011",
  3005=>"000000000",
  3006=>"001001000",
  3007=>"001011000",
  3008=>"111100000",
  3009=>"001000000",
  3010=>"001001000",
  3011=>"000000000",
  3012=>"000000111",
  3013=>"011010111",
  3014=>"001001000",
  3015=>"111111111",
  3016=>"101000000",
  3017=>"011011001",
  3018=>"001000000",
  3019=>"100100000",
  3020=>"110110111",
  3021=>"000000000",
  3022=>"011000000",
  3023=>"111010111",
  3024=>"000000111",
  3025=>"010010000",
  3026=>"101101100",
  3027=>"000000001",
  3028=>"100000000",
  3029=>"111111100",
  3030=>"111111111",
  3031=>"001011011",
  3032=>"000000000",
  3033=>"111000000",
  3034=>"100100100",
  3035=>"000000000",
  3036=>"011000000",
  3037=>"011011000",
  3038=>"100110000",
  3039=>"000000001",
  3040=>"000111111",
  3041=>"100000000",
  3042=>"000000011",
  3043=>"001001000",
  3044=>"000110111",
  3045=>"001111111",
  3046=>"111001001",
  3047=>"111111111",
  3048=>"111111110",
  3049=>"011011011",
  3050=>"000000011",
  3051=>"010010000",
  3052=>"000000000",
  3053=>"000100011",
  3054=>"001111011",
  3055=>"000000111",
  3056=>"000000000",
  3057=>"000000000",
  3058=>"000000000",
  3059=>"001000000",
  3060=>"111111100",
  3061=>"000000000",
  3062=>"000000000",
  3063=>"000000000",
  3064=>"000000000",
  3065=>"001001111",
  3066=>"111111111",
  3067=>"111111111",
  3068=>"000000000",
  3069=>"000100000",
  3070=>"000000000",
  3071=>"000000100",
  3072=>"110111111",
  3073=>"000000000",
  3074=>"000000000",
  3075=>"111111111",
  3076=>"111111000",
  3077=>"000000000",
  3078=>"111000101",
  3079=>"111111111",
  3080=>"000001111",
  3081=>"111111000",
  3082=>"001000000",
  3083=>"000000001",
  3084=>"111111111",
  3085=>"111111111",
  3086=>"010101111",
  3087=>"001111011",
  3088=>"111100000",
  3089=>"000000001",
  3090=>"111101111",
  3091=>"111111001",
  3092=>"111111000",
  3093=>"111111000",
  3094=>"011000000",
  3095=>"111111001",
  3096=>"100011100",
  3097=>"001001000",
  3098=>"110111111",
  3099=>"000000011",
  3100=>"111100100",
  3101=>"000100111",
  3102=>"011111111",
  3103=>"000000001",
  3104=>"000001001",
  3105=>"111110111",
  3106=>"111111110",
  3107=>"110111111",
  3108=>"000011111",
  3109=>"000000000",
  3110=>"111110000",
  3111=>"111100000",
  3112=>"111111111",
  3113=>"110111000",
  3114=>"001000000",
  3115=>"101111000",
  3116=>"001000000",
  3117=>"110000000",
  3118=>"111100000",
  3119=>"000111110",
  3120=>"000000000",
  3121=>"000000001",
  3122=>"001100100",
  3123=>"110111101",
  3124=>"110000000",
  3125=>"111011000",
  3126=>"000000111",
  3127=>"000101001",
  3128=>"001101001",
  3129=>"001000111",
  3130=>"000000100",
  3131=>"000110111",
  3132=>"000100111",
  3133=>"000000101",
  3134=>"000000000",
  3135=>"000000000",
  3136=>"101100111",
  3137=>"100001011",
  3138=>"000000001",
  3139=>"111111100",
  3140=>"000000000",
  3141=>"101001000",
  3142=>"111111010",
  3143=>"111111111",
  3144=>"000100110",
  3145=>"000000111",
  3146=>"010111111",
  3147=>"000000000",
  3148=>"111111100",
  3149=>"000000111",
  3150=>"011000000",
  3151=>"000010111",
  3152=>"000000010",
  3153=>"101000000",
  3154=>"000111111",
  3155=>"000001011",
  3156=>"000000101",
  3157=>"000000111",
  3158=>"111001000",
  3159=>"000000000",
  3160=>"000010000",
  3161=>"000000010",
  3162=>"000011000",
  3163=>"001000000",
  3164=>"101111100",
  3165=>"011001000",
  3166=>"110111000",
  3167=>"010000110",
  3168=>"111110000",
  3169=>"111111100",
  3170=>"011111111",
  3171=>"111111110",
  3172=>"000111000",
  3173=>"000000111",
  3174=>"111000011",
  3175=>"100000111",
  3176=>"000000000",
  3177=>"111010010",
  3178=>"111011000",
  3179=>"000000111",
  3180=>"000001000",
  3181=>"000001111",
  3182=>"000000111",
  3183=>"111000000",
  3184=>"111000000",
  3185=>"000000111",
  3186=>"010111111",
  3187=>"111111111",
  3188=>"000000100",
  3189=>"011011000",
  3190=>"101000000",
  3191=>"000000000",
  3192=>"000000000",
  3193=>"110111111",
  3194=>"111111101",
  3195=>"001001000",
  3196=>"111011001",
  3197=>"111111011",
  3198=>"111100110",
  3199=>"111111000",
  3200=>"000001000",
  3201=>"000101111",
  3202=>"110000011",
  3203=>"000110111",
  3204=>"110110111",
  3205=>"000000000",
  3206=>"000000110",
  3207=>"111111100",
  3208=>"010111111",
  3209=>"111111000",
  3210=>"100111111",
  3211=>"000110110",
  3212=>"000000111",
  3213=>"111000010",
  3214=>"100000110",
  3215=>"000000110",
  3216=>"111111111",
  3217=>"000010010",
  3218=>"000000000",
  3219=>"000000000",
  3220=>"100000000",
  3221=>"000111111",
  3222=>"111100010",
  3223=>"000111000",
  3224=>"000000100",
  3225=>"111111110",
  3226=>"000000111",
  3227=>"000000000",
  3228=>"111111101",
  3229=>"101100000",
  3230=>"000000001",
  3231=>"000000001",
  3232=>"111111000",
  3233=>"000000110",
  3234=>"000000111",
  3235=>"000111111",
  3236=>"110110000",
  3237=>"111111111",
  3238=>"110111010",
  3239=>"001000000",
  3240=>"000000000",
  3241=>"111001001",
  3242=>"000000000",
  3243=>"000000000",
  3244=>"011000000",
  3245=>"000000010",
  3246=>"110111000",
  3247=>"111111111",
  3248=>"111111000",
  3249=>"111111110",
  3250=>"111111111",
  3251=>"010000000",
  3252=>"111110000",
  3253=>"000000100",
  3254=>"000000000",
  3255=>"001111111",
  3256=>"111101111",
  3257=>"000000111",
  3258=>"000110111",
  3259=>"011100111",
  3260=>"111111111",
  3261=>"000000000",
  3262=>"100100111",
  3263=>"111111111",
  3264=>"001010111",
  3265=>"111010100",
  3266=>"000010011",
  3267=>"000000000",
  3268=>"000000000",
  3269=>"111111000",
  3270=>"000111111",
  3271=>"000001001",
  3272=>"010011000",
  3273=>"000000101",
  3274=>"011111111",
  3275=>"111000000",
  3276=>"111000000",
  3277=>"111111111",
  3278=>"000000000",
  3279=>"000100101",
  3280=>"000000000",
  3281=>"011111110",
  3282=>"000111000",
  3283=>"111111111",
  3284=>"001000000",
  3285=>"111100000",
  3286=>"010000000",
  3287=>"000111111",
  3288=>"111111000",
  3289=>"000110000",
  3290=>"011001000",
  3291=>"111000000",
  3292=>"000000000",
  3293=>"110000000",
  3294=>"010111111",
  3295=>"000111111",
  3296=>"010000000",
  3297=>"000000111",
  3298=>"110111111",
  3299=>"000000000",
  3300=>"111100000",
  3301=>"001000100",
  3302=>"111111111",
  3303=>"111111111",
  3304=>"001111111",
  3305=>"111101000",
  3306=>"111111000",
  3307=>"000000011",
  3308=>"111000000",
  3309=>"000010011",
  3310=>"110001111",
  3311=>"111000000",
  3312=>"111111000",
  3313=>"000111111",
  3314=>"111111000",
  3315=>"000010101",
  3316=>"001000001",
  3317=>"000001001",
  3318=>"000110000",
  3319=>"111000101",
  3320=>"111000111",
  3321=>"000000011",
  3322=>"001000110",
  3323=>"101001111",
  3324=>"110100100",
  3325=>"001001001",
  3326=>"111111111",
  3327=>"000011000",
  3328=>"001111111",
  3329=>"100110110",
  3330=>"111111111",
  3331=>"001101000",
  3332=>"000000111",
  3333=>"000001000",
  3334=>"000000000",
  3335=>"000000000",
  3336=>"111111111",
  3337=>"000000001",
  3338=>"000101101",
  3339=>"011011111",
  3340=>"111111111",
  3341=>"000000000",
  3342=>"000000000",
  3343=>"100111111",
  3344=>"101001101",
  3345=>"011111111",
  3346=>"000000001",
  3347=>"000111111",
  3348=>"001011000",
  3349=>"110000000",
  3350=>"010000111",
  3351=>"000000101",
  3352=>"111111001",
  3353=>"101111000",
  3354=>"111111111",
  3355=>"110111000",
  3356=>"011111111",
  3357=>"111000000",
  3358=>"000000000",
  3359=>"000000000",
  3360=>"010110000",
  3361=>"110110000",
  3362=>"111111111",
  3363=>"000001111",
  3364=>"111111111",
  3365=>"111010001",
  3366=>"000000000",
  3367=>"110100111",
  3368=>"111111000",
  3369=>"110100111",
  3370=>"000110111",
  3371=>"000111110",
  3372=>"110110000",
  3373=>"110111001",
  3374=>"000000000",
  3375=>"000000000",
  3376=>"011011111",
  3377=>"111110000",
  3378=>"111101000",
  3379=>"111000000",
  3380=>"100000000",
  3381=>"111111111",
  3382=>"010000001",
  3383=>"111001001",
  3384=>"010000000",
  3385=>"000000111",
  3386=>"111100101",
  3387=>"110100100",
  3388=>"011111111",
  3389=>"000001000",
  3390=>"111111111",
  3391=>"111111000",
  3392=>"011000000",
  3393=>"111111001",
  3394=>"000000111",
  3395=>"000100101",
  3396=>"000000111",
  3397=>"000010111",
  3398=>"000101111",
  3399=>"110100111",
  3400=>"111000010",
  3401=>"111111000",
  3402=>"000011000",
  3403=>"110100001",
  3404=>"001111111",
  3405=>"000001111",
  3406=>"000000100",
  3407=>"110111111",
  3408=>"111100110",
  3409=>"000111000",
  3410=>"000000111",
  3411=>"111000000",
  3412=>"110110111",
  3413=>"111001001",
  3414=>"000000000",
  3415=>"111000000",
  3416=>"111000011",
  3417=>"100000011",
  3418=>"000111111",
  3419=>"111000111",
  3420=>"000000000",
  3421=>"011111111",
  3422=>"111111000",
  3423=>"000111111",
  3424=>"001000111",
  3425=>"000111111",
  3426=>"110110111",
  3427=>"000000000",
  3428=>"110110110",
  3429=>"000000100",
  3430=>"111110000",
  3431=>"000000111",
  3432=>"111111110",
  3433=>"000000001",
  3434=>"111111000",
  3435=>"111110101",
  3436=>"010010011",
  3437=>"011000000",
  3438=>"000000000",
  3439=>"001111111",
  3440=>"000000000",
  3441=>"111111011",
  3442=>"111000111",
  3443=>"101111100",
  3444=>"000110111",
  3445=>"000000000",
  3446=>"001111111",
  3447=>"000000000",
  3448=>"011111011",
  3449=>"000000011",
  3450=>"001000000",
  3451=>"111101000",
  3452=>"001000111",
  3453=>"111111000",
  3454=>"000001000",
  3455=>"011111111",
  3456=>"111011010",
  3457=>"111000000",
  3458=>"111000000",
  3459=>"100000111",
  3460=>"111111111",
  3461=>"111111111",
  3462=>"111111000",
  3463=>"010011010",
  3464=>"000011000",
  3465=>"000001111",
  3466=>"011000000",
  3467=>"001111000",
  3468=>"111001111",
  3469=>"111110100",
  3470=>"000001101",
  3471=>"110110010",
  3472=>"011011111",
  3473=>"000100000",
  3474=>"000110100",
  3475=>"100110011",
  3476=>"111111111",
  3477=>"111101000",
  3478=>"111111111",
  3479=>"111111110",
  3480=>"000000100",
  3481=>"111000111",
  3482=>"011001001",
  3483=>"011011011",
  3484=>"000101101",
  3485=>"110000000",
  3486=>"011011111",
  3487=>"000000000",
  3488=>"010000000",
  3489=>"111111100",
  3490=>"000100001",
  3491=>"000111111",
  3492=>"001000000",
  3493=>"000000000",
  3494=>"000000000",
  3495=>"011011001",
  3496=>"111110011",
  3497=>"111111111",
  3498=>"111111111",
  3499=>"000000100",
  3500=>"000100111",
  3501=>"000000000",
  3502=>"000000001",
  3503=>"111111111",
  3504=>"111111000",
  3505=>"111000000",
  3506=>"110110111",
  3507=>"000000011",
  3508=>"111111111",
  3509=>"111111111",
  3510=>"011111111",
  3511=>"000000000",
  3512=>"111000000",
  3513=>"110000000",
  3514=>"111111111",
  3515=>"101111000",
  3516=>"000000000",
  3517=>"000000100",
  3518=>"111111100",
  3519=>"000011111",
  3520=>"111111010",
  3521=>"010010000",
  3522=>"010111111",
  3523=>"110111110",
  3524=>"111111111",
  3525=>"011001000",
  3526=>"000000001",
  3527=>"000011111",
  3528=>"111110111",
  3529=>"000111111",
  3530=>"000000000",
  3531=>"111110000",
  3532=>"001000000",
  3533=>"000111111",
  3534=>"110111111",
  3535=>"111111011",
  3536=>"111110000",
  3537=>"001011011",
  3538=>"110111111",
  3539=>"111000111",
  3540=>"000110111",
  3541=>"111000000",
  3542=>"000000000",
  3543=>"000000011",
  3544=>"111111000",
  3545=>"011000000",
  3546=>"111111111",
  3547=>"000000111",
  3548=>"000000001",
  3549=>"000000011",
  3550=>"000000000",
  3551=>"111111111",
  3552=>"000010010",
  3553=>"000000111",
  3554=>"000000000",
  3555=>"000010111",
  3556=>"110110100",
  3557=>"111001011",
  3558=>"000000010",
  3559=>"111111000",
  3560=>"110111001",
  3561=>"000000111",
  3562=>"000011011",
  3563=>"000000000",
  3564=>"011011000",
  3565=>"000100000",
  3566=>"110111110",
  3567=>"000000100",
  3568=>"000000000",
  3569=>"001000000",
  3570=>"001111111",
  3571=>"010011010",
  3572=>"000001101",
  3573=>"111011000",
  3574=>"111111110",
  3575=>"000011111",
  3576=>"001010111",
  3577=>"001001001",
  3578=>"000000000",
  3579=>"110000000",
  3580=>"000111000",
  3581=>"011111111",
  3582=>"000000011",
  3583=>"111111111",
  3584=>"111110111",
  3585=>"000001000",
  3586=>"000000000",
  3587=>"000000000",
  3588=>"111111111",
  3589=>"000100000",
  3590=>"000000000",
  3591=>"111000000",
  3592=>"000000000",
  3593=>"000110110",
  3594=>"001111110",
  3595=>"000010010",
  3596=>"100000000",
  3597=>"001000000",
  3598=>"001001111",
  3599=>"001101111",
  3600=>"000000000",
  3601=>"000000000",
  3602=>"001001111",
  3603=>"101000001",
  3604=>"011011111",
  3605=>"000000000",
  3606=>"110111111",
  3607=>"001000000",
  3608=>"111011001",
  3609=>"100000000",
  3610=>"000000010",
  3611=>"000111011",
  3612=>"111011111",
  3613=>"000011100",
  3614=>"111111111",
  3615=>"111111111",
  3616=>"111111111",
  3617=>"111111111",
  3618=>"000000000",
  3619=>"111110111",
  3620=>"111111111",
  3621=>"000000001",
  3622=>"111111111",
  3623=>"000000000",
  3624=>"000000000",
  3625=>"000000000",
  3626=>"111111111",
  3627=>"110110111",
  3628=>"111111111",
  3629=>"111100100",
  3630=>"000000000",
  3631=>"000000010",
  3632=>"111111111",
  3633=>"111111111",
  3634=>"001000000",
  3635=>"010110000",
  3636=>"111111001",
  3637=>"001011110",
  3638=>"000000000",
  3639=>"111111111",
  3640=>"000100111",
  3641=>"010000000",
  3642=>"000000000",
  3643=>"001100000",
  3644=>"111001111",
  3645=>"111100101",
  3646=>"111111111",
  3647=>"000000000",
  3648=>"000110111",
  3649=>"000000001",
  3650=>"000000000",
  3651=>"110111111",
  3652=>"010010000",
  3653=>"100111111",
  3654=>"000101100",
  3655=>"000000000",
  3656=>"100100100",
  3657=>"111111111",
  3658=>"000001011",
  3659=>"100100111",
  3660=>"001001110",
  3661=>"111100100",
  3662=>"111110000",
  3663=>"000000000",
  3664=>"100100000",
  3665=>"000000000",
  3666=>"000001001",
  3667=>"001011111",
  3668=>"111101101",
  3669=>"000000111",
  3670=>"100000110",
  3671=>"100100110",
  3672=>"011011111",
  3673=>"101001111",
  3674=>"000000100",
  3675=>"110011001",
  3676=>"111001001",
  3677=>"111111000",
  3678=>"010000000",
  3679=>"011110110",
  3680=>"111001001",
  3681=>"111111100",
  3682=>"011000000",
  3683=>"111111111",
  3684=>"111010000",
  3685=>"011111111",
  3686=>"110110111",
  3687=>"000000000",
  3688=>"111111000",
  3689=>"000110110",
  3690=>"000000000",
  3691=>"010110110",
  3692=>"110110100",
  3693=>"111111111",
  3694=>"000000100",
  3695=>"110110100",
  3696=>"011000111",
  3697=>"000000000",
  3698=>"011011111",
  3699=>"011111111",
  3700=>"111101100",
  3701=>"000000000",
  3702=>"111000000",
  3703=>"111101000",
  3704=>"111111111",
  3705=>"011111111",
  3706=>"000000011",
  3707=>"101100101",
  3708=>"011011010",
  3709=>"000000000",
  3710=>"000000000",
  3711=>"111111111",
  3712=>"111111111",
  3713=>"111111110",
  3714=>"100100100",
  3715=>"111111111",
  3716=>"110000100",
  3717=>"011101101",
  3718=>"101000000",
  3719=>"000000000",
  3720=>"011000000",
  3721=>"000000000",
  3722=>"000000000",
  3723=>"000000000",
  3724=>"000000000",
  3725=>"110111000",
  3726=>"000001000",
  3727=>"111101000",
  3728=>"000000000",
  3729=>"111111111",
  3730=>"000110111",
  3731=>"111111001",
  3732=>"010000001",
  3733=>"111111111",
  3734=>"111111111",
  3735=>"000000000",
  3736=>"000000000",
  3737=>"111111111",
  3738=>"111110110",
  3739=>"111111111",
  3740=>"100000000",
  3741=>"001000100",
  3742=>"100000000",
  3743=>"111111101",
  3744=>"000000000",
  3745=>"111100000",
  3746=>"111111111",
  3747=>"111111111",
  3748=>"000000000",
  3749=>"111111111",
  3750=>"011010000",
  3751=>"111111110",
  3752=>"111111110",
  3753=>"111111111",
  3754=>"000000000",
  3755=>"111011000",
  3756=>"111111111",
  3757=>"000000001",
  3758=>"100100111",
  3759=>"000001001",
  3760=>"100110111",
  3761=>"111111101",
  3762=>"011000000",
  3763=>"111111111",
  3764=>"111110011",
  3765=>"000001101",
  3766=>"111000000",
  3767=>"000000001",
  3768=>"111111111",
  3769=>"100001100",
  3770=>"000001010",
  3771=>"110000001",
  3772=>"110011111",
  3773=>"111111001",
  3774=>"000101100",
  3775=>"000000001",
  3776=>"001001000",
  3777=>"111000000",
  3778=>"101111110",
  3779=>"000000000",
  3780=>"111000000",
  3781=>"000000000",
  3782=>"111111111",
  3783=>"001111111",
  3784=>"000000000",
  3785=>"111111101",
  3786=>"000000001",
  3787=>"000000100",
  3788=>"111001101",
  3789=>"101000000",
  3790=>"111111111",
  3791=>"100100111",
  3792=>"000000001",
  3793=>"000000000",
  3794=>"111000000",
  3795=>"111000000",
  3796=>"111111111",
  3797=>"011011001",
  3798=>"100100110",
  3799=>"001001000",
  3800=>"011111100",
  3801=>"110000001",
  3802=>"111111111",
  3803=>"011111111",
  3804=>"111111011",
  3805=>"000000011",
  3806=>"001101111",
  3807=>"000000000",
  3808=>"000000000",
  3809=>"000000000",
  3810=>"000000000",
  3811=>"000001111",
  3812=>"111101111",
  3813=>"000000000",
  3814=>"111111111",
  3815=>"110110000",
  3816=>"000000000",
  3817=>"100000110",
  3818=>"000000000",
  3819=>"000000000",
  3820=>"011111110",
  3821=>"000000000",
  3822=>"000000111",
  3823=>"110110110",
  3824=>"001000011",
  3825=>"011100100",
  3826=>"111111111",
  3827=>"000000000",
  3828=>"000000000",
  3829=>"110100100",
  3830=>"000000000",
  3831=>"111000000",
  3832=>"000000000",
  3833=>"000000000",
  3834=>"000000001",
  3835=>"101000000",
  3836=>"011011011",
  3837=>"100000111",
  3838=>"000000000",
  3839=>"111000000",
  3840=>"000000000",
  3841=>"011011011",
  3842=>"111111111",
  3843=>"000001101",
  3844=>"111111111",
  3845=>"111010000",
  3846=>"111111111",
  3847=>"000000111",
  3848=>"111111111",
  3849=>"000000100",
  3850=>"000000000",
  3851=>"111111111",
  3852=>"100110110",
  3853=>"000000111",
  3854=>"000111111",
  3855=>"000000000",
  3856=>"000000000",
  3857=>"001000000",
  3858=>"111000000",
  3859=>"011000000",
  3860=>"111001001",
  3861=>"101111000",
  3862=>"001001001",
  3863=>"111111101",
  3864=>"101111111",
  3865=>"011111111",
  3866=>"111111111",
  3867=>"001000000",
  3868=>"100100111",
  3869=>"000000000",
  3870=>"111111111",
  3871=>"011100100",
  3872=>"000001011",
  3873=>"111111111",
  3874=>"000000000",
  3875=>"111110110",
  3876=>"011000000",
  3877=>"111111111",
  3878=>"110110111",
  3879=>"111000111",
  3880=>"111111111",
  3881=>"111111111",
  3882=>"000100100",
  3883=>"011000000",
  3884=>"001001001",
  3885=>"100100100",
  3886=>"111111000",
  3887=>"010010010",
  3888=>"011001001",
  3889=>"111111111",
  3890=>"111111111",
  3891=>"111000000",
  3892=>"111111000",
  3893=>"111000000",
  3894=>"111111100",
  3895=>"000000000",
  3896=>"110111111",
  3897=>"110100000",
  3898=>"000000100",
  3899=>"111111100",
  3900=>"110100100",
  3901=>"100111110",
  3902=>"000000000",
  3903=>"110000011",
  3904=>"000111111",
  3905=>"111111111",
  3906=>"000000000",
  3907=>"111111100",
  3908=>"000111111",
  3909=>"001111111",
  3910=>"111111111",
  3911=>"100100111",
  3912=>"111000000",
  3913=>"111111111",
  3914=>"001000000",
  3915=>"111011000",
  3916=>"000000000",
  3917=>"000000111",
  3918=>"111000000",
  3919=>"111111111",
  3920=>"111110110",
  3921=>"000000101",
  3922=>"111111000",
  3923=>"000001111",
  3924=>"000000000",
  3925=>"000000100",
  3926=>"110111111",
  3927=>"111101111",
  3928=>"000000000",
  3929=>"000000000",
  3930=>"111111111",
  3931=>"111111111",
  3932=>"000000000",
  3933=>"111111111",
  3934=>"000000000",
  3935=>"000110000",
  3936=>"111111111",
  3937=>"111111111",
  3938=>"111111111",
  3939=>"111011000",
  3940=>"111111100",
  3941=>"001000011",
  3942=>"000000000",
  3943=>"111111111",
  3944=>"010010000",
  3945=>"000000000",
  3946=>"100000111",
  3947=>"010001010",
  3948=>"000000000",
  3949=>"000000000",
  3950=>"000000000",
  3951=>"111111111",
  3952=>"111110111",
  3953=>"110111111",
  3954=>"000111111",
  3955=>"100100110",
  3956=>"000000000",
  3957=>"000001011",
  3958=>"011111111",
  3959=>"000000111",
  3960=>"111111111",
  3961=>"001011110",
  3962=>"111000100",
  3963=>"000000001",
  3964=>"101100100",
  3965=>"110111111",
  3966=>"110000000",
  3967=>"000000001",
  3968=>"000000100",
  3969=>"000000111",
  3970=>"110111111",
  3971=>"111111111",
  3972=>"111110001",
  3973=>"000000110",
  3974=>"111111111",
  3975=>"111110000",
  3976=>"111001010",
  3977=>"000111111",
  3978=>"100111111",
  3979=>"110100110",
  3980=>"111111111",
  3981=>"000100000",
  3982=>"000000111",
  3983=>"000010010",
  3984=>"111111111",
  3985=>"010000000",
  3986=>"100000000",
  3987=>"101000001",
  3988=>"000000010",
  3989=>"111110000",
  3990=>"111011001",
  3991=>"001111111",
  3992=>"110000001",
  3993=>"011011011",
  3994=>"111111111",
  3995=>"000000000",
  3996=>"111111111",
  3997=>"111010111",
  3998=>"000000000",
  3999=>"000000000",
  4000=>"000000110",
  4001=>"000000000",
  4002=>"110110111",
  4003=>"100100111",
  4004=>"000111111",
  4005=>"111111110",
  4006=>"111111000",
  4007=>"100000011",
  4008=>"111111111",
  4009=>"111111011",
  4010=>"000000111",
  4011=>"000000000",
  4012=>"001001001",
  4013=>"110100101",
  4014=>"000001000",
  4015=>"111111111",
  4016=>"000001011",
  4017=>"000011000",
  4018=>"100000001",
  4019=>"111000000",
  4020=>"000111001",
  4021=>"000000001",
  4022=>"111111011",
  4023=>"000000001",
  4024=>"111111011",
  4025=>"100000010",
  4026=>"000000000",
  4027=>"111111111",
  4028=>"111111110",
  4029=>"111111111",
  4030=>"100100000",
  4031=>"001011001",
  4032=>"000000001",
  4033=>"000001111",
  4034=>"000000000",
  4035=>"111111110",
  4036=>"101100111",
  4037=>"000000110",
  4038=>"000001111",
  4039=>"011100100",
  4040=>"010000000",
  4041=>"001111111",
  4042=>"111111111",
  4043=>"000000000",
  4044=>"100001001",
  4045=>"111111111",
  4046=>"000111111",
  4047=>"111111111",
  4048=>"011000000",
  4049=>"000100100",
  4050=>"111111111",
  4051=>"000010000",
  4052=>"001001011",
  4053=>"111101111",
  4054=>"111000000",
  4055=>"011001001",
  4056=>"100001001",
  4057=>"111101111",
  4058=>"000000000",
  4059=>"111000000",
  4060=>"000000000",
  4061=>"000000010",
  4062=>"000110000",
  4063=>"011011111",
  4064=>"111111110",
  4065=>"111111101",
  4066=>"010111111",
  4067=>"111111110",
  4068=>"110110100",
  4069=>"111100100",
  4070=>"001111111",
  4071=>"110111111",
  4072=>"111000001",
  4073=>"111111001",
  4074=>"000000000",
  4075=>"111111111",
  4076=>"000000000",
  4077=>"100111110",
  4078=>"011011000",
  4079=>"000000000",
  4080=>"000000000",
  4081=>"000001111",
  4082=>"101000000",
  4083=>"000011111",
  4084=>"000000000",
  4085=>"111111111",
  4086=>"000111111",
  4087=>"100100000",
  4088=>"000110000",
  4089=>"000110110",
  4090=>"111011000",
  4091=>"000111010",
  4092=>"110000000",
  4093=>"011000011",
  4094=>"110111001",
  4095=>"000000000",
  4096=>"111111101",
  4097=>"000000100",
  4098=>"001001101",
  4099=>"000000000",
  4100=>"000000111",
  4101=>"000101000",
  4102=>"001011011",
  4103=>"111111111",
  4104=>"110111111",
  4105=>"000000000",
  4106=>"000000000",
  4107=>"000000111",
  4108=>"000000110",
  4109=>"000100110",
  4110=>"111000000",
  4111=>"111111111",
  4112=>"111011011",
  4113=>"011111111",
  4114=>"000000000",
  4115=>"111000001",
  4116=>"111111110",
  4117=>"000000100",
  4118=>"111111111",
  4119=>"111111111",
  4120=>"110000000",
  4121=>"011001011",
  4122=>"100000000",
  4123=>"010110110",
  4124=>"000000000",
  4125=>"000111111",
  4126=>"101011011",
  4127=>"000111111",
  4128=>"001001111",
  4129=>"000000000",
  4130=>"000000000",
  4131=>"000000000",
  4132=>"100000001",
  4133=>"001000000",
  4134=>"000100000",
  4135=>"111111111",
  4136=>"000000111",
  4137=>"100000000",
  4138=>"111111100",
  4139=>"000100100",
  4140=>"111110110",
  4141=>"111101101",
  4142=>"101101111",
  4143=>"010110000",
  4144=>"000000111",
  4145=>"111111001",
  4146=>"001000000",
  4147=>"000000000",
  4148=>"111111101",
  4149=>"100100010",
  4150=>"000000011",
  4151=>"110100100",
  4152=>"001000000",
  4153=>"100100111",
  4154=>"000111111",
  4155=>"111111111",
  4156=>"100000000",
  4157=>"011011111",
  4158=>"000000011",
  4159=>"000000000",
  4160=>"000000000",
  4161=>"111111000",
  4162=>"111111111",
  4163=>"100111111",
  4164=>"000000000",
  4165=>"100000000",
  4166=>"000000000",
  4167=>"001001001",
  4168=>"111111111",
  4169=>"000000001",
  4170=>"111100000",
  4171=>"000001101",
  4172=>"100111111",
  4173=>"111111111",
  4174=>"011011010",
  4175=>"111111111",
  4176=>"111111000",
  4177=>"000000000",
  4178=>"000000000",
  4179=>"000010010",
  4180=>"000000000",
  4181=>"010000000",
  4182=>"000000000",
  4183=>"000000000",
  4184=>"000001001",
  4185=>"000000111",
  4186=>"110111010",
  4187=>"010110011",
  4188=>"111111010",
  4189=>"000000000",
  4190=>"000001011",
  4191=>"000000000",
  4192=>"000000111",
  4193=>"010010001",
  4194=>"011001100",
  4195=>"111110111",
  4196=>"000000000",
  4197=>"001001001",
  4198=>"000000000",
  4199=>"000100000",
  4200=>"000000000",
  4201=>"000000001",
  4202=>"001000000",
  4203=>"100110111",
  4204=>"000010110",
  4205=>"000000000",
  4206=>"111000000",
  4207=>"000000111",
  4208=>"111111000",
  4209=>"000001111",
  4210=>"100000000",
  4211=>"000100100",
  4212=>"011111111",
  4213=>"111111111",
  4214=>"000000000",
  4215=>"011000000",
  4216=>"000000000",
  4217=>"110111101",
  4218=>"011011001",
  4219=>"001001001",
  4220=>"110100110",
  4221=>"110111111",
  4222=>"111111001",
  4223=>"001001101",
  4224=>"010000000",
  4225=>"100110111",
  4226=>"000000000",
  4227=>"001101100",
  4228=>"111111111",
  4229=>"100100111",
  4230=>"110111111",
  4231=>"010100111",
  4232=>"000011111",
  4233=>"000001001",
  4234=>"000000000",
  4235=>"111101111",
  4236=>"000000000",
  4237=>"010000000",
  4238=>"100110111",
  4239=>"000000001",
  4240=>"111111111",
  4241=>"111111111",
  4242=>"000100100",
  4243=>"000000000",
  4244=>"001111111",
  4245=>"100100100",
  4246=>"000001011",
  4247=>"000100100",
  4248=>"000000000",
  4249=>"011111111",
  4250=>"000000001",
  4251=>"000000000",
  4252=>"111111111",
  4253=>"001011000",
  4254=>"001001000",
  4255=>"111111111",
  4256=>"010010000",
  4257=>"000000100",
  4258=>"000000000",
  4259=>"000100110",
  4260=>"000000000",
  4261=>"111111111",
  4262=>"000000000",
  4263=>"001001000",
  4264=>"010110010",
  4265=>"001000000",
  4266=>"111010000",
  4267=>"111111111",
  4268=>"001001011",
  4269=>"000000100",
  4270=>"000000000",
  4271=>"111111111",
  4272=>"011111011",
  4273=>"111001101",
  4274=>"011111011",
  4275=>"111111111",
  4276=>"111101111",
  4277=>"000000000",
  4278=>"000000000",
  4279=>"111111111",
  4280=>"001111111",
  4281=>"111011111",
  4282=>"010000000",
  4283=>"000101100",
  4284=>"000000000",
  4285=>"111111111",
  4286=>"111111111",
  4287=>"111111111",
  4288=>"101000000",
  4289=>"000000000",
  4290=>"001001001",
  4291=>"000000000",
  4292=>"100100100",
  4293=>"000000000",
  4294=>"111111000",
  4295=>"111000000",
  4296=>"000100000",
  4297=>"011001101",
  4298=>"000000000",
  4299=>"111000000",
  4300=>"000000000",
  4301=>"111110110",
  4302=>"111111111",
  4303=>"000000000",
  4304=>"111111111",
  4305=>"011100100",
  4306=>"011011111",
  4307=>"111111111",
  4308=>"100000000",
  4309=>"000001011",
  4310=>"001000000",
  4311=>"000000101",
  4312=>"111000000",
  4313=>"111111111",
  4314=>"000010000",
  4315=>"110111111",
  4316=>"000110111",
  4317=>"000000110",
  4318=>"000000000",
  4319=>"000000000",
  4320=>"000000000",
  4321=>"100110000",
  4322=>"000000000",
  4323=>"000000000",
  4324=>"111011001",
  4325=>"000000110",
  4326=>"101101000",
  4327=>"111110000",
  4328=>"101111110",
  4329=>"011001001",
  4330=>"101001000",
  4331=>"000000000",
  4332=>"000000000",
  4333=>"010010000",
  4334=>"111111101",
  4335=>"000010010",
  4336=>"001000100",
  4337=>"111110110",
  4338=>"000001111",
  4339=>"000000001",
  4340=>"000000111",
  4341=>"000000000",
  4342=>"111111111",
  4343=>"000000000",
  4344=>"011011111",
  4345=>"000000000",
  4346=>"000000000",
  4347=>"000001011",
  4348=>"000000000",
  4349=>"000000000",
  4350=>"010000111",
  4351=>"011111111",
  4352=>"000110000",
  4353=>"111101001",
  4354=>"100100100",
  4355=>"111111110",
  4356=>"111111111",
  4357=>"011111111",
  4358=>"111111111",
  4359=>"000000000",
  4360=>"000100111",
  4361=>"000000100",
  4362=>"111111111",
  4363=>"000000000",
  4364=>"110111110",
  4365=>"000000011",
  4366=>"000110000",
  4367=>"000000011",
  4368=>"000000000",
  4369=>"011100111",
  4370=>"000000111",
  4371=>"011000111",
  4372=>"111111001",
  4373=>"000000000",
  4374=>"100101001",
  4375=>"101001111",
  4376=>"111111111",
  4377=>"111001001",
  4378=>"000100100",
  4379=>"110110111",
  4380=>"000100000",
  4381=>"000000110",
  4382=>"000000000",
  4383=>"001101111",
  4384=>"100100010",
  4385=>"100111111",
  4386=>"111111010",
  4387=>"100100111",
  4388=>"111110100",
  4389=>"000000000",
  4390=>"110110000",
  4391=>"000111001",
  4392=>"111111100",
  4393=>"000000000",
  4394=>"111111111",
  4395=>"000110100",
  4396=>"000011011",
  4397=>"110000001",
  4398=>"000000000",
  4399=>"000000000",
  4400=>"100000000",
  4401=>"000000000",
  4402=>"000000000",
  4403=>"111001000",
  4404=>"000000000",
  4405=>"111101111",
  4406=>"000000000",
  4407=>"110110110",
  4408=>"001001000",
  4409=>"100000000",
  4410=>"110110111",
  4411=>"000000100",
  4412=>"100000000",
  4413=>"000000000",
  4414=>"110000000",
  4415=>"110000000",
  4416=>"000000000",
  4417=>"000110110",
  4418=>"000000000",
  4419=>"100100110",
  4420=>"111111111",
  4421=>"010110111",
  4422=>"110100000",
  4423=>"000010111",
  4424=>"111001000",
  4425=>"100100111",
  4426=>"111111100",
  4427=>"111110110",
  4428=>"111111111",
  4429=>"000011000",
  4430=>"110111110",
  4431=>"111011100",
  4432=>"100111111",
  4433=>"000000000",
  4434=>"000111111",
  4435=>"111111111",
  4436=>"001000000",
  4437=>"001001001",
  4438=>"000000001",
  4439=>"111111111",
  4440=>"111111111",
  4441=>"110110111",
  4442=>"000010011",
  4443=>"000010110",
  4444=>"000100111",
  4445=>"111111000",
  4446=>"000000000",
  4447=>"110110000",
  4448=>"111110000",
  4449=>"110111111",
  4450=>"000000110",
  4451=>"000000000",
  4452=>"111110111",
  4453=>"111111001",
  4454=>"100100011",
  4455=>"000000110",
  4456=>"101001001",
  4457=>"011001000",
  4458=>"111111111",
  4459=>"111011001",
  4460=>"111001001",
  4461=>"000000000",
  4462=>"000000000",
  4463=>"000010000",
  4464=>"111111011",
  4465=>"011111011",
  4466=>"111111111",
  4467=>"001001000",
  4468=>"000000000",
  4469=>"000000111",
  4470=>"000000000",
  4471=>"000000000",
  4472=>"110100111",
  4473=>"111111010",
  4474=>"000110111",
  4475=>"110110000",
  4476=>"011111100",
  4477=>"101101101",
  4478=>"000000000",
  4479=>"111111000",
  4480=>"100100010",
  4481=>"110000000",
  4482=>"110110110",
  4483=>"000100110",
  4484=>"000000111",
  4485=>"000001001",
  4486=>"111110000",
  4487=>"000001001",
  4488=>"000000000",
  4489=>"111111111",
  4490=>"000000111",
  4491=>"000001001",
  4492=>"000000111",
  4493=>"111111111",
  4494=>"000000000",
  4495=>"000000000",
  4496=>"000000000",
  4497=>"010111111",
  4498=>"000000001",
  4499=>"000000000",
  4500=>"000110110",
  4501=>"000000000",
  4502=>"000000000",
  4503=>"000001111",
  4504=>"000000000",
  4505=>"000011111",
  4506=>"000111111",
  4507=>"111000100",
  4508=>"011011011",
  4509=>"000000000",
  4510=>"011010000",
  4511=>"111111101",
  4512=>"111010000",
  4513=>"111110100",
  4514=>"000100111",
  4515=>"000010010",
  4516=>"111111111",
  4517=>"000000000",
  4518=>"111111111",
  4519=>"000111111",
  4520=>"011011111",
  4521=>"100000000",
  4522=>"000011111",
  4523=>"011001000",
  4524=>"110111111",
  4525=>"000000000",
  4526=>"111110100",
  4527=>"111111111",
  4528=>"000000000",
  4529=>"000000000",
  4530=>"111100101",
  4531=>"000111111",
  4532=>"000110100",
  4533=>"010000000",
  4534=>"001000000",
  4535=>"000001110",
  4536=>"111111110",
  4537=>"111111111",
  4538=>"000000100",
  4539=>"000000110",
  4540=>"011011000",
  4541=>"001000001",
  4542=>"111001000",
  4543=>"111111111",
  4544=>"000000000",
  4545=>"000000001",
  4546=>"001001000",
  4547=>"000100111",
  4548=>"000000111",
  4549=>"011000011",
  4550=>"101101111",
  4551=>"000001001",
  4552=>"000000000",
  4553=>"001001000",
  4554=>"000000001",
  4555=>"000000001",
  4556=>"111000000",
  4557=>"000000000",
  4558=>"011111100",
  4559=>"110000001",
  4560=>"011011000",
  4561=>"110111111",
  4562=>"111111001",
  4563=>"110110111",
  4564=>"111111001",
  4565=>"110111111",
  4566=>"000000000",
  4567=>"001001000",
  4568=>"000000000",
  4569=>"000000010",
  4570=>"000100100",
  4571=>"000000011",
  4572=>"000000000",
  4573=>"000000000",
  4574=>"001000000",
  4575=>"111000011",
  4576=>"111001000",
  4577=>"111000000",
  4578=>"000100110",
  4579=>"111111100",
  4580=>"111111111",
  4581=>"111111111",
  4582=>"101100000",
  4583=>"000000100",
  4584=>"111111100",
  4585=>"110100101",
  4586=>"111110110",
  4587=>"111111111",
  4588=>"000010000",
  4589=>"001001000",
  4590=>"000000000",
  4591=>"000000111",
  4592=>"011001000",
  4593=>"000000000",
  4594=>"000000000",
  4595=>"000001000",
  4596=>"000000000",
  4597=>"110110010",
  4598=>"000000000",
  4599=>"111111110",
  4600=>"111101000",
  4601=>"011011011",
  4602=>"001000000",
  4603=>"100000000",
  4604=>"110111111",
  4605=>"111111000",
  4606=>"111111111",
  4607=>"001001011",
  4608=>"110010101",
  4609=>"010000110",
  4610=>"000000111",
  4611=>"000000110",
  4612=>"011011001",
  4613=>"010010000",
  4614=>"000000111",
  4615=>"111111111",
  4616=>"010000011",
  4617=>"100000000",
  4618=>"000000000",
  4619=>"000100100",
  4620=>"101001010",
  4621=>"100111100",
  4622=>"111000000",
  4623=>"000000000",
  4624=>"111000000",
  4625=>"000000011",
  4626=>"110000000",
  4627=>"000111011",
  4628=>"000100001",
  4629=>"011000000",
  4630=>"111111011",
  4631=>"000111111",
  4632=>"111110110",
  4633=>"000110100",
  4634=>"101001111",
  4635=>"000011000",
  4636=>"001001111",
  4637=>"111111111",
  4638=>"101111011",
  4639=>"111010000",
  4640=>"000000001",
  4641=>"001001001",
  4642=>"111111111",
  4643=>"101000111",
  4644=>"111111111",
  4645=>"001001101",
  4646=>"110010010",
  4647=>"000010000",
  4648=>"100000000",
  4649=>"000000000",
  4650=>"000101101",
  4651=>"000001111",
  4652=>"110110000",
  4653=>"100101001",
  4654=>"000000000",
  4655=>"111010000",
  4656=>"110101000",
  4657=>"000000010",
  4658=>"011111101",
  4659=>"011111110",
  4660=>"000110000",
  4661=>"101101001",
  4662=>"000110000",
  4663=>"000001000",
  4664=>"000000000",
  4665=>"000001111",
  4666=>"001101000",
  4667=>"000111111",
  4668=>"000000000",
  4669=>"001001000",
  4670=>"100101111",
  4671=>"000001000",
  4672=>"000000000",
  4673=>"000110000",
  4674=>"000011111",
  4675=>"111010000",
  4676=>"100100111",
  4677=>"011000000",
  4678=>"001000111",
  4679=>"000000000",
  4680=>"111111000",
  4681=>"101000001",
  4682=>"011111100",
  4683=>"010111111",
  4684=>"110110110",
  4685=>"111010000",
  4686=>"000000010",
  4687=>"111111111",
  4688=>"011111011",
  4689=>"111000100",
  4690=>"000110000",
  4691=>"001001001",
  4692=>"000001000",
  4693=>"000000000",
  4694=>"000000000",
  4695=>"000000000",
  4696=>"110110111",
  4697=>"101000101",
  4698=>"001011001",
  4699=>"111111010",
  4700=>"000000111",
  4701=>"000111010",
  4702=>"011111010",
  4703=>"000111111",
  4704=>"110000000",
  4705=>"111111111",
  4706=>"110000000",
  4707=>"000000111",
  4708=>"010000110",
  4709=>"000000111",
  4710=>"111111111",
  4711=>"000000000",
  4712=>"111000000",
  4713=>"000001111",
  4714=>"000000000",
  4715=>"000110111",
  4716=>"111111111",
  4717=>"000000010",
  4718=>"111010000",
  4719=>"000000000",
  4720=>"100100100",
  4721=>"101000010",
  4722=>"111100100",
  4723=>"111001000",
  4724=>"100000100",
  4725=>"001000111",
  4726=>"011001111",
  4727=>"000000110",
  4728=>"111100101",
  4729=>"111111111",
  4730=>"111001001",
  4731=>"111001111",
  4732=>"000110100",
  4733=>"110111011",
  4734=>"110100111",
  4735=>"110111101",
  4736=>"101000111",
  4737=>"111101100",
  4738=>"001000000",
  4739=>"000000110",
  4740=>"000111101",
  4741=>"110110110",
  4742=>"000110001",
  4743=>"110000111",
  4744=>"111000000",
  4745=>"110110000",
  4746=>"100100000",
  4747=>"100100111",
  4748=>"010010001",
  4749=>"100000100",
  4750=>"001000111",
  4751=>"000000001",
  4752=>"101101111",
  4753=>"110000000",
  4754=>"011111110",
  4755=>"110110111",
  4756=>"110110000",
  4757=>"111001000",
  4758=>"000001111",
  4759=>"101000000",
  4760=>"000000111",
  4761=>"111101101",
  4762=>"111100110",
  4763=>"010111111",
  4764=>"010010111",
  4765=>"000000001",
  4766=>"000111000",
  4767=>"000101111",
  4768=>"101101001",
  4769=>"101111011",
  4770=>"000000111",
  4771=>"010111011",
  4772=>"001001001",
  4773=>"000000000",
  4774=>"010111111",
  4775=>"101111100",
  4776=>"000010000",
  4777=>"110000111",
  4778=>"000000011",
  4779=>"111010110",
  4780=>"010111111",
  4781=>"000100001",
  4782=>"100000101",
  4783=>"000000000",
  4784=>"000011110",
  4785=>"000011001",
  4786=>"110111111",
  4787=>"111111111",
  4788=>"010111111",
  4789=>"100011011",
  4790=>"111010000",
  4791=>"001001001",
  4792=>"100100101",
  4793=>"111111111",
  4794=>"111001111",
  4795=>"111111111",
  4796=>"010111110",
  4797=>"111110110",
  4798=>"000110111",
  4799=>"011000011",
  4800=>"000000000",
  4801=>"010110010",
  4802=>"000000111",
  4803=>"000010000",
  4804=>"111000000",
  4805=>"000000101",
  4806=>"011111000",
  4807=>"010010011",
  4808=>"000000000",
  4809=>"101101000",
  4810=>"111111010",
  4811=>"110011011",
  4812=>"111111110",
  4813=>"000111110",
  4814=>"000100110",
  4815=>"000001000",
  4816=>"000010110",
  4817=>"000000000",
  4818=>"111110110",
  4819=>"000000101",
  4820=>"111101001",
  4821=>"101101111",
  4822=>"000011000",
  4823=>"000000000",
  4824=>"000000000",
  4825=>"001111000",
  4826=>"000111011",
  4827=>"000000111",
  4828=>"111111100",
  4829=>"110111111",
  4830=>"111111000",
  4831=>"000011111",
  4832=>"111111111",
  4833=>"000010010",
  4834=>"111001000",
  4835=>"111111111",
  4836=>"000111001",
  4837=>"111111110",
  4838=>"010110010",
  4839=>"010010111",
  4840=>"111111101",
  4841=>"000100100",
  4842=>"000000000",
  4843=>"111111100",
  4844=>"000000100",
  4845=>"111000000",
  4846=>"010010111",
  4847=>"000000111",
  4848=>"111011001",
  4849=>"000000001",
  4850=>"001001000",
  4851=>"101001101",
  4852=>"111111010",
  4853=>"000001111",
  4854=>"101111111",
  4855=>"000011011",
  4856=>"101000001",
  4857=>"000000001",
  4858=>"001101100",
  4859=>"000000110",
  4860=>"100111000",
  4861=>"111111111",
  4862=>"111000000",
  4863=>"100110110",
  4864=>"100001010",
  4865=>"011110000",
  4866=>"111001011",
  4867=>"011001001",
  4868=>"100101111",
  4869=>"110000011",
  4870=>"010111111",
  4871=>"011111111",
  4872=>"100100000",
  4873=>"110000000",
  4874=>"110110010",
  4875=>"000111011",
  4876=>"111000001",
  4877=>"001000110",
  4878=>"000000100",
  4879=>"111001110",
  4880=>"000011111",
  4881=>"110000110",
  4882=>"000000000",
  4883=>"010010000",
  4884=>"101111111",
  4885=>"110000000",
  4886=>"000100111",
  4887=>"000000000",
  4888=>"000000100",
  4889=>"111011000",
  4890=>"000000000",
  4891=>"000000111",
  4892=>"111111111",
  4893=>"010000010",
  4894=>"111111111",
  4895=>"001101111",
  4896=>"101111011",
  4897=>"010110111",
  4898=>"111010000",
  4899=>"101101111",
  4900=>"010010000",
  4901=>"110110011",
  4902=>"000001111",
  4903=>"000000001",
  4904=>"100101111",
  4905=>"111011000",
  4906=>"010000001",
  4907=>"001000011",
  4908=>"111111000",
  4909=>"000001001",
  4910=>"110000111",
  4911=>"000000100",
  4912=>"000100100",
  4913=>"011111010",
  4914=>"100100000",
  4915=>"111000000",
  4916=>"000000000",
  4917=>"000000000",
  4918=>"000000111",
  4919=>"000000111",
  4920=>"101101000",
  4921=>"101001111",
  4922=>"111111010",
  4923=>"001001000",
  4924=>"000000100",
  4925=>"111010000",
  4926=>"100000001",
  4927=>"100100111",
  4928=>"111000100",
  4929=>"111110000",
  4930=>"000000001",
  4931=>"000100100",
  4932=>"100111010",
  4933=>"010000100",
  4934=>"000001000",
  4935=>"111000000",
  4936=>"100000000",
  4937=>"010010111",
  4938=>"011110000",
  4939=>"000100000",
  4940=>"010000011",
  4941=>"110000000",
  4942=>"000011111",
  4943=>"111000100",
  4944=>"000000000",
  4945=>"000000101",
  4946=>"100101000",
  4947=>"110101101",
  4948=>"000000000",
  4949=>"011011000",
  4950=>"010010000",
  4951=>"111010000",
  4952=>"111001000",
  4953=>"000010011",
  4954=>"111000100",
  4955=>"101101000",
  4956=>"000000000",
  4957=>"111000111",
  4958=>"110000100",
  4959=>"011000011",
  4960=>"111111111",
  4961=>"000111111",
  4962=>"100110100",
  4963=>"011111111",
  4964=>"000100110",
  4965=>"000000001",
  4966=>"111100000",
  4967=>"001001001",
  4968=>"000100100",
  4969=>"111001000",
  4970=>"100000111",
  4971=>"000110000",
  4972=>"000110110",
  4973=>"001011111",
  4974=>"111100100",
  4975=>"000000111",
  4976=>"100100111",
  4977=>"000110110",
  4978=>"000111111",
  4979=>"111111111",
  4980=>"000000000",
  4981=>"111110110",
  4982=>"011111100",
  4983=>"000000000",
  4984=>"000111111",
  4985=>"000000010",
  4986=>"000100100",
  4987=>"000000001",
  4988=>"111111111",
  4989=>"000000000",
  4990=>"000000000",
  4991=>"000000000",
  4992=>"011011000",
  4993=>"111111000",
  4994=>"110000000",
  4995=>"111111110",
  4996=>"000000000",
  4997=>"000000000",
  4998=>"110111000",
  4999=>"000110100",
  5000=>"110100111",
  5001=>"111111000",
  5002=>"010010000",
  5003=>"111010000",
  5004=>"110111111",
  5005=>"000111001",
  5006=>"000000000",
  5007=>"000000000",
  5008=>"000110010",
  5009=>"111111011",
  5010=>"111110100",
  5011=>"000000001",
  5012=>"000000010",
  5013=>"111010000",
  5014=>"000000111",
  5015=>"101111011",
  5016=>"100000111",
  5017=>"011011011",
  5018=>"001111111",
  5019=>"111000000",
  5020=>"000000000",
  5021=>"111001011",
  5022=>"000111111",
  5023=>"000111111",
  5024=>"101001011",
  5025=>"011110111",
  5026=>"111111001",
  5027=>"111000000",
  5028=>"111111011",
  5029=>"000000000",
  5030=>"111111111",
  5031=>"011000110",
  5032=>"100110000",
  5033=>"111011111",
  5034=>"000000001",
  5035=>"011011000",
  5036=>"000000000",
  5037=>"100000000",
  5038=>"000000001",
  5039=>"111011000",
  5040=>"000000001",
  5041=>"111111010",
  5042=>"000000111",
  5043=>"111100000",
  5044=>"010000110",
  5045=>"100000111",
  5046=>"101001101",
  5047=>"011111111",
  5048=>"001010000",
  5049=>"011011011",
  5050=>"000000011",
  5051=>"010110000",
  5052=>"000000111",
  5053=>"100000000",
  5054=>"000001111",
  5055=>"000000000",
  5056=>"010010000",
  5057=>"111101111",
  5058=>"100000001",
  5059=>"000111010",
  5060=>"110100000",
  5061=>"000001100",
  5062=>"111111001",
  5063=>"000010000",
  5064=>"100100000",
  5065=>"100000000",
  5066=>"000000000",
  5067=>"110111111",
  5068=>"010000000",
  5069=>"111111111",
  5070=>"000010010",
  5071=>"001101111",
  5072=>"000110100",
  5073=>"000110000",
  5074=>"111111110",
  5075=>"110100100",
  5076=>"110111111",
  5077=>"011111111",
  5078=>"110010000",
  5079=>"100000000",
  5080=>"010111101",
  5081=>"000000110",
  5082=>"000001011",
  5083=>"000000000",
  5084=>"001000000",
  5085=>"000000111",
  5086=>"011011111",
  5087=>"111010000",
  5088=>"100100111",
  5089=>"000000000",
  5090=>"111001001",
  5091=>"111111000",
  5092=>"111010011",
  5093=>"000000001",
  5094=>"111000000",
  5095=>"010000111",
  5096=>"011101001",
  5097=>"000010011",
  5098=>"000010011",
  5099=>"000001111",
  5100=>"000010111",
  5101=>"001000000",
  5102=>"100100111",
  5103=>"000000100",
  5104=>"101000101",
  5105=>"001001001",
  5106=>"000111111",
  5107=>"000000000",
  5108=>"111111111",
  5109=>"111000000",
  5110=>"110110000",
  5111=>"111101111",
  5112=>"110111111",
  5113=>"001001000",
  5114=>"000000111",
  5115=>"011000111",
  5116=>"110011111",
  5117=>"111110000",
  5118=>"010110111",
  5119=>"111101111",
  5120=>"000000110",
  5121=>"011010010",
  5122=>"111111111",
  5123=>"000000000",
  5124=>"011000000",
  5125=>"111111111",
  5126=>"000111111",
  5127=>"001111111",
  5128=>"111111100",
  5129=>"111000000",
  5130=>"000000000",
  5131=>"000011011",
  5132=>"000110000",
  5133=>"000000101",
  5134=>"111111111",
  5135=>"100100100",
  5136=>"011011111",
  5137=>"000000011",
  5138=>"000100111",
  5139=>"110111110",
  5140=>"110000000",
  5141=>"010111110",
  5142=>"111000001",
  5143=>"001001000",
  5144=>"110110000",
  5145=>"000100111",
  5146=>"000000111",
  5147=>"000001011",
  5148=>"110110000",
  5149=>"000001001",
  5150=>"000000111",
  5151=>"010111000",
  5152=>"000000111",
  5153=>"000111001",
  5154=>"111111111",
  5155=>"111000000",
  5156=>"000000000",
  5157=>"111111011",
  5158=>"000000100",
  5159=>"110000001",
  5160=>"110110111",
  5161=>"000110111",
  5162=>"001001000",
  5163=>"111111111",
  5164=>"001000111",
  5165=>"110111110",
  5166=>"001011111",
  5167=>"000100110",
  5168=>"000001011",
  5169=>"000000111",
  5170=>"001111110",
  5171=>"111111000",
  5172=>"001000111",
  5173=>"000111111",
  5174=>"100000000",
  5175=>"101110110",
  5176=>"001111110",
  5177=>"111111000",
  5178=>"000111111",
  5179=>"011001111",
  5180=>"000000001",
  5181=>"111111110",
  5182=>"000000001",
  5183=>"000001111",
  5184=>"110111111",
  5185=>"100000101",
  5186=>"111111100",
  5187=>"110000100",
  5188=>"010000000",
  5189=>"001001001",
  5190=>"000000011",
  5191=>"101100101",
  5192=>"011100101",
  5193=>"000000111",
  5194=>"000000000",
  5195=>"111111111",
  5196=>"111111100",
  5197=>"111111000",
  5198=>"000010011",
  5199=>"000000110",
  5200=>"100110110",
  5201=>"111001111",
  5202=>"110111111",
  5203=>"110110110",
  5204=>"000000000",
  5205=>"000110100",
  5206=>"000000000",
  5207=>"000000000",
  5208=>"111001100",
  5209=>"000000111",
  5210=>"010000110",
  5211=>"010011100",
  5212=>"111111111",
  5213=>"111111001",
  5214=>"111110100",
  5215=>"010110000",
  5216=>"000111000",
  5217=>"001100111",
  5218=>"000000111",
  5219=>"000101111",
  5220=>"111111000",
  5221=>"000000111",
  5222=>"000000000",
  5223=>"111000111",
  5224=>"111111111",
  5225=>"111111111",
  5226=>"111111110",
  5227=>"010000000",
  5228=>"111011001",
  5229=>"111111000",
  5230=>"111111111",
  5231=>"111111100",
  5232=>"000000000",
  5233=>"000000100",
  5234=>"000000111",
  5235=>"000000000",
  5236=>"000101111",
  5237=>"111010000",
  5238=>"100100101",
  5239=>"001100111",
  5240=>"000000111",
  5241=>"000001000",
  5242=>"111000000",
  5243=>"001000011",
  5244=>"100110110",
  5245=>"111111111",
  5246=>"101111000",
  5247=>"111111111",
  5248=>"111000000",
  5249=>"111010110",
  5250=>"110111000",
  5251=>"011011011",
  5252=>"000111111",
  5253=>"001001111",
  5254=>"111111111",
  5255=>"100101111",
  5256=>"001000000",
  5257=>"110001000",
  5258=>"111111111",
  5259=>"111111111",
  5260=>"000000000",
  5261=>"000000000",
  5262=>"111100000",
  5263=>"000111111",
  5264=>"000000111",
  5265=>"000000111",
  5266=>"111010110",
  5267=>"000111111",
  5268=>"111010000",
  5269=>"000000111",
  5270=>"111110111",
  5271=>"111000000",
  5272=>"000000000",
  5273=>"000000111",
  5274=>"010011111",
  5275=>"111000110",
  5276=>"001001000",
  5277=>"001000110",
  5278=>"011011011",
  5279=>"100100101",
  5280=>"000100110",
  5281=>"111111111",
  5282=>"111111111",
  5283=>"111111111",
  5284=>"101001111",
  5285=>"100100111",
  5286=>"000000000",
  5287=>"000111111",
  5288=>"000001011",
  5289=>"000000100",
  5290=>"010111001",
  5291=>"100111111",
  5292=>"111111011",
  5293=>"100000001",
  5294=>"000100111",
  5295=>"000000000",
  5296=>"000101111",
  5297=>"000111111",
  5298=>"000011010",
  5299=>"111111000",
  5300=>"000010111",
  5301=>"000000000",
  5302=>"000000111",
  5303=>"101011111",
  5304=>"111111111",
  5305=>"000000000",
  5306=>"001000000",
  5307=>"101011111",
  5308=>"000000000",
  5309=>"111111100",
  5310=>"111111111",
  5311=>"000000001",
  5312=>"111100110",
  5313=>"111001001",
  5314=>"011111111",
  5315=>"000000001",
  5316=>"000100111",
  5317=>"011000000",
  5318=>"111110000",
  5319=>"000000010",
  5320=>"000111111",
  5321=>"000000000",
  5322=>"110010000",
  5323=>"010111111",
  5324=>"111111110",
  5325=>"000000000",
  5326=>"000110100",
  5327=>"010000010",
  5328=>"110101111",
  5329=>"000011011",
  5330=>"110010111",
  5331=>"100100100",
  5332=>"111000100",
  5333=>"000011111",
  5334=>"000000101",
  5335=>"111111111",
  5336=>"000000011",
  5337=>"111111000",
  5338=>"110110000",
  5339=>"000000000",
  5340=>"111110000",
  5341=>"000000111",
  5342=>"111001000",
  5343=>"000011001",
  5344=>"000000000",
  5345=>"000000111",
  5346=>"011011011",
  5347=>"111111111",
  5348=>"000011000",
  5349=>"110110001",
  5350=>"011111111",
  5351=>"111111111",
  5352=>"111111111",
  5353=>"111111000",
  5354=>"000000000",
  5355=>"000110111",
  5356=>"100001001",
  5357=>"000000110",
  5358=>"000100111",
  5359=>"000000111",
  5360=>"000001011",
  5361=>"000000000",
  5362=>"000000000",
  5363=>"000000000",
  5364=>"001011111",
  5365=>"000001001",
  5366=>"111111000",
  5367=>"000000010",
  5368=>"100000000",
  5369=>"000110011",
  5370=>"111111001",
  5371=>"001111110",
  5372=>"000000110",
  5373=>"000000001",
  5374=>"111000000",
  5375=>"100111111",
  5376=>"111101000",
  5377=>"001000111",
  5378=>"011111111",
  5379=>"111000001",
  5380=>"001111110",
  5381=>"101111101",
  5382=>"110100111",
  5383=>"000000001",
  5384=>"111111111",
  5385=>"111010000",
  5386=>"000000000",
  5387=>"111111110",
  5388=>"100111111",
  5389=>"000000111",
  5390=>"111000000",
  5391=>"011111111",
  5392=>"000000000",
  5393=>"000000011",
  5394=>"000010011",
  5395=>"000000000",
  5396=>"000001011",
  5397=>"111110000",
  5398=>"010111111",
  5399=>"000111000",
  5400=>"111111110",
  5401=>"000000101",
  5402=>"010000000",
  5403=>"100100110",
  5404=>"000000000",
  5405=>"000000110",
  5406=>"000000100",
  5407=>"111111011",
  5408=>"011010000",
  5409=>"000111010",
  5410=>"110111111",
  5411=>"111111111",
  5412=>"010000011",
  5413=>"111000000",
  5414=>"000011000",
  5415=>"001011010",
  5416=>"000111011",
  5417=>"010011011",
  5418=>"111010000",
  5419=>"000000111",
  5420=>"111111111",
  5421=>"111111111",
  5422=>"000111111",
  5423=>"101111000",
  5424=>"000011000",
  5425=>"111111111",
  5426=>"110111111",
  5427=>"000000000",
  5428=>"111010001",
  5429=>"111110010",
  5430=>"000000001",
  5431=>"000001001",
  5432=>"111111000",
  5433=>"111111111",
  5434=>"111011001",
  5435=>"111111111",
  5436=>"111111111",
  5437=>"000000000",
  5438=>"001001111",
  5439=>"100000110",
  5440=>"111001111",
  5441=>"111111110",
  5442=>"001001000",
  5443=>"001001111",
  5444=>"111010000",
  5445=>"000000000",
  5446=>"000110000",
  5447=>"000000000",
  5448=>"111111111",
  5449=>"111111111",
  5450=>"001000000",
  5451=>"001000000",
  5452=>"000010010",
  5453=>"111110000",
  5454=>"111001110",
  5455=>"111111110",
  5456=>"111111000",
  5457=>"001000000",
  5458=>"111111111",
  5459=>"000000111",
  5460=>"000010010",
  5461=>"011011011",
  5462=>"111111111",
  5463=>"001000000",
  5464=>"000000100",
  5465=>"011011111",
  5466=>"000000000",
  5467=>"000000000",
  5468=>"010110110",
  5469=>"000011000",
  5470=>"000010110",
  5471=>"000000000",
  5472=>"111001000",
  5473=>"010111000",
  5474=>"000000111",
  5475=>"000000000",
  5476=>"000000011",
  5477=>"000000000",
  5478=>"110000000",
  5479=>"111111000",
  5480=>"000000100",
  5481=>"111000000",
  5482=>"000000000",
  5483=>"111101111",
  5484=>"000111111",
  5485=>"001000000",
  5486=>"000000000",
  5487=>"100101111",
  5488=>"111111111",
  5489=>"010010110",
  5490=>"000000111",
  5491=>"100011111",
  5492=>"111111111",
  5493=>"000000000",
  5494=>"111000111",
  5495=>"111111000",
  5496=>"111000100",
  5497=>"000000111",
  5498=>"000000000",
  5499=>"001000001",
  5500=>"100000111",
  5501=>"111111111",
  5502=>"110000000",
  5503=>"000000000",
  5504=>"001001001",
  5505=>"001001111",
  5506=>"000100110",
  5507=>"000100111",
  5508=>"100011011",
  5509=>"010000000",
  5510=>"111111111",
  5511=>"111111111",
  5512=>"000000000",
  5513=>"011111111",
  5514=>"000000110",
  5515=>"000111000",
  5516=>"110111111",
  5517=>"100110111",
  5518=>"110000111",
  5519=>"000000000",
  5520=>"000000000",
  5521=>"001101111",
  5522=>"100111110",
  5523=>"111111111",
  5524=>"011111111",
  5525=>"000110000",
  5526=>"000000111",
  5527=>"000110110",
  5528=>"111101111",
  5529=>"000100110",
  5530=>"001000000",
  5531=>"111111111",
  5532=>"000000000",
  5533=>"000000111",
  5534=>"000000000",
  5535=>"000111001",
  5536=>"100111100",
  5537=>"111111111",
  5538=>"110111111",
  5539=>"111111000",
  5540=>"111011000",
  5541=>"111000000",
  5542=>"111111111",
  5543=>"111000000",
  5544=>"000000111",
  5545=>"000000111",
  5546=>"110101111",
  5547=>"111111000",
  5548=>"000000011",
  5549=>"000000001",
  5550=>"110010111",
  5551=>"101111111",
  5552=>"010000111",
  5553=>"000000000",
  5554=>"101111111",
  5555=>"110111110",
  5556=>"000000000",
  5557=>"011000000",
  5558=>"111111101",
  5559=>"010010000",
  5560=>"111111000",
  5561=>"010010000",
  5562=>"000000111",
  5563=>"001011111",
  5564=>"000111111",
  5565=>"000001001",
  5566=>"011000000",
  5567=>"000110000",
  5568=>"100111000",
  5569=>"000010000",
  5570=>"001011111",
  5571=>"000001001",
  5572=>"000000001",
  5573=>"011001000",
  5574=>"111111000",
  5575=>"010001000",
  5576=>"000000000",
  5577=>"100100100",
  5578=>"000000011",
  5579=>"000000000",
  5580=>"000000000",
  5581=>"111111100",
  5582=>"000000000",
  5583=>"011111111",
  5584=>"101111111",
  5585=>"101111001",
  5586=>"110110110",
  5587=>"011000011",
  5588=>"000000010",
  5589=>"000000101",
  5590=>"000000111",
  5591=>"001111111",
  5592=>"100111111",
  5593=>"100111100",
  5594=>"000001011",
  5595=>"000000111",
  5596=>"000000001",
  5597=>"000000111",
  5598=>"111000000",
  5599=>"100100000",
  5600=>"110000100",
  5601=>"010000000",
  5602=>"000000000",
  5603=>"110110110",
  5604=>"000001111",
  5605=>"110000000",
  5606=>"111111111",
  5607=>"000000000",
  5608=>"111111010",
  5609=>"110000000",
  5610=>"101000001",
  5611=>"111011000",
  5612=>"100000010",
  5613=>"000011011",
  5614=>"001111111",
  5615=>"001000000",
  5616=>"111111101",
  5617=>"000000001",
  5618=>"000000000",
  5619=>"111011111",
  5620=>"111111000",
  5621=>"000100110",
  5622=>"111011000",
  5623=>"010011000",
  5624=>"011011000",
  5625=>"000001111",
  5626=>"000011011",
  5627=>"111101111",
  5628=>"000011111",
  5629=>"111111111",
  5630=>"000000011",
  5631=>"001000000",
  5632=>"001000111",
  5633=>"111111001",
  5634=>"111111111",
  5635=>"000111111",
  5636=>"111001100",
  5637=>"000000001",
  5638=>"000110100",
  5639=>"001001111",
  5640=>"100110001",
  5641=>"000011111",
  5642=>"111110010",
  5643=>"011111010",
  5644=>"000000000",
  5645=>"001011111",
  5646=>"111110000",
  5647=>"111110110",
  5648=>"111101100",
  5649=>"000000111",
  5650=>"000000110",
  5651=>"010111111",
  5652=>"000000101",
  5653=>"111000000",
  5654=>"010100100",
  5655=>"111111111",
  5656=>"100000000",
  5657=>"001000100",
  5658=>"111000101",
  5659=>"000000000",
  5660=>"111000111",
  5661=>"100111000",
  5662=>"010100000",
  5663=>"111111000",
  5664=>"000000000",
  5665=>"100000001",
  5666=>"110000001",
  5667=>"111111000",
  5668=>"000000000",
  5669=>"001000000",
  5670=>"111111011",
  5671=>"111000111",
  5672=>"000000111",
  5673=>"111000000",
  5674=>"000001001",
  5675=>"000000111",
  5676=>"111100000",
  5677=>"110111010",
  5678=>"111111111",
  5679=>"000000000",
  5680=>"000000000",
  5681=>"000111011",
  5682=>"111110000",
  5683=>"110000111",
  5684=>"111111110",
  5685=>"010110100",
  5686=>"100110000",
  5687=>"000000000",
  5688=>"000000111",
  5689=>"000001011",
  5690=>"011001000",
  5691=>"000000000",
  5692=>"111111111",
  5693=>"000000000",
  5694=>"111100111",
  5695=>"000000000",
  5696=>"000000110",
  5697=>"011001000",
  5698=>"111011000",
  5699=>"000001000",
  5700=>"110000000",
  5701=>"000110011",
  5702=>"111111000",
  5703=>"000000000",
  5704=>"000000111",
  5705=>"000101111",
  5706=>"000011000",
  5707=>"111111111",
  5708=>"110110110",
  5709=>"000000110",
  5710=>"001000011",
  5711=>"111111111",
  5712=>"011001001",
  5713=>"111111111",
  5714=>"101001111",
  5715=>"100110100",
  5716=>"110111000",
  5717=>"000010111",
  5718=>"111001001",
  5719=>"111111111",
  5720=>"100100000",
  5721=>"111000001",
  5722=>"000000111",
  5723=>"000000100",
  5724=>"111111111",
  5725=>"011111111",
  5726=>"000000000",
  5727=>"111110010",
  5728=>"000111111",
  5729=>"100000111",
  5730=>"000000111",
  5731=>"000000000",
  5732=>"100000000",
  5733=>"000111111",
  5734=>"000001000",
  5735=>"100000000",
  5736=>"000000000",
  5737=>"111000000",
  5738=>"010000110",
  5739=>"111001000",
  5740=>"011111111",
  5741=>"000111111",
  5742=>"000000100",
  5743=>"000000000",
  5744=>"111011000",
  5745=>"111111000",
  5746=>"000001001",
  5747=>"100110111",
  5748=>"110111011",
  5749=>"000100110",
  5750=>"000110111",
  5751=>"000000000",
  5752=>"000000000",
  5753=>"111101000",
  5754=>"000111111",
  5755=>"000000000",
  5756=>"000000000",
  5757=>"111111000",
  5758=>"111111111",
  5759=>"111111111",
  5760=>"000000100",
  5761=>"000111111",
  5762=>"111111111",
  5763=>"000011011",
  5764=>"111111000",
  5765=>"111011000",
  5766=>"100000110",
  5767=>"111111111",
  5768=>"111111111",
  5769=>"000011111",
  5770=>"000000000",
  5771=>"111111111",
  5772=>"100100111",
  5773=>"001011111",
  5774=>"000000001",
  5775=>"000000000",
  5776=>"111111000",
  5777=>"011011000",
  5778=>"111100000",
  5779=>"111111000",
  5780=>"000000000",
  5781=>"000100111",
  5782=>"110011000",
  5783=>"000111000",
  5784=>"000100111",
  5785=>"110110110",
  5786=>"000110111",
  5787=>"111110000",
  5788=>"111100100",
  5789=>"111110010",
  5790=>"111011111",
  5791=>"000000011",
  5792=>"000000111",
  5793=>"011111111",
  5794=>"000111111",
  5795=>"000000000",
  5796=>"000010110",
  5797=>"110111111",
  5798=>"000110010",
  5799=>"001001001",
  5800=>"111111001",
  5801=>"001011000",
  5802=>"111111111",
  5803=>"111000111",
  5804=>"111000000",
  5805=>"000010011",
  5806=>"010011111",
  5807=>"101111000",
  5808=>"000001111",
  5809=>"111001111",
  5810=>"010000010",
  5811=>"011010111",
  5812=>"001100000",
  5813=>"011111111",
  5814=>"001000000",
  5815=>"000001111",
  5816=>"000000000",
  5817=>"000000000",
  5818=>"000000000",
  5819=>"000001101",
  5820=>"111100110",
  5821=>"000000000",
  5822=>"111111111",
  5823=>"101100100",
  5824=>"000000111",
  5825=>"000110111",
  5826=>"011010111",
  5827=>"111111111",
  5828=>"111111111",
  5829=>"000111111",
  5830=>"000001111",
  5831=>"001001001",
  5832=>"011001000",
  5833=>"111000000",
  5834=>"111111111",
  5835=>"010011000",
  5836=>"000011111",
  5837=>"000000111",
  5838=>"110111000",
  5839=>"000010011",
  5840=>"000111110",
  5841=>"111111111",
  5842=>"000000000",
  5843=>"000000111",
  5844=>"001111000",
  5845=>"100111111",
  5846=>"000000110",
  5847=>"111110111",
  5848=>"111101000",
  5849=>"111000000",
  5850=>"000100000",
  5851=>"111000101",
  5852=>"010111111",
  5853=>"111111001",
  5854=>"100111111",
  5855=>"000000000",
  5856=>"000111000",
  5857=>"111000000",
  5858=>"010000000",
  5859=>"111111111",
  5860=>"011111111",
  5861=>"100100100",
  5862=>"000001000",
  5863=>"000000011",
  5864=>"000000101",
  5865=>"000010011",
  5866=>"101111111",
  5867=>"000000000",
  5868=>"111111111",
  5869=>"111110111",
  5870=>"000100000",
  5871=>"011111111",
  5872=>"000011000",
  5873=>"011111111",
  5874=>"000001011",
  5875=>"110000000",
  5876=>"111111111",
  5877=>"111111100",
  5878=>"111111001",
  5879=>"111111111",
  5880=>"111011001",
  5881=>"000000000",
  5882=>"111011000",
  5883=>"000001000",
  5884=>"000011000",
  5885=>"000001111",
  5886=>"111000111",
  5887=>"000111100",
  5888=>"000010000",
  5889=>"110110101",
  5890=>"110100000",
  5891=>"000100101",
  5892=>"000101111",
  5893=>"011111111",
  5894=>"111111001",
  5895=>"110000000",
  5896=>"111000000",
  5897=>"000000100",
  5898=>"111111111",
  5899=>"110111110",
  5900=>"001111110",
  5901=>"000000000",
  5902=>"110110000",
  5903=>"111111010",
  5904=>"000110000",
  5905=>"001011001",
  5906=>"011011001",
  5907=>"000000101",
  5908=>"111000000",
  5909=>"111100100",
  5910=>"110111111",
  5911=>"111111001",
  5912=>"000100000",
  5913=>"001011000",
  5914=>"110111000",
  5915=>"000010011",
  5916=>"001000000",
  5917=>"000111111",
  5918=>"000000111",
  5919=>"111111111",
  5920=>"000000001",
  5921=>"111111100",
  5922=>"111010000",
  5923=>"000000010",
  5924=>"111011111",
  5925=>"001001000",
  5926=>"111111111",
  5927=>"000000000",
  5928=>"000000101",
  5929=>"111000000",
  5930=>"111111111",
  5931=>"111110100",
  5932=>"000000000",
  5933=>"011111110",
  5934=>"101111110",
  5935=>"111000000",
  5936=>"000000100",
  5937=>"110110110",
  5938=>"111111111",
  5939=>"100100111",
  5940=>"000000000",
  5941=>"101101111",
  5942=>"000000000",
  5943=>"100100111",
  5944=>"111111000",
  5945=>"111000000",
  5946=>"000000000",
  5947=>"111111111",
  5948=>"000000000",
  5949=>"000111000",
  5950=>"000001111",
  5951=>"010111111",
  5952=>"000000000",
  5953=>"111111100",
  5954=>"111111111",
  5955=>"111101001",
  5956=>"001000000",
  5957=>"100100000",
  5958=>"100000000",
  5959=>"001011011",
  5960=>"111111000",
  5961=>"000000000",
  5962=>"000111110",
  5963=>"111100100",
  5964=>"000000100",
  5965=>"001000111",
  5966=>"110011000",
  5967=>"001001001",
  5968=>"100110100",
  5969=>"111111111",
  5970=>"111000000",
  5971=>"000000001",
  5972=>"000111111",
  5973=>"001001000",
  5974=>"111100000",
  5975=>"111001011",
  5976=>"111111111",
  5977=>"000111010",
  5978=>"111111000",
  5979=>"000000000",
  5980=>"000000000",
  5981=>"111111000",
  5982=>"110000000",
  5983=>"111111000",
  5984=>"000000000",
  5985=>"000000000",
  5986=>"000001010",
  5987=>"111111111",
  5988=>"111110110",
  5989=>"000110111",
  5990=>"111000111",
  5991=>"100110111",
  5992=>"111000001",
  5993=>"101000000",
  5994=>"100000100",
  5995=>"111111111",
  5996=>"000000000",
  5997=>"110100000",
  5998=>"000000000",
  5999=>"000001000",
  6000=>"000011111",
  6001=>"100110100",
  6002=>"000111110",
  6003=>"111111000",
  6004=>"100000111",
  6005=>"111111111",
  6006=>"110111100",
  6007=>"000000000",
  6008=>"111001011",
  6009=>"000001001",
  6010=>"111000000",
  6011=>"000000000",
  6012=>"111101000",
  6013=>"000000000",
  6014=>"000000000",
  6015=>"111111111",
  6016=>"001001000",
  6017=>"010111000",
  6018=>"001011000",
  6019=>"111111111",
  6020=>"111000000",
  6021=>"110000000",
  6022=>"000010111",
  6023=>"000100111",
  6024=>"000010000",
  6025=>"100110110",
  6026=>"111011111",
  6027=>"011000111",
  6028=>"111111110",
  6029=>"000000000",
  6030=>"111111111",
  6031=>"100100100",
  6032=>"000000000",
  6033=>"110111111",
  6034=>"010010000",
  6035=>"000001001",
  6036=>"000000000",
  6037=>"000000000",
  6038=>"100111111",
  6039=>"010111110",
  6040=>"111000000",
  6041=>"110111000",
  6042=>"000000110",
  6043=>"100100111",
  6044=>"111101111",
  6045=>"000001000",
  6046=>"010000000",
  6047=>"100111110",
  6048=>"000111110",
  6049=>"110100100",
  6050=>"101111000",
  6051=>"111111010",
  6052=>"111111111",
  6053=>"000000000",
  6054=>"000111111",
  6055=>"001101111",
  6056=>"010000000",
  6057=>"010011011",
  6058=>"111111111",
  6059=>"111111111",
  6060=>"000000000",
  6061=>"000001001",
  6062=>"111000000",
  6063=>"011000000",
  6064=>"000111111",
  6065=>"111111111",
  6066=>"000001001",
  6067=>"010111111",
  6068=>"001101111",
  6069=>"100000001",
  6070=>"000111111",
  6071=>"000110000",
  6072=>"001001001",
  6073=>"101100100",
  6074=>"111111100",
  6075=>"001001000",
  6076=>"000111111",
  6077=>"000110111",
  6078=>"111001000",
  6079=>"000011011",
  6080=>"111001111",
  6081=>"000000000",
  6082=>"011000011",
  6083=>"000000000",
  6084=>"111110111",
  6085=>"011001111",
  6086=>"001111111",
  6087=>"110110000",
  6088=>"111111000",
  6089=>"001000000",
  6090=>"000000000",
  6091=>"000010000",
  6092=>"001001000",
  6093=>"111111000",
  6094=>"111111101",
  6095=>"100111111",
  6096=>"111111011",
  6097=>"001000100",
  6098=>"101111111",
  6099=>"111111111",
  6100=>"111111100",
  6101=>"111111110",
  6102=>"000000011",
  6103=>"001001001",
  6104=>"000111001",
  6105=>"010010011",
  6106=>"111101111",
  6107=>"000000111",
  6108=>"111000000",
  6109=>"111111000",
  6110=>"101111000",
  6111=>"111001001",
  6112=>"000110010",
  6113=>"111100000",
  6114=>"111111111",
  6115=>"111111011",
  6116=>"000000000",
  6117=>"111000000",
  6118=>"100110101",
  6119=>"000000101",
  6120=>"001001011",
  6121=>"101001111",
  6122=>"000101111",
  6123=>"011001001",
  6124=>"111000000",
  6125=>"000100110",
  6126=>"111011010",
  6127=>"010000000",
  6128=>"001001001",
  6129=>"000111111",
  6130=>"001000111",
  6131=>"111111010",
  6132=>"111111111",
  6133=>"000011000",
  6134=>"111111111",
  6135=>"000111111",
  6136=>"011011000",
  6137=>"011100100",
  6138=>"000000000",
  6139=>"000111000",
  6140=>"000000000",
  6141=>"100100111",
  6142=>"010111111",
  6143=>"000000000",
  6144=>"000000000",
  6145=>"111111111",
  6146=>"000000100",
  6147=>"101111111",
  6148=>"000100100",
  6149=>"001001001",
  6150=>"000000000",
  6151=>"111001001",
  6152=>"000000001",
  6153=>"000111111",
  6154=>"111110000",
  6155=>"000000000",
  6156=>"110111111",
  6157=>"000000001",
  6158=>"001101101",
  6159=>"111111111",
  6160=>"111011000",
  6161=>"000000000",
  6162=>"111100111",
  6163=>"000000000",
  6164=>"101111111",
  6165=>"000111111",
  6166=>"000000000",
  6167=>"000000000",
  6168=>"000000000",
  6169=>"110000010",
  6170=>"000000000",
  6171=>"000000000",
  6172=>"000000100",
  6173=>"111111111",
  6174=>"111000000",
  6175=>"000000011",
  6176=>"110110111",
  6177=>"110100000",
  6178=>"001001111",
  6179=>"111111111",
  6180=>"000000001",
  6181=>"000000000",
  6182=>"111111111",
  6183=>"111110011",
  6184=>"101111111",
  6185=>"011011111",
  6186=>"000000000",
  6187=>"111101000",
  6188=>"111111000",
  6189=>"000001000",
  6190=>"111110110",
  6191=>"000011000",
  6192=>"001001001",
  6193=>"111001011",
  6194=>"100100100",
  6195=>"000111111",
  6196=>"110110011",
  6197=>"110111111",
  6198=>"111111000",
  6199=>"000000000",
  6200=>"111111111",
  6201=>"111100000",
  6202=>"111111111",
  6203=>"000000000",
  6204=>"111111111",
  6205=>"111111000",
  6206=>"111000001",
  6207=>"111111101",
  6208=>"111101111",
  6209=>"110110110",
  6210=>"101110111",
  6211=>"000000101",
  6212=>"100111111",
  6213=>"101000110",
  6214=>"000000111",
  6215=>"110111111",
  6216=>"111100110",
  6217=>"001001001",
  6218=>"010010110",
  6219=>"000111011",
  6220=>"111111111",
  6221=>"111111111",
  6222=>"000000100",
  6223=>"111111010",
  6224=>"011000000",
  6225=>"000000110",
  6226=>"111111111",
  6227=>"001001111",
  6228=>"111111111",
  6229=>"011111111",
  6230=>"111000000",
  6231=>"001000000",
  6232=>"000001111",
  6233=>"111000000",
  6234=>"111111111",
  6235=>"110011011",
  6236=>"111111001",
  6237=>"111111111",
  6238=>"011000000",
  6239=>"111111000",
  6240=>"111001000",
  6241=>"111111111",
  6242=>"011001001",
  6243=>"111001111",
  6244=>"001101111",
  6245=>"100111111",
  6246=>"000000000",
  6247=>"111111111",
  6248=>"000000000",
  6249=>"000000000",
  6250=>"000000000",
  6251=>"000000000",
  6252=>"011011000",
  6253=>"000000000",
  6254=>"111110000",
  6255=>"000101001",
  6256=>"000000000",
  6257=>"111111111",
  6258=>"110111111",
  6259=>"111000000",
  6260=>"011001000",
  6261=>"111011010",
  6262=>"010010000",
  6263=>"110110110",
  6264=>"111110110",
  6265=>"001000110",
  6266=>"000000000",
  6267=>"000000000",
  6268=>"110110110",
  6269=>"101000000",
  6270=>"000100111",
  6271=>"010110000",
  6272=>"000000000",
  6273=>"111111000",
  6274=>"000000000",
  6275=>"000000001",
  6276=>"000000000",
  6277=>"111111111",
  6278=>"011111110",
  6279=>"111001000",
  6280=>"110100000",
  6281=>"110110100",
  6282=>"000001111",
  6283=>"111100000",
  6284=>"111111111",
  6285=>"001000000",
  6286=>"001011100",
  6287=>"011001001",
  6288=>"101111111",
  6289=>"000000000",
  6290=>"000000111",
  6291=>"110111111",
  6292=>"000000000",
  6293=>"111111110",
  6294=>"000000111",
  6295=>"000100000",
  6296=>"000000000",
  6297=>"111101111",
  6298=>"000000000",
  6299=>"110111011",
  6300=>"000000000",
  6301=>"111110000",
  6302=>"111111111",
  6303=>"000011011",
  6304=>"000111111",
  6305=>"111010000",
  6306=>"000000011",
  6307=>"111110100",
  6308=>"000000000",
  6309=>"111111111",
  6310=>"111111001",
  6311=>"111111111",
  6312=>"001011111",
  6313=>"111101101",
  6314=>"000000000",
  6315=>"111111111",
  6316=>"000000100",
  6317=>"110111111",
  6318=>"000001111",
  6319=>"111101001",
  6320=>"111111000",
  6321=>"011101110",
  6322=>"111111111",
  6323=>"100100100",
  6324=>"110110011",
  6325=>"001111111",
  6326=>"111111111",
  6327=>"111000000",
  6328=>"111110111",
  6329=>"111111111",
  6330=>"000000000",
  6331=>"100000000",
  6332=>"000000000",
  6333=>"000100000",
  6334=>"000000000",
  6335=>"000000000",
  6336=>"000000000",
  6337=>"000000111",
  6338=>"000000100",
  6339=>"000000000",
  6340=>"111111111",
  6341=>"000000000",
  6342=>"000001000",
  6343=>"110111111",
  6344=>"000000000",
  6345=>"111111111",
  6346=>"001001101",
  6347=>"010000000",
  6348=>"111111111",
  6349=>"111111111",
  6350=>"110000000",
  6351=>"000000000",
  6352=>"111111111",
  6353=>"100000000",
  6354=>"111001101",
  6355=>"000000000",
  6356=>"001000000",
  6357=>"100100100",
  6358=>"111101111",
  6359=>"001000001",
  6360=>"111100111",
  6361=>"100100111",
  6362=>"001000111",
  6363=>"111111111",
  6364=>"001011010",
  6365=>"111111011",
  6366=>"111101000",
  6367=>"000000000",
  6368=>"000000000",
  6369=>"000010000",
  6370=>"000000001",
  6371=>"111000000",
  6372=>"111111101",
  6373=>"010011010",
  6374=>"100000111",
  6375=>"111111111",
  6376=>"111101111",
  6377=>"011011001",
  6378=>"000100111",
  6379=>"001000000",
  6380=>"111111111",
  6381=>"000000000",
  6382=>"000000100",
  6383=>"111111100",
  6384=>"000000000",
  6385=>"000000111",
  6386=>"000000000",
  6387=>"000000000",
  6388=>"111111010",
  6389=>"111111111",
  6390=>"000000001",
  6391=>"000111111",
  6392=>"000000000",
  6393=>"111101101",
  6394=>"001001111",
  6395=>"111111111",
  6396=>"000000000",
  6397=>"001001001",
  6398=>"111111111",
  6399=>"111001001",
  6400=>"000011000",
  6401=>"100000100",
  6402=>"000000000",
  6403=>"000000000",
  6404=>"000110100",
  6405=>"000000101",
  6406=>"001001001",
  6407=>"000001001",
  6408=>"000000000",
  6409=>"111111111",
  6410=>"011001011",
  6411=>"000000000",
  6412=>"111111011",
  6413=>"011011011",
  6414=>"100111111",
  6415=>"111111111",
  6416=>"111111111",
  6417=>"000000001",
  6418=>"111000111",
  6419=>"111111111",
  6420=>"000000000",
  6421=>"111111111",
  6422=>"011011001",
  6423=>"000000000",
  6424=>"000110110",
  6425=>"111110111",
  6426=>"101000000",
  6427=>"111111110",
  6428=>"111111111",
  6429=>"000000000",
  6430=>"110111111",
  6431=>"000101000",
  6432=>"111111001",
  6433=>"011011011",
  6434=>"111111111",
  6435=>"001001111",
  6436=>"000000000",
  6437=>"000000000",
  6438=>"111101111",
  6439=>"010111000",
  6440=>"111100100",
  6441=>"111111111",
  6442=>"111111101",
  6443=>"011011001",
  6444=>"001111111",
  6445=>"111111100",
  6446=>"000000000",
  6447=>"111111011",
  6448=>"000000000",
  6449=>"111111100",
  6450=>"000000000",
  6451=>"111001111",
  6452=>"000000000",
  6453=>"000000000",
  6454=>"001111010",
  6455=>"100100001",
  6456=>"000110000",
  6457=>"000000000",
  6458=>"011101111",
  6459=>"111111110",
  6460=>"000000000",
  6461=>"000101101",
  6462=>"111111111",
  6463=>"111111100",
  6464=>"111110111",
  6465=>"000010011",
  6466=>"100000000",
  6467=>"111011001",
  6468=>"111111111",
  6469=>"001111101",
  6470=>"000111111",
  6471=>"000000100",
  6472=>"100000000",
  6473=>"100000111",
  6474=>"110000000",
  6475=>"111111111",
  6476=>"001000000",
  6477=>"111111101",
  6478=>"011111111",
  6479=>"100000000",
  6480=>"111111111",
  6481=>"111111111",
  6482=>"000011111",
  6483=>"110100100",
  6484=>"000000000",
  6485=>"011011001",
  6486=>"111100111",
  6487=>"111111111",
  6488=>"111111111",
  6489=>"111111111",
  6490=>"000000101",
  6491=>"011010110",
  6492=>"000000001",
  6493=>"111111111",
  6494=>"111011111",
  6495=>"000000001",
  6496=>"000000010",
  6497=>"111111111",
  6498=>"111100011",
  6499=>"000000000",
  6500=>"000000010",
  6501=>"000000000",
  6502=>"100000100",
  6503=>"000100100",
  6504=>"111001101",
  6505=>"110000100",
  6506=>"000000000",
  6507=>"111101111",
  6508=>"110110100",
  6509=>"000110000",
  6510=>"111111111",
  6511=>"000000001",
  6512=>"000000100",
  6513=>"110000000",
  6514=>"111111111",
  6515=>"000100000",
  6516=>"111111000",
  6517=>"100100000",
  6518=>"110100100",
  6519=>"000111000",
  6520=>"111111111",
  6521=>"000000000",
  6522=>"111000000",
  6523=>"000000000",
  6524=>"000000000",
  6525=>"111111111",
  6526=>"000000000",
  6527=>"001000000",
  6528=>"000000000",
  6529=>"111111111",
  6530=>"000000001",
  6531=>"111011001",
  6532=>"001101100",
  6533=>"011111111",
  6534=>"001000110",
  6535=>"101001111",
  6536=>"001001111",
  6537=>"000000000",
  6538=>"011001000",
  6539=>"000000000",
  6540=>"111111111",
  6541=>"000110100",
  6542=>"000001001",
  6543=>"011011000",
  6544=>"000000001",
  6545=>"000000000",
  6546=>"111111111",
  6547=>"000000001",
  6548=>"000110110",
  6549=>"111111000",
  6550=>"101111111",
  6551=>"000100000",
  6552=>"111101000",
  6553=>"010011111",
  6554=>"110111111",
  6555=>"111111111",
  6556=>"000000000",
  6557=>"000110111",
  6558=>"000000111",
  6559=>"000110111",
  6560=>"110110110",
  6561=>"011111111",
  6562=>"001001111",
  6563=>"000111111",
  6564=>"001001111",
  6565=>"111111110",
  6566=>"111111111",
  6567=>"001111111",
  6568=>"110110000",
  6569=>"000000110",
  6570=>"111101111",
  6571=>"111111111",
  6572=>"010000111",
  6573=>"000010010",
  6574=>"110111111",
  6575=>"111111001",
  6576=>"110100101",
  6577=>"000111110",
  6578=>"111111001",
  6579=>"000000100",
  6580=>"000000000",
  6581=>"000001011",
  6582=>"100000101",
  6583=>"111111111",
  6584=>"110100111",
  6585=>"111111111",
  6586=>"000000110",
  6587=>"111001001",
  6588=>"000011000",
  6589=>"000111111",
  6590=>"010001000",
  6591=>"111111111",
  6592=>"111111011",
  6593=>"111110000",
  6594=>"000000000",
  6595=>"111111111",
  6596=>"111111111",
  6597=>"000000000",
  6598=>"000110110",
  6599=>"000101111",
  6600=>"000000000",
  6601=>"000111011",
  6602=>"000000000",
  6603=>"000000011",
  6604=>"000000000",
  6605=>"001000000",
  6606=>"100111101",
  6607=>"000000000",
  6608=>"110100000",
  6609=>"000000000",
  6610=>"000000000",
  6611=>"101000000",
  6612=>"110100100",
  6613=>"011001000",
  6614=>"001000111",
  6615=>"011010010",
  6616=>"111111111",
  6617=>"001000010",
  6618=>"011011000",
  6619=>"111111100",
  6620=>"000000001",
  6621=>"000001001",
  6622=>"000000010",
  6623=>"001001000",
  6624=>"111110110",
  6625=>"000000000",
  6626=>"111111110",
  6627=>"000100111",
  6628=>"001001001",
  6629=>"110110010",
  6630=>"011001001",
  6631=>"000000000",
  6632=>"000000110",
  6633=>"000010111",
  6634=>"000000000",
  6635=>"111100111",
  6636=>"101101011",
  6637=>"100110101",
  6638=>"001000100",
  6639=>"111111101",
  6640=>"000001000",
  6641=>"100111111",
  6642=>"000001000",
  6643=>"000000100",
  6644=>"000000000",
  6645=>"111111111",
  6646=>"000000000",
  6647=>"111100000",
  6648=>"000000111",
  6649=>"000100111",
  6650=>"111001001",
  6651=>"000000000",
  6652=>"000000000",
  6653=>"000111111",
  6654=>"111110100",
  6655=>"001111111",
  6656=>"000000000",
  6657=>"000000111",
  6658=>"111010111",
  6659=>"111111101",
  6660=>"011011000",
  6661=>"110111111",
  6662=>"111001001",
  6663=>"111111111",
  6664=>"000111110",
  6665=>"111111110",
  6666=>"111111111",
  6667=>"000111111",
  6668=>"100101101",
  6669=>"100111111",
  6670=>"000101001",
  6671=>"111111111",
  6672=>"001011111",
  6673=>"000111101",
  6674=>"000000000",
  6675=>"001001000",
  6676=>"000000100",
  6677=>"100100111",
  6678=>"000011111",
  6679=>"111111110",
  6680=>"111111101",
  6681=>"001101000",
  6682=>"000000110",
  6683=>"000100111",
  6684=>"001001111",
  6685=>"110111010",
  6686=>"111100110",
  6687=>"000000111",
  6688=>"011111011",
  6689=>"000111111",
  6690=>"011101111",
  6691=>"111000000",
  6692=>"111111111",
  6693=>"111111100",
  6694=>"000000000",
  6695=>"011001000",
  6696=>"000000000",
  6697=>"111000000",
  6698=>"011001101",
  6699=>"000000111",
  6700=>"100101101",
  6701=>"111111111",
  6702=>"110110010",
  6703=>"100000000",
  6704=>"111110000",
  6705=>"100101000",
  6706=>"100101111",
  6707=>"111010111",
  6708=>"101000000",
  6709=>"110110000",
  6710=>"000000101",
  6711=>"010000110",
  6712=>"000001001",
  6713=>"001001000",
  6714=>"111111000",
  6715=>"000001000",
  6716=>"001000000",
  6717=>"011011000",
  6718=>"111111111",
  6719=>"011111000",
  6720=>"111011111",
  6721=>"111111100",
  6722=>"101000100",
  6723=>"000000000",
  6724=>"001000000",
  6725=>"110110000",
  6726=>"111000111",
  6727=>"000010000",
  6728=>"000000110",
  6729=>"000000101",
  6730=>"111111111",
  6731=>"001001101",
  6732=>"110110110",
  6733=>"000000001",
  6734=>"011011001",
  6735=>"001111111",
  6736=>"110111111",
  6737=>"000000000",
  6738=>"011011111",
  6739=>"110110110",
  6740=>"000010000",
  6741=>"101100000",
  6742=>"001001001",
  6743=>"111111110",
  6744=>"100100000",
  6745=>"000000111",
  6746=>"010110000",
  6747=>"111111111",
  6748=>"000000000",
  6749=>"000000000",
  6750=>"001101001",
  6751=>"011110100",
  6752=>"001001111",
  6753=>"001001000",
  6754=>"000000011",
  6755=>"000000000",
  6756=>"011000000",
  6757=>"111001001",
  6758=>"111111000",
  6759=>"101000000",
  6760=>"101000000",
  6761=>"111111111",
  6762=>"000000111",
  6763=>"111101101",
  6764=>"111101011",
  6765=>"111111111",
  6766=>"001001001",
  6767=>"111111111",
  6768=>"001001001",
  6769=>"010110111",
  6770=>"111110000",
  6771=>"111011011",
  6772=>"011011011",
  6773=>"111111111",
  6774=>"101111111",
  6775=>"001001000",
  6776=>"011011000",
  6777=>"000000000",
  6778=>"111111000",
  6779=>"000000000",
  6780=>"100101100",
  6781=>"111111000",
  6782=>"010100110",
  6783=>"110111110",
  6784=>"100000100",
  6785=>"111101010",
  6786=>"111000111",
  6787=>"100000000",
  6788=>"001000011",
  6789=>"000000000",
  6790=>"000000000",
  6791=>"111111011",
  6792=>"101111111",
  6793=>"110110110",
  6794=>"000000111",
  6795=>"000001111",
  6796=>"011000000",
  6797=>"000000000",
  6798=>"111111111",
  6799=>"011111111",
  6800=>"000000000",
  6801=>"110110110",
  6802=>"001011001",
  6803=>"111111111",
  6804=>"000000100",
  6805=>"001111111",
  6806=>"111111111",
  6807=>"000110111",
  6808=>"011111111",
  6809=>"101101111",
  6810=>"011111111",
  6811=>"110000000",
  6812=>"000000000",
  6813=>"011001001",
  6814=>"000000000",
  6815=>"000000000",
  6816=>"111111111",
  6817=>"000000000",
  6818=>"000000000",
  6819=>"110110110",
  6820=>"110110000",
  6821=>"110111111",
  6822=>"000110000",
  6823=>"100110110",
  6824=>"110101111",
  6825=>"111001001",
  6826=>"111111111",
  6827=>"111111010",
  6828=>"110010000",
  6829=>"111110111",
  6830=>"111100000",
  6831=>"000000111",
  6832=>"010110000",
  6833=>"111111111",
  6834=>"110111110",
  6835=>"111111111",
  6836=>"111111110",
  6837=>"111001001",
  6838=>"000000000",
  6839=>"111100000",
  6840=>"001000000",
  6841=>"101001000",
  6842=>"111011000",
  6843=>"000001001",
  6844=>"101100101",
  6845=>"011100101",
  6846=>"001000101",
  6847=>"000000000",
  6848=>"001000000",
  6849=>"001001001",
  6850=>"111111111",
  6851=>"000000110",
  6852=>"011000011",
  6853=>"111011011",
  6854=>"000000000",
  6855=>"001100000",
  6856=>"000000111",
  6857=>"000000001",
  6858=>"001000001",
  6859=>"111100000",
  6860=>"000100110",
  6861=>"000011110",
  6862=>"111101000",
  6863=>"011000000",
  6864=>"111001000",
  6865=>"011101111",
  6866=>"111110010",
  6867=>"110101000",
  6868=>"101110110",
  6869=>"100000001",
  6870=>"100100000",
  6871=>"101100100",
  6872=>"111111111",
  6873=>"000000101",
  6874=>"001000000",
  6875=>"000111111",
  6876=>"111001000",
  6877=>"110111110",
  6878=>"010110010",
  6879=>"010000000",
  6880=>"001001000",
  6881=>"000000000",
  6882=>"111111000",
  6883=>"110000000",
  6884=>"100000100",
  6885=>"101101100",
  6886=>"001101000",
  6887=>"000111111",
  6888=>"000000001",
  6889=>"000000000",
  6890=>"111001111",
  6891=>"000000001",
  6892=>"111111100",
  6893=>"111110111",
  6894=>"101110111",
  6895=>"000011111",
  6896=>"111111111",
  6897=>"001000001",
  6898=>"000000111",
  6899=>"010010000",
  6900=>"000110000",
  6901=>"011000110",
  6902=>"001000000",
  6903=>"011110110",
  6904=>"101000000",
  6905=>"000000101",
  6906=>"110110000",
  6907=>"000101111",
  6908=>"011000000",
  6909=>"110011011",
  6910=>"000000000",
  6911=>"001001000",
  6912=>"110111011",
  6913=>"101001011",
  6914=>"011001111",
  6915=>"111000000",
  6916=>"001001001",
  6917=>"000000110",
  6918=>"000000111",
  6919=>"111111111",
  6920=>"000000000",
  6921=>"001101101",
  6922=>"111000000",
  6923=>"000000001",
  6924=>"000000000",
  6925=>"010111110",
  6926=>"000000000",
  6927=>"001001010",
  6928=>"111011111",
  6929=>"110000000",
  6930=>"000010000",
  6931=>"000011011",
  6932=>"100000100",
  6933=>"000000011",
  6934=>"100110111",
  6935=>"111111100",
  6936=>"111000000",
  6937=>"111110111",
  6938=>"011000000",
  6939=>"011111111",
  6940=>"000100100",
  6941=>"011000110",
  6942=>"101100111",
  6943=>"000010111",
  6944=>"100110000",
  6945=>"000000000",
  6946=>"000110111",
  6947=>"111111011",
  6948=>"000000011",
  6949=>"010000111",
  6950=>"000001110",
  6951=>"000011000",
  6952=>"110111001",
  6953=>"111111111",
  6954=>"011111001",
  6955=>"001001000",
  6956=>"011011110",
  6957=>"110110110",
  6958=>"111111111",
  6959=>"000000001",
  6960=>"110110110",
  6961=>"000110000",
  6962=>"000000000",
  6963=>"111111000",
  6964=>"000000010",
  6965=>"011011001",
  6966=>"110111111",
  6967=>"111001101",
  6968=>"111110110",
  6969=>"001000000",
  6970=>"000001001",
  6971=>"000011011",
  6972=>"111111100",
  6973=>"000000000",
  6974=>"110111110",
  6975=>"111111111",
  6976=>"000000000",
  6977=>"000000000",
  6978=>"001011000",
  6979=>"111001001",
  6980=>"111000000",
  6981=>"000100101",
  6982=>"000000000",
  6983=>"111111111",
  6984=>"000000000",
  6985=>"001101111",
  6986=>"111111111",
  6987=>"111000000",
  6988=>"011001000",
  6989=>"101000111",
  6990=>"000101111",
  6991=>"111110100",
  6992=>"000000000",
  6993=>"000111111",
  6994=>"110100000",
  6995=>"000000000",
  6996=>"000000000",
  6997=>"011011011",
  6998=>"111110000",
  6999=>"111001001",
  7000=>"001011010",
  7001=>"000110111",
  7002=>"001000000",
  7003=>"010000000",
  7004=>"110110110",
  7005=>"010000001",
  7006=>"110000111",
  7007=>"000101001",
  7008=>"111111001",
  7009=>"000000000",
  7010=>"111101001",
  7011=>"000000000",
  7012=>"111111111",
  7013=>"000000000",
  7014=>"111111111",
  7015=>"000000000",
  7016=>"001000000",
  7017=>"001001001",
  7018=>"000000001",
  7019=>"000000000",
  7020=>"111110110",
  7021=>"111111000",
  7022=>"001000000",
  7023=>"110000001",
  7024=>"000001011",
  7025=>"000000000",
  7026=>"010000000",
  7027=>"111111110",
  7028=>"000000001",
  7029=>"111111111",
  7030=>"000000111",
  7031=>"111000010",
  7032=>"111011111",
  7033=>"000000000",
  7034=>"000000000",
  7035=>"111111111",
  7036=>"111011000",
  7037=>"000000001",
  7038=>"010000010",
  7039=>"100000101",
  7040=>"011011111",
  7041=>"001000000",
  7042=>"111100100",
  7043=>"000000001",
  7044=>"111111111",
  7045=>"000111010",
  7046=>"000001111",
  7047=>"111111011",
  7048=>"110000000",
  7049=>"111111111",
  7050=>"110111110",
  7051=>"000000111",
  7052=>"110110111",
  7053=>"111101100",
  7054=>"110110000",
  7055=>"001000000",
  7056=>"000110000",
  7057=>"111111111",
  7058=>"111111110",
  7059=>"000001001",
  7060=>"111111111",
  7061=>"010011000",
  7062=>"111111111",
  7063=>"111110000",
  7064=>"000000001",
  7065=>"111111011",
  7066=>"001000100",
  7067=>"111000000",
  7068=>"000000000",
  7069=>"000000000",
  7070=>"100110100",
  7071=>"000000101",
  7072=>"000100011",
  7073=>"011011111",
  7074=>"000000000",
  7075=>"100110110",
  7076=>"111111101",
  7077=>"000000110",
  7078=>"101001001",
  7079=>"001111111",
  7080=>"101000100",
  7081=>"000000111",
  7082=>"111111111",
  7083=>"000000100",
  7084=>"000010110",
  7085=>"011111111",
  7086=>"000000000",
  7087=>"000000000",
  7088=>"011011111",
  7089=>"000001011",
  7090=>"000000001",
  7091=>"000000000",
  7092=>"001001001",
  7093=>"111000000",
  7094=>"001111111",
  7095=>"001001101",
  7096=>"111111000",
  7097=>"111111111",
  7098=>"011011111",
  7099=>"000000011",
  7100=>"111100000",
  7101=>"111111111",
  7102=>"001000111",
  7103=>"000000000",
  7104=>"111110010",
  7105=>"110110110",
  7106=>"001101111",
  7107=>"000000000",
  7108=>"000000111",
  7109=>"001000100",
  7110=>"001000001",
  7111=>"101100110",
  7112=>"010000000",
  7113=>"010010011",
  7114=>"111000000",
  7115=>"000000000",
  7116=>"111111000",
  7117=>"101101000",
  7118=>"111000000",
  7119=>"000011011",
  7120=>"000000111",
  7121=>"111111000",
  7122=>"101101101",
  7123=>"011000101",
  7124=>"111110111",
  7125=>"000100111",
  7126=>"000100110",
  7127=>"100000000",
  7128=>"111111000",
  7129=>"001001000",
  7130=>"000001001",
  7131=>"010011111",
  7132=>"110111111",
  7133=>"001001101",
  7134=>"111111111",
  7135=>"000000010",
  7136=>"000111111",
  7137=>"111001001",
  7138=>"111001111",
  7139=>"001000000",
  7140=>"001111111",
  7141=>"000000110",
  7142=>"000010000",
  7143=>"111011011",
  7144=>"001000000",
  7145=>"000000000",
  7146=>"000000010",
  7147=>"110110110",
  7148=>"000000000",
  7149=>"111111100",
  7150=>"000000111",
  7151=>"110111110",
  7152=>"110111101",
  7153=>"000100111",
  7154=>"111000100",
  7155=>"111111000",
  7156=>"110000000",
  7157=>"000000111",
  7158=>"001001001",
  7159=>"000000000",
  7160=>"000000000",
  7161=>"100000000",
  7162=>"111001001",
  7163=>"001000000",
  7164=>"001001000",
  7165=>"001001000",
  7166=>"010000000",
  7167=>"001000100",
  7168=>"001111111",
  7169=>"111111011",
  7170=>"000000111",
  7171=>"111111111",
  7172=>"110111110",
  7173=>"011110010",
  7174=>"010111111",
  7175=>"000000111",
  7176=>"000000000",
  7177=>"010010010",
  7178=>"111111111",
  7179=>"011010010",
  7180=>"100110110",
  7181=>"111111011",
  7182=>"111111001",
  7183=>"000000000",
  7184=>"111111111",
  7185=>"000111111",
  7186=>"010111000",
  7187=>"010111111",
  7188=>"001101111",
  7189=>"011000111",
  7190=>"111111111",
  7191=>"010010111",
  7192=>"110110110",
  7193=>"001110110",
  7194=>"000001000",
  7195=>"111011000",
  7196=>"111110000",
  7197=>"010111111",
  7198=>"100000000",
  7199=>"000111111",
  7200=>"110110110",
  7201=>"110110111",
  7202=>"110110110",
  7203=>"110111010",
  7204=>"001000000",
  7205=>"111111000",
  7206=>"111111000",
  7207=>"000111000",
  7208=>"000000000",
  7209=>"000000000",
  7210=>"110111011",
  7211=>"000000111",
  7212=>"000110110",
  7213=>"011111111",
  7214=>"101001001",
  7215=>"111111111",
  7216=>"000000000",
  7217=>"000000111",
  7218=>"111111001",
  7219=>"111111111",
  7220=>"001001000",
  7221=>"000000000",
  7222=>"000000001",
  7223=>"001000000",
  7224=>"111111011",
  7225=>"000010000",
  7226=>"010000000",
  7227=>"001111111",
  7228=>"000000000",
  7229=>"000000000",
  7230=>"111111111",
  7231=>"000000100",
  7232=>"101111110",
  7233=>"000111001",
  7234=>"000000111",
  7235=>"000000001",
  7236=>"100110100",
  7237=>"100100111",
  7238=>"111000000",
  7239=>"000000111",
  7240=>"011111001",
  7241=>"010010010",
  7242=>"010111101",
  7243=>"010110111",
  7244=>"000000111",
  7245=>"111001001",
  7246=>"001000100",
  7247=>"000000000",
  7248=>"000000000",
  7249=>"101111110",
  7250=>"111111000",
  7251=>"001000000",
  7252=>"001001111",
  7253=>"100111111",
  7254=>"100000000",
  7255=>"111111100",
  7256=>"001000001",
  7257=>"000000101",
  7258=>"110111111",
  7259=>"100011001",
  7260=>"001001001",
  7261=>"111001111",
  7262=>"010110111",
  7263=>"000000001",
  7264=>"001001101",
  7265=>"111001000",
  7266=>"111111111",
  7267=>"111101111",
  7268=>"110110010",
  7269=>"001000000",
  7270=>"111110000",
  7271=>"111111000",
  7272=>"111111111",
  7273=>"111000000",
  7274=>"000000000",
  7275=>"000000000",
  7276=>"110110000",
  7277=>"000000000",
  7278=>"111111111",
  7279=>"000010000",
  7280=>"111000010",
  7281=>"000000001",
  7282=>"111111011",
  7283=>"000000111",
  7284=>"111111000",
  7285=>"100001001",
  7286=>"000000111",
  7287=>"111111111",
  7288=>"111000010",
  7289=>"000000000",
  7290=>"101000001",
  7291=>"000000000",
  7292=>"011001001",
  7293=>"111111111",
  7294=>"000000000",
  7295=>"000000000",
  7296=>"111111101",
  7297=>"111111011",
  7298=>"000000000",
  7299=>"000111010",
  7300=>"111111010",
  7301=>"000000000",
  7302=>"000000111",
  7303=>"111101111",
  7304=>"000010111",
  7305=>"000111111",
  7306=>"110111110",
  7307=>"111111000",
  7308=>"111111110",
  7309=>"110000000",
  7310=>"110111001",
  7311=>"000100100",
  7312=>"000000101",
  7313=>"001000001",
  7314=>"111111111",
  7315=>"111001000",
  7316=>"110001000",
  7317=>"001000001",
  7318=>"110110110",
  7319=>"000000000",
  7320=>"101001111",
  7321=>"000000111",
  7322=>"000010111",
  7323=>"111111111",
  7324=>"010011000",
  7325=>"011000001",
  7326=>"000110111",
  7327=>"000001000",
  7328=>"111111110",
  7329=>"000111111",
  7330=>"011111111",
  7331=>"111001011",
  7332=>"011000001",
  7333=>"000111011",
  7334=>"001001000",
  7335=>"100100100",
  7336=>"000000111",
  7337=>"101000001",
  7338=>"100100111",
  7339=>"111000101",
  7340=>"101000000",
  7341=>"100101111",
  7342=>"000001111",
  7343=>"000000001",
  7344=>"000000001",
  7345=>"011011000",
  7346=>"010111010",
  7347=>"101001100",
  7348=>"100000110",
  7349=>"101101111",
  7350=>"000101100",
  7351=>"100010000",
  7352=>"000000000",
  7353=>"110111110",
  7354=>"111000000",
  7355=>"000101111",
  7356=>"111100000",
  7357=>"111111111",
  7358=>"101100100",
  7359=>"000000000",
  7360=>"000000000",
  7361=>"001000000",
  7362=>"111100110",
  7363=>"010110000",
  7364=>"001001101",
  7365=>"000000110",
  7366=>"111000111",
  7367=>"100000001",
  7368=>"000000000",
  7369=>"000000101",
  7370=>"000000100",
  7371=>"000000000",
  7372=>"000000101",
  7373=>"001101000",
  7374=>"000000001",
  7375=>"000000000",
  7376=>"111000000",
  7377=>"001001000",
  7378=>"111100100",
  7379=>"001001001",
  7380=>"000000000",
  7381=>"001000000",
  7382=>"101001111",
  7383=>"000000001",
  7384=>"000000111",
  7385=>"111110111",
  7386=>"111111110",
  7387=>"000010111",
  7388=>"111101101",
  7389=>"001001001",
  7390=>"101000000",
  7391=>"000001111",
  7392=>"000001011",
  7393=>"010010000",
  7394=>"011111111",
  7395=>"000000110",
  7396=>"000100111",
  7397=>"100110100",
  7398=>"101111111",
  7399=>"111111010",
  7400=>"111111000",
  7401=>"000000000",
  7402=>"000101111",
  7403=>"111010000",
  7404=>"000000000",
  7405=>"111011001",
  7406=>"111111111",
  7407=>"111111111",
  7408=>"110011001",
  7409=>"101100100",
  7410=>"010000001",
  7411=>"101001011",
  7412=>"111111110",
  7413=>"001000100",
  7414=>"011000000",
  7415=>"011000000",
  7416=>"110110000",
  7417=>"000010000",
  7418=>"000001101",
  7419=>"001001111",
  7420=>"000110111",
  7421=>"001001000",
  7422=>"101111011",
  7423=>"000000000",
  7424=>"110111110",
  7425=>"101000000",
  7426=>"111111111",
  7427=>"110110000",
  7428=>"000000101",
  7429=>"010100000",
  7430=>"110000010",
  7431=>"000000001",
  7432=>"000000000",
  7433=>"111001001",
  7434=>"000000000",
  7435=>"110011111",
  7436=>"000000100",
  7437=>"111110111",
  7438=>"000000111",
  7439=>"010010000",
  7440=>"000100100",
  7441=>"000111111",
  7442=>"000000000",
  7443=>"001000000",
  7444=>"010000111",
  7445=>"010111111",
  7446=>"111101101",
  7447=>"000001001",
  7448=>"000000111",
  7449=>"000100111",
  7450=>"000000000",
  7451=>"111000000",
  7452=>"110110000",
  7453=>"111111111",
  7454=>"000000000",
  7455=>"000000100",
  7456=>"000000000",
  7457=>"011111111",
  7458=>"000010111",
  7459=>"111110110",
  7460=>"011011001",
  7461=>"000100111",
  7462=>"011111011",
  7463=>"100000101",
  7464=>"000000101",
  7465=>"110111010",
  7466=>"001000000",
  7467=>"000000111",
  7468=>"111101111",
  7469=>"000000001",
  7470=>"011111110",
  7471=>"000101111",
  7472=>"000000111",
  7473=>"100100000",
  7474=>"001000000",
  7475=>"111111111",
  7476=>"111111111",
  7477=>"011011001",
  7478=>"011011111",
  7479=>"001001001",
  7480=>"010010011",
  7481=>"101000000",
  7482=>"000000101",
  7483=>"111000000",
  7484=>"000011111",
  7485=>"110001000",
  7486=>"000100101",
  7487=>"000000100",
  7488=>"100100100",
  7489=>"000000011",
  7490=>"000110010",
  7491=>"001001011",
  7492=>"000000000",
  7493=>"000000111",
  7494=>"000111111",
  7495=>"110110000",
  7496=>"111101101",
  7497=>"111000000",
  7498=>"000111111",
  7499=>"000000000",
  7500=>"111011111",
  7501=>"111001001",
  7502=>"111000000",
  7503=>"100110110",
  7504=>"111110110",
  7505=>"111111001",
  7506=>"111010000",
  7507=>"110010010",
  7508=>"111111110",
  7509=>"001011001",
  7510=>"001000001",
  7511=>"111111111",
  7512=>"110110111",
  7513=>"111111111",
  7514=>"100111111",
  7515=>"000000101",
  7516=>"110001000",
  7517=>"100000000",
  7518=>"110110100",
  7519=>"000110110",
  7520=>"101111101",
  7521=>"100000000",
  7522=>"100000000",
  7523=>"101000000",
  7524=>"110110000",
  7525=>"001000000",
  7526=>"011010111",
  7527=>"111111000",
  7528=>"111101111",
  7529=>"000000011",
  7530=>"111001000",
  7531=>"011000110",
  7532=>"000000000",
  7533=>"111111110",
  7534=>"110111010",
  7535=>"111101111",
  7536=>"011111111",
  7537=>"101001001",
  7538=>"101000001",
  7539=>"000110111",
  7540=>"000000000",
  7541=>"111111000",
  7542=>"001111001",
  7543=>"111111000",
  7544=>"101000000",
  7545=>"001001000",
  7546=>"000000101",
  7547=>"111000000",
  7548=>"000100111",
  7549=>"000000000",
  7550=>"111110110",
  7551=>"000000101",
  7552=>"000000100",
  7553=>"001010101",
  7554=>"100111111",
  7555=>"000000100",
  7556=>"101111111",
  7557=>"010010010",
  7558=>"100001001",
  7559=>"011111111",
  7560=>"111111111",
  7561=>"000000000",
  7562=>"000100110",
  7563=>"111110010",
  7564=>"001000001",
  7565=>"100110100",
  7566=>"111111110",
  7567=>"000000000",
  7568=>"110010000",
  7569=>"000000111",
  7570=>"100101111",
  7571=>"000000001",
  7572=>"000000110",
  7573=>"000000000",
  7574=>"000000001",
  7575=>"001001011",
  7576=>"110111111",
  7577=>"111100100",
  7578=>"001010000",
  7579=>"000001111",
  7580=>"110111111",
  7581=>"000000000",
  7582=>"101001001",
  7583=>"111000000",
  7584=>"001000000",
  7585=>"110000111",
  7586=>"010110010",
  7587=>"000000111",
  7588=>"000000001",
  7589=>"001001001",
  7590=>"111101100",
  7591=>"110000000",
  7592=>"111111000",
  7593=>"111110011",
  7594=>"110111110",
  7595=>"001001011",
  7596=>"000000000",
  7597=>"000000000",
  7598=>"101001101",
  7599=>"000000000",
  7600=>"101100111",
  7601=>"000000000",
  7602=>"111111101",
  7603=>"000000110",
  7604=>"101111011",
  7605=>"000100111",
  7606=>"111011111",
  7607=>"110110000",
  7608=>"000001011",
  7609=>"111110110",
  7610=>"111111110",
  7611=>"000000111",
  7612=>"111111101",
  7613=>"110111111",
  7614=>"011111111",
  7615=>"111111111",
  7616=>"100110110",
  7617=>"100110100",
  7618=>"110111111",
  7619=>"001001000",
  7620=>"000000000",
  7621=>"000000000",
  7622=>"000000001",
  7623=>"000000111",
  7624=>"000000111",
  7625=>"000000100",
  7626=>"111111011",
  7627=>"111111111",
  7628=>"111001111",
  7629=>"010110110",
  7630=>"000111111",
  7631=>"001001011",
  7632=>"111111111",
  7633=>"000000000",
  7634=>"010000110",
  7635=>"111111111",
  7636=>"001000000",
  7637=>"100101001",
  7638=>"111111111",
  7639=>"010111011",
  7640=>"000111111",
  7641=>"000000010",
  7642=>"101000000",
  7643=>"001111010",
  7644=>"000000000",
  7645=>"100100001",
  7646=>"000011011",
  7647=>"000001111",
  7648=>"110110111",
  7649=>"000000000",
  7650=>"000000000",
  7651=>"111111000",
  7652=>"111100100",
  7653=>"100111111",
  7654=>"000000000",
  7655=>"001000111",
  7656=>"101111001",
  7657=>"000111111",
  7658=>"111000000",
  7659=>"110011011",
  7660=>"010111111",
  7661=>"011011001",
  7662=>"111111111",
  7663=>"001010110",
  7664=>"111000100",
  7665=>"011110111",
  7666=>"000011011",
  7667=>"111111111",
  7668=>"010110010",
  7669=>"001101000",
  7670=>"111111100",
  7671=>"111100100",
  7672=>"110111111",
  7673=>"100110110",
  7674=>"000000000",
  7675=>"000000001",
  7676=>"110110000",
  7677=>"111011011",
  7678=>"011000100",
  7679=>"001111111",
  7680=>"000100110",
  7681=>"000000000",
  7682=>"111000000",
  7683=>"000000111",
  7684=>"011000000",
  7685=>"111000000",
  7686=>"111001000",
  7687=>"111000111",
  7688=>"011010010",
  7689=>"111110100",
  7690=>"001000000",
  7691=>"000111100",
  7692=>"001001001",
  7693=>"101001100",
  7694=>"000000100",
  7695=>"101001001",
  7696=>"100111000",
  7697=>"110000000",
  7698=>"001000110",
  7699=>"000000000",
  7700=>"110111111",
  7701=>"001001000",
  7702=>"001000000",
  7703=>"011111111",
  7704=>"110110110",
  7705=>"111000000",
  7706=>"001101101",
  7707=>"111011011",
  7708=>"111111111",
  7709=>"111000001",
  7710=>"000000100",
  7711=>"000000000",
  7712=>"000001001",
  7713=>"111001101",
  7714=>"011111111",
  7715=>"110111111",
  7716=>"000111111",
  7717=>"000000100",
  7718=>"011001000",
  7719=>"011011001",
  7720=>"111100100",
  7721=>"111000100",
  7722=>"000000000",
  7723=>"001001000",
  7724=>"000111100",
  7725=>"111010000",
  7726=>"011001000",
  7727=>"011001001",
  7728=>"000000011",
  7729=>"111100000",
  7730=>"111111111",
  7731=>"000000000",
  7732=>"000001001",
  7733=>"111001000",
  7734=>"111111001",
  7735=>"000100000",
  7736=>"001100111",
  7737=>"101000111",
  7738=>"001000001",
  7739=>"111000000",
  7740=>"111101101",
  7741=>"001000000",
  7742=>"001001000",
  7743=>"101001000",
  7744=>"111111111",
  7745=>"001001001",
  7746=>"000111111",
  7747=>"000001011",
  7748=>"100000011",
  7749=>"000011000",
  7750=>"000000110",
  7751=>"000000111",
  7752=>"001000000",
  7753=>"001000001",
  7754=>"111111111",
  7755=>"111111011",
  7756=>"000000000",
  7757=>"110111111",
  7758=>"011000000",
  7759=>"111110100",
  7760=>"001000010",
  7761=>"011000000",
  7762=>"100000000",
  7763=>"001000000",
  7764=>"001001000",
  7765=>"111101000",
  7766=>"111100000",
  7767=>"110111110",
  7768=>"011001001",
  7769=>"001001001",
  7770=>"011010010",
  7771=>"000000011",
  7772=>"110111111",
  7773=>"111111111",
  7774=>"110101010",
  7775=>"111111101",
  7776=>"111001001",
  7777=>"001001100",
  7778=>"000000000",
  7779=>"100100000",
  7780=>"001000111",
  7781=>"111001001",
  7782=>"111111111",
  7783=>"001001001",
  7784=>"000001111",
  7785=>"100100001",
  7786=>"000000100",
  7787=>"000000000",
  7788=>"000000001",
  7789=>"001001101",
  7790=>"111001000",
  7791=>"110110100",
  7792=>"000000000",
  7793=>"011101111",
  7794=>"011000000",
  7795=>"100100100",
  7796=>"000110000",
  7797=>"100111111",
  7798=>"111001111",
  7799=>"000000010",
  7800=>"000000000",
  7801=>"010111111",
  7802=>"110010000",
  7803=>"111001000",
  7804=>"000001000",
  7805=>"110001000",
  7806=>"111110000",
  7807=>"000000000",
  7808=>"111000000",
  7809=>"111111000",
  7810=>"111000000",
  7811=>"111111111",
  7812=>"101111111",
  7813=>"001001111",
  7814=>"001111111",
  7815=>"111110111",
  7816=>"111111111",
  7817=>"000111111",
  7818=>"000000000",
  7819=>"001001001",
  7820=>"111111111",
  7821=>"001001000",
  7822=>"011001101",
  7823=>"000000000",
  7824=>"000000000",
  7825=>"001000000",
  7826=>"100110011",
  7827=>"101111111",
  7828=>"101111100",
  7829=>"011011001",
  7830=>"110111111",
  7831=>"000000001",
  7832=>"111001101",
  7833=>"001111111",
  7834=>"011011011",
  7835=>"000000000",
  7836=>"001111111",
  7837=>"110100000",
  7838=>"001000100",
  7839=>"000010111",
  7840=>"111111111",
  7841=>"011010100",
  7842=>"101101101",
  7843=>"000010110",
  7844=>"111110010",
  7845=>"001001000",
  7846=>"001111101",
  7847=>"001000001",
  7848=>"011011001",
  7849=>"001000000",
  7850=>"010111111",
  7851=>"111001001",
  7852=>"000000001",
  7853=>"000000011",
  7854=>"011001001",
  7855=>"000011111",
  7856=>"000011111",
  7857=>"001111110",
  7858=>"010111011",
  7859=>"111111011",
  7860=>"011110000",
  7861=>"001000000",
  7862=>"111101111",
  7863=>"000000100",
  7864=>"011111011",
  7865=>"000000100",
  7866=>"110000001",
  7867=>"000000000",
  7868=>"000000000",
  7869=>"111111111",
  7870=>"110000000",
  7871=>"110110111",
  7872=>"001001001",
  7873=>"111111111",
  7874=>"000000000",
  7875=>"111111010",
  7876=>"101111101",
  7877=>"111111001",
  7878=>"101000000",
  7879=>"001000001",
  7880=>"111111111",
  7881=>"000000000",
  7882=>"000000000",
  7883=>"011011010",
  7884=>"111111111",
  7885=>"000000000",
  7886=>"000010111",
  7887=>"000000000",
  7888=>"000000000",
  7889=>"000010000",
  7890=>"100111111",
  7891=>"000000000",
  7892=>"001000101",
  7893=>"110110110",
  7894=>"010010000",
  7895=>"111011000",
  7896=>"000000001",
  7897=>"111011001",
  7898=>"000000111",
  7899=>"100001001",
  7900=>"001000000",
  7901=>"110111110",
  7902=>"011011111",
  7903=>"101100111",
  7904=>"000111001",
  7905=>"000000110",
  7906=>"011111111",
  7907=>"001001000",
  7908=>"010010000",
  7909=>"001000001",
  7910=>"101111111",
  7911=>"011001000",
  7912=>"000000010",
  7913=>"110000000",
  7914=>"000000111",
  7915=>"000000000",
  7916=>"110000001",
  7917=>"100110111",
  7918=>"110111111",
  7919=>"000000001",
  7920=>"000111111",
  7921=>"111111111",
  7922=>"100111011",
  7923=>"000000000",
  7924=>"000000100",
  7925=>"100100111",
  7926=>"001000000",
  7927=>"000000000",
  7928=>"111101111",
  7929=>"000011000",
  7930=>"111111101",
  7931=>"000100001",
  7932=>"010111110",
  7933=>"101001000",
  7934=>"111110110",
  7935=>"011011111",
  7936=>"000000100",
  7937=>"000001001",
  7938=>"001000101",
  7939=>"110110111",
  7940=>"110100110",
  7941=>"001001111",
  7942=>"000000001",
  7943=>"111000000",
  7944=>"000000010",
  7945=>"000001000",
  7946=>"111101000",
  7947=>"000001111",
  7948=>"000000100",
  7949=>"010111111",
  7950=>"111010010",
  7951=>"010011011",
  7952=>"111110010",
  7953=>"101000100",
  7954=>"111111111",
  7955=>"000000000",
  7956=>"011111110",
  7957=>"110000000",
  7958=>"001001101",
  7959=>"111111110",
  7960=>"011111101",
  7961=>"100000000",
  7962=>"011000000",
  7963=>"011111111",
  7964=>"000001001",
  7965=>"111001101",
  7966=>"000000000",
  7967=>"111011101",
  7968=>"111001001",
  7969=>"010111110",
  7970=>"010010000",
  7971=>"100110111",
  7972=>"100110110",
  7973=>"000000000",
  7974=>"000000100",
  7975=>"011111000",
  7976=>"110110010",
  7977=>"000011010",
  7978=>"000001100",
  7979=>"110110000",
  7980=>"001000110",
  7981=>"010000000",
  7982=>"000010010",
  7983=>"011001001",
  7984=>"011001101",
  7985=>"000000000",
  7986=>"000000000",
  7987=>"000000000",
  7988=>"000000110",
  7989=>"001001001",
  7990=>"011111111",
  7991=>"000000101",
  7992=>"011000000",
  7993=>"101000000",
  7994=>"111000011",
  7995=>"110000001",
  7996=>"010000001",
  7997=>"001000000",
  7998=>"100010011",
  7999=>"111111011",
  8000=>"000101111",
  8001=>"111110111",
  8002=>"000000001",
  8003=>"111111110",
  8004=>"001101000",
  8005=>"000110111",
  8006=>"000000010",
  8007=>"000000000",
  8008=>"000000000",
  8009=>"000110111",
  8010=>"000000000",
  8011=>"011011001",
  8012=>"000100000",
  8013=>"000111111",
  8014=>"011011111",
  8015=>"110111111",
  8016=>"011011011",
  8017=>"111000000",
  8018=>"100010000",
  8019=>"001001001",
  8020=>"001001000",
  8021=>"011011011",
  8022=>"000000000",
  8023=>"111101101",
  8024=>"001000000",
  8025=>"111111001",
  8026=>"111111010",
  8027=>"110000000",
  8028=>"110111111",
  8029=>"001001000",
  8030=>"010000011",
  8031=>"000000000",
  8032=>"010110111",
  8033=>"111111111",
  8034=>"111011011",
  8035=>"000111111",
  8036=>"000111100",
  8037=>"000000000",
  8038=>"110111111",
  8039=>"000000000",
  8040=>"000000000",
  8041=>"111111111",
  8042=>"001001001",
  8043=>"111111101",
  8044=>"000100001",
  8045=>"111111111",
  8046=>"000000000",
  8047=>"011011111",
  8048=>"000000000",
  8049=>"100100110",
  8050=>"000000000",
  8051=>"101100100",
  8052=>"110111111",
  8053=>"011000000",
  8054=>"100100000",
  8055=>"100000010",
  8056=>"101000111",
  8057=>"000001001",
  8058=>"011000000",
  8059=>"111110111",
  8060=>"100000000",
  8061=>"000000000",
  8062=>"110011011",
  8063=>"011111111",
  8064=>"100100100",
  8065=>"001101011",
  8066=>"111111111",
  8067=>"000000110",
  8068=>"111001000",
  8069=>"010110000",
  8070=>"100110110",
  8071=>"111100000",
  8072=>"111111111",
  8073=>"011111011",
  8074=>"011011000",
  8075=>"000000111",
  8076=>"111101111",
  8077=>"100100110",
  8078=>"011111111",
  8079=>"010111111",
  8080=>"011000000",
  8081=>"001001000",
  8082=>"011001000",
  8083=>"111101001",
  8084=>"000111111",
  8085=>"000010010",
  8086=>"000000000",
  8087=>"000001000",
  8088=>"011001001",
  8089=>"100110110",
  8090=>"100100101",
  8091=>"111001111",
  8092=>"000000001",
  8093=>"100110100",
  8094=>"000000011",
  8095=>"001000111",
  8096=>"111111000",
  8097=>"001001011",
  8098=>"011011011",
  8099=>"010111111",
  8100=>"000000101",
  8101=>"011111011",
  8102=>"111111001",
  8103=>"000010000",
  8104=>"001011011",
  8105=>"000000110",
  8106=>"000100111",
  8107=>"011001001",
  8108=>"010111000",
  8109=>"101001111",
  8110=>"100000000",
  8111=>"001000000",
  8112=>"110110000",
  8113=>"000001111",
  8114=>"000000110",
  8115=>"111111111",
  8116=>"000000010",
  8117=>"001000000",
  8118=>"001001101",
  8119=>"100000000",
  8120=>"101100110",
  8121=>"000011111",
  8122=>"000000000",
  8123=>"011111111",
  8124=>"111001001",
  8125=>"001001000",
  8126=>"001001001",
  8127=>"000000000",
  8128=>"000000110",
  8129=>"101111111",
  8130=>"000000001",
  8131=>"000111110",
  8132=>"001001001",
  8133=>"001000111",
  8134=>"000111111",
  8135=>"111111011",
  8136=>"100000001",
  8137=>"011011000",
  8138=>"000000000",
  8139=>"000010000",
  8140=>"000000000",
  8141=>"011111011",
  8142=>"101001001",
  8143=>"010110111",
  8144=>"000111110",
  8145=>"110111111",
  8146=>"000001011",
  8147=>"000000110",
  8148=>"111111100",
  8149=>"101000000",
  8150=>"011001001",
  8151=>"001001001",
  8152=>"001001111",
  8153=>"011111111",
  8154=>"100111000",
  8155=>"111001000",
  8156=>"110111111",
  8157=>"111111111",
  8158=>"111111011",
  8159=>"000001011",
  8160=>"111111111",
  8161=>"110111110",
  8162=>"111111010",
  8163=>"011111111",
  8164=>"111110110",
  8165=>"111111111",
  8166=>"111111110",
  8167=>"000000010",
  8168=>"101101000",
  8169=>"010000000",
  8170=>"110001111",
  8171=>"101110000",
  8172=>"100101111",
  8173=>"011000000",
  8174=>"000000000",
  8175=>"111101001",
  8176=>"111000000",
  8177=>"000110000",
  8178=>"000111111",
  8179=>"111010000",
  8180=>"000000000",
  8181=>"000000000",
  8182=>"010110110",
  8183=>"101100110",
  8184=>"000000000",
  8185=>"011001000",
  8186=>"000000000",
  8187=>"111000000",
  8188=>"000000100",
  8189=>"100000000",
  8190=>"111100100",
  8191=>"000000001",
  8192=>"010110010",
  8193=>"000000000",
  8194=>"000000111",
  8195=>"100111111",
  8196=>"001000000",
  8197=>"110100100",
  8198=>"111100110",
  8199=>"000000000",
  8200=>"011000000",
  8201=>"100101111",
  8202=>"111111111",
  8203=>"000111010",
  8204=>"100110110",
  8205=>"011000101",
  8206=>"000001111",
  8207=>"111111110",
  8208=>"100111111",
  8209=>"100100001",
  8210=>"011111000",
  8211=>"000001111",
  8212=>"111000000",
  8213=>"111111011",
  8214=>"111110111",
  8215=>"111001001",
  8216=>"000000000",
  8217=>"000011111",
  8218=>"010000000",
  8219=>"000000011",
  8220=>"000000000",
  8221=>"001111000",
  8222=>"000000110",
  8223=>"100000000",
  8224=>"110111011",
  8225=>"111111111",
  8226=>"010111000",
  8227=>"010111110",
  8228=>"001000000",
  8229=>"011111111",
  8230=>"111000000",
  8231=>"011011000",
  8232=>"000100111",
  8233=>"100110110",
  8234=>"011111111",
  8235=>"111001000",
  8236=>"000001111",
  8237=>"000010000",
  8238=>"000011111",
  8239=>"010111101",
  8240=>"000000001",
  8241=>"111011000",
  8242=>"000110000",
  8243=>"000001111",
  8244=>"000011011",
  8245=>"011011110",
  8246=>"111001011",
  8247=>"000101111",
  8248=>"111111110",
  8249=>"010000111",
  8250=>"111111111",
  8251=>"111011011",
  8252=>"111111111",
  8253=>"111111000",
  8254=>"010110000",
  8255=>"101111011",
  8256=>"111111001",
  8257=>"000111111",
  8258=>"000111111",
  8259=>"111001001",
  8260=>"011000000",
  8261=>"001000000",
  8262=>"011000000",
  8263=>"111111111",
  8264=>"011011011",
  8265=>"000000111",
  8266=>"111001100",
  8267=>"100100110",
  8268=>"110011111",
  8269=>"110010000",
  8270=>"000000100",
  8271=>"100111111",
  8272=>"111000000",
  8273=>"001111011",
  8274=>"001001001",
  8275=>"000110110",
  8276=>"000000000",
  8277=>"000111101",
  8278=>"111110111",
  8279=>"000000000",
  8280=>"111111011",
  8281=>"000000000",
  8282=>"111000111",
  8283=>"000001001",
  8284=>"110000101",
  8285=>"111111000",
  8286=>"110110000",
  8287=>"111011001",
  8288=>"111111110",
  8289=>"000111111",
  8290=>"000000011",
  8291=>"110111111",
  8292=>"000000000",
  8293=>"110000001",
  8294=>"110100111",
  8295=>"101100101",
  8296=>"000110000",
  8297=>"111000000",
  8298=>"111100110",
  8299=>"000111111",
  8300=>"111110000",
  8301=>"111111111",
  8302=>"111001001",
  8303=>"011001101",
  8304=>"000000111",
  8305=>"110100100",
  8306=>"001101101",
  8307=>"111000000",
  8308=>"000000100",
  8309=>"110111111",
  8310=>"100111111",
  8311=>"100001000",
  8312=>"010100000",
  8313=>"111011001",
  8314=>"100000100",
  8315=>"111111001",
  8316=>"000011010",
  8317=>"000001011",
  8318=>"000000000",
  8319=>"100000000",
  8320=>"111011011",
  8321=>"111110111",
  8322=>"111111000",
  8323=>"111111000",
  8324=>"111001001",
  8325=>"110000111",
  8326=>"000000000",
  8327=>"101001001",
  8328=>"111111111",
  8329=>"000001001",
  8330=>"111111001",
  8331=>"000110100",
  8332=>"000000000",
  8333=>"000111111",
  8334=>"111111000",
  8335=>"111111000",
  8336=>"000000000",
  8337=>"001000001",
  8338=>"000111111",
  8339=>"110110011",
  8340=>"011100100",
  8341=>"001001001",
  8342=>"111111111",
  8343=>"001000001",
  8344=>"001000000",
  8345=>"011011000",
  8346=>"111111111",
  8347=>"000000001",
  8348=>"011000000",
  8349=>"111100100",
  8350=>"000110111",
  8351=>"000000000",
  8352=>"111111111",
  8353=>"101001001",
  8354=>"111111111",
  8355=>"111000010",
  8356=>"100001011",
  8357=>"101101111",
  8358=>"001001101",
  8359=>"100101001",
  8360=>"110111110",
  8361=>"101001001",
  8362=>"100000000",
  8363=>"000001111",
  8364=>"001000000",
  8365=>"001000001",
  8366=>"001000000",
  8367=>"101111111",
  8368=>"000011111",
  8369=>"001101001",
  8370=>"001101001",
  8371=>"100101000",
  8372=>"111111000",
  8373=>"000000001",
  8374=>"000000001",
  8375=>"000000010",
  8376=>"001000001",
  8377=>"000001111",
  8378=>"110010000",
  8379=>"110110111",
  8380=>"001111111",
  8381=>"000101111",
  8382=>"110111100",
  8383=>"000000001",
  8384=>"111111000",
  8385=>"111101111",
  8386=>"111111111",
  8387=>"001000000",
  8388=>"000000000",
  8389=>"000000001",
  8390=>"000000110",
  8391=>"010110110",
  8392=>"111111111",
  8393=>"111000100",
  8394=>"100110111",
  8395=>"111111111",
  8396=>"000001001",
  8397=>"000111111",
  8398=>"111111000",
  8399=>"110000000",
  8400=>"001001000",
  8401=>"110110111",
  8402=>"111111001",
  8403=>"000000000",
  8404=>"101000100",
  8405=>"110010111",
  8406=>"101100101",
  8407=>"000000000",
  8408=>"001111111",
  8409=>"011111000",
  8410=>"000110111",
  8411=>"001000100",
  8412=>"110111111",
  8413=>"001000000",
  8414=>"111111111",
  8415=>"000111101",
  8416=>"001011011",
  8417=>"000000110",
  8418=>"111111111",
  8419=>"101100110",
  8420=>"010000000",
  8421=>"001000000",
  8422=>"110111111",
  8423=>"000000111",
  8424=>"111111111",
  8425=>"001000000",
  8426=>"111111011",
  8427=>"110000000",
  8428=>"101101000",
  8429=>"000100110",
  8430=>"101000000",
  8431=>"000000111",
  8432=>"011111000",
  8433=>"110000000",
  8434=>"111000000",
  8435=>"110000000",
  8436=>"000000111",
  8437=>"111100000",
  8438=>"000000111",
  8439=>"111111110",
  8440=>"110000000",
  8441=>"101111111",
  8442=>"111111111",
  8443=>"000001000",
  8444=>"100110000",
  8445=>"100110011",
  8446=>"111000000",
  8447=>"111100000",
  8448=>"101000111",
  8449=>"011011111",
  8450=>"111110110",
  8451=>"101000000",
  8452=>"111111110",
  8453=>"000111111",
  8454=>"000000000",
  8455=>"111101001",
  8456=>"101000000",
  8457=>"011111111",
  8458=>"000000000",
  8459=>"111100000",
  8460=>"000000000",
  8461=>"000000000",
  8462=>"000000111",
  8463=>"111111011",
  8464=>"110110111",
  8465=>"111011001",
  8466=>"000000000",
  8467=>"000110111",
  8468=>"000000000",
  8469=>"111111110",
  8470=>"000101001",
  8471=>"111111111",
  8472=>"111111111",
  8473=>"111111000",
  8474=>"000000000",
  8475=>"000000000",
  8476=>"111111111",
  8477=>"100110110",
  8478=>"000000111",
  8479=>"101001111",
  8480=>"000000000",
  8481=>"111000000",
  8482=>"000111011",
  8483=>"111111000",
  8484=>"001011111",
  8485=>"111000000",
  8486=>"000000000",
  8487=>"111111000",
  8488=>"000000000",
  8489=>"000000101",
  8490=>"010000000",
  8491=>"011000000",
  8492=>"011011000",
  8493=>"010011001",
  8494=>"101000000",
  8495=>"000000000",
  8496=>"000000000",
  8497=>"000000000",
  8498=>"011111111",
  8499=>"000000110",
  8500=>"111111110",
  8501=>"001011001",
  8502=>"111111010",
  8503=>"010111111",
  8504=>"000000000",
  8505=>"000000010",
  8506=>"111100000",
  8507=>"111001000",
  8508=>"001000000",
  8509=>"011111111",
  8510=>"110111111",
  8511=>"111111010",
  8512=>"000000110",
  8513=>"110111001",
  8514=>"000000001",
  8515=>"000000000",
  8516=>"011010000",
  8517=>"100000000",
  8518=>"000111111",
  8519=>"000000000",
  8520=>"001000000",
  8521=>"111000000",
  8522=>"001001000",
  8523=>"111111001",
  8524=>"111111010",
  8525=>"000111111",
  8526=>"111011011",
  8527=>"000000101",
  8528=>"011001100",
  8529=>"111011000",
  8530=>"000111100",
  8531=>"111111010",
  8532=>"110000000",
  8533=>"010011111",
  8534=>"111111111",
  8535=>"101000001",
  8536=>"000011101",
  8537=>"001000000",
  8538=>"110110010",
  8539=>"000000110",
  8540=>"111111111",
  8541=>"110111111",
  8542=>"111111011",
  8543=>"000000110",
  8544=>"111111111",
  8545=>"000000000",
  8546=>"000011011",
  8547=>"001001001",
  8548=>"000011011",
  8549=>"001000000",
  8550=>"111111111",
  8551=>"001001011",
  8552=>"000001000",
  8553=>"100000000",
  8554=>"000000000",
  8555=>"001000000",
  8556=>"111001000",
  8557=>"110000111",
  8558=>"000000001",
  8559=>"001001111",
  8560=>"111111111",
  8561=>"111100100",
  8562=>"111111111",
  8563=>"111111001",
  8564=>"100000100",
  8565=>"111111111",
  8566=>"101000000",
  8567=>"101111011",
  8568=>"111100000",
  8569=>"100110100",
  8570=>"011000000",
  8571=>"111111110",
  8572=>"100000111",
  8573=>"000000001",
  8574=>"000111111",
  8575=>"111111111",
  8576=>"000000000",
  8577=>"000000000",
  8578=>"110000000",
  8579=>"100101111",
  8580=>"100000000",
  8581=>"000000000",
  8582=>"001000100",
  8583=>"000000001",
  8584=>"000001011",
  8585=>"011001000",
  8586=>"000000000",
  8587=>"000001000",
  8588=>"000000111",
  8589=>"000101111",
  8590=>"111001000",
  8591=>"000000110",
  8592=>"000000110",
  8593=>"001001001",
  8594=>"000000000",
  8595=>"111100000",
  8596=>"000000111",
  8597=>"000110000",
  8598=>"000000000",
  8599=>"010010000",
  8600=>"000110110",
  8601=>"010110111",
  8602=>"011010110",
  8603=>"000110110",
  8604=>"000110111",
  8605=>"110010000",
  8606=>"000110110",
  8607=>"111111001",
  8608=>"111111100",
  8609=>"111110111",
  8610=>"111000010",
  8611=>"100110111",
  8612=>"001001111",
  8613=>"110100000",
  8614=>"110101000",
  8615=>"001000000",
  8616=>"000000000",
  8617=>"000000010",
  8618=>"111000000",
  8619=>"000110110",
  8620=>"111111100",
  8621=>"000000000",
  8622=>"111000100",
  8623=>"111111000",
  8624=>"110110111",
  8625=>"100000101",
  8626=>"101100100",
  8627=>"111111101",
  8628=>"000100101",
  8629=>"111111111",
  8630=>"111111010",
  8631=>"001111011",
  8632=>"101110000",
  8633=>"000000111",
  8634=>"110100010",
  8635=>"001000101",
  8636=>"000110111",
  8637=>"001011111",
  8638=>"000001001",
  8639=>"000011011",
  8640=>"000111111",
  8641=>"100100111",
  8642=>"111000111",
  8643=>"000000000",
  8644=>"000000111",
  8645=>"001000010",
  8646=>"000000010",
  8647=>"000111011",
  8648=>"111000111",
  8649=>"011000100",
  8650=>"110110100",
  8651=>"111111000",
  8652=>"000111000",
  8653=>"000000111",
  8654=>"000110110",
  8655=>"110110100",
  8656=>"000000000",
  8657=>"000000000",
  8658=>"111111000",
  8659=>"101000111",
  8660=>"111011001",
  8661=>"100100100",
  8662=>"000000011",
  8663=>"111111000",
  8664=>"000000110",
  8665=>"110110110",
  8666=>"000000001",
  8667=>"000000000",
  8668=>"000000000",
  8669=>"010000001",
  8670=>"111111000",
  8671=>"000000001",
  8672=>"001000000",
  8673=>"111001000",
  8674=>"000000001",
  8675=>"101101111",
  8676=>"101100100",
  8677=>"000000110",
  8678=>"001000000",
  8679=>"111000000",
  8680=>"111111111",
  8681=>"100101111",
  8682=>"000000000",
  8683=>"111111111",
  8684=>"010010111",
  8685=>"111000000",
  8686=>"101101100",
  8687=>"001001111",
  8688=>"000000100",
  8689=>"000111111",
  8690=>"000000111",
  8691=>"100000000",
  8692=>"001111111",
  8693=>"001001111",
  8694=>"010001000",
  8695=>"011111111",
  8696=>"011001000",
  8697=>"001001000",
  8698=>"111111001",
  8699=>"000000011",
  8700=>"100000101",
  8701=>"111000000",
  8702=>"011110100",
  8703=>"011010011",
  8704=>"000000000",
  8705=>"100110111",
  8706=>"111111111",
  8707=>"111111111",
  8708=>"100000111",
  8709=>"111110000",
  8710=>"000000000",
  8711=>"110000000",
  8712=>"000000110",
  8713=>"110110111",
  8714=>"111111111",
  8715=>"111000000",
  8716=>"000100100",
  8717=>"011111110",
  8718=>"110110110",
  8719=>"000000000",
  8720=>"000000000",
  8721=>"000000100",
  8722=>"011111011",
  8723=>"100000000",
  8724=>"000000000",
  8725=>"110111111",
  8726=>"000110111",
  8727=>"000111100",
  8728=>"111100000",
  8729=>"000011011",
  8730=>"011011000",
  8731=>"000000000",
  8732=>"000000000",
  8733=>"111111011",
  8734=>"111110000",
  8735=>"011000000",
  8736=>"000000001",
  8737=>"000000001",
  8738=>"000000001",
  8739=>"111111011",
  8740=>"001001010",
  8741=>"111111111",
  8742=>"000000111",
  8743=>"111111011",
  8744=>"000000000",
  8745=>"111000101",
  8746=>"111000111",
  8747=>"111111011",
  8748=>"000011111",
  8749=>"000111111",
  8750=>"110011001",
  8751=>"111011000",
  8752=>"111111111",
  8753=>"000000000",
  8754=>"000000000",
  8755=>"001111000",
  8756=>"000000001",
  8757=>"010000010",
  8758=>"001000000",
  8759=>"111111111",
  8760=>"111101000",
  8761=>"010000111",
  8762=>"111111111",
  8763=>"111111111",
  8764=>"111100000",
  8765=>"111111111",
  8766=>"000000000",
  8767=>"000001001",
  8768=>"011111111",
  8769=>"000000110",
  8770=>"111001001",
  8771=>"000001000",
  8772=>"000000000",
  8773=>"001000001",
  8774=>"000000000",
  8775=>"110111111",
  8776=>"111111111",
  8777=>"111111110",
  8778=>"111110100",
  8779=>"000000110",
  8780=>"111011111",
  8781=>"111111110",
  8782=>"000000000",
  8783=>"000000000",
  8784=>"000000001",
  8785=>"111111111",
  8786=>"000000000",
  8787=>"110011111",
  8788=>"000000000",
  8789=>"011111000",
  8790=>"011111111",
  8791=>"111111000",
  8792=>"001111011",
  8793=>"000000000",
  8794=>"010110111",
  8795=>"000000100",
  8796=>"111111111",
  8797=>"111111111",
  8798=>"000000000",
  8799=>"000000011",
  8800=>"000000000",
  8801=>"111111111",
  8802=>"110111111",
  8803=>"100000100",
  8804=>"001111010",
  8805=>"000100111",
  8806=>"000000000",
  8807=>"010000000",
  8808=>"111101111",
  8809=>"000000000",
  8810=>"000100111",
  8811=>"110111111",
  8812=>"111101101",
  8813=>"111111111",
  8814=>"010010010",
  8815=>"111110100",
  8816=>"111111111",
  8817=>"111101111",
  8818=>"000000011",
  8819=>"111111111",
  8820=>"111011111",
  8821=>"000000110",
  8822=>"100000000",
  8823=>"111111000",
  8824=>"000011110",
  8825=>"001000110",
  8826=>"000001000",
  8827=>"110000000",
  8828=>"110100100",
  8829=>"011000000",
  8830=>"000000000",
  8831=>"000000000",
  8832=>"000000100",
  8833=>"000000000",
  8834=>"000110111",
  8835=>"111101110",
  8836=>"000111111",
  8837=>"000100111",
  8838=>"111111111",
  8839=>"000000000",
  8840=>"000000000",
  8841=>"000000000",
  8842=>"111111111",
  8843=>"111111111",
  8844=>"101101111",
  8845=>"001001001",
  8846=>"000000000",
  8847=>"011111100",
  8848=>"000000000",
  8849=>"101000000",
  8850=>"000000000",
  8851=>"101111111",
  8852=>"000110100",
  8853=>"111111111",
  8854=>"000000111",
  8855=>"001000000",
  8856=>"000110000",
  8857=>"110111111",
  8858=>"001111111",
  8859=>"111111111",
  8860=>"000000111",
  8861=>"111100000",
  8862=>"010010000",
  8863=>"000000000",
  8864=>"000000000",
  8865=>"000101001",
  8866=>"001001000",
  8867=>"000000000",
  8868=>"000000110",
  8869=>"110111011",
  8870=>"111001000",
  8871=>"111111111",
  8872=>"011001110",
  8873=>"111111111",
  8874=>"110101101",
  8875=>"111111111",
  8876=>"111111111",
  8877=>"001001001",
  8878=>"001111111",
  8879=>"101001001",
  8880=>"000000000",
  8881=>"000000000",
  8882=>"111111111",
  8883=>"001000000",
  8884=>"000000000",
  8885=>"010000000",
  8886=>"000001001",
  8887=>"111111101",
  8888=>"010000000",
  8889=>"010000010",
  8890=>"000000000",
  8891=>"010011111",
  8892=>"001001000",
  8893=>"000000111",
  8894=>"111111000",
  8895=>"101000101",
  8896=>"100000001",
  8897=>"000000000",
  8898=>"000000000",
  8899=>"000000000",
  8900=>"000001111",
  8901=>"011011001",
  8902=>"010111111",
  8903=>"110100000",
  8904=>"111111111",
  8905=>"011001001",
  8906=>"111101111",
  8907=>"000000010",
  8908=>"111111011",
  8909=>"000000100",
  8910=>"000000001",
  8911=>"010111000",
  8912=>"100000000",
  8913=>"111110000",
  8914=>"001000000",
  8915=>"010011101",
  8916=>"101101000",
  8917=>"000000001",
  8918=>"001000000",
  8919=>"101100000",
  8920=>"000000000",
  8921=>"111001101",
  8922=>"000000000",
  8923=>"111111111",
  8924=>"011001001",
  8925=>"100000111",
  8926=>"000000111",
  8927=>"010011011",
  8928=>"111011001",
  8929=>"110111110",
  8930=>"000010111",
  8931=>"111111111",
  8932=>"111111001",
  8933=>"111100000",
  8934=>"000000111",
  8935=>"111111000",
  8936=>"000001000",
  8937=>"001101100",
  8938=>"000000000",
  8939=>"000000000",
  8940=>"001000001",
  8941=>"001000000",
  8942=>"011111100",
  8943=>"111111111",
  8944=>"111111111",
  8945=>"000000001",
  8946=>"110100111",
  8947=>"001001001",
  8948=>"111111100",
  8949=>"000000000",
  8950=>"110111111",
  8951=>"001000000",
  8952=>"111111111",
  8953=>"000000000",
  8954=>"000000001",
  8955=>"111111111",
  8956=>"111110100",
  8957=>"000000000",
  8958=>"010011001",
  8959=>"100111111",
  8960=>"010011000",
  8961=>"011000000",
  8962=>"000000111",
  8963=>"010111111",
  8964=>"000000001",
  8965=>"111111111",
  8966=>"111111111",
  8967=>"000000000",
  8968=>"000000100",
  8969=>"000000000",
  8970=>"000000001",
  8971=>"111111111",
  8972=>"000000111",
  8973=>"111111111",
  8974=>"000000000",
  8975=>"000000000",
  8976=>"000000000",
  8977=>"000111111",
  8978=>"111100001",
  8979=>"000100111",
  8980=>"000000000",
  8981=>"000000000",
  8982=>"001011011",
  8983=>"111101001",
  8984=>"100100001",
  8985=>"111111000",
  8986=>"001000000",
  8987=>"000111111",
  8988=>"000000000",
  8989=>"111111111",
  8990=>"000000000",
  8991=>"001100000",
  8992=>"000000010",
  8993=>"001111111",
  8994=>"101111111",
  8995=>"000000111",
  8996=>"100100000",
  8997=>"000000000",
  8998=>"000101111",
  8999=>"101101111",
  9000=>"000011111",
  9001=>"001001000",
  9002=>"100000101",
  9003=>"111111111",
  9004=>"001011011",
  9005=>"000001111",
  9006=>"000000000",
  9007=>"011010000",
  9008=>"000000111",
  9009=>"000000000",
  9010=>"111111011",
  9011=>"111111111",
  9012=>"101000101",
  9013=>"001001011",
  9014=>"011110000",
  9015=>"000000000",
  9016=>"000000000",
  9017=>"000000111",
  9018=>"000000111",
  9019=>"000110111",
  9020=>"000000000",
  9021=>"101101000",
  9022=>"011000000",
  9023=>"000000001",
  9024=>"000000000",
  9025=>"101100000",
  9026=>"001011101",
  9027=>"101101100",
  9028=>"111111111",
  9029=>"001011111",
  9030=>"000011000",
  9031=>"000100110",
  9032=>"000000000",
  9033=>"100000000",
  9034=>"111111111",
  9035=>"111000000",
  9036=>"010111110",
  9037=>"100100110",
  9038=>"111111111",
  9039=>"011001000",
  9040=>"110010111",
  9041=>"111111111",
  9042=>"111111111",
  9043=>"000000101",
  9044=>"011000000",
  9045=>"011011001",
  9046=>"111101101",
  9047=>"111111111",
  9048=>"111111111",
  9049=>"111111010",
  9050=>"000010110",
  9051=>"100100000",
  9052=>"100101101",
  9053=>"000000000",
  9054=>"101111111",
  9055=>"111011001",
  9056=>"001101100",
  9057=>"111111111",
  9058=>"101001001",
  9059=>"000000000",
  9060=>"101111010",
  9061=>"000000000",
  9062=>"110110001",
  9063=>"111111111",
  9064=>"110110011",
  9065=>"000001011",
  9066=>"000000000",
  9067=>"111111111",
  9068=>"000000000",
  9069=>"000111111",
  9070=>"111000111",
  9071=>"000000000",
  9072=>"111000100",
  9073=>"000000000",
  9074=>"000000000",
  9075=>"111111000",
  9076=>"101111111",
  9077=>"101000000",
  9078=>"000000111",
  9079=>"001011000",
  9080=>"000000000",
  9081=>"111111111",
  9082=>"111111111",
  9083=>"010010000",
  9084=>"000000000",
  9085=>"110110000",
  9086=>"010000000",
  9087=>"000000000",
  9088=>"000000001",
  9089=>"111111111",
  9090=>"000000011",
  9091=>"111100100",
  9092=>"111111000",
  9093=>"111111111",
  9094=>"000000000",
  9095=>"111110101",
  9096=>"111111111",
  9097=>"000000110",
  9098=>"000000000",
  9099=>"100100100",
  9100=>"101000001",
  9101=>"000000000",
  9102=>"000100110",
  9103=>"111111111",
  9104=>"000000110",
  9105=>"111000000",
  9106=>"000000000",
  9107=>"000000000",
  9108=>"000000000",
  9109=>"000000110",
  9110=>"000000111",
  9111=>"100111111",
  9112=>"100111011",
  9113=>"000010110",
  9114=>"111110100",
  9115=>"111111111",
  9116=>"011011000",
  9117=>"000000000",
  9118=>"000000010",
  9119=>"000000000",
  9120=>"000000000",
  9121=>"110111111",
  9122=>"000000111",
  9123=>"000011000",
  9124=>"111111111",
  9125=>"000011111",
  9126=>"111111111",
  9127=>"111011000",
  9128=>"110111111",
  9129=>"111011011",
  9130=>"111111111",
  9131=>"000000000",
  9132=>"111101000",
  9133=>"111101111",
  9134=>"000111111",
  9135=>"111111011",
  9136=>"110111111",
  9137=>"111000000",
  9138=>"011100000",
  9139=>"100001111",
  9140=>"000000000",
  9141=>"111110000",
  9142=>"100001001",
  9143=>"111101111",
  9144=>"001000000",
  9145=>"111111111",
  9146=>"111111000",
  9147=>"001000001",
  9148=>"000000000",
  9149=>"111011000",
  9150=>"000000000",
  9151=>"011111111",
  9152=>"111111001",
  9153=>"111111111",
  9154=>"000011111",
  9155=>"111111111",
  9156=>"100111111",
  9157=>"111011010",
  9158=>"000111111",
  9159=>"000000100",
  9160=>"001000000",
  9161=>"000000100",
  9162=>"000101001",
  9163=>"000000001",
  9164=>"100000000",
  9165=>"100111111",
  9166=>"010111000",
  9167=>"010011111",
  9168=>"111100000",
  9169=>"100000000",
  9170=>"000000000",
  9171=>"000000000",
  9172=>"000000000",
  9173=>"110111000",
  9174=>"111001011",
  9175=>"000000010",
  9176=>"000000000",
  9177=>"000000011",
  9178=>"110000000",
  9179=>"000000000",
  9180=>"000000011",
  9181=>"001011011",
  9182=>"000000000",
  9183=>"001011011",
  9184=>"000000111",
  9185=>"000000000",
  9186=>"000000111",
  9187=>"001000000",
  9188=>"100110111",
  9189=>"000000000",
  9190=>"000001111",
  9191=>"000001000",
  9192=>"101111111",
  9193=>"011001001",
  9194=>"111111111",
  9195=>"000000000",
  9196=>"110110000",
  9197=>"000100100",
  9198=>"000000000",
  9199=>"000000011",
  9200=>"000000000",
  9201=>"000000000",
  9202=>"001001000",
  9203=>"000000000",
  9204=>"000000000",
  9205=>"111111111",
  9206=>"000110011",
  9207=>"110111011",
  9208=>"011011000",
  9209=>"010111111",
  9210=>"000000000",
  9211=>"111111110",
  9212=>"000000000",
  9213=>"111111111",
  9214=>"111110000",
  9215=>"000001001",
  9216=>"111111110",
  9217=>"001001000",
  9218=>"000000000",
  9219=>"111001011",
  9220=>"000001111",
  9221=>"010111000",
  9222=>"111111111",
  9223=>"000000000",
  9224=>"001100000",
  9225=>"111111111",
  9226=>"001101000",
  9227=>"111111000",
  9228=>"000000000",
  9229=>"000100001",
  9230=>"000000000",
  9231=>"010000110",
  9232=>"000111000",
  9233=>"111001111",
  9234=>"111000000",
  9235=>"000110110",
  9236=>"000111000",
  9237=>"110111000",
  9238=>"110111111",
  9239=>"111000000",
  9240=>"110110110",
  9241=>"111000101",
  9242=>"010011111",
  9243=>"100111011",
  9244=>"010000000",
  9245=>"011000001",
  9246=>"011001011",
  9247=>"000000000",
  9248=>"111111000",
  9249=>"110111000",
  9250=>"001001001",
  9251=>"000000000",
  9252=>"111111111",
  9253=>"000001000",
  9254=>"001100110",
  9255=>"000001000",
  9256=>"111111100",
  9257=>"101111111",
  9258=>"000111111",
  9259=>"000011010",
  9260=>"000000001",
  9261=>"111111010",
  9262=>"110111111",
  9263=>"011000000",
  9264=>"011001000",
  9265=>"111000100",
  9266=>"000100110",
  9267=>"001111011",
  9268=>"111001111",
  9269=>"111001111",
  9270=>"000011000",
  9271=>"110011101",
  9272=>"000111111",
  9273=>"001001100",
  9274=>"111111111",
  9275=>"111111011",
  9276=>"000000000",
  9277=>"000011001",
  9278=>"110100010",
  9279=>"001110001",
  9280=>"100001111",
  9281=>"001111111",
  9282=>"000000000",
  9283=>"001111111",
  9284=>"001111010",
  9285=>"011111110",
  9286=>"000000000",
  9287=>"111111100",
  9288=>"001111111",
  9289=>"101000000",
  9290=>"000000000",
  9291=>"000111000",
  9292=>"111111011",
  9293=>"111000101",
  9294=>"000001000",
  9295=>"101111101",
  9296=>"000111101",
  9297=>"111110011",
  9298=>"111110000",
  9299=>"011011000",
  9300=>"000000001",
  9301=>"011000110",
  9302=>"000011111",
  9303=>"111111111",
  9304=>"000111000",
  9305=>"000111000",
  9306=>"000111000",
  9307=>"000101001",
  9308=>"110111000",
  9309=>"001101100",
  9310=>"000000000",
  9311=>"101111011",
  9312=>"000110000",
  9313=>"000111000",
  9314=>"110110111",
  9315=>"111111000",
  9316=>"001011011",
  9317=>"110001000",
  9318=>"001111111",
  9319=>"111101111",
  9320=>"010000010",
  9321=>"000110010",
  9322=>"000000111",
  9323=>"111111111",
  9324=>"010000000",
  9325=>"110111111",
  9326=>"111110100",
  9327=>"111111011",
  9328=>"001011000",
  9329=>"001000000",
  9330=>"111001111",
  9331=>"001111110",
  9332=>"001111111",
  9333=>"111111101",
  9334=>"001111111",
  9335=>"010111111",
  9336=>"000111110",
  9337=>"000100111",
  9338=>"110110100",
  9339=>"000011000",
  9340=>"100100110",
  9341=>"110011000",
  9342=>"110110100",
  9343=>"111000000",
  9344=>"000000001",
  9345=>"010100000",
  9346=>"111001000",
  9347=>"000001000",
  9348=>"101101111",
  9349=>"111111000",
  9350=>"000111000",
  9351=>"111011001",
  9352=>"011111010",
  9353=>"110110111",
  9354=>"000001000",
  9355=>"000000000",
  9356=>"000111011",
  9357=>"011111100",
  9358=>"101111111",
  9359=>"111111101",
  9360=>"110110110",
  9361=>"111000000",
  9362=>"001001111",
  9363=>"000110010",
  9364=>"111111111",
  9365=>"110011011",
  9366=>"000000000",
  9367=>"001101000",
  9368=>"001101000",
  9369=>"000111111",
  9370=>"111111000",
  9371=>"111111000",
  9372=>"000100001",
  9373=>"000111000",
  9374=>"000001000",
  9375=>"000110111",
  9376=>"100000000",
  9377=>"000111000",
  9378=>"000111111",
  9379=>"000111111",
  9380=>"111000110",
  9381=>"000111111",
  9382=>"000000000",
  9383=>"011010111",
  9384=>"000011010",
  9385=>"111111000",
  9386=>"111111101",
  9387=>"000011001",
  9388=>"000100111",
  9389=>"101111011",
  9390=>"111101001",
  9391=>"000111111",
  9392=>"000000000",
  9393=>"001001101",
  9394=>"111010111",
  9395=>"000000000",
  9396=>"110110010",
  9397=>"000000000",
  9398=>"111111011",
  9399=>"110000000",
  9400=>"001111111",
  9401=>"000001111",
  9402=>"110000111",
  9403=>"110001101",
  9404=>"000111111",
  9405=>"000000100",
  9406=>"000000000",
  9407=>"110010111",
  9408=>"111111111",
  9409=>"000110100",
  9410=>"011011000",
  9411=>"000000000",
  9412=>"001001111",
  9413=>"100101111",
  9414=>"111101101",
  9415=>"010001011",
  9416=>"000000000",
  9417=>"011111110",
  9418=>"001111010",
  9419=>"111111111",
  9420=>"001111010",
  9421=>"111001111",
  9422=>"111111111",
  9423=>"010000100",
  9424=>"111111000",
  9425=>"111111000",
  9426=>"110111000",
  9427=>"111111111",
  9428=>"111111111",
  9429=>"001111100",
  9430=>"011000000",
  9431=>"000111011",
  9432=>"000000000",
  9433=>"000011001",
  9434=>"111111111",
  9435=>"000111000",
  9436=>"000111110",
  9437=>"000000000",
  9438=>"111000000",
  9439=>"011111000",
  9440=>"001010000",
  9441=>"001000100",
  9442=>"000000000",
  9443=>"000100111",
  9444=>"111100110",
  9445=>"011001001",
  9446=>"000000000",
  9447=>"111111000",
  9448=>"000000111",
  9449=>"111110010",
  9450=>"000000001",
  9451=>"000001111",
  9452=>"111111111",
  9453=>"111000001",
  9454=>"001111000",
  9455=>"000111000",
  9456=>"111000110",
  9457=>"110000000",
  9458=>"110100000",
  9459=>"000001000",
  9460=>"000001001",
  9461=>"111111111",
  9462=>"010110111",
  9463=>"000000011",
  9464=>"011001000",
  9465=>"111111111",
  9466=>"000111111",
  9467=>"111111001",
  9468=>"110000111",
  9469=>"110011110",
  9470=>"000111111",
  9471=>"100110111",
  9472=>"000001111",
  9473=>"010010010",
  9474=>"111111111",
  9475=>"000000000",
  9476=>"111110000",
  9477=>"100111111",
  9478=>"011111000",
  9479=>"000111011",
  9480=>"111111000",
  9481=>"110111111",
  9482=>"000000000",
  9483=>"000101111",
  9484=>"111111111",
  9485=>"000111111",
  9486=>"000001000",
  9487=>"111111000",
  9488=>"110111110",
  9489=>"011011000",
  9490=>"000000001",
  9491=>"110111111",
  9492=>"111001000",
  9493=>"111111000",
  9494=>"110111101",
  9495=>"111111111",
  9496=>"111100111",
  9497=>"111111111",
  9498=>"000000000",
  9499=>"111111001",
  9500=>"110111111",
  9501=>"001101000",
  9502=>"111111111",
  9503=>"111001000",
  9504=>"111111100",
  9505=>"001101000",
  9506=>"111101100",
  9507=>"000111111",
  9508=>"001111001",
  9509=>"110110100",
  9510=>"110100100",
  9511=>"100000000",
  9512=>"111001111",
  9513=>"111111111",
  9514=>"000111001",
  9515=>"000000000",
  9516=>"111111111",
  9517=>"111000001",
  9518=>"000000000",
  9519=>"111001000",
  9520=>"011111110",
  9521=>"110111111",
  9522=>"000000000",
  9523=>"111111111",
  9524=>"000000000",
  9525=>"101111100",
  9526=>"000000000",
  9527=>"000111000",
  9528=>"111000011",
  9529=>"000110111",
  9530=>"111111111",
  9531=>"111001000",
  9532=>"000000000",
  9533=>"000000000",
  9534=>"000000111",
  9535=>"000111000",
  9536=>"000111001",
  9537=>"000000000",
  9538=>"000011111",
  9539=>"000100101",
  9540=>"111011000",
  9541=>"000000000",
  9542=>"011001111",
  9543=>"111111111",
  9544=>"000101001",
  9545=>"000011000",
  9546=>"000000000",
  9547=>"110110111",
  9548=>"111101000",
  9549=>"111111011",
  9550=>"000111111",
  9551=>"000000000",
  9552=>"111001111",
  9553=>"100011110",
  9554=>"000000100",
  9555=>"111000110",
  9556=>"111000000",
  9557=>"111011011",
  9558=>"111111111",
  9559=>"111111110",
  9560=>"000000111",
  9561=>"000111000",
  9562=>"001100100",
  9563=>"111101000",
  9564=>"000111010",
  9565=>"001111111",
  9566=>"111111000",
  9567=>"111100100",
  9568=>"110100000",
  9569=>"000000111",
  9570=>"110100100",
  9571=>"000000011",
  9572=>"000001101",
  9573=>"000011001",
  9574=>"111001111",
  9575=>"000000111",
  9576=>"111111111",
  9577=>"010111000",
  9578=>"111010000",
  9579=>"010110000",
  9580=>"000110110",
  9581=>"110000111",
  9582=>"110010000",
  9583=>"000011010",
  9584=>"111100000",
  9585=>"000000111",
  9586=>"111100000",
  9587=>"111111111",
  9588=>"100111111",
  9589=>"111111000",
  9590=>"000011000",
  9591=>"111001001",
  9592=>"000000100",
  9593=>"000000000",
  9594=>"000000000",
  9595=>"000001111",
  9596=>"100000000",
  9597=>"011111111",
  9598=>"010111110",
  9599=>"001000000",
  9600=>"111111000",
  9601=>"111001111",
  9602=>"110111111",
  9603=>"000000000",
  9604=>"010111111",
  9605=>"000000100",
  9606=>"011001000",
  9607=>"000111111",
  9608=>"000110000",
  9609=>"100000111",
  9610=>"001110000",
  9611=>"000000000",
  9612=>"001000000",
  9613=>"111000111",
  9614=>"000000110",
  9615=>"111111111",
  9616=>"000011011",
  9617=>"000111000",
  9618=>"010010000",
  9619=>"000000000",
  9620=>"111111010",
  9621=>"111000111",
  9622=>"100100110",
  9623=>"100000000",
  9624=>"111111000",
  9625=>"010110110",
  9626=>"010111111",
  9627=>"111000100",
  9628=>"000001111",
  9629=>"111111010",
  9630=>"111110111",
  9631=>"111111000",
  9632=>"110100111",
  9633=>"010001000",
  9634=>"000111110",
  9635=>"000110110",
  9636=>"000110110",
  9637=>"000110111",
  9638=>"000000000",
  9639=>"000000000",
  9640=>"010010000",
  9641=>"000001001",
  9642=>"000001000",
  9643=>"111000000",
  9644=>"000010000",
  9645=>"000001000",
  9646=>"000111100",
  9647=>"010010000",
  9648=>"111100110",
  9649=>"000111111",
  9650=>"011001001",
  9651=>"000000110",
  9652=>"111000000",
  9653=>"011001011",
  9654=>"000000010",
  9655=>"000110100",
  9656=>"000000000",
  9657=>"100011111",
  9658=>"001110111",
  9659=>"000000000",
  9660=>"000000010",
  9661=>"000010000",
  9662=>"111110000",
  9663=>"111011111",
  9664=>"000110111",
  9665=>"000000000",
  9666=>"000000000",
  9667=>"000000000",
  9668=>"000110100",
  9669=>"000110111",
  9670=>"101111111",
  9671=>"001001000",
  9672=>"000001111",
  9673=>"111000111",
  9674=>"001111000",
  9675=>"000000000",
  9676=>"011111000",
  9677=>"000000000",
  9678=>"110000000",
  9679=>"100110111",
  9680=>"000000000",
  9681=>"010010011",
  9682=>"111110110",
  9683=>"001111000",
  9684=>"100111001",
  9685=>"000000110",
  9686=>"010000010",
  9687=>"111001111",
  9688=>"000100000",
  9689=>"000001001",
  9690=>"111011000",
  9691=>"100111111",
  9692=>"010001000",
  9693=>"000011011",
  9694=>"011111000",
  9695=>"110101100",
  9696=>"000111111",
  9697=>"101000101",
  9698=>"110110111",
  9699=>"000111101",
  9700=>"000000001",
  9701=>"110111000",
  9702=>"001110000",
  9703=>"000111001",
  9704=>"000101001",
  9705=>"011000000",
  9706=>"000000000",
  9707=>"111110011",
  9708=>"111111000",
  9709=>"011000010",
  9710=>"111101001",
  9711=>"011110110",
  9712=>"111111111",
  9713=>"111000000",
  9714=>"010111111",
  9715=>"000111001",
  9716=>"110111011",
  9717=>"111000000",
  9718=>"000001111",
  9719=>"110001001",
  9720=>"000000000",
  9721=>"111100110",
  9722=>"111111111",
  9723=>"000000000",
  9724=>"001010110",
  9725=>"011011111",
  9726=>"110111110",
  9727=>"111111011",
  9728=>"111111111",
  9729=>"111001001",
  9730=>"111111111",
  9731=>"011000000",
  9732=>"111100100",
  9733=>"100100111",
  9734=>"011111111",
  9735=>"101111111",
  9736=>"000000000",
  9737=>"111011111",
  9738=>"000000000",
  9739=>"000011011",
  9740=>"001000000",
  9741=>"000000001",
  9742=>"111111111",
  9743=>"111111111",
  9744=>"000000000",
  9745=>"111111100",
  9746=>"111111111",
  9747=>"001000000",
  9748=>"111111000",
  9749=>"000000000",
  9750=>"111111111",
  9751=>"011001011",
  9752=>"101100111",
  9753=>"000000000",
  9754=>"000001000",
  9755=>"110110110",
  9756=>"000000001",
  9757=>"111111000",
  9758=>"011011111",
  9759=>"010000000",
  9760=>"110111111",
  9761=>"111111111",
  9762=>"100100111",
  9763=>"000000000",
  9764=>"011011011",
  9765=>"000100111",
  9766=>"001000101",
  9767=>"000000000",
  9768=>"001000000",
  9769=>"100100100",
  9770=>"000000000",
  9771=>"000000010",
  9772=>"110111111",
  9773=>"110110000",
  9774=>"011011110",
  9775=>"000110000",
  9776=>"111110111",
  9777=>"011011111",
  9778=>"011011111",
  9779=>"111111011",
  9780=>"000000000",
  9781=>"000000000",
  9782=>"000100100",
  9783=>"000101111",
  9784=>"011011001",
  9785=>"111011111",
  9786=>"111111110",
  9787=>"000000000",
  9788=>"101101000",
  9789=>"100111111",
  9790=>"111111111",
  9791=>"000000000",
  9792=>"000001111",
  9793=>"001000111",
  9794=>"000000000",
  9795=>"000000111",
  9796=>"000000010",
  9797=>"000000000",
  9798=>"000000000",
  9799=>"111111111",
  9800=>"111110110",
  9801=>"000000100",
  9802=>"000000010",
  9803=>"111111010",
  9804=>"010011000",
  9805=>"000000111",
  9806=>"111011111",
  9807=>"011011001",
  9808=>"000101111",
  9809=>"000000000",
  9810=>"111101000",
  9811=>"001111111",
  9812=>"000000000",
  9813=>"111111011",
  9814=>"100100111",
  9815=>"000000000",
  9816=>"111111111",
  9817=>"000000000",
  9818=>"111111111",
  9819=>"000000000",
  9820=>"101100010",
  9821=>"000000000",
  9822=>"011111111",
  9823=>"100110100",
  9824=>"100111111",
  9825=>"000100100",
  9826=>"111111111",
  9827=>"111111101",
  9828=>"100000011",
  9829=>"011000000",
  9830=>"111000110",
  9831=>"111111000",
  9832=>"000000000",
  9833=>"010000000",
  9834=>"000000010",
  9835=>"010011011",
  9836=>"111111111",
  9837=>"100000000",
  9838=>"000001000",
  9839=>"001101111",
  9840=>"000000000",
  9841=>"111111111",
  9842=>"110100110",
  9843=>"101111111",
  9844=>"111111111",
  9845=>"000100110",
  9846=>"000000000",
  9847=>"011111111",
  9848=>"000000000",
  9849=>"011000000",
  9850=>"000010010",
  9851=>"111111000",
  9852=>"000100000",
  9853=>"011011011",
  9854=>"111111111",
  9855=>"110111111",
  9856=>"111111111",
  9857=>"110110011",
  9858=>"111011001",
  9859=>"011011111",
  9860=>"111010000",
  9861=>"100000111",
  9862=>"110110110",
  9863=>"000000000",
  9864=>"000000000",
  9865=>"010001001",
  9866=>"000000001",
  9867=>"001011001",
  9868=>"111111111",
  9869=>"000110111",
  9870=>"000000000",
  9871=>"001000000",
  9872=>"111111111",
  9873=>"111111111",
  9874=>"000000000",
  9875=>"000111111",
  9876=>"000000111",
  9877=>"011011011",
  9878=>"000000000",
  9879=>"000000000",
  9880=>"000111000",
  9881=>"100100000",
  9882=>"000000000",
  9883=>"111100100",
  9884=>"100010011",
  9885=>"011001001",
  9886=>"011011111",
  9887=>"001001001",
  9888=>"000000101",
  9889=>"000000000",
  9890=>"111111111",
  9891=>"111111111",
  9892=>"000000000",
  9893=>"001001111",
  9894=>"111111111",
  9895=>"000000000",
  9896=>"000000000",
  9897=>"111111111",
  9898=>"000000000",
  9899=>"111000111",
  9900=>"111111110",
  9901=>"111111111",
  9902=>"000000000",
  9903=>"000000111",
  9904=>"000111111",
  9905=>"000001000",
  9906=>"111111111",
  9907=>"001100000",
  9908=>"001000000",
  9909=>"000000000",
  9910=>"001000000",
  9911=>"000001001",
  9912=>"100111111",
  9913=>"000000000",
  9914=>"000000011",
  9915=>"000000010",
  9916=>"000000000",
  9917=>"101111111",
  9918=>"111000000",
  9919=>"000010110",
  9920=>"111100111",
  9921=>"011111011",
  9922=>"110110000",
  9923=>"000000000",
  9924=>"111111111",
  9925=>"111111111",
  9926=>"111110100",
  9927=>"111111111",
  9928=>"000000100",
  9929=>"001000000",
  9930=>"111101111",
  9931=>"111111111",
  9932=>"000000001",
  9933=>"111111111",
  9934=>"000011101",
  9935=>"000000000",
  9936=>"000000000",
  9937=>"001100111",
  9938=>"001000111",
  9939=>"000000000",
  9940=>"111111111",
  9941=>"110100000",
  9942=>"100000000",
  9943=>"111101111",
  9944=>"111111111",
  9945=>"001101111",
  9946=>"000000000",
  9947=>"000000000",
  9948=>"010000000",
  9949=>"000010000",
  9950=>"000000111",
  9951=>"000000011",
  9952=>"111111111",
  9953=>"100000111",
  9954=>"111111010",
  9955=>"110000011",
  9956=>"111100110",
  9957=>"000000000",
  9958=>"000110110",
  9959=>"011001001",
  9960=>"000000001",
  9961=>"011000111",
  9962=>"111110111",
  9963=>"000000000",
  9964=>"000000000",
  9965=>"111111111",
  9966=>"111111001",
  9967=>"000000001",
  9968=>"111011011",
  9969=>"000000000",
  9970=>"000000110",
  9971=>"000000000",
  9972=>"111111111",
  9973=>"000000000",
  9974=>"111111000",
  9975=>"000000111",
  9976=>"111110000",
  9977=>"000000000",
  9978=>"000000000",
  9979=>"000000000",
  9980=>"010110110",
  9981=>"111111111",
  9982=>"000000000",
  9983=>"100110111",
  9984=>"000000000",
  9985=>"111111110",
  9986=>"000000000",
  9987=>"000000000",
  9988=>"000000000",
  9989=>"000000000",
  9990=>"000000111",
  9991=>"111100111",
  9992=>"111111111",
  9993=>"001000000",
  9994=>"000000001",
  9995=>"100000111",
  9996=>"110000000",
  9997=>"111111111",
  9998=>"000000000",
  9999=>"111110111",
  10000=>"001011000",
  10001=>"111000000",
  10002=>"011001001",
  10003=>"110000000",
  10004=>"111111111",
  10005=>"000000000",
  10006=>"010110111",
  10007=>"000010000",
  10008=>"111111111",
  10009=>"000000000",
  10010=>"011000011",
  10011=>"000000000",
  10012=>"101100101",
  10013=>"111111111",
  10014=>"000110000",
  10015=>"111000000",
  10016=>"000000000",
  10017=>"111000000",
  10018=>"100100111",
  10019=>"111111111",
  10020=>"000000000",
  10021=>"000000100",
  10022=>"000000001",
  10023=>"111011111",
  10024=>"000100100",
  10025=>"000111111",
  10026=>"111100000",
  10027=>"111111111",
  10028=>"000011000",
  10029=>"111110110",
  10030=>"111111111",
  10031=>"010000000",
  10032=>"001001001",
  10033=>"011011011",
  10034=>"110111111",
  10035=>"111111010",
  10036=>"000000000",
  10037=>"000011001",
  10038=>"000100111",
  10039=>"000100110",
  10040=>"000000010",
  10041=>"111100100",
  10042=>"110110110",
  10043=>"000000000",
  10044=>"000010000",
  10045=>"110110000",
  10046=>"111111111",
  10047=>"111111111",
  10048=>"000000010",
  10049=>"101101111",
  10050=>"100000000",
  10051=>"111111111",
  10052=>"000000111",
  10053=>"111111111",
  10054=>"111111111",
  10055=>"110110110",
  10056=>"111111111",
  10057=>"111001101",
  10058=>"100100110",
  10059=>"000000000",
  10060=>"000011011",
  10061=>"111111111",
  10062=>"000000000",
  10063=>"111111110",
  10064=>"000000000",
  10065=>"000000000",
  10066=>"000000000",
  10067=>"100000000",
  10068=>"000000000",
  10069=>"010010011",
  10070=>"011011001",
  10071=>"111100100",
  10072=>"000000001",
  10073=>"000111111",
  10074=>"111100111",
  10075=>"000000111",
  10076=>"111011110",
  10077=>"111111111",
  10078=>"000000001",
  10079=>"110111111",
  10080=>"111111111",
  10081=>"101001111",
  10082=>"100100111",
  10083=>"000000000",
  10084=>"000000101",
  10085=>"000000100",
  10086=>"011010110",
  10087=>"000000000",
  10088=>"001001000",
  10089=>"000000111",
  10090=>"000000001",
  10091=>"001110110",
  10092=>"011001001",
  10093=>"010111111",
  10094=>"000010010",
  10095=>"111111111",
  10096=>"000000100",
  10097=>"111101000",
  10098=>"111000000",
  10099=>"110110110",
  10100=>"000000000",
  10101=>"111111111",
  10102=>"000000000",
  10103=>"100111111",
  10104=>"000011111",
  10105=>"000000000",
  10106=>"111111110",
  10107=>"110001000",
  10108=>"111111010",
  10109=>"111100000",
  10110=>"000001111",
  10111=>"111000000",
  10112=>"111111001",
  10113=>"111111111",
  10114=>"001011010",
  10115=>"111111111",
  10116=>"000000000",
  10117=>"000000000",
  10118=>"001001000",
  10119=>"111111111",
  10120=>"001011000",
  10121=>"000000001",
  10122=>"111111001",
  10123=>"000000111",
  10124=>"111111111",
  10125=>"001101111",
  10126=>"100000000",
  10127=>"010011010",
  10128=>"101000000",
  10129=>"100000001",
  10130=>"011000000",
  10131=>"011011000",
  10132=>"110101101",
  10133=>"000000111",
  10134=>"111111111",
  10135=>"000000000",
  10136=>"000000000",
  10137=>"000000000",
  10138=>"100000001",
  10139=>"111111111",
  10140=>"000011111",
  10141=>"000000001",
  10142=>"000000000",
  10143=>"111111111",
  10144=>"000010000",
  10145=>"111001111",
  10146=>"100000000",
  10147=>"000000000",
  10148=>"111110010",
  10149=>"000000101",
  10150=>"111111111",
  10151=>"011011000",
  10152=>"000100100",
  10153=>"001111111",
  10154=>"111111111",
  10155=>"011111111",
  10156=>"111100000",
  10157=>"110111101",
  10158=>"001111000",
  10159=>"111111001",
  10160=>"100001000",
  10161=>"000000000",
  10162=>"111110111",
  10163=>"011001011",
  10164=>"011111111",
  10165=>"000000000",
  10166=>"111101101",
  10167=>"000000011",
  10168=>"000000000",
  10169=>"000000000",
  10170=>"001001001",
  10171=>"111111111",
  10172=>"000011111",
  10173=>"011001000",
  10174=>"000000000",
  10175=>"000000000",
  10176=>"110111011",
  10177=>"000000100",
  10178=>"000000000",
  10179=>"111111111",
  10180=>"000000011",
  10181=>"111011011",
  10182=>"000000000",
  10183=>"110000000",
  10184=>"000000000",
  10185=>"001011011",
  10186=>"000100111",
  10187=>"000110111",
  10188=>"000000000",
  10189=>"011011111",
  10190=>"011000000",
  10191=>"000000000",
  10192=>"000000000",
  10193=>"111111011",
  10194=>"111101111",
  10195=>"111111111",
  10196=>"000000100",
  10197=>"000111111",
  10198=>"111111111",
  10199=>"000010110",
  10200=>"000000000",
  10201=>"111011111",
  10202=>"000000011",
  10203=>"000000000",
  10204=>"000001111",
  10205=>"111111111",
  10206=>"001000111",
  10207=>"010000001",
  10208=>"000000000",
  10209=>"001111111",
  10210=>"111111011",
  10211=>"000001101",
  10212=>"001101001",
  10213=>"101100000",
  10214=>"000010000",
  10215=>"010000010",
  10216=>"111011101",
  10217=>"111111110",
  10218=>"000001011",
  10219=>"111111111",
  10220=>"001000011",
  10221=>"000000000",
  10222=>"111111111",
  10223=>"000000001",
  10224=>"000000000",
  10225=>"001001111",
  10226=>"111000000",
  10227=>"000000000",
  10228=>"100100111",
  10229=>"100000111",
  10230=>"000000000",
  10231=>"000000000",
  10232=>"000000110",
  10233=>"010010010",
  10234=>"111111011",
  10235=>"110110111",
  10236=>"001001001",
  10237=>"000000100",
  10238=>"111111101",
  10239=>"001000000",
  10240=>"010000010",
  10241=>"110111111",
  10242=>"000001011",
  10243=>"000100100",
  10244=>"111111111",
  10245=>"000000000",
  10246=>"011011011",
  10247=>"111111111",
  10248=>"111111111",
  10249=>"111111011",
  10250=>"111111111",
  10251=>"000110110",
  10252=>"111101111",
  10253=>"101000000",
  10254=>"011001100",
  10255=>"111001000",
  10256=>"000100000",
  10257=>"001100000",
  10258=>"111111111",
  10259=>"110111111",
  10260=>"111111111",
  10261=>"111101001",
  10262=>"000000111",
  10263=>"000000000",
  10264=>"111001100",
  10265=>"100000000",
  10266=>"000000000",
  10267=>"000000000",
  10268=>"011011111",
  10269=>"111010010",
  10270=>"000000111",
  10271=>"111100100",
  10272=>"010010000",
  10273=>"000000000",
  10274=>"110111111",
  10275=>"000000100",
  10276=>"001000011",
  10277=>"001001000",
  10278=>"000000000",
  10279=>"111111101",
  10280=>"111111111",
  10281=>"000000000",
  10282=>"111111101",
  10283=>"011000000",
  10284=>"000000000",
  10285=>"000110110",
  10286=>"011111111",
  10287=>"000000000",
  10288=>"000000000",
  10289=>"111000000",
  10290=>"111001111",
  10291=>"100110100",
  10292=>"000000001",
  10293=>"001001001",
  10294=>"111111100",
  10295=>"100001000",
  10296=>"000000001",
  10297=>"011011111",
  10298=>"111111111",
  10299=>"110100100",
  10300=>"000000000",
  10301=>"000000100",
  10302=>"100110000",
  10303=>"111111111",
  10304=>"010000000",
  10305=>"000000000",
  10306=>"000000101",
  10307=>"000000000",
  10308=>"111111101",
  10309=>"000000000",
  10310=>"111111110",
  10311=>"111111111",
  10312=>"000000100",
  10313=>"000000000",
  10314=>"000110110",
  10315=>"011000101",
  10316=>"011011111",
  10317=>"001111111",
  10318=>"010110110",
  10319=>"000000110",
  10320=>"111110110",
  10321=>"000011000",
  10322=>"111101100",
  10323=>"110100111",
  10324=>"000000001",
  10325=>"101001000",
  10326=>"010011000",
  10327=>"001001001",
  10328=>"111111111",
  10329=>"000000000",
  10330=>"111111111",
  10331=>"000000000",
  10332=>"000000001",
  10333=>"000000110",
  10334=>"001000000",
  10335=>"111111001",
  10336=>"000000000",
  10337=>"000111111",
  10338=>"000010000",
  10339=>"000000000",
  10340=>"101101111",
  10341=>"011001111",
  10342=>"000000000",
  10343=>"111100000",
  10344=>"000000111",
  10345=>"011111111",
  10346=>"111001011",
  10347=>"111010010",
  10348=>"111111100",
  10349=>"011011011",
  10350=>"111111001",
  10351=>"000000000",
  10352=>"000000000",
  10353=>"010000111",
  10354=>"111111111",
  10355=>"100100110",
  10356=>"011000000",
  10357=>"111111111",
  10358=>"000000000",
  10359=>"001000001",
  10360=>"100000010",
  10361=>"011011010",
  10362=>"011000111",
  10363=>"111111111",
  10364=>"010001000",
  10365=>"111001001",
  10366=>"000100100",
  10367=>"111011000",
  10368=>"000000000",
  10369=>"101111110",
  10370=>"000010011",
  10371=>"110110111",
  10372=>"011011000",
  10373=>"010011011",
  10374=>"100001100",
  10375=>"101111111",
  10376=>"111111000",
  10377=>"100100000",
  10378=>"000001001",
  10379=>"111011011",
  10380=>"010000100",
  10381=>"000011111",
  10382=>"111111000",
  10383=>"111111011",
  10384=>"111111111",
  10385=>"000111101",
  10386=>"001011011",
  10387=>"011001001",
  10388=>"001001001",
  10389=>"000010100",
  10390=>"111111111",
  10391=>"000000000",
  10392=>"011111111",
  10393=>"010100100",
  10394=>"011011000",
  10395=>"111111111",
  10396=>"000000000",
  10397=>"011000001",
  10398=>"000101101",
  10399=>"111111111",
  10400=>"000110100",
  10401=>"111011000",
  10402=>"111001001",
  10403=>"100000100",
  10404=>"001001001",
  10405=>"001000000",
  10406=>"111111111",
  10407=>"110100100",
  10408=>"110000000",
  10409=>"110100000",
  10410=>"011111011",
  10411=>"000000100",
  10412=>"001011111",
  10413=>"001001000",
  10414=>"000101111",
  10415=>"100100110",
  10416=>"111100001",
  10417=>"000000000",
  10418=>"000000000",
  10419=>"000000101",
  10420=>"011011111",
  10421=>"000000000",
  10422=>"110100111",
  10423=>"111011111",
  10424=>"100100100",
  10425=>"111111011",
  10426=>"001001001",
  10427=>"000011111",
  10428=>"000010000",
  10429=>"000000111",
  10430=>"000000000",
  10431=>"111111111",
  10432=>"111111101",
  10433=>"001001111",
  10434=>"111011011",
  10435=>"000000000",
  10436=>"000000000",
  10437=>"011011001",
  10438=>"001001001",
  10439=>"111111111",
  10440=>"000000000",
  10441=>"111111010",
  10442=>"010000100",
  10443=>"111111111",
  10444=>"100000100",
  10445=>"110110100",
  10446=>"100110100",
  10447=>"000000000",
  10448=>"000000000",
  10449=>"000000000",
  10450=>"000000000",
  10451=>"001000000",
  10452=>"111111111",
  10453=>"000000000",
  10454=>"110111010",
  10455=>"101101100",
  10456=>"111111111",
  10457=>"000001101",
  10458=>"100100100",
  10459=>"011111111",
  10460=>"100111111",
  10461=>"100000111",
  10462=>"111111110",
  10463=>"000001001",
  10464=>"000000000",
  10465=>"000001000",
  10466=>"111111110",
  10467=>"011011111",
  10468=>"111001000",
  10469=>"100110110",
  10470=>"011001000",
  10471=>"000000110",
  10472=>"000100111",
  10473=>"111100000",
  10474=>"011111111",
  10475=>"111111111",
  10476=>"000000000",
  10477=>"100000000",
  10478=>"000100111",
  10479=>"000011011",
  10480=>"111111111",
  10481=>"111100111",
  10482=>"010000010",
  10483=>"010010100",
  10484=>"011011111",
  10485=>"111111111",
  10486=>"111100100",
  10487=>"000000010",
  10488=>"010111111",
  10489=>"001000000",
  10490=>"100000010",
  10491=>"000000000",
  10492=>"111110111",
  10493=>"000000000",
  10494=>"001001111",
  10495=>"111111111",
  10496=>"011000111",
  10497=>"001000001",
  10498=>"111111111",
  10499=>"100100110",
  10500=>"000000000",
  10501=>"111111111",
  10502=>"100100001",
  10503=>"111010011",
  10504=>"000000101",
  10505=>"000000000",
  10506=>"001000000",
  10507=>"011001101",
  10508=>"000111111",
  10509=>"111111111",
  10510=>"000101111",
  10511=>"111001000",
  10512=>"010001111",
  10513=>"011000000",
  10514=>"000000111",
  10515=>"111011011",
  10516=>"010010000",
  10517=>"111100000",
  10518=>"001001001",
  10519=>"111101101",
  10520=>"100001101",
  10521=>"000111100",
  10522=>"000000000",
  10523=>"000111111",
  10524=>"111000000",
  10525=>"000000111",
  10526=>"011001001",
  10527=>"000000000",
  10528=>"111000011",
  10529=>"110111000",
  10530=>"010010111",
  10531=>"010000000",
  10532=>"111011111",
  10533=>"111100000",
  10534=>"100110100",
  10535=>"111011111",
  10536=>"001111011",
  10537=>"111110110",
  10538=>"110100000",
  10539=>"000000000",
  10540=>"000000010",
  10541=>"111110000",
  10542=>"000001000",
  10543=>"001000111",
  10544=>"111001111",
  10545=>"000000100",
  10546=>"101101111",
  10547=>"001100000",
  10548=>"111111111",
  10549=>"000000000",
  10550=>"111111111",
  10551=>"111111111",
  10552=>"000000110",
  10553=>"011001011",
  10554=>"000000000",
  10555=>"100000000",
  10556=>"011011000",
  10557=>"111111111",
  10558=>"011011111",
  10559=>"001001001",
  10560=>"000110110",
  10561=>"110111111",
  10562=>"000000111",
  10563=>"000000000",
  10564=>"111101111",
  10565=>"100100111",
  10566=>"000000000",
  10567=>"001111111",
  10568=>"111111111",
  10569=>"000100000",
  10570=>"111010110",
  10571=>"100000101",
  10572=>"100000000",
  10573=>"111111111",
  10574=>"001111111",
  10575=>"111101111",
  10576=>"100000000",
  10577=>"111000001",
  10578=>"000000111",
  10579=>"011111111",
  10580=>"000101001",
  10581=>"001011111",
  10582=>"111111111",
  10583=>"000000000",
  10584=>"000000000",
  10585=>"011111111",
  10586=>"110111111",
  10587=>"111111110",
  10588=>"000000000",
  10589=>"000000111",
  10590=>"000000000",
  10591=>"110000100",
  10592=>"111111111",
  10593=>"000010111",
  10594=>"100100101",
  10595=>"111111111",
  10596=>"111111110",
  10597=>"000000001",
  10598=>"000000000",
  10599=>"000000000",
  10600=>"011001001",
  10601=>"000000000",
  10602=>"001000011",
  10603=>"000110111",
  10604=>"001011001",
  10605=>"011111111",
  10606=>"011001000",
  10607=>"100111111",
  10608=>"000000001",
  10609=>"110111111",
  10610=>"000000110",
  10611=>"110111111",
  10612=>"011010010",
  10613=>"011001101",
  10614=>"111111111",
  10615=>"111111111",
  10616=>"000100100",
  10617=>"111110000",
  10618=>"100000100",
  10619=>"011011111",
  10620=>"000000000",
  10621=>"111111111",
  10622=>"110000000",
  10623=>"000000000",
  10624=>"000000001",
  10625=>"010000101",
  10626=>"011000000",
  10627=>"111100111",
  10628=>"011000000",
  10629=>"000000000",
  10630=>"101101111",
  10631=>"011011011",
  10632=>"101111111",
  10633=>"111111111",
  10634=>"000000100",
  10635=>"111111111",
  10636=>"111001101",
  10637=>"000100100",
  10638=>"101100101",
  10639=>"111110111",
  10640=>"000110111",
  10641=>"110111111",
  10642=>"111000000",
  10643=>"000000001",
  10644=>"010011111",
  10645=>"011011111",
  10646=>"000110110",
  10647=>"001001111",
  10648=>"111111111",
  10649=>"000000011",
  10650=>"011111111",
  10651=>"111101101",
  10652=>"000000000",
  10653=>"111111111",
  10654=>"110111111",
  10655=>"101100000",
  10656=>"011000110",
  10657=>"111110110",
  10658=>"110110000",
  10659=>"100110110",
  10660=>"111111001",
  10661=>"000000000",
  10662=>"000000000",
  10663=>"111101111",
  10664=>"111111111",
  10665=>"000000000",
  10666=>"111111110",
  10667=>"000100110",
  10668=>"000000000",
  10669=>"000111111",
  10670=>"111001100",
  10671=>"011011111",
  10672=>"000000111",
  10673=>"011011010",
  10674=>"011111111",
  10675=>"110111110",
  10676=>"111111001",
  10677=>"000100110",
  10678=>"101111111",
  10679=>"000000000",
  10680=>"111000000",
  10681=>"110111111",
  10682=>"000000000",
  10683=>"000100111",
  10684=>"000000010",
  10685=>"111010111",
  10686=>"010110000",
  10687=>"101000100",
  10688=>"111010110",
  10689=>"000000000",
  10690=>"111111111",
  10691=>"001001000",
  10692=>"000010110",
  10693=>"000111011",
  10694=>"111111111",
  10695=>"000111011",
  10696=>"001111111",
  10697=>"001001011",
  10698=>"010000000",
  10699=>"001001011",
  10700=>"000000000",
  10701=>"001000000",
  10702=>"111111111",
  10703=>"100100100",
  10704=>"010000000",
  10705=>"000111111",
  10706=>"000000000",
  10707=>"110000000",
  10708=>"111011011",
  10709=>"111111111",
  10710=>"000110110",
  10711=>"110000001",
  10712=>"111111111",
  10713=>"000100100",
  10714=>"001000000",
  10715=>"000000000",
  10716=>"001000000",
  10717=>"010111111",
  10718=>"111111111",
  10719=>"111111111",
  10720=>"100000000",
  10721=>"111011011",
  10722=>"000000000",
  10723=>"111111111",
  10724=>"000000000",
  10725=>"000011111",
  10726=>"100100100",
  10727=>"000000000",
  10728=>"011001000",
  10729=>"000000000",
  10730=>"111110000",
  10731=>"011011001",
  10732=>"010010011",
  10733=>"100000000",
  10734=>"000000000",
  10735=>"110111111",
  10736=>"001001001",
  10737=>"000011111",
  10738=>"000011001",
  10739=>"111011011",
  10740=>"011110110",
  10741=>"000000000",
  10742=>"000000000",
  10743=>"001001111",
  10744=>"000000000",
  10745=>"000000000",
  10746=>"011011111",
  10747=>"111100000",
  10748=>"000000001",
  10749=>"100000100",
  10750=>"000000000",
  10751=>"001000110",
  10752=>"001001000",
  10753=>"000111111",
  10754=>"000111111",
  10755=>"000000000",
  10756=>"010110110",
  10757=>"100100000",
  10758=>"000000000",
  10759=>"111111111",
  10760=>"111001000",
  10761=>"111111111",
  10762=>"001111111",
  10763=>"111001000",
  10764=>"000100110",
  10765=>"110100111",
  10766=>"111001000",
  10767=>"010000111",
  10768=>"010000000",
  10769=>"000000001",
  10770=>"111010010",
  10771=>"001001011",
  10772=>"000000111",
  10773=>"111000000",
  10774=>"111111000",
  10775=>"111111111",
  10776=>"000001001",
  10777=>"001111111",
  10778=>"000000000",
  10779=>"100110110",
  10780=>"110111111",
  10781=>"111111001",
  10782=>"011011011",
  10783=>"111111111",
  10784=>"000010000",
  10785=>"100111000",
  10786=>"000000000",
  10787=>"001011000",
  10788=>"111111111",
  10789=>"111000001",
  10790=>"000000000",
  10791=>"100000100",
  10792=>"000000000",
  10793=>"011000000",
  10794=>"111111111",
  10795=>"000000011",
  10796=>"111111111",
  10797=>"000000000",
  10798=>"000000011",
  10799=>"111111111",
  10800=>"000011000",
  10801=>"011111111",
  10802=>"001011111",
  10803=>"111101111",
  10804=>"000000000",
  10805=>"000000000",
  10806=>"111111111",
  10807=>"000000000",
  10808=>"110110111",
  10809=>"111011001",
  10810=>"000000000",
  10811=>"011111111",
  10812=>"000000000",
  10813=>"010000000",
  10814=>"111100111",
  10815=>"000100111",
  10816=>"011011000",
  10817=>"000000000",
  10818=>"000000001",
  10819=>"111111111",
  10820=>"111111011",
  10821=>"011111111",
  10822=>"111111000",
  10823=>"000000000",
  10824=>"011011111",
  10825=>"111111111",
  10826=>"000000000",
  10827=>"111001001",
  10828=>"111111010",
  10829=>"000100111",
  10830=>"001000000",
  10831=>"111111000",
  10832=>"000110100",
  10833=>"101000000",
  10834=>"111000000",
  10835=>"010001001",
  10836=>"000000000",
  10837=>"000000000",
  10838=>"001011000",
  10839=>"000010000",
  10840=>"000011111",
  10841=>"001001111",
  10842=>"111100000",
  10843=>"100000000",
  10844=>"000001001",
  10845=>"001001111",
  10846=>"000100111",
  10847=>"111111111",
  10848=>"111111111",
  10849=>"111011011",
  10850=>"011111111",
  10851=>"000000000",
  10852=>"000000111",
  10853=>"100100111",
  10854=>"110111111",
  10855=>"000000000",
  10856=>"000101110",
  10857=>"111111111",
  10858=>"111101100",
  10859=>"000000000",
  10860=>"000110111",
  10861=>"000000000",
  10862=>"101001000",
  10863=>"000000000",
  10864=>"011011001",
  10865=>"000000101",
  10866=>"000000000",
  10867=>"000000000",
  10868=>"100010000",
  10869=>"000000100",
  10870=>"000000111",
  10871=>"111111001",
  10872=>"000000000",
  10873=>"111100111",
  10874=>"000000000",
  10875=>"111000011",
  10876=>"000000000",
  10877=>"000100111",
  10878=>"011111011",
  10879=>"111111111",
  10880=>"000000000",
  10881=>"000000000",
  10882=>"111111111",
  10883=>"111100100",
  10884=>"111111111",
  10885=>"000000110",
  10886=>"111000000",
  10887=>"111000000",
  10888=>"111001000",
  10889=>"111111110",
  10890=>"000000000",
  10891=>"110111111",
  10892=>"000000000",
  10893=>"111110111",
  10894=>"000000000",
  10895=>"111111111",
  10896=>"001000001",
  10897=>"000000101",
  10898=>"000000000",
  10899=>"111111111",
  10900=>"111111110",
  10901=>"011011110",
  10902=>"110100111",
  10903=>"000000000",
  10904=>"000000000",
  10905=>"110110111",
  10906=>"111111111",
  10907=>"111111010",
  10908=>"100000011",
  10909=>"000000000",
  10910=>"111111100",
  10911=>"111101001",
  10912=>"000000000",
  10913=>"001000000",
  10914=>"111111111",
  10915=>"110110011",
  10916=>"000111010",
  10917=>"111111111",
  10918=>"000111000",
  10919=>"000000001",
  10920=>"000000000",
  10921=>"001001111",
  10922=>"111111111",
  10923=>"111111000",
  10924=>"110010000",
  10925=>"110000000",
  10926=>"111011111",
  10927=>"001001011",
  10928=>"111111000",
  10929=>"111101111",
  10930=>"000001000",
  10931=>"111111000",
  10932=>"000110111",
  10933=>"111111111",
  10934=>"000111111",
  10935=>"111101111",
  10936=>"000000110",
  10937=>"111111001",
  10938=>"000010000",
  10939=>"110001111",
  10940=>"000000000",
  10941=>"111001001",
  10942=>"111110110",
  10943=>"001101111",
  10944=>"000000000",
  10945=>"100000101",
  10946=>"000101111",
  10947=>"001111111",
  10948=>"010000111",
  10949=>"000000000",
  10950=>"000000000",
  10951=>"111011111",
  10952=>"000000000",
  10953=>"101001011",
  10954=>"010100000",
  10955=>"000110000",
  10956=>"001000000",
  10957=>"001001011",
  10958=>"111001111",
  10959=>"000000001",
  10960=>"111111000",
  10961=>"000000000",
  10962=>"001001001",
  10963=>"111111110",
  10964=>"111111111",
  10965=>"111111111",
  10966=>"000000000",
  10967=>"011001100",
  10968=>"001001111",
  10969=>"110110111",
  10970=>"000000000",
  10971=>"111111111",
  10972=>"011000000",
  10973=>"000101111",
  10974=>"111111100",
  10975=>"000110111",
  10976=>"000000000",
  10977=>"000000110",
  10978=>"100110010",
  10979=>"000000000",
  10980=>"000110111",
  10981=>"000000000",
  10982=>"110110111",
  10983=>"111010000",
  10984=>"000000000",
  10985=>"101101111",
  10986=>"111111111",
  10987=>"111111111",
  10988=>"111101101",
  10989=>"111111111",
  10990=>"000001001",
  10991=>"010000000",
  10992=>"000000111",
  10993=>"110111111",
  10994=>"001001000",
  10995=>"101101111",
  10996=>"110110111",
  10997=>"110100111",
  10998=>"101101111",
  10999=>"011000000",
  11000=>"100000000",
  11001=>"111111101",
  11002=>"110110110",
  11003=>"000000000",
  11004=>"100000000",
  11005=>"110111111",
  11006=>"000001001",
  11007=>"111111111",
  11008=>"111111111",
  11009=>"001001001",
  11010=>"111000010",
  11011=>"000000000",
  11012=>"111000000",
  11013=>"100000000",
  11014=>"111110000",
  11015=>"000000000",
  11016=>"111011000",
  11017=>"000000101",
  11018=>"111111111",
  11019=>"001001100",
  11020=>"100100000",
  11021=>"000000000",
  11022=>"111111111",
  11023=>"111111000",
  11024=>"000000001",
  11025=>"100000000",
  11026=>"000110000",
  11027=>"111111011",
  11028=>"111011000",
  11029=>"110010111",
  11030=>"111000001",
  11031=>"000000101",
  11032=>"001001000",
  11033=>"101000000",
  11034=>"000000001",
  11035=>"000000000",
  11036=>"111111111",
  11037=>"110100101",
  11038=>"100111111",
  11039=>"000000000",
  11040=>"111111111",
  11041=>"111111111",
  11042=>"100110000",
  11043=>"111111100",
  11044=>"000000000",
  11045=>"111111111",
  11046=>"111111100",
  11047=>"000000000",
  11048=>"000000000",
  11049=>"111111111",
  11050=>"000000000",
  11051=>"000000000",
  11052=>"011000000",
  11053=>"000001111",
  11054=>"111111000",
  11055=>"111101000",
  11056=>"000000010",
  11057=>"111111000",
  11058=>"110110100",
  11059=>"000100100",
  11060=>"111111111",
  11061=>"110111111",
  11062=>"000000000",
  11063=>"010111011",
  11064=>"110111111",
  11065=>"111111111",
  11066=>"000111111",
  11067=>"100111111",
  11068=>"000000001",
  11069=>"101001000",
  11070=>"000000111",
  11071=>"000000000",
  11072=>"000000000",
  11073=>"101111111",
  11074=>"100000111",
  11075=>"111000101",
  11076=>"111111111",
  11077=>"111111111",
  11078=>"111111111",
  11079=>"000000000",
  11080=>"011000001",
  11081=>"111111111",
  11082=>"111000001",
  11083=>"001001000",
  11084=>"100111111",
  11085=>"111110100",
  11086=>"000000000",
  11087=>"000000000",
  11088=>"011000000",
  11089=>"100100101",
  11090=>"101100000",
  11091=>"000001000",
  11092=>"000000000",
  11093=>"001001001",
  11094=>"111111111",
  11095=>"111111111",
  11096=>"111101111",
  11097=>"000001000",
  11098=>"010110101",
  11099=>"111111111",
  11100=>"100000000",
  11101=>"000000000",
  11102=>"101001000",
  11103=>"000000001",
  11104=>"111111111",
  11105=>"111111111",
  11106=>"101101111",
  11107=>"000000000",
  11108=>"111110110",
  11109=>"000100001",
  11110=>"000000000",
  11111=>"111110000",
  11112=>"100000000",
  11113=>"000000000",
  11114=>"111111111",
  11115=>"000111111",
  11116=>"001001000",
  11117=>"011000000",
  11118=>"111111111",
  11119=>"000000001",
  11120=>"000100011",
  11121=>"000000011",
  11122=>"001001001",
  11123=>"111111000",
  11124=>"111111111",
  11125=>"011111111",
  11126=>"000000000",
  11127=>"000000000",
  11128=>"000000111",
  11129=>"111011010",
  11130=>"000000000",
  11131=>"010010111",
  11132=>"010111110",
  11133=>"000011011",
  11134=>"000000000",
  11135=>"001001111",
  11136=>"111011011",
  11137=>"000011011",
  11138=>"110110110",
  11139=>"000000100",
  11140=>"111111111",
  11141=>"000000000",
  11142=>"000000000",
  11143=>"000000000",
  11144=>"111111000",
  11145=>"111001000",
  11146=>"111111000",
  11147=>"111111111",
  11148=>"111111111",
  11149=>"111101111",
  11150=>"001000001",
  11151=>"000000000",
  11152=>"000000101",
  11153=>"000000000",
  11154=>"111111111",
  11155=>"000000100",
  11156=>"111011000",
  11157=>"000010010",
  11158=>"111111111",
  11159=>"000001011",
  11160=>"000000111",
  11161=>"111111111",
  11162=>"000000111",
  11163=>"000001111",
  11164=>"001111111",
  11165=>"111000111",
  11166=>"111111011",
  11167=>"111000000",
  11168=>"110101111",
  11169=>"001000000",
  11170=>"001000001",
  11171=>"000101000",
  11172=>"100100111",
  11173=>"010000000",
  11174=>"000000000",
  11175=>"001111111",
  11176=>"000000000",
  11177=>"000000000",
  11178=>"111111111",
  11179=>"101111010",
  11180=>"111111101",
  11181=>"111001100",
  11182=>"001000000",
  11183=>"000000011",
  11184=>"000000000",
  11185=>"111111001",
  11186=>"100100000",
  11187=>"111111111",
  11188=>"000111111",
  11189=>"111111111",
  11190=>"111111111",
  11191=>"011111001",
  11192=>"111111110",
  11193=>"011000000",
  11194=>"010000000",
  11195=>"111111111",
  11196=>"110100000",
  11197=>"001111111",
  11198=>"001000000",
  11199=>"101000001",
  11200=>"111111111",
  11201=>"000100111",
  11202=>"011011011",
  11203=>"000000000",
  11204=>"000010010",
  11205=>"010000000",
  11206=>"000000001",
  11207=>"000001011",
  11208=>"111110000",
  11209=>"000000000",
  11210=>"000001000",
  11211=>"011000000",
  11212=>"111000000",
  11213=>"001011011",
  11214=>"011001001",
  11215=>"111111111",
  11216=>"001001000",
  11217=>"111110110",
  11218=>"111111101",
  11219=>"000011011",
  11220=>"111101111",
  11221=>"000100110",
  11222=>"100000000",
  11223=>"001101001",
  11224=>"101111101",
  11225=>"100100110",
  11226=>"111111111",
  11227=>"000111111",
  11228=>"111111111",
  11229=>"001001111",
  11230=>"111111111",
  11231=>"000000000",
  11232=>"000000000",
  11233=>"000000001",
  11234=>"111111111",
  11235=>"111111011",
  11236=>"100111111",
  11237=>"000100110",
  11238=>"000000000",
  11239=>"000000100",
  11240=>"111001001",
  11241=>"111111111",
  11242=>"000000000",
  11243=>"111111001",
  11244=>"111001001",
  11245=>"111111111",
  11246=>"110111110",
  11247=>"010011011",
  11248=>"000000000",
  11249=>"011011111",
  11250=>"111000000",
  11251=>"000000000",
  11252=>"111000000",
  11253=>"110100101",
  11254=>"000000000",
  11255=>"110010010",
  11256=>"001011011",
  11257=>"111111111",
  11258=>"000000000",
  11259=>"000000000",
  11260=>"111111011",
  11261=>"111011011",
  11262=>"001000000",
  11263=>"001000000",
  11264=>"010000111",
  11265=>"111111111",
  11266=>"111111110",
  11267=>"000101000",
  11268=>"111001001",
  11269=>"111111000",
  11270=>"111000000",
  11271=>"011000111",
  11272=>"100111111",
  11273=>"111100111",
  11274=>"111110001",
  11275=>"101100100",
  11276=>"100000110",
  11277=>"111011111",
  11278=>"111000000",
  11279=>"000000000",
  11280=>"100111111",
  11281=>"111001011",
  11282=>"001000001",
  11283=>"010101110",
  11284=>"000111000",
  11285=>"010111111",
  11286=>"000100000",
  11287=>"110000111",
  11288=>"101000111",
  11289=>"100110000",
  11290=>"110111000",
  11291=>"101001000",
  11292=>"111111111",
  11293=>"000000111",
  11294=>"011000111",
  11295=>"000110111",
  11296=>"000011000",
  11297=>"100000111",
  11298=>"000000000",
  11299=>"100101000",
  11300=>"000000000",
  11301=>"000111001",
  11302=>"000111011",
  11303=>"101100111",
  11304=>"100111111",
  11305=>"010000111",
  11306=>"000101000",
  11307=>"110111111",
  11308=>"111110111",
  11309=>"100111111",
  11310=>"110000001",
  11311=>"100100000",
  11312=>"000000111",
  11313=>"011111000",
  11314=>"111101111",
  11315=>"101000000",
  11316=>"111000110",
  11317=>"111000111",
  11318=>"111111011",
  11319=>"101111111",
  11320=>"111011011",
  11321=>"000110111",
  11322=>"111000010",
  11323=>"000000000",
  11324=>"111111000",
  11325=>"001001111",
  11326=>"111100111",
  11327=>"111111111",
  11328=>"000000000",
  11329=>"110000010",
  11330=>"000110000",
  11331=>"000000111",
  11332=>"110000100",
  11333=>"001011001",
  11334=>"110000111",
  11335=>"111111111",
  11336=>"111000011",
  11337=>"111111011",
  11338=>"000000000",
  11339=>"111111101",
  11340=>"000100110",
  11341=>"011001011",
  11342=>"010110111",
  11343=>"111111110",
  11344=>"000000100",
  11345=>"110000000",
  11346=>"111000000",
  11347=>"100001111",
  11348=>"001001111",
  11349=>"011101101",
  11350=>"100100100",
  11351=>"000000000",
  11352=>"000110110",
  11353=>"000111000",
  11354=>"100100000",
  11355=>"100111101",
  11356=>"000111101",
  11357=>"000000111",
  11358=>"111110100",
  11359=>"111111111",
  11360=>"100000111",
  11361=>"000011000",
  11362=>"000111111",
  11363=>"000000000",
  11364=>"100111000",
  11365=>"111101000",
  11366=>"000100000",
  11367=>"000111110",
  11368=>"101111111",
  11369=>"000111000",
  11370=>"111110111",
  11371=>"000000000",
  11372=>"001111111",
  11373=>"000001000",
  11374=>"000110000",
  11375=>"111111110",
  11376=>"010000000",
  11377=>"010110111",
  11378=>"011010000",
  11379=>"011011011",
  11380=>"101001000",
  11381=>"111110010",
  11382=>"000000000",
  11383=>"000001101",
  11384=>"000000000",
  11385=>"100000000",
  11386=>"111101001",
  11387=>"000000000",
  11388=>"111000111",
  11389=>"111101101",
  11390=>"111001110",
  11391=>"010000000",
  11392=>"000111111",
  11393=>"000111000",
  11394=>"111010111",
  11395=>"001000110",
  11396=>"011000100",
  11397=>"000000111",
  11398=>"000000001",
  11399=>"000111010",
  11400=>"110011000",
  11401=>"111111000",
  11402=>"000000101",
  11403=>"111000000",
  11404=>"011111111",
  11405=>"111111111",
  11406=>"110000000",
  11407=>"000110000",
  11408=>"001111011",
  11409=>"000100000",
  11410=>"111111000",
  11411=>"111000001",
  11412=>"001000111",
  11413=>"101000111",
  11414=>"000000111",
  11415=>"000000110",
  11416=>"000111110",
  11417=>"011111001",
  11418=>"000001111",
  11419=>"110110111",
  11420=>"000100000",
  11421=>"111110100",
  11422=>"101101111",
  11423=>"000000101",
  11424=>"011000100",
  11425=>"111011110",
  11426=>"000011010",
  11427=>"110111111",
  11428=>"111011111",
  11429=>"010111100",
  11430=>"110111000",
  11431=>"000000010",
  11432=>"000101101",
  11433=>"000010111",
  11434=>"000111111",
  11435=>"000100111",
  11436=>"111111000",
  11437=>"111000111",
  11438=>"101001111",
  11439=>"000000000",
  11440=>"000000000",
  11441=>"011110110",
  11442=>"000000000",
  11443=>"111000000",
  11444=>"111101101",
  11445=>"000000000",
  11446=>"111000111",
  11447=>"100101000",
  11448=>"000101001",
  11449=>"110111111",
  11450=>"111111110",
  11451=>"100101111",
  11452=>"111011111",
  11453=>"000000001",
  11454=>"111000000",
  11455=>"101100111",
  11456=>"100000000",
  11457=>"001011111",
  11458=>"111101011",
  11459=>"111111111",
  11460=>"000000000",
  11461=>"111000110",
  11462=>"010011111",
  11463=>"000000111",
  11464=>"000110111",
  11465=>"110000111",
  11466=>"111000111",
  11467=>"011100100",
  11468=>"000011001",
  11469=>"111111001",
  11470=>"111111111",
  11471=>"111111111",
  11472=>"000010000",
  11473=>"011000000",
  11474=>"111011000",
  11475=>"000001000",
  11476=>"111110010",
  11477=>"000000011",
  11478=>"000011011",
  11479=>"111111111",
  11480=>"111111111",
  11481=>"111111110",
  11482=>"000111000",
  11483=>"000110111",
  11484=>"001001111",
  11485=>"000111011",
  11486=>"111000000",
  11487=>"010011000",
  11488=>"000010011",
  11489=>"111111111",
  11490=>"000000000",
  11491=>"001111111",
  11492=>"111000111",
  11493=>"000000100",
  11494=>"111001000",
  11495=>"111011111",
  11496=>"111111000",
  11497=>"011111110",
  11498=>"011011000",
  11499=>"000001111",
  11500=>"101111010",
  11501=>"000111000",
  11502=>"000011110",
  11503=>"010111000",
  11504=>"111111110",
  11505=>"111111110",
  11506=>"000000111",
  11507=>"000000000",
  11508=>"001000000",
  11509=>"110011111",
  11510=>"101000111",
  11511=>"100110100",
  11512=>"111111000",
  11513=>"001000000",
  11514=>"000111111",
  11515=>"000010111",
  11516=>"111000111",
  11517=>"111100111",
  11518=>"000000101",
  11519=>"011001111",
  11520=>"000001001",
  11521=>"111001111",
  11522=>"110111011",
  11523=>"110110111",
  11524=>"100000000",
  11525=>"110110110",
  11526=>"111111111",
  11527=>"011110100",
  11528=>"100000111",
  11529=>"111111110",
  11530=>"000001000",
  11531=>"001000110",
  11532=>"100000100",
  11533=>"111110111",
  11534=>"111000000",
  11535=>"000000000",
  11536=>"001001000",
  11537=>"000000101",
  11538=>"111111000",
  11539=>"111011010",
  11540=>"011001001",
  11541=>"000000111",
  11542=>"111000111",
  11543=>"111100111",
  11544=>"010000111",
  11545=>"111110101",
  11546=>"000000111",
  11547=>"000011000",
  11548=>"000000110",
  11549=>"000000000",
  11550=>"000000000",
  11551=>"111010010",
  11552=>"011001111",
  11553=>"000111001",
  11554=>"000001111",
  11555=>"011001111",
  11556=>"110111101",
  11557=>"010000110",
  11558=>"010000000",
  11559=>"100111000",
  11560=>"000000010",
  11561=>"111000000",
  11562=>"010111110",
  11563=>"000111000",
  11564=>"000000000",
  11565=>"001100101",
  11566=>"000000001",
  11567=>"000111000",
  11568=>"000000111",
  11569=>"011001111",
  11570=>"001000100",
  11571=>"100100000",
  11572=>"000111000",
  11573=>"111000000",
  11574=>"010011111",
  11575=>"001100000",
  11576=>"110000010",
  11577=>"000000010",
  11578=>"111111000",
  11579=>"110010000",
  11580=>"000000001",
  11581=>"011000000",
  11582=>"111001000",
  11583=>"011000100",
  11584=>"000111111",
  11585=>"100011111",
  11586=>"000000100",
  11587=>"011111011",
  11588=>"010000000",
  11589=>"000100110",
  11590=>"001001111",
  11591=>"000000000",
  11592=>"000010011",
  11593=>"111000000",
  11594=>"000111111",
  11595=>"111000100",
  11596=>"011000001",
  11597=>"000111111",
  11598=>"000111111",
  11599=>"100100110",
  11600=>"001000100",
  11601=>"111011101",
  11602=>"000110111",
  11603=>"011001011",
  11604=>"100111001",
  11605=>"011000011",
  11606=>"000110110",
  11607=>"110111100",
  11608=>"000000001",
  11609=>"111111001",
  11610=>"111000111",
  11611=>"000111000",
  11612=>"111000111",
  11613=>"111000000",
  11614=>"010000000",
  11615=>"111101111",
  11616=>"000111000",
  11617=>"111000011",
  11618=>"110000111",
  11619=>"000111000",
  11620=>"111000111",
  11621=>"011000001",
  11622=>"000111000",
  11623=>"111011111",
  11624=>"000000000",
  11625=>"111010111",
  11626=>"000000111",
  11627=>"111111000",
  11628=>"000000000",
  11629=>"111110111",
  11630=>"111000000",
  11631=>"010111111",
  11632=>"000000111",
  11633=>"111111111",
  11634=>"001011000",
  11635=>"111111110",
  11636=>"111111111",
  11637=>"111111001",
  11638=>"100100101",
  11639=>"110110111",
  11640=>"000111000",
  11641=>"000101001",
  11642=>"000011000",
  11643=>"000000001",
  11644=>"110111010",
  11645=>"100111111",
  11646=>"111111000",
  11647=>"000000000",
  11648=>"100100011",
  11649=>"001011111",
  11650=>"101100100",
  11651=>"010110110",
  11652=>"000111000",
  11653=>"010000110",
  11654=>"111111000",
  11655=>"000000100",
  11656=>"010000000",
  11657=>"000000111",
  11658=>"001001000",
  11659=>"110111110",
  11660=>"111111000",
  11661=>"100000111",
  11662=>"111101111",
  11663=>"110011000",
  11664=>"000000110",
  11665=>"011111000",
  11666=>"000000000",
  11667=>"101111001",
  11668=>"111000111",
  11669=>"001000011",
  11670=>"111111001",
  11671=>"100100110",
  11672=>"001111111",
  11673=>"111000111",
  11674=>"111111000",
  11675=>"111111110",
  11676=>"001000111",
  11677=>"010001000",
  11678=>"001000000",
  11679=>"000000000",
  11680=>"111000000",
  11681=>"101000110",
  11682=>"100100100",
  11683=>"000111101",
  11684=>"110110110",
  11685=>"100000111",
  11686=>"111111000",
  11687=>"000011011",
  11688=>"000000001",
  11689=>"000111111",
  11690=>"000000010",
  11691=>"100111111",
  11692=>"111111000",
  11693=>"111111110",
  11694=>"010111111",
  11695=>"111000111",
  11696=>"010111111",
  11697=>"000111111",
  11698=>"000110100",
  11699=>"101000011",
  11700=>"101001111",
  11701=>"001011011",
  11702=>"000000011",
  11703=>"001000000",
  11704=>"111111111",
  11705=>"111111000",
  11706=>"111111001",
  11707=>"100100111",
  11708=>"111000100",
  11709=>"111111000",
  11710=>"000011111",
  11711=>"000000000",
  11712=>"000111110",
  11713=>"000000000",
  11714=>"010000000",
  11715=>"111111111",
  11716=>"000100111",
  11717=>"000110111",
  11718=>"111001111",
  11719=>"111111111",
  11720=>"000000011",
  11721=>"000111110",
  11722=>"000100101",
  11723=>"000011000",
  11724=>"000111110",
  11725=>"000001000",
  11726=>"011111100",
  11727=>"000000000",
  11728=>"000000111",
  11729=>"100110011",
  11730=>"111001001",
  11731=>"001011001",
  11732=>"010111100",
  11733=>"010110111",
  11734=>"111110110",
  11735=>"000000001",
  11736=>"000000100",
  11737=>"001100111",
  11738=>"000000000",
  11739=>"100101000",
  11740=>"111000001",
  11741=>"011010000",
  11742=>"000001000",
  11743=>"100110110",
  11744=>"000000111",
  11745=>"100111011",
  11746=>"111010000",
  11747=>"111111010",
  11748=>"000110000",
  11749=>"111111011",
  11750=>"110111000",
  11751=>"000111000",
  11752=>"011111101",
  11753=>"000110001",
  11754=>"111010000",
  11755=>"100100111",
  11756=>"000110000",
  11757=>"001001001",
  11758=>"000000000",
  11759=>"111011000",
  11760=>"111111111",
  11761=>"111111100",
  11762=>"111000111",
  11763=>"111011000",
  11764=>"000001011",
  11765=>"001000000",
  11766=>"000011000",
  11767=>"101000011",
  11768=>"000000011",
  11769=>"000000000",
  11770=>"010000000",
  11771=>"000000000",
  11772=>"000000000",
  11773=>"100010111",
  11774=>"011000101",
  11775=>"100111111",
  11776=>"001011111",
  11777=>"110000000",
  11778=>"111111101",
  11779=>"111111111",
  11780=>"111111111",
  11781=>"111111001",
  11782=>"000000000",
  11783=>"100000000",
  11784=>"111111110",
  11785=>"111111111",
  11786=>"111001111",
  11787=>"111111110",
  11788=>"100100100",
  11789=>"000000000",
  11790=>"000100100",
  11791=>"000000110",
  11792=>"000000000",
  11793=>"111111111",
  11794=>"000000000",
  11795=>"000000000",
  11796=>"000100100",
  11797=>"111111000",
  11798=>"111110000",
  11799=>"000000001",
  11800=>"111111111",
  11801=>"111111111",
  11802=>"100100100",
  11803=>"111111111",
  11804=>"100111111",
  11805=>"111111001",
  11806=>"110000000",
  11807=>"000110111",
  11808=>"110100000",
  11809=>"110110111",
  11810=>"000000000",
  11811=>"111111000",
  11812=>"110100100",
  11813=>"011111111",
  11814=>"011011000",
  11815=>"000100000",
  11816=>"101111111",
  11817=>"000100001",
  11818=>"000000000",
  11819=>"111111000",
  11820=>"111001000",
  11821=>"000110000",
  11822=>"110111110",
  11823=>"000101111",
  11824=>"010111111",
  11825=>"010111111",
  11826=>"000001001",
  11827=>"000000000",
  11828=>"000000000",
  11829=>"111111111",
  11830=>"000000000",
  11831=>"111110110",
  11832=>"111111111",
  11833=>"001101100",
  11834=>"001001001",
  11835=>"111110111",
  11836=>"111111101",
  11837=>"111111111",
  11838=>"111110100",
  11839=>"101100100",
  11840=>"111000000",
  11841=>"111111000",
  11842=>"000111111",
  11843=>"111011111",
  11844=>"100100110",
  11845=>"000000000",
  11846=>"111101111",
  11847=>"000000000",
  11848=>"111001011",
  11849=>"111101101",
  11850=>"110110111",
  11851=>"111011000",
  11852=>"000000000",
  11853=>"000000111",
  11854=>"000000000",
  11855=>"000000000",
  11856=>"111111111",
  11857=>"000000000",
  11858=>"111110000",
  11859=>"000000110",
  11860=>"001001011",
  11861=>"000000000",
  11862=>"110100101",
  11863=>"000000000",
  11864=>"001000000",
  11865=>"101100101",
  11866=>"110001001",
  11867=>"111110110",
  11868=>"000111111",
  11869=>"000100111",
  11870=>"101111111",
  11871=>"111110110",
  11872=>"111001001",
  11873=>"111001000",
  11874=>"000000100",
  11875=>"111000000",
  11876=>"111100100",
  11877=>"111110100",
  11878=>"111111111",
  11879=>"111111111",
  11880=>"111000000",
  11881=>"111111001",
  11882=>"000000000",
  11883=>"100100000",
  11884=>"001001001",
  11885=>"111111111",
  11886=>"111111111",
  11887=>"111111011",
  11888=>"110111111",
  11889=>"111111111",
  11890=>"111111111",
  11891=>"001001001",
  11892=>"111111001",
  11893=>"111111110",
  11894=>"110111111",
  11895=>"011011000",
  11896=>"001001001",
  11897=>"000000101",
  11898=>"001000000",
  11899=>"111001001",
  11900=>"110100111",
  11901=>"000111111",
  11902=>"000000000",
  11903=>"111010000",
  11904=>"111111001",
  11905=>"001001000",
  11906=>"000000000",
  11907=>"111011111",
  11908=>"111111001",
  11909=>"111101111",
  11910=>"000000101",
  11911=>"110000000",
  11912=>"100000000",
  11913=>"110000011",
  11914=>"000010010",
  11915=>"000000100",
  11916=>"111101101",
  11917=>"000000000",
  11918=>"111101101",
  11919=>"111111111",
  11920=>"000000000",
  11921=>"001000001",
  11922=>"110100111",
  11923=>"000000011",
  11924=>"001011001",
  11925=>"111111111",
  11926=>"001000000",
  11927=>"111111111",
  11928=>"001001000",
  11929=>"000000000",
  11930=>"001000001",
  11931=>"000000110",
  11932=>"010000000",
  11933=>"100000000",
  11934=>"001000000",
  11935=>"000000000",
  11936=>"111101101",
  11937=>"110111111",
  11938=>"111110000",
  11939=>"000000000",
  11940=>"000000000",
  11941=>"110111111",
  11942=>"111111111",
  11943=>"111011011",
  11944=>"110110000",
  11945=>"000111111",
  11946=>"000000000",
  11947=>"111010000",
  11948=>"111111000",
  11949=>"100000100",
  11950=>"111111111",
  11951=>"000000111",
  11952=>"010010110",
  11953=>"111111111",
  11954=>"111111111",
  11955=>"010000111",
  11956=>"110111111",
  11957=>"000000000",
  11958=>"000000000",
  11959=>"111111011",
  11960=>"000000100",
  11961=>"100111111",
  11962=>"000001000",
  11963=>"110111111",
  11964=>"000000000",
  11965=>"111101100",
  11966=>"110010000",
  11967=>"001000000",
  11968=>"000000000",
  11969=>"111111111",
  11970=>"111000000",
  11971=>"001111111",
  11972=>"111011000",
  11973=>"000000000",
  11974=>"000000000",
  11975=>"100100100",
  11976=>"001101111",
  11977=>"000000111",
  11978=>"011111111",
  11979=>"000011011",
  11980=>"111011001",
  11981=>"100111111",
  11982=>"000000000",
  11983=>"000000000",
  11984=>"000000000",
  11985=>"111111111",
  11986=>"111000000",
  11987=>"010000010",
  11988=>"111111111",
  11989=>"110000000",
  11990=>"100000001",
  11991=>"000000101",
  11992=>"000000000",
  11993=>"000110110",
  11994=>"000000000",
  11995=>"110110110",
  11996=>"100000001",
  11997=>"110111111",
  11998=>"111011000",
  11999=>"000000001",
  12000=>"111111111",
  12001=>"100111011",
  12002=>"100000001",
  12003=>"111010000",
  12004=>"000000000",
  12005=>"011111111",
  12006=>"000100100",
  12007=>"000000000",
  12008=>"000000010",
  12009=>"000000010",
  12010=>"111111110",
  12011=>"100100000",
  12012=>"000000000",
  12013=>"111100000",
  12014=>"110001001",
  12015=>"111111111",
  12016=>"111100001",
  12017=>"000000000",
  12018=>"011011111",
  12019=>"000000000",
  12020=>"100000111",
  12021=>"110000010",
  12022=>"111111100",
  12023=>"110111111",
  12024=>"111111110",
  12025=>"111111111",
  12026=>"000111111",
  12027=>"111111100",
  12028=>"000100110",
  12029=>"001000000",
  12030=>"110110110",
  12031=>"000000001",
  12032=>"000100100",
  12033=>"110110111",
  12034=>"000000000",
  12035=>"011001000",
  12036=>"000000000",
  12037=>"111111111",
  12038=>"100000101",
  12039=>"000000000",
  12040=>"000000100",
  12041=>"011111001",
  12042=>"000000000",
  12043=>"111111100",
  12044=>"001001001",
  12045=>"100000000",
  12046=>"000111111",
  12047=>"011001001",
  12048=>"000100100",
  12049=>"000000000",
  12050=>"000000000",
  12051=>"100000000",
  12052=>"000100110",
  12053=>"111101111",
  12054=>"001000001",
  12055=>"000000000",
  12056=>"010010010",
  12057=>"010000000",
  12058=>"111111111",
  12059=>"010000000",
  12060=>"111110100",
  12061=>"111101111",
  12062=>"000111000",
  12063=>"100000001",
  12064=>"000000000",
  12065=>"111111111",
  12066=>"111111111",
  12067=>"100000111",
  12068=>"111000100",
  12069=>"000110101",
  12070=>"011011011",
  12071=>"111111111",
  12072=>"111111111",
  12073=>"110000000",
  12074=>"110000010",
  12075=>"000000111",
  12076=>"011011111",
  12077=>"111111100",
  12078=>"000010110",
  12079=>"000000000",
  12080=>"111111111",
  12081=>"000000000",
  12082=>"000000001",
  12083=>"000000000",
  12084=>"110000000",
  12085=>"000110111",
  12086=>"100000000",
  12087=>"110111111",
  12088=>"000000000",
  12089=>"111001011",
  12090=>"000000010",
  12091=>"111111110",
  12092=>"000000000",
  12093=>"000000000",
  12094=>"001011000",
  12095=>"111011011",
  12096=>"111101000",
  12097=>"111111111",
  12098=>"000000000",
  12099=>"000000000",
  12100=>"000011101",
  12101=>"010000000",
  12102=>"000000011",
  12103=>"001001101",
  12104=>"010111010",
  12105=>"111000000",
  12106=>"000000000",
  12107=>"000000000",
  12108=>"111001011",
  12109=>"111111111",
  12110=>"001000000",
  12111=>"110111111",
  12112=>"111111110",
  12113=>"000000000",
  12114=>"000111011",
  12115=>"000000000",
  12116=>"000001011",
  12117=>"001011001",
  12118=>"010000010",
  12119=>"001000000",
  12120=>"000001111",
  12121=>"000000110",
  12122=>"001111111",
  12123=>"111100100",
  12124=>"000000000",
  12125=>"001000010",
  12126=>"111111111",
  12127=>"011011111",
  12128=>"110000000",
  12129=>"111111101",
  12130=>"111111110",
  12131=>"110100100",
  12132=>"000000000",
  12133=>"000000000",
  12134=>"111100000",
  12135=>"111111000",
  12136=>"000000000",
  12137=>"000000000",
  12138=>"100111111",
  12139=>"111100110",
  12140=>"110110000",
  12141=>"000000000",
  12142=>"000010000",
  12143=>"011111111",
  12144=>"000000000",
  12145=>"000000000",
  12146=>"000000010",
  12147=>"111111111",
  12148=>"110111010",
  12149=>"001001101",
  12150=>"000111111",
  12151=>"010111111",
  12152=>"100001011",
  12153=>"010000000",
  12154=>"111001001",
  12155=>"011011001",
  12156=>"010000000",
  12157=>"110000111",
  12158=>"111111001",
  12159=>"111011111",
  12160=>"111111011",
  12161=>"011111111",
  12162=>"000000000",
  12163=>"000000000",
  12164=>"111111111",
  12165=>"000000000",
  12166=>"100100000",
  12167=>"000000000",
  12168=>"000000000",
  12169=>"000000000",
  12170=>"111111111",
  12171=>"000000000",
  12172=>"101111111",
  12173=>"000000001",
  12174=>"010000100",
  12175=>"111111111",
  12176=>"000000000",
  12177=>"000000000",
  12178=>"000000100",
  12179=>"000000000",
  12180=>"011111000",
  12181=>"000010000",
  12182=>"111111111",
  12183=>"101111001",
  12184=>"111111011",
  12185=>"110100110",
  12186=>"000100000",
  12187=>"111000000",
  12188=>"000111111",
  12189=>"110000000",
  12190=>"001011011",
  12191=>"011011111",
  12192=>"000111111",
  12193=>"000101101",
  12194=>"100000100",
  12195=>"000000111",
  12196=>"000000100",
  12197=>"111111111",
  12198=>"111111111",
  12199=>"000000001",
  12200=>"010010000",
  12201=>"000000000",
  12202=>"000000111",
  12203=>"000000001",
  12204=>"000000000",
  12205=>"100001001",
  12206=>"100111111",
  12207=>"000000000",
  12208=>"100111110",
  12209=>"000000000",
  12210=>"111111000",
  12211=>"110100111",
  12212=>"111100100",
  12213=>"111110000",
  12214=>"011010100",
  12215=>"111111111",
  12216=>"111110000",
  12217=>"000000110",
  12218=>"000000000",
  12219=>"111111111",
  12220=>"101100000",
  12221=>"110000011",
  12222=>"000000111",
  12223=>"000000100",
  12224=>"111011111",
  12225=>"111111111",
  12226=>"100100101",
  12227=>"000000000",
  12228=>"111011000",
  12229=>"111111010",
  12230=>"110100100",
  12231=>"000000111",
  12232=>"000000000",
  12233=>"111111111",
  12234=>"111111111",
  12235=>"011000000",
  12236=>"000001001",
  12237=>"111000111",
  12238=>"000000000",
  12239=>"110111111",
  12240=>"000000000",
  12241=>"111111111",
  12242=>"000000000",
  12243=>"100000000",
  12244=>"111111111",
  12245=>"000000000",
  12246=>"111001111",
  12247=>"001011011",
  12248=>"111111111",
  12249=>"000010011",
  12250=>"111111111",
  12251=>"111111111",
  12252=>"010111111",
  12253=>"100001111",
  12254=>"000000100",
  12255=>"011011111",
  12256=>"010000000",
  12257=>"000000000",
  12258=>"000001100",
  12259=>"101111111",
  12260=>"000000000",
  12261=>"111111111",
  12262=>"000000101",
  12263=>"000110110",
  12264=>"000000000",
  12265=>"000000100",
  12266=>"100100010",
  12267=>"111110110",
  12268=>"000000000",
  12269=>"110010000",
  12270=>"000000100",
  12271=>"101000000",
  12272=>"000011001",
  12273=>"000000000",
  12274=>"111000111",
  12275=>"000000000",
  12276=>"110110000",
  12277=>"011001011",
  12278=>"111010000",
  12279=>"000000000",
  12280=>"000000100",
  12281=>"001001001",
  12282=>"111000010",
  12283=>"110001101",
  12284=>"100100000",
  12285=>"000000000",
  12286=>"101111111",
  12287=>"111111111",
  12288=>"111101100",
  12289=>"000000011",
  12290=>"000101101",
  12291=>"000010000",
  12292=>"000000111",
  12293=>"000000000",
  12294=>"111110110",
  12295=>"000000000",
  12296=>"000000111",
  12297=>"000001000",
  12298=>"000000000",
  12299=>"111111110",
  12300=>"001011000",
  12301=>"001000101",
  12302=>"100000011",
  12303=>"000000000",
  12304=>"000111111",
  12305=>"011111000",
  12306=>"000111111",
  12307=>"000000001",
  12308=>"000000000",
  12309=>"111111000",
  12310=>"000000000",
  12311=>"100000111",
  12312=>"111111000",
  12313=>"111111110",
  12314=>"111111110",
  12315=>"011110111",
  12316=>"111111110",
  12317=>"100111111",
  12318=>"001000001",
  12319=>"100100000",
  12320=>"000000000",
  12321=>"111110000",
  12322=>"111111110",
  12323=>"111000000",
  12324=>"001111111",
  12325=>"111101111",
  12326=>"000000000",
  12327=>"111010100",
  12328=>"000000000",
  12329=>"111111001",
  12330=>"100111111",
  12331=>"111001000",
  12332=>"111100001",
  12333=>"000001000",
  12334=>"000000000",
  12335=>"110101000",
  12336=>"111000110",
  12337=>"000111111",
  12338=>"000000000",
  12339=>"000000010",
  12340=>"001001101",
  12341=>"000011111",
  12342=>"001000000",
  12343=>"111100000",
  12344=>"000000111",
  12345=>"100101000",
  12346=>"100100111",
  12347=>"011111101",
  12348=>"001000100",
  12349=>"111111000",
  12350=>"010111111",
  12351=>"111111111",
  12352=>"111101111",
  12353=>"111111000",
  12354=>"111111000",
  12355=>"111000000",
  12356=>"011011011",
  12357=>"000000000",
  12358=>"001000000",
  12359=>"111111000",
  12360=>"111101100",
  12361=>"111000000",
  12362=>"111111111",
  12363=>"111111111",
  12364=>"111111111",
  12365=>"000111111",
  12366=>"000100001",
  12367=>"000000100",
  12368=>"111110000",
  12369=>"111111111",
  12370=>"111110000",
  12371=>"000000111",
  12372=>"111111111",
  12373=>"110000000",
  12374=>"111000000",
  12375=>"000000100",
  12376=>"001000111",
  12377=>"111000100",
  12378=>"000011111",
  12379=>"111110110",
  12380=>"000001011",
  12381=>"001000111",
  12382=>"111111000",
  12383=>"000000000",
  12384=>"000111111",
  12385=>"111010000",
  12386=>"001000000",
  12387=>"001001111",
  12388=>"001011100",
  12389=>"111110000",
  12390=>"111111111",
  12391=>"111111011",
  12392=>"000000000",
  12393=>"111111111",
  12394=>"000000000",
  12395=>"000110000",
  12396=>"000000111",
  12397=>"000001111",
  12398=>"000111111",
  12399=>"000000000",
  12400=>"001111000",
  12401=>"000000011",
  12402=>"000001001",
  12403=>"111111000",
  12404=>"000000011",
  12405=>"000111111",
  12406=>"000011111",
  12407=>"000100111",
  12408=>"000000000",
  12409=>"111111000",
  12410=>"000111111",
  12411=>"000000000",
  12412=>"110110100",
  12413=>"111111011",
  12414=>"010111111",
  12415=>"111011111",
  12416=>"000000100",
  12417=>"000111111",
  12418=>"111000000",
  12419=>"000111111",
  12420=>"000000110",
  12421=>"000010010",
  12422=>"111100000",
  12423=>"011001000",
  12424=>"000000111",
  12425=>"111111000",
  12426=>"000111011",
  12427=>"000000110",
  12428=>"111111100",
  12429=>"111111001",
  12430=>"100011011",
  12431=>"111000111",
  12432=>"000000111",
  12433=>"000000001",
  12434=>"000000100",
  12435=>"111111111",
  12436=>"100100000",
  12437=>"101000100",
  12438=>"000000111",
  12439=>"111111101",
  12440=>"000000101",
  12441=>"000000111",
  12442=>"011000100",
  12443=>"000000000",
  12444=>"111111110",
  12445=>"000001111",
  12446=>"000100111",
  12447=>"000110110",
  12448=>"000001101",
  12449=>"011001000",
  12450=>"111000101",
  12451=>"000100111",
  12452=>"000111111",
  12453=>"111001001",
  12454=>"100000000",
  12455=>"000011001",
  12456=>"111110010",
  12457=>"011000000",
  12458=>"000000000",
  12459=>"000000100",
  12460=>"010111011",
  12461=>"110000000",
  12462=>"111111000",
  12463=>"111111111",
  12464=>"111111000",
  12465=>"110110100",
  12466=>"111111111",
  12467=>"011000110",
  12468=>"000000101",
  12469=>"101111111",
  12470=>"000000000",
  12471=>"000000110",
  12472=>"100100111",
  12473=>"111111111",
  12474=>"000111110",
  12475=>"111000000",
  12476=>"001011000",
  12477=>"101100111",
  12478=>"000111111",
  12479=>"111111000",
  12480=>"011000000",
  12481=>"011010111",
  12482=>"111111110",
  12483=>"000000111",
  12484=>"111000000",
  12485=>"000000000",
  12486=>"001000000",
  12487=>"000001110",
  12488=>"010111111",
  12489=>"111000000",
  12490=>"000000000",
  12491=>"000000111",
  12492=>"101000000",
  12493=>"000011000",
  12494=>"111001111",
  12495=>"000111111",
  12496=>"111111000",
  12497=>"111111111",
  12498=>"111111111",
  12499=>"011111011",
  12500=>"111111000",
  12501=>"000100110",
  12502=>"111111000",
  12503=>"000000000",
  12504=>"000000000",
  12505=>"001000000",
  12506=>"000100000",
  12507=>"111111000",
  12508=>"001000000",
  12509=>"000000100",
  12510=>"000000100",
  12511=>"100000001",
  12512=>"000111000",
  12513=>"000000000",
  12514=>"000000000",
  12515=>"100001111",
  12516=>"000111111",
  12517=>"111111111",
  12518=>"000010111",
  12519=>"111111100",
  12520=>"000000111",
  12521=>"111110111",
  12522=>"101101111",
  12523=>"001001111",
  12524=>"000000101",
  12525=>"000000000",
  12526=>"000000111",
  12527=>"111111000",
  12528=>"111111000",
  12529=>"000000111",
  12530=>"111111111",
  12531=>"001001001",
  12532=>"000000000",
  12533=>"000000000",
  12534=>"000000011",
  12535=>"011101111",
  12536=>"000000111",
  12537=>"111100000",
  12538=>"111001111",
  12539=>"100000000",
  12540=>"000000000",
  12541=>"111110100",
  12542=>"010001111",
  12543=>"111111100",
  12544=>"111111000",
  12545=>"000100101",
  12546=>"000000111",
  12547=>"110000000",
  12548=>"011011111",
  12549=>"110101100",
  12550=>"000000111",
  12551=>"011000001",
  12552=>"001011111",
  12553=>"000000010",
  12554=>"111111111",
  12555=>"000110111",
  12556=>"111000101",
  12557=>"000011000",
  12558=>"000000000",
  12559=>"111111111",
  12560=>"000000111",
  12561=>"001001000",
  12562=>"111000000",
  12563=>"000000000",
  12564=>"111010000",
  12565=>"000000100",
  12566=>"110100111",
  12567=>"111000000",
  12568=>"000111101",
  12569=>"111000000",
  12570=>"000000101",
  12571=>"111000111",
  12572=>"001001001",
  12573=>"000011111",
  12574=>"010000000",
  12575=>"001000111",
  12576=>"000011110",
  12577=>"001000000",
  12578=>"000000101",
  12579=>"101000000",
  12580=>"111000000",
  12581=>"111111111",
  12582=>"111100100",
  12583=>"000000000",
  12584=>"111111111",
  12585=>"111111000",
  12586=>"111111101",
  12587=>"000111111",
  12588=>"111111010",
  12589=>"000000111",
  12590=>"000011111",
  12591=>"000000000",
  12592=>"000100000",
  12593=>"000000010",
  12594=>"000000000",
  12595=>"000000001",
  12596=>"001000000",
  12597=>"010111101",
  12598=>"000000011",
  12599=>"000110110",
  12600=>"000000111",
  12601=>"111000101",
  12602=>"110000000",
  12603=>"100000000",
  12604=>"000000000",
  12605=>"000000101",
  12606=>"010000000",
  12607=>"000000000",
  12608=>"000000111",
  12609=>"000011000",
  12610=>"110111000",
  12611=>"001111111",
  12612=>"111000100",
  12613=>"000111111",
  12614=>"000100110",
  12615=>"000000111",
  12616=>"001000001",
  12617=>"111000000",
  12618=>"000000100",
  12619=>"011011001",
  12620=>"000100110",
  12621=>"000000000",
  12622=>"000000000",
  12623=>"000000000",
  12624=>"000000111",
  12625=>"001000100",
  12626=>"111011111",
  12627=>"000000111",
  12628=>"001111111",
  12629=>"011011001",
  12630=>"111001000",
  12631=>"111111111",
  12632=>"111111100",
  12633=>"111110111",
  12634=>"111010000",
  12635=>"111111110",
  12636=>"111000000",
  12637=>"001011011",
  12638=>"000000111",
  12639=>"111000000",
  12640=>"111110001",
  12641=>"111111111",
  12642=>"100100100",
  12643=>"111111000",
  12644=>"000011111",
  12645=>"101100111",
  12646=>"000000001",
  12647=>"111000000",
  12648=>"110000000",
  12649=>"000000111",
  12650=>"000001111",
  12651=>"111111110",
  12652=>"000000010",
  12653=>"000111111",
  12654=>"000000000",
  12655=>"001000000",
  12656=>"111111011",
  12657=>"101011111",
  12658=>"000000100",
  12659=>"011011011",
  12660=>"000111111",
  12661=>"011010111",
  12662=>"111001111",
  12663=>"000101111",
  12664=>"111111111",
  12665=>"000111111",
  12666=>"000000000",
  12667=>"000001000",
  12668=>"000000100",
  12669=>"000010111",
  12670=>"000000000",
  12671=>"111111111",
  12672=>"100100100",
  12673=>"000000000",
  12674=>"100000000",
  12675=>"111100000",
  12676=>"000000011",
  12677=>"000111111",
  12678=>"110010000",
  12679=>"001000000",
  12680=>"111000000",
  12681=>"111111001",
  12682=>"111111111",
  12683=>"111111000",
  12684=>"101000111",
  12685=>"001011111",
  12686=>"001000110",
  12687=>"011111111",
  12688=>"000001000",
  12689=>"111111110",
  12690=>"111111111",
  12691=>"000000001",
  12692=>"000111111",
  12693=>"000000010",
  12694=>"111010100",
  12695=>"111111000",
  12696=>"000000011",
  12697=>"000100111",
  12698=>"110000111",
  12699=>"011111111",
  12700=>"111111111",
  12701=>"000000000",
  12702=>"000000111",
  12703=>"000000111",
  12704=>"000011111",
  12705=>"000000101",
  12706=>"001000001",
  12707=>"000000011",
  12708=>"001001101",
  12709=>"000100111",
  12710=>"000111111",
  12711=>"000000011",
  12712=>"000000000",
  12713=>"100110111",
  12714=>"111101000",
  12715=>"111111101",
  12716=>"000000000",
  12717=>"000000001",
  12718=>"000000011",
  12719=>"111000000",
  12720=>"111111000",
  12721=>"000000000",
  12722=>"101100101",
  12723=>"000000000",
  12724=>"111111111",
  12725=>"111000111",
  12726=>"111000001",
  12727=>"000001111",
  12728=>"111111100",
  12729=>"111110110",
  12730=>"010000001",
  12731=>"111111111",
  12732=>"000000000",
  12733=>"000000000",
  12734=>"101001111",
  12735=>"110110100",
  12736=>"001001111",
  12737=>"111100101",
  12738=>"111101111",
  12739=>"010010100",
  12740=>"111111000",
  12741=>"111000000",
  12742=>"111111000",
  12743=>"000111011",
  12744=>"000000001",
  12745=>"100111000",
  12746=>"100000000",
  12747=>"111101100",
  12748=>"000000111",
  12749=>"000000000",
  12750=>"100000000",
  12751=>"110111000",
  12752=>"000011001",
  12753=>"111111011",
  12754=>"000111111",
  12755=>"111111111",
  12756=>"000000000",
  12757=>"110110000",
  12758=>"000110000",
  12759=>"100100000",
  12760=>"100100100",
  12761=>"001111111",
  12762=>"001111100",
  12763=>"000000101",
  12764=>"001111111",
  12765=>"001000101",
  12766=>"101000000",
  12767=>"110000001",
  12768=>"011001000",
  12769=>"000010010",
  12770=>"111111111",
  12771=>"001001000",
  12772=>"111000000",
  12773=>"100111111",
  12774=>"000000000",
  12775=>"000000000",
  12776=>"111101000",
  12777=>"111000000",
  12778=>"111001001",
  12779=>"111111000",
  12780=>"001111111",
  12781=>"011011000",
  12782=>"000000000",
  12783=>"111111111",
  12784=>"111011000",
  12785=>"111111111",
  12786=>"001000001",
  12787=>"000000111",
  12788=>"111111010",
  12789=>"000011111",
  12790=>"000000100",
  12791=>"000000000",
  12792=>"111111000",
  12793=>"110010000",
  12794=>"000000100",
  12795=>"111101111",
  12796=>"000011111",
  12797=>"001000100",
  12798=>"000000000",
  12799=>"000000111",
  12800=>"111000001",
  12801=>"101000000",
  12802=>"111111111",
  12803=>"000111111",
  12804=>"111000000",
  12805=>"000110000",
  12806=>"000000000",
  12807=>"101100111",
  12808=>"011010000",
  12809=>"000000100",
  12810=>"101000000",
  12811=>"000000000",
  12812=>"111111111",
  12813=>"000000000",
  12814=>"000100101",
  12815=>"111111111",
  12816=>"010010010",
  12817=>"111000000",
  12818=>"000000000",
  12819=>"011001000",
  12820=>"000000000",
  12821=>"000000000",
  12822=>"111111111",
  12823=>"001000001",
  12824=>"000000000",
  12825=>"110101001",
  12826=>"111110100",
  12827=>"110010000",
  12828=>"111111111",
  12829=>"111100111",
  12830=>"111011000",
  12831=>"111111111",
  12832=>"111111111",
  12833=>"111111110",
  12834=>"000110110",
  12835=>"000000000",
  12836=>"111111111",
  12837=>"000101101",
  12838=>"000000000",
  12839=>"000000000",
  12840=>"000000000",
  12841=>"111111111",
  12842=>"001000001",
  12843=>"111111111",
  12844=>"010110111",
  12845=>"011000000",
  12846=>"001000111",
  12847=>"101000100",
  12848=>"000000000",
  12849=>"111111111",
  12850=>"001001000",
  12851=>"100000101",
  12852=>"111111111",
  12853=>"001001111",
  12854=>"101000000",
  12855=>"110110000",
  12856=>"111011011",
  12857=>"000000000",
  12858=>"111100101",
  12859=>"000000000",
  12860=>"101000000",
  12861=>"111111011",
  12862=>"111111011",
  12863=>"000100000",
  12864=>"100000111",
  12865=>"000000101",
  12866=>"111111110",
  12867=>"000001000",
  12868=>"111100111",
  12869=>"111011011",
  12870=>"000001000",
  12871=>"111111111",
  12872=>"011000000",
  12873=>"000000000",
  12874=>"111111111",
  12875=>"000000000",
  12876=>"001111111",
  12877=>"000000111",
  12878=>"000110110",
  12879=>"010111111",
  12880=>"000000000",
  12881=>"000001101",
  12882=>"101000000",
  12883=>"000000000",
  12884=>"111111011",
  12885=>"000000000",
  12886=>"000000000",
  12887=>"110000000",
  12888=>"111111111",
  12889=>"111101111",
  12890=>"000000110",
  12891=>"110010000",
  12892=>"000110110",
  12893=>"011011011",
  12894=>"111000000",
  12895=>"000000001",
  12896=>"100110110",
  12897=>"000000000",
  12898=>"111111111",
  12899=>"111111111",
  12900=>"000000001",
  12901=>"001000110",
  12902=>"000001111",
  12903=>"001001101",
  12904=>"111111111",
  12905=>"000110111",
  12906=>"111111110",
  12907=>"111111111",
  12908=>"111110001",
  12909=>"111111111",
  12910=>"011111111",
  12911=>"111111111",
  12912=>"000000000",
  12913=>"010010000",
  12914=>"110100111",
  12915=>"111000010",
  12916=>"000000000",
  12917=>"111111111",
  12918=>"111111001",
  12919=>"111101000",
  12920=>"011011100",
  12921=>"101000000",
  12922=>"000000000",
  12923=>"111111111",
  12924=>"000100001",
  12925=>"000110110",
  12926=>"000000111",
  12927=>"111100100",
  12928=>"111111100",
  12929=>"111000000",
  12930=>"000000111",
  12931=>"110111011",
  12932=>"000000000",
  12933=>"010000000",
  12934=>"000000000",
  12935=>"000000000",
  12936=>"000000011",
  12937=>"000000111",
  12938=>"000000111",
  12939=>"000101111",
  12940=>"101000000",
  12941=>"000000111",
  12942=>"110000000",
  12943=>"111111111",
  12944=>"100100000",
  12945=>"000001000",
  12946=>"000111011",
  12947=>"111110000",
  12948=>"000000111",
  12949=>"000100111",
  12950=>"000000000",
  12951=>"000000000",
  12952=>"000000111",
  12953=>"111111111",
  12954=>"111111111",
  12955=>"000100000",
  12956=>"111000100",
  12957=>"101000000",
  12958=>"111111111",
  12959=>"100000000",
  12960=>"000011111",
  12961=>"101010000",
  12962=>"111111111",
  12963=>"110111111",
  12964=>"000000100",
  12965=>"111111111",
  12966=>"000000000",
  12967=>"111110111",
  12968=>"000111011",
  12969=>"000000010",
  12970=>"111111111",
  12971=>"011111111",
  12972=>"100110110",
  12973=>"000000001",
  12974=>"000000111",
  12975=>"000000100",
  12976=>"111111111",
  12977=>"111111111",
  12978=>"011011011",
  12979=>"111000000",
  12980=>"111101101",
  12981=>"000010000",
  12982=>"000000100",
  12983=>"000000001",
  12984=>"101000000",
  12985=>"000111000",
  12986=>"000000000",
  12987=>"000111111",
  12988=>"111111111",
  12989=>"111101010",
  12990=>"111111111",
  12991=>"000000000",
  12992=>"111101111",
  12993=>"111001001",
  12994=>"111111100",
  12995=>"001000000",
  12996=>"011000000",
  12997=>"000000000",
  12998=>"001111111",
  12999=>"011011001",
  13000=>"100100000",
  13001=>"110110110",
  13002=>"100110000",
  13003=>"000000000",
  13004=>"000000100",
  13005=>"111111111",
  13006=>"111000000",
  13007=>"000000000",
  13008=>"111111111",
  13009=>"111000100",
  13010=>"101100111",
  13011=>"100000000",
  13012=>"001000001",
  13013=>"100000000",
  13014=>"000000000",
  13015=>"100001001",
  13016=>"111011000",
  13017=>"000000100",
  13018=>"111110000",
  13019=>"111111111",
  13020=>"000000001",
  13021=>"000000110",
  13022=>"011011111",
  13023=>"111111000",
  13024=>"000000000",
  13025=>"100100111",
  13026=>"000000111",
  13027=>"111111010",
  13028=>"110000001",
  13029=>"011001000",
  13030=>"110010000",
  13031=>"000000000",
  13032=>"001000011",
  13033=>"111111110",
  13034=>"111111111",
  13035=>"111011000",
  13036=>"101000101",
  13037=>"011000110",
  13038=>"000001011",
  13039=>"000000000",
  13040=>"101000000",
  13041=>"000000100",
  13042=>"000000000",
  13043=>"000110111",
  13044=>"111111111",
  13045=>"100000000",
  13046=>"001011111",
  13047=>"111111111",
  13048=>"011111111",
  13049=>"111101101",
  13050=>"111111111",
  13051=>"000000111",
  13052=>"111100000",
  13053=>"000000000",
  13054=>"100001111",
  13055=>"101001111",
  13056=>"101101111",
  13057=>"010011011",
  13058=>"000000000",
  13059=>"000000000",
  13060=>"111111111",
  13061=>"000111111",
  13062=>"111111111",
  13063=>"100000101",
  13064=>"111111111",
  13065=>"110110110",
  13066=>"000010000",
  13067=>"111100000",
  13068=>"111111011",
  13069=>"000001111",
  13070=>"000010110",
  13071=>"001000011",
  13072=>"000000011",
  13073=>"111111111",
  13074=>"000000111",
  13075=>"110111111",
  13076=>"110000000",
  13077=>"111111111",
  13078=>"111111011",
  13079=>"110000000",
  13080=>"111011001",
  13081=>"111111000",
  13082=>"001111111",
  13083=>"111010010",
  13084=>"000000000",
  13085=>"111111111",
  13086=>"000000000",
  13087=>"000110111",
  13088=>"011010100",
  13089=>"011111000",
  13090=>"110100100",
  13091=>"111111110",
  13092=>"110111110",
  13093=>"000000000",
  13094=>"000010010",
  13095=>"110110110",
  13096=>"000100100",
  13097=>"111111101",
  13098=>"010010000",
  13099=>"000111111",
  13100=>"011011001",
  13101=>"110110110",
  13102=>"000000000",
  13103=>"000000000",
  13104=>"010011011",
  13105=>"111011001",
  13106=>"000111000",
  13107=>"111111111",
  13108=>"011111010",
  13109=>"111111111",
  13110=>"000000000",
  13111=>"001000000",
  13112=>"010111110",
  13113=>"000000101",
  13114=>"000000000",
  13115=>"011011110",
  13116=>"110000001",
  13117=>"001111100",
  13118=>"111111111",
  13119=>"101100100",
  13120=>"000111110",
  13121=>"000000001",
  13122=>"111111100",
  13123=>"001000000",
  13124=>"000000001",
  13125=>"000000100",
  13126=>"111000000",
  13127=>"000000000",
  13128=>"000000000",
  13129=>"000100000",
  13130=>"001100100",
  13131=>"111111100",
  13132=>"000010110",
  13133=>"100111111",
  13134=>"111111100",
  13135=>"111100100",
  13136=>"111101111",
  13137=>"000000111",
  13138=>"110000000",
  13139=>"001000011",
  13140=>"000000000",
  13141=>"001001001",
  13142=>"111111010",
  13143=>"000101111",
  13144=>"111111000",
  13145=>"010010000",
  13146=>"000000000",
  13147=>"000000000",
  13148=>"000000101",
  13149=>"111111111",
  13150=>"111111100",
  13151=>"000100111",
  13152=>"001001111",
  13153=>"001001111",
  13154=>"100100100",
  13155=>"000000000",
  13156=>"111111100",
  13157=>"000000000",
  13158=>"001001001",
  13159=>"000000000",
  13160=>"110000000",
  13161=>"111111111",
  13162=>"111010111",
  13163=>"000001111",
  13164=>"111100001",
  13165=>"001000000",
  13166=>"111111111",
  13167=>"000000001",
  13168=>"110111111",
  13169=>"111111111",
  13170=>"011111111",
  13171=>"111110110",
  13172=>"111111111",
  13173=>"001000001",
  13174=>"011000000",
  13175=>"100111111",
  13176=>"111100001",
  13177=>"000111111",
  13178=>"000111111",
  13179=>"101111111",
  13180=>"001010000",
  13181=>"111111111",
  13182=>"001000101",
  13183=>"111111111",
  13184=>"111001001",
  13185=>"000000000",
  13186=>"111110110",
  13187=>"100000001",
  13188=>"111110110",
  13189=>"000000001",
  13190=>"111111111",
  13191=>"000000000",
  13192=>"000111111",
  13193=>"000111111",
  13194=>"000000000",
  13195=>"000010000",
  13196=>"000111111",
  13197=>"000000100",
  13198=>"101011000",
  13199=>"000000000",
  13200=>"000000000",
  13201=>"000000001",
  13202=>"110111111",
  13203=>"111100110",
  13204=>"000000000",
  13205=>"111111111",
  13206=>"100000011",
  13207=>"010110010",
  13208=>"111111100",
  13209=>"000000111",
  13210=>"000000111",
  13211=>"111111101",
  13212=>"000000001",
  13213=>"111110111",
  13214=>"000000111",
  13215=>"001111111",
  13216=>"011001011",
  13217=>"011011111",
  13218=>"011000000",
  13219=>"110111111",
  13220=>"000000000",
  13221=>"010000000",
  13222=>"000001010",
  13223=>"000000111",
  13224=>"000000000",
  13225=>"000100100",
  13226=>"100110110",
  13227=>"000111011",
  13228=>"000000000",
  13229=>"000001111",
  13230=>"000000110",
  13231=>"111111111",
  13232=>"111110111",
  13233=>"111111000",
  13234=>"110110010",
  13235=>"000001111",
  13236=>"011010111",
  13237=>"110000000",
  13238=>"111111111",
  13239=>"000000000",
  13240=>"100111100",
  13241=>"000100000",
  13242=>"111001111",
  13243=>"111111111",
  13244=>"000000010",
  13245=>"000011111",
  13246=>"000010110",
  13247=>"000011011",
  13248=>"110000011",
  13249=>"111111111",
  13250=>"000000000",
  13251=>"111111010",
  13252=>"111110010",
  13253=>"000000100",
  13254=>"010010010",
  13255=>"000101111",
  13256=>"000000101",
  13257=>"111111111",
  13258=>"100100000",
  13259=>"000110000",
  13260=>"111111000",
  13261=>"111111111",
  13262=>"000100110",
  13263=>"111110100",
  13264=>"100000000",
  13265=>"000100101",
  13266=>"111111111",
  13267=>"011011011",
  13268=>"000011111",
  13269=>"000001000",
  13270=>"011111111",
  13271=>"111101101",
  13272=>"100000000",
  13273=>"000001111",
  13274=>"101101111",
  13275=>"001101111",
  13276=>"001000000",
  13277=>"000000111",
  13278=>"011111001",
  13279=>"111101001",
  13280=>"111011000",
  13281=>"111000000",
  13282=>"001111111",
  13283=>"000000011",
  13284=>"000001001",
  13285=>"111101111",
  13286=>"000000010",
  13287=>"001000101",
  13288=>"101000100",
  13289=>"111110000",
  13290=>"111000000",
  13291=>"000000100",
  13292=>"001000000",
  13293=>"110100100",
  13294=>"011111111",
  13295=>"000000100",
  13296=>"000000000",
  13297=>"000111111",
  13298=>"000000000",
  13299=>"110010011",
  13300=>"000111111",
  13301=>"000000101",
  13302=>"111111101",
  13303=>"001110110",
  13304=>"000000000",
  13305=>"111100100",
  13306=>"111000000",
  13307=>"110111000",
  13308=>"111000000",
  13309=>"000000101",
  13310=>"000011011",
  13311=>"000000001",
  13312=>"110110111",
  13313=>"111001000",
  13314=>"101000101",
  13315=>"011111111",
  13316=>"001001001",
  13317=>"111100100",
  13318=>"111000000",
  13319=>"000000101",
  13320=>"000000111",
  13321=>"110101001",
  13322=>"111111101",
  13323=>"000101101",
  13324=>"110111111",
  13325=>"000000011",
  13326=>"110001000",
  13327=>"111111100",
  13328=>"111001001",
  13329=>"011000000",
  13330=>"101000011",
  13331=>"011000000",
  13332=>"111010000",
  13333=>"000001111",
  13334=>"110111110",
  13335=>"011000000",
  13336=>"001001111",
  13337=>"000000000",
  13338=>"110000000",
  13339=>"101100100",
  13340=>"000111111",
  13341=>"111111000",
  13342=>"111110110",
  13343=>"000000111",
  13344=>"000000000",
  13345=>"111111010",
  13346=>"011011111",
  13347=>"111110000",
  13348=>"101001100",
  13349=>"111000000",
  13350=>"111100001",
  13351=>"000010000",
  13352=>"000001000",
  13353=>"000000000",
  13354=>"111011000",
  13355=>"100000000",
  13356=>"000111101",
  13357=>"101111100",
  13358=>"011011111",
  13359=>"000000011",
  13360=>"111111110",
  13361=>"000000111",
  13362=>"110000000",
  13363=>"111000000",
  13364=>"111111000",
  13365=>"011011111",
  13366=>"111111100",
  13367=>"101100110",
  13368=>"000001111",
  13369=>"110010000",
  13370=>"111000000",
  13371=>"000000000",
  13372=>"010111111",
  13373=>"111000000",
  13374=>"000000001",
  13375=>"111110111",
  13376=>"111110000",
  13377=>"111111001",
  13378=>"000001010",
  13379=>"110111000",
  13380=>"111000000",
  13381=>"110110110",
  13382=>"111111101",
  13383=>"000100000",
  13384=>"111010011",
  13385=>"000000001",
  13386=>"111111101",
  13387=>"000111111",
  13388=>"111110111",
  13389=>"111111000",
  13390=>"111000000",
  13391=>"010000101",
  13392=>"111000000",
  13393=>"000111100",
  13394=>"111111000",
  13395=>"110000111",
  13396=>"111111111",
  13397=>"011000000",
  13398=>"111000000",
  13399=>"010111010",
  13400=>"111000100",
  13401=>"000000000",
  13402=>"110000111",
  13403=>"111110101",
  13404=>"111000000",
  13405=>"000000110",
  13406=>"000000111",
  13407=>"000100100",
  13408=>"000001001",
  13409=>"010000000",
  13410=>"111110111",
  13411=>"000001111",
  13412=>"000000000",
  13413=>"000111111",
  13414=>"000000000",
  13415=>"000000100",
  13416=>"111000000",
  13417=>"111110110",
  13418=>"000000111",
  13419=>"000000111",
  13420=>"000000111",
  13421=>"111000000",
  13422=>"000000111",
  13423=>"000000000",
  13424=>"101001100",
  13425=>"000000111",
  13426=>"000110000",
  13427=>"001000001",
  13428=>"000000000",
  13429=>"111111111",
  13430=>"000000000",
  13431=>"000000001",
  13432=>"000000000",
  13433=>"000001000",
  13434=>"100111000",
  13435=>"111001001",
  13436=>"001011011",
  13437=>"000011111",
  13438=>"001000000",
  13439=>"000000000",
  13440=>"111100000",
  13441=>"100000111",
  13442=>"111101111",
  13443=>"111011000",
  13444=>"111101111",
  13445=>"101001000",
  13446=>"000000000",
  13447=>"111001001",
  13448=>"111010001",
  13449=>"000000011",
  13450=>"111000000",
  13451=>"000000000",
  13452=>"000000111",
  13453=>"111111011",
  13454=>"111111111",
  13455=>"111111000",
  13456=>"000011011",
  13457=>"000100111",
  13458=>"000001101",
  13459=>"111111110",
  13460=>"110000000",
  13461=>"000000111",
  13462=>"000000000",
  13463=>"000100110",
  13464=>"001000100",
  13465=>"001111111",
  13466=>"111000000",
  13467=>"001001101",
  13468=>"111110110",
  13469=>"000000000",
  13470=>"110010111",
  13471=>"110110110",
  13472=>"111111111",
  13473=>"111000000",
  13474=>"000000000",
  13475=>"111000000",
  13476=>"001111000",
  13477=>"111010101",
  13478=>"010010010",
  13479=>"100100111",
  13480=>"000000011",
  13481=>"111111000",
  13482=>"110111111",
  13483=>"101000000",
  13484=>"000000000",
  13485=>"111100000",
  13486=>"111001000",
  13487=>"110000000",
  13488=>"000000001",
  13489=>"001000011",
  13490=>"010111111",
  13491=>"010000000",
  13492=>"000000111",
  13493=>"000111000",
  13494=>"111001001",
  13495=>"111111110",
  13496=>"111000000",
  13497=>"000000000",
  13498=>"000000111",
  13499=>"010010111",
  13500=>"000000111",
  13501=>"000000100",
  13502=>"111111101",
  13503=>"000010110",
  13504=>"011000111",
  13505=>"111110000",
  13506=>"111000000",
  13507=>"111111000",
  13508=>"000101000",
  13509=>"111111111",
  13510=>"110111111",
  13511=>"000000110",
  13512=>"111111111",
  13513=>"000111111",
  13514=>"001111111",
  13515=>"100001011",
  13516=>"110111011",
  13517=>"011111111",
  13518=>"000000000",
  13519=>"010000000",
  13520=>"101101000",
  13521=>"011011010",
  13522=>"011000011",
  13523=>"111000111",
  13524=>"000000111",
  13525=>"000000011",
  13526=>"000011001",
  13527=>"011111111",
  13528=>"111111111",
  13529=>"010000001",
  13530=>"000000001",
  13531=>"111111000",
  13532=>"010000110",
  13533=>"100000010",
  13534=>"000010111",
  13535=>"111111111",
  13536=>"111111000",
  13537=>"000000111",
  13538=>"111000000",
  13539=>"111111111",
  13540=>"000111111",
  13541=>"111001100",
  13542=>"000000101",
  13543=>"000001101",
  13544=>"111111111",
  13545=>"101101000",
  13546=>"111111111",
  13547=>"111000011",
  13548=>"111000000",
  13549=>"000000111",
  13550=>"111000000",
  13551=>"111111010",
  13552=>"011000000",
  13553=>"000000001",
  13554=>"000000111",
  13555=>"111100110",
  13556=>"101000000",
  13557=>"001111001",
  13558=>"111110111",
  13559=>"010111111",
  13560=>"111110000",
  13561=>"111111110",
  13562=>"111000000",
  13563=>"000100000",
  13564=>"001011111",
  13565=>"111111111",
  13566=>"111011011",
  13567=>"000100100",
  13568=>"111000000",
  13569=>"000111110",
  13570=>"111111000",
  13571=>"000000000",
  13572=>"000001001",
  13573=>"101001111",
  13574=>"111111000",
  13575=>"111000000",
  13576=>"110000000",
  13577=>"000111001",
  13578=>"100000111",
  13579=>"111000000",
  13580=>"111000110",
  13581=>"111111111",
  13582=>"110111111",
  13583=>"000111111",
  13584=>"011011011",
  13585=>"111000000",
  13586=>"000001111",
  13587=>"000000000",
  13588=>"000000000",
  13589=>"000001111",
  13590=>"000000010",
  13591=>"000000111",
  13592=>"010100010",
  13593=>"000110110",
  13594=>"001001111",
  13595=>"110010000",
  13596=>"001000000",
  13597=>"000011000",
  13598=>"111111111",
  13599=>"111100001",
  13600=>"000000100",
  13601=>"110110000",
  13602=>"001001111",
  13603=>"111111111",
  13604=>"101111111",
  13605=>"111001111",
  13606=>"000111111",
  13607=>"100000111",
  13608=>"000000011",
  13609=>"111000000",
  13610=>"010000000",
  13611=>"001000110",
  13612=>"000111111",
  13613=>"000000011",
  13614=>"000000010",
  13615=>"000000000",
  13616=>"111000001",
  13617=>"000010010",
  13618=>"111011111",
  13619=>"000111111",
  13620=>"111000000",
  13621=>"011111111",
  13622=>"111101001",
  13623=>"000000110",
  13624=>"111100000",
  13625=>"100000111",
  13626=>"111000000",
  13627=>"111111000",
  13628=>"111110011",
  13629=>"110101000",
  13630=>"000000000",
  13631=>"111111100",
  13632=>"111000000",
  13633=>"000110111",
  13634=>"000000111",
  13635=>"010111111",
  13636=>"000000000",
  13637=>"111111000",
  13638=>"011011111",
  13639=>"000111111",
  13640=>"000000000",
  13641=>"111000000",
  13642=>"111001000",
  13643=>"000111111",
  13644=>"000000000",
  13645=>"011000111",
  13646=>"111010000",
  13647=>"000001111",
  13648=>"111111000",
  13649=>"000111001",
  13650=>"011001111",
  13651=>"000110111",
  13652=>"000000000",
  13653=>"000101000",
  13654=>"111111111",
  13655=>"100100111",
  13656=>"100111111",
  13657=>"010000000",
  13658=>"111010000",
  13659=>"000000100",
  13660=>"001111001",
  13661=>"000000011",
  13662=>"000000111",
  13663=>"110111111",
  13664=>"111111111",
  13665=>"010111000",
  13666=>"111001011",
  13667=>"000111000",
  13668=>"000111111",
  13669=>"111000111",
  13670=>"000000000",
  13671=>"000000111",
  13672=>"000001111",
  13673=>"000001000",
  13674=>"000000000",
  13675=>"010100101",
  13676=>"100000011",
  13677=>"101000111",
  13678=>"000000000",
  13679=>"111111000",
  13680=>"000000000",
  13681=>"110000001",
  13682=>"000001111",
  13683=>"111011001",
  13684=>"111111111",
  13685=>"101101111",
  13686=>"100001000",
  13687=>"010000100",
  13688=>"000111000",
  13689=>"111111000",
  13690=>"110111110",
  13691=>"111110000",
  13692=>"000000000",
  13693=>"011000111",
  13694=>"111111000",
  13695=>"111111000",
  13696=>"010111111",
  13697=>"010011000",
  13698=>"000000000",
  13699=>"000000000",
  13700=>"001000001",
  13701=>"100111000",
  13702=>"000000011",
  13703=>"100000111",
  13704=>"111111111",
  13705=>"111111000",
  13706=>"000000111",
  13707=>"101001100",
  13708=>"111101001",
  13709=>"111100100",
  13710=>"111000100",
  13711=>"010000000",
  13712=>"111111000",
  13713=>"111000110",
  13714=>"000001000",
  13715=>"111100000",
  13716=>"110111100",
  13717=>"111111011",
  13718=>"000000000",
  13719=>"011111110",
  13720=>"111000000",
  13721=>"111111011",
  13722=>"011111111",
  13723=>"010000110",
  13724=>"111111111",
  13725=>"111011010",
  13726=>"000111111",
  13727=>"000000000",
  13728=>"001111110",
  13729=>"011111111",
  13730=>"011011011",
  13731=>"111111000",
  13732=>"111001001",
  13733=>"111111000",
  13734=>"000000111",
  13735=>"110000000",
  13736=>"000000000",
  13737=>"000000000",
  13738=>"000000100",
  13739=>"000000111",
  13740=>"000100111",
  13741=>"110000010",
  13742=>"111101000",
  13743=>"000000001",
  13744=>"000000001",
  13745=>"000000001",
  13746=>"000000001",
  13747=>"000000000",
  13748=>"000000011",
  13749=>"001000111",
  13750=>"100101111",
  13751=>"111001001",
  13752=>"111000000",
  13753=>"000000010",
  13754=>"000001111",
  13755=>"000011101",
  13756=>"000000000",
  13757=>"111111111",
  13758=>"111000000",
  13759=>"101000000",
  13760=>"111001001",
  13761=>"000000111",
  13762=>"111110110",
  13763=>"110000000",
  13764=>"111001010",
  13765=>"111011000",
  13766=>"111111000",
  13767=>"111111000",
  13768=>"111010110",
  13769=>"000000111",
  13770=>"111000000",
  13771=>"111110000",
  13772=>"111000000",
  13773=>"111011000",
  13774=>"111000011",
  13775=>"110111111",
  13776=>"111001000",
  13777=>"000100111",
  13778=>"000111111",
  13779=>"000000010",
  13780=>"000000111",
  13781=>"111000001",
  13782=>"000001111",
  13783=>"011011111",
  13784=>"000001000",
  13785=>"000000000",
  13786=>"111110111",
  13787=>"111100111",
  13788=>"111111111",
  13789=>"111111000",
  13790=>"011001000",
  13791=>"000000011",
  13792=>"111111001",
  13793=>"100000000",
  13794=>"100000111",
  13795=>"111111111",
  13796=>"000000110",
  13797=>"111000000",
  13798=>"001100111",
  13799=>"000000101",
  13800=>"111000111",
  13801=>"111111000",
  13802=>"000000010",
  13803=>"000000000",
  13804=>"111000000",
  13805=>"100110111",
  13806=>"000010110",
  13807=>"000000100",
  13808=>"000000000",
  13809=>"111111111",
  13810=>"110111111",
  13811=>"000111111",
  13812=>"011111111",
  13813=>"000000000",
  13814=>"111111111",
  13815=>"000011111",
  13816=>"111010000",
  13817=>"000000100",
  13818=>"111000110",
  13819=>"111000111",
  13820=>"000000000",
  13821=>"000000110",
  13822=>"000010011",
  13823=>"011001000",
  13824=>"000000110",
  13825=>"111001111",
  13826=>"011000000",
  13827=>"110110000",
  13828=>"001000000",
  13829=>"000000001",
  13830=>"111111100",
  13831=>"000000000",
  13832=>"000100100",
  13833=>"000000110",
  13834=>"000000000",
  13835=>"000110000",
  13836=>"010010010",
  13837=>"001000100",
  13838=>"101111111",
  13839=>"111111111",
  13840=>"000000001",
  13841=>"011111001",
  13842=>"111111111",
  13843=>"000000000",
  13844=>"111111111",
  13845=>"000000101",
  13846=>"101100100",
  13847=>"111011101",
  13848=>"111000101",
  13849=>"111100100",
  13850=>"001000110",
  13851=>"000010010",
  13852=>"111101101",
  13853=>"111111111",
  13854=>"111011111",
  13855=>"111111000",
  13856=>"000000000",
  13857=>"111110010",
  13858=>"111110100",
  13859=>"001001101",
  13860=>"001001011",
  13861=>"101100000",
  13862=>"000011011",
  13863=>"000111111",
  13864=>"000000001",
  13865=>"000011111",
  13866=>"010110000",
  13867=>"111110110",
  13868=>"111111101",
  13869=>"111111111",
  13870=>"000000000",
  13871=>"111111111",
  13872=>"110100111",
  13873=>"100100000",
  13874=>"011001011",
  13875=>"111110111",
  13876=>"000000000",
  13877=>"110000000",
  13878=>"000000000",
  13879=>"001111111",
  13880=>"011011011",
  13881=>"100110100",
  13882=>"000000000",
  13883=>"111000000",
  13884=>"111001111",
  13885=>"001000000",
  13886=>"001011111",
  13887=>"111111100",
  13888=>"000000000",
  13889=>"000000000",
  13890=>"000101111",
  13891=>"000000111",
  13892=>"000000000",
  13893=>"100100100",
  13894=>"111111000",
  13895=>"111111111",
  13896=>"011000000",
  13897=>"111101110",
  13898=>"000000000",
  13899=>"111011111",
  13900=>"000110110",
  13901=>"011110000",
  13902=>"000000000",
  13903=>"110111111",
  13904=>"111111000",
  13905=>"111111111",
  13906=>"000000000",
  13907=>"000000000",
  13908=>"101111110",
  13909=>"111111110",
  13910=>"000001001",
  13911=>"000000100",
  13912=>"000000000",
  13913=>"000000000",
  13914=>"000100111",
  13915=>"000000001",
  13916=>"001001001",
  13917=>"111111111",
  13918=>"000000000",
  13919=>"000000010",
  13920=>"000000100",
  13921=>"111111111",
  13922=>"000000000",
  13923=>"111111111",
  13924=>"000000000",
  13925=>"000000000",
  13926=>"110110000",
  13927=>"000000000",
  13928=>"000010111",
  13929=>"000000000",
  13930=>"000010000",
  13931=>"000000000",
  13932=>"010011111",
  13933=>"111101000",
  13934=>"110110111",
  13935=>"000100100",
  13936=>"000001111",
  13937=>"110011000",
  13938=>"000001001",
  13939=>"000100001",
  13940=>"101101100",
  13941=>"111111111",
  13942=>"011111000",
  13943=>"000000000",
  13944=>"010000000",
  13945=>"110111111",
  13946=>"101101111",
  13947=>"000000001",
  13948=>"110110110",
  13949=>"111111111",
  13950=>"111111111",
  13951=>"000001011",
  13952=>"111111010",
  13953=>"111110100",
  13954=>"101000000",
  13955=>"010000111",
  13956=>"111111111",
  13957=>"111111111",
  13958=>"011111111",
  13959=>"001000000",
  13960=>"110111111",
  13961=>"111110000",
  13962=>"000000000",
  13963=>"000000000",
  13964=>"011111010",
  13965=>"100000000",
  13966=>"100111111",
  13967=>"000000000",
  13968=>"000000111",
  13969=>"000001000",
  13970=>"111111111",
  13971=>"101001000",
  13972=>"100100110",
  13973=>"000000000",
  13974=>"100100000",
  13975=>"000000000",
  13976=>"001001000",
  13977=>"111011011",
  13978=>"111111111",
  13979=>"000000000",
  13980=>"111101101",
  13981=>"000000000",
  13982=>"111111100",
  13983=>"000000000",
  13984=>"000000110",
  13985=>"000001001",
  13986=>"111011111",
  13987=>"100110111",
  13988=>"001001000",
  13989=>"010110111",
  13990=>"011111111",
  13991=>"111111011",
  13992=>"111110011",
  13993=>"111111111",
  13994=>"000000000",
  13995=>"100000000",
  13996=>"111111111",
  13997=>"110100111",
  13998=>"001001001",
  13999=>"110010001",
  14000=>"011011011",
  14001=>"010011001",
  14002=>"101101101",
  14003=>"100000111",
  14004=>"111111111",
  14005=>"000100100",
  14006=>"000000000",
  14007=>"001100101",
  14008=>"001000000",
  14009=>"111001000",
  14010=>"000000000",
  14011=>"111100000",
  14012=>"000000000",
  14013=>"111110000",
  14014=>"111001000",
  14015=>"000000100",
  14016=>"111001111",
  14017=>"001000000",
  14018=>"111111011",
  14019=>"111111111",
  14020=>"000000000",
  14021=>"111001010",
  14022=>"000000000",
  14023=>"011111111",
  14024=>"111111111",
  14025=>"110111011",
  14026=>"110111111",
  14027=>"011111111",
  14028=>"111111011",
  14029=>"001110000",
  14030=>"100001000",
  14031=>"000000000",
  14032=>"011000000",
  14033=>"110111111",
  14034=>"101100101",
  14035=>"000000000",
  14036=>"000000000",
  14037=>"110000000",
  14038=>"111111111",
  14039=>"011110110",
  14040=>"111110111",
  14041=>"011110110",
  14042=>"000010000",
  14043=>"000000000",
  14044=>"010000000",
  14045=>"111111111",
  14046=>"111111011",
  14047=>"011111010",
  14048=>"001111111",
  14049=>"011111111",
  14050=>"000001001",
  14051=>"111111111",
  14052=>"111111001",
  14053=>"101001000",
  14054=>"111111111",
  14055=>"011111111",
  14056=>"111000000",
  14057=>"000000000",
  14058=>"000111111",
  14059=>"000100010",
  14060=>"010010000",
  14061=>"100100000",
  14062=>"100111111",
  14063=>"000011111",
  14064=>"101000000",
  14065=>"000110111",
  14066=>"000001001",
  14067=>"000000000",
  14068=>"111111111",
  14069=>"000000110",
  14070=>"001011011",
  14071=>"000000000",
  14072=>"111111111",
  14073=>"000000000",
  14074=>"111111111",
  14075=>"000000000",
  14076=>"111111110",
  14077=>"001000010",
  14078=>"000000000",
  14079=>"111111111",
  14080=>"000000000",
  14081=>"100101001",
  14082=>"000000111",
  14083=>"000110111",
  14084=>"100000000",
  14085=>"111111011",
  14086=>"111111111",
  14087=>"000000000",
  14088=>"111111111",
  14089=>"000000000",
  14090=>"110110100",
  14091=>"001000000",
  14092=>"001011001",
  14093=>"000000110",
  14094=>"000110110",
  14095=>"010010000",
  14096=>"100110110",
  14097=>"111111111",
  14098=>"111111111",
  14099=>"000001111",
  14100=>"011110000",
  14101=>"100100101",
  14102=>"011011011",
  14103=>"000110111",
  14104=>"111111110",
  14105=>"110110111",
  14106=>"110110100",
  14107=>"011001100",
  14108=>"110100000",
  14109=>"110000100",
  14110=>"011111011",
  14111=>"000000001",
  14112=>"000001100",
  14113=>"001001111",
  14114=>"000100000",
  14115=>"111111000",
  14116=>"001100100",
  14117=>"111110111",
  14118=>"000000000",
  14119=>"100001100",
  14120=>"111111001",
  14121=>"000100100",
  14122=>"111111111",
  14123=>"010000000",
  14124=>"011010000",
  14125=>"000000000",
  14126=>"000000000",
  14127=>"000000001",
  14128=>"100101111",
  14129=>"111011100",
  14130=>"011000111",
  14131=>"110110100",
  14132=>"111111111",
  14133=>"100000000",
  14134=>"011111011",
  14135=>"111000001",
  14136=>"111111111",
  14137=>"000000111",
  14138=>"010110110",
  14139=>"000000000",
  14140=>"100000000",
  14141=>"011111011",
  14142=>"111110100",
  14143=>"111001111",
  14144=>"111111111",
  14145=>"011001001",
  14146=>"111100110",
  14147=>"111111111",
  14148=>"001111111",
  14149=>"011000000",
  14150=>"100100000",
  14151=>"110111110",
  14152=>"111111111",
  14153=>"111111111",
  14154=>"111001001",
  14155=>"110011111",
  14156=>"101100000",
  14157=>"111111001",
  14158=>"001100000",
  14159=>"000000000",
  14160=>"111011000",
  14161=>"010000000",
  14162=>"111110111",
  14163=>"010000111",
  14164=>"000000110",
  14165=>"111011001",
  14166=>"111111111",
  14167=>"111111111",
  14168=>"111111111",
  14169=>"111111111",
  14170=>"100000000",
  14171=>"001011111",
  14172=>"110110111",
  14173=>"000000000",
  14174=>"111111110",
  14175=>"111111111",
  14176=>"001101111",
  14177=>"001000000",
  14178=>"110110011",
  14179=>"110111011",
  14180=>"000000010",
  14181=>"000000000",
  14182=>"011000100",
  14183=>"111111110",
  14184=>"000100101",
  14185=>"000111111",
  14186=>"111101001",
  14187=>"000001111",
  14188=>"000001000",
  14189=>"000000000",
  14190=>"000000000",
  14191=>"110111111",
  14192=>"001100001",
  14193=>"000000111",
  14194=>"110111000",
  14195=>"110111110",
  14196=>"000000000",
  14197=>"111101101",
  14198=>"111000111",
  14199=>"000010111",
  14200=>"111111110",
  14201=>"111010111",
  14202=>"110110000",
  14203=>"011110110",
  14204=>"011011111",
  14205=>"111111111",
  14206=>"110100110",
  14207=>"000001001",
  14208=>"011111010",
  14209=>"011111111",
  14210=>"100100000",
  14211=>"111111111",
  14212=>"111111110",
  14213=>"000000000",
  14214=>"101111000",
  14215=>"000000001",
  14216=>"100111000",
  14217=>"110000001",
  14218=>"111011011",
  14219=>"111111011",
  14220=>"111111111",
  14221=>"001101101",
  14222=>"011011000",
  14223=>"000000000",
  14224=>"111111111",
  14225=>"111111100",
  14226=>"000111111",
  14227=>"111101101",
  14228=>"111111011",
  14229=>"001000111",
  14230=>"111100111",
  14231=>"110110010",
  14232=>"111111111",
  14233=>"101100111",
  14234=>"011111110",
  14235=>"111111111",
  14236=>"100000000",
  14237=>"100111110",
  14238=>"001001000",
  14239=>"111111111",
  14240=>"111111001",
  14241=>"100000000",
  14242=>"010010100",
  14243=>"000000001",
  14244=>"111111010",
  14245=>"000000000",
  14246=>"101000000",
  14247=>"000111000",
  14248=>"100001001",
  14249=>"011011010",
  14250=>"000000001",
  14251=>"110000000",
  14252=>"100010010",
  14253=>"001110010",
  14254=>"000100000",
  14255=>"011011011",
  14256=>"001001001",
  14257=>"111111111",
  14258=>"101001000",
  14259=>"010111000",
  14260=>"001101101",
  14261=>"111111110",
  14262=>"110000001",
  14263=>"100001000",
  14264=>"101100111",
  14265=>"000011011",
  14266=>"000101001",
  14267=>"100110101",
  14268=>"001111111",
  14269=>"000000000",
  14270=>"001011011",
  14271=>"111000000",
  14272=>"111111100",
  14273=>"000001100",
  14274=>"000000000",
  14275=>"111111111",
  14276=>"000101111",
  14277=>"000000110",
  14278=>"001100111",
  14279=>"001001111",
  14280=>"111111111",
  14281=>"101100111",
  14282=>"000000111",
  14283=>"000000111",
  14284=>"100110000",
  14285=>"000000100",
  14286=>"001111111",
  14287=>"111110100",
  14288=>"111011000",
  14289=>"001011011",
  14290=>"000000111",
  14291=>"111111000",
  14292=>"011111010",
  14293=>"000000101",
  14294=>"100000000",
  14295=>"001000011",
  14296=>"111000001",
  14297=>"000000000",
  14298=>"000000000",
  14299=>"110110100",
  14300=>"001000111",
  14301=>"111111010",
  14302=>"000000000",
  14303=>"011110000",
  14304=>"000000101",
  14305=>"000000100",
  14306=>"100000001",
  14307=>"111111111",
  14308=>"111111111",
  14309=>"110100111",
  14310=>"011011001",
  14311=>"000000100",
  14312=>"011011111",
  14313=>"000100110",
  14314=>"001100110",
  14315=>"111111111",
  14316=>"101101001",
  14317=>"001011011",
  14318=>"110100000",
  14319=>"011111110",
  14320=>"000000000",
  14321=>"001111111",
  14322=>"000000101",
  14323=>"000000000",
  14324=>"011001000",
  14325=>"111000000",
  14326=>"110100000",
  14327=>"111011010",
  14328=>"111111011",
  14329=>"001001001",
  14330=>"111111111",
  14331=>"000000000",
  14332=>"111111100",
  14333=>"001000100",
  14334=>"000111011",
  14335=>"111111111",
  14336=>"011011001",
  14337=>"000000000",
  14338=>"000000111",
  14339=>"101000000",
  14340=>"111111111",
  14341=>"011111000",
  14342=>"101101111",
  14343=>"000000111",
  14344=>"111000111",
  14345=>"111111110",
  14346=>"001001000",
  14347=>"000100110",
  14348=>"000111000",
  14349=>"011100100",
  14350=>"111111111",
  14351=>"011000111",
  14352=>"011000000",
  14353=>"101001111",
  14354=>"011001110",
  14355=>"111111111",
  14356=>"100100111",
  14357=>"000000111",
  14358=>"000000000",
  14359=>"000000000",
  14360=>"111010000",
  14361=>"000010111",
  14362=>"100000000",
  14363=>"000000100",
  14364=>"111000001",
  14365=>"010010000",
  14366=>"000000100",
  14367=>"111000000",
  14368=>"001001111",
  14369=>"000000111",
  14370=>"001000000",
  14371=>"001111110",
  14372=>"111111011",
  14373=>"000000111",
  14374=>"000000111",
  14375=>"100000000",
  14376=>"101111111",
  14377=>"011000000",
  14378=>"111110001",
  14379=>"100100011",
  14380=>"000010111",
  14381=>"111001111",
  14382=>"001111111",
  14383=>"000010000",
  14384=>"000001111",
  14385=>"011011111",
  14386=>"000000000",
  14387=>"111111111",
  14388=>"000000000",
  14389=>"111111001",
  14390=>"001000111",
  14391=>"111101101",
  14392=>"000000111",
  14393=>"000000000",
  14394=>"111111000",
  14395=>"111000110",
  14396=>"000101111",
  14397=>"001001111",
  14398=>"011010000",
  14399=>"001000111",
  14400=>"001000001",
  14401=>"000111111",
  14402=>"100110110",
  14403=>"111111111",
  14404=>"011000000",
  14405=>"110000000",
  14406=>"000000011",
  14407=>"100010011",
  14408=>"000000111",
  14409=>"111111111",
  14410=>"000000000",
  14411=>"000000011",
  14412=>"000010110",
  14413=>"111111111",
  14414=>"111101001",
  14415=>"000000000",
  14416=>"100111100",
  14417=>"111111000",
  14418=>"111111000",
  14419=>"001000011",
  14420=>"111111011",
  14421=>"111111000",
  14422=>"000000000",
  14423=>"000000000",
  14424=>"011000000",
  14425=>"100100101",
  14426=>"011011000",
  14427=>"000100100",
  14428=>"111111000",
  14429=>"001011011",
  14430=>"111110110",
  14431=>"000000000",
  14432=>"111011000",
  14433=>"000000000",
  14434=>"111000100",
  14435=>"111000100",
  14436=>"011110110",
  14437=>"100011011",
  14438=>"111010000",
  14439=>"110110100",
  14440=>"000000000",
  14441=>"001000000",
  14442=>"100000000",
  14443=>"000000000",
  14444=>"000000101",
  14445=>"101111111",
  14446=>"111111010",
  14447=>"000000000",
  14448=>"101111000",
  14449=>"000000000",
  14450=>"111111000",
  14451=>"011011011",
  14452=>"100111111",
  14453=>"011000110",
  14454=>"001000010",
  14455=>"111000011",
  14456=>"111111111",
  14457=>"100111111",
  14458=>"111000000",
  14459=>"111001000",
  14460=>"010010000",
  14461=>"011011011",
  14462=>"111000000",
  14463=>"000000011",
  14464=>"001111110",
  14465=>"000000110",
  14466=>"111111111",
  14467=>"000000000",
  14468=>"110110100",
  14469=>"111111111",
  14470=>"111101100",
  14471=>"000000111",
  14472=>"000000111",
  14473=>"000000000",
  14474=>"111111000",
  14475=>"001111111",
  14476=>"001001100",
  14477=>"001001001",
  14478=>"011110111",
  14479=>"111111000",
  14480=>"111111111",
  14481=>"011011111",
  14482=>"001000000",
  14483=>"000110000",
  14484=>"110111111",
  14485=>"100000110",
  14486=>"011000000",
  14487=>"111001111",
  14488=>"100001001",
  14489=>"000000000",
  14490=>"100000000",
  14491=>"111111111",
  14492=>"100111100",
  14493=>"111111001",
  14494=>"000000111",
  14495=>"111111111",
  14496=>"000000100",
  14497=>"100111100",
  14498=>"111110000",
  14499=>"111111000",
  14500=>"111001100",
  14501=>"100000000",
  14502=>"011000000",
  14503=>"111111100",
  14504=>"110000111",
  14505=>"000000000",
  14506=>"111111111",
  14507=>"000000000",
  14508=>"001001001",
  14509=>"000110111",
  14510=>"101000100",
  14511=>"100011110",
  14512=>"111111111",
  14513=>"000000111",
  14514=>"110110111",
  14515=>"001000100",
  14516=>"001001110",
  14517=>"111111111",
  14518=>"000000000",
  14519=>"111111000",
  14520=>"001100111",
  14521=>"000000111",
  14522=>"111101111",
  14523=>"100101011",
  14524=>"000100101",
  14525=>"000011000",
  14526=>"000110111",
  14527=>"111000000",
  14528=>"111110110",
  14529=>"111111110",
  14530=>"000000001",
  14531=>"111100000",
  14532=>"011111111",
  14533=>"000000111",
  14534=>"000000111",
  14535=>"101111111",
  14536=>"001000111",
  14537=>"000000111",
  14538=>"111111000",
  14539=>"110111110",
  14540=>"101111111",
  14541=>"000111000",
  14542=>"110000100",
  14543=>"111101000",
  14544=>"111111111",
  14545=>"000000000",
  14546=>"111111110",
  14547=>"110111111",
  14548=>"111111000",
  14549=>"111011000",
  14550=>"000000111",
  14551=>"000000000",
  14552=>"111000000",
  14553=>"000000001",
  14554=>"000000000",
  14555=>"100000000",
  14556=>"001000101",
  14557=>"110110000",
  14558=>"000000110",
  14559=>"000000111",
  14560=>"000001111",
  14561=>"000000111",
  14562=>"000111111",
  14563=>"101001001",
  14564=>"111010000",
  14565=>"001001011",
  14566=>"111110111",
  14567=>"111001000",
  14568=>"111111111",
  14569=>"111111111",
  14570=>"001111111",
  14571=>"000000100",
  14572=>"111111000",
  14573=>"010010000",
  14574=>"011111111",
  14575=>"010000000",
  14576=>"100110111",
  14577=>"111101000",
  14578=>"111111110",
  14579=>"000000111",
  14580=>"101111111",
  14581=>"000000010",
  14582=>"100011010",
  14583=>"000111111",
  14584=>"000100110",
  14585=>"000000000",
  14586=>"000110111",
  14587=>"011011000",
  14588=>"001001000",
  14589=>"000000111",
  14590=>"110000000",
  14591=>"000000100",
  14592=>"001111111",
  14593=>"111111100",
  14594=>"000000000",
  14595=>"111111000",
  14596=>"100111111",
  14597=>"110100000",
  14598=>"111111001",
  14599=>"111111000",
  14600=>"000110100",
  14601=>"111111111",
  14602=>"000111110",
  14603=>"000001111",
  14604=>"111101000",
  14605=>"101111110",
  14606=>"111111111",
  14607=>"000111111",
  14608=>"100100100",
  14609=>"001111101",
  14610=>"011011000",
  14611=>"001111111",
  14612=>"111111001",
  14613=>"111100100",
  14614=>"010001111",
  14615=>"000000000",
  14616=>"000111111",
  14617=>"001000000",
  14618=>"000001111",
  14619=>"010000111",
  14620=>"000000011",
  14621=>"011011010",
  14622=>"000000000",
  14623=>"000000100",
  14624=>"100110100",
  14625=>"111111010",
  14626=>"000101111",
  14627=>"000000111",
  14628=>"110000101",
  14629=>"111111111",
  14630=>"001101111",
  14631=>"110100000",
  14632=>"000000000",
  14633=>"111111101",
  14634=>"001000000",
  14635=>"000010111",
  14636=>"000000111",
  14637=>"100000000",
  14638=>"000110110",
  14639=>"110000000",
  14640=>"111111111",
  14641=>"001101111",
  14642=>"000010110",
  14643=>"111110011",
  14644=>"001001000",
  14645=>"001001011",
  14646=>"010000000",
  14647=>"000111111",
  14648=>"000111111",
  14649=>"111111111",
  14650=>"011111111",
  14651=>"100100000",
  14652=>"000110111",
  14653=>"111110000",
  14654=>"101000110",
  14655=>"111111000",
  14656=>"011111000",
  14657=>"100000000",
  14658=>"000000000",
  14659=>"000001111",
  14660=>"111111111",
  14661=>"000000110",
  14662=>"100100111",
  14663=>"100000100",
  14664=>"000000111",
  14665=>"111000111",
  14666=>"111110111",
  14667=>"011010011",
  14668=>"111100111",
  14669=>"000110111",
  14670=>"110100111",
  14671=>"111111000",
  14672=>"001001011",
  14673=>"000000110",
  14674=>"111111111",
  14675=>"111100000",
  14676=>"001000000",
  14677=>"001011001",
  14678=>"111010000",
  14679=>"001010010",
  14680=>"111111100",
  14681=>"111111000",
  14682=>"000000000",
  14683=>"111111110",
  14684=>"000100101",
  14685=>"001001000",
  14686=>"111110000",
  14687=>"111111001",
  14688=>"000000000",
  14689=>"111000000",
  14690=>"100000000",
  14691=>"111111000",
  14692=>"111111011",
  14693=>"000000111",
  14694=>"000000110",
  14695=>"111111111",
  14696=>"001000001",
  14697=>"000110111",
  14698=>"111111111",
  14699=>"000000000",
  14700=>"000111111",
  14701=>"000000110",
  14702=>"000000000",
  14703=>"111000000",
  14704=>"101000100",
  14705=>"010111111",
  14706=>"000000001",
  14707=>"001111011",
  14708=>"110100100",
  14709=>"000000000",
  14710=>"001111000",
  14711=>"111111111",
  14712=>"110101111",
  14713=>"011011000",
  14714=>"000000110",
  14715=>"101111110",
  14716=>"100100111",
  14717=>"101000000",
  14718=>"100000000",
  14719=>"001001000",
  14720=>"000000000",
  14721=>"000000100",
  14722=>"111111000",
  14723=>"110110100",
  14724=>"010011001",
  14725=>"111101011",
  14726=>"000000000",
  14727=>"000000011",
  14728=>"111111000",
  14729=>"000100111",
  14730=>"100111111",
  14731=>"110000000",
  14732=>"111111101",
  14733=>"000000000",
  14734=>"111111110",
  14735=>"111000000",
  14736=>"100010000",
  14737=>"011101111",
  14738=>"111111111",
  14739=>"001001011",
  14740=>"000000000",
  14741=>"000011111",
  14742=>"111110110",
  14743=>"000011011",
  14744=>"001000100",
  14745=>"000000000",
  14746=>"101111111",
  14747=>"001011111",
  14748=>"111111111",
  14749=>"000000011",
  14750=>"000101111",
  14751=>"111111111",
  14752=>"111000000",
  14753=>"011011000",
  14754=>"001000111",
  14755=>"111111000",
  14756=>"001000100",
  14757=>"011111111",
  14758=>"011000100",
  14759=>"000111111",
  14760=>"000000000",
  14761=>"000100111",
  14762=>"111110000",
  14763=>"000000101",
  14764=>"100111100",
  14765=>"000000000",
  14766=>"000110111",
  14767=>"100000110",
  14768=>"011110111",
  14769=>"000000011",
  14770=>"111111111",
  14771=>"001000011",
  14772=>"111111011",
  14773=>"001000000",
  14774=>"111011000",
  14775=>"010000110",
  14776=>"000000000",
  14777=>"110000011",
  14778=>"101001011",
  14779=>"111111111",
  14780=>"111111111",
  14781=>"111111111",
  14782=>"110111110",
  14783=>"100100111",
  14784=>"000000110",
  14785=>"111110000",
  14786=>"111110111",
  14787=>"000110110",
  14788=>"000000000",
  14789=>"111111000",
  14790=>"000000001",
  14791=>"001001000",
  14792=>"100000011",
  14793=>"101000100",
  14794=>"000000000",
  14795=>"111111010",
  14796=>"000111000",
  14797=>"111111001",
  14798=>"101100000",
  14799=>"000000000",
  14800=>"111111111",
  14801=>"111100000",
  14802=>"100000000",
  14803=>"110110111",
  14804=>"000000000",
  14805=>"111111111",
  14806=>"000000000",
  14807=>"100000000",
  14808=>"000111111",
  14809=>"001011111",
  14810=>"000000000",
  14811=>"111111111",
  14812=>"111110111",
  14813=>"111111000",
  14814=>"010000111",
  14815=>"100000011",
  14816=>"111100111",
  14817=>"100000110",
  14818=>"111000000",
  14819=>"000100000",
  14820=>"001000000",
  14821=>"111111000",
  14822=>"111111111",
  14823=>"100110110",
  14824=>"000111111",
  14825=>"000001111",
  14826=>"111001000",
  14827=>"000100111",
  14828=>"011000000",
  14829=>"000000111",
  14830=>"111001111",
  14831=>"111111111",
  14832=>"111000000",
  14833=>"111100000",
  14834=>"000000000",
  14835=>"000000111",
  14836=>"001000001",
  14837=>"111111011",
  14838=>"000000111",
  14839=>"000010111",
  14840=>"111111111",
  14841=>"001011111",
  14842=>"011011110",
  14843=>"000111111",
  14844=>"100111111",
  14845=>"111000000",
  14846=>"100100000",
  14847=>"111111111",
  14848=>"101101000",
  14849=>"100000001",
  14850=>"111111111",
  14851=>"111101111",
  14852=>"100110010",
  14853=>"000000000",
  14854=>"011011011",
  14855=>"100100000",
  14856=>"011100000",
  14857=>"111111101",
  14858=>"111100000",
  14859=>"110000001",
  14860=>"111001000",
  14861=>"110111000",
  14862=>"100100110",
  14863=>"000000111",
  14864=>"000000100",
  14865=>"111111000",
  14866=>"000011011",
  14867=>"111111011",
  14868=>"000100110",
  14869=>"111111111",
  14870=>"111011000",
  14871=>"000011111",
  14872=>"001000000",
  14873=>"010111001",
  14874=>"111111111",
  14875=>"000000001",
  14876=>"011000000",
  14877=>"111111111",
  14878=>"111111011",
  14879=>"011111111",
  14880=>"000000000",
  14881=>"100110110",
  14882=>"000001111",
  14883=>"111111111",
  14884=>"000001111",
  14885=>"111110111",
  14886=>"111111111",
  14887=>"100110110",
  14888=>"000100001",
  14889=>"111101000",
  14890=>"100101111",
  14891=>"101000000",
  14892=>"001000000",
  14893=>"111011000",
  14894=>"111010000",
  14895=>"000011010",
  14896=>"000011001",
  14897=>"011001011",
  14898=>"111111111",
  14899=>"000000000",
  14900=>"111111111",
  14901=>"110000111",
  14902=>"000001011",
  14903=>"011000000",
  14904=>"000000000",
  14905=>"000000100",
  14906=>"000000100",
  14907=>"000000000",
  14908=>"000000000",
  14909=>"111111111",
  14910=>"111111111",
  14911=>"000000000",
  14912=>"111100111",
  14913=>"101101111",
  14914=>"011110000",
  14915=>"111111100",
  14916=>"000000000",
  14917=>"000000000",
  14918=>"000111000",
  14919=>"111111111",
  14920=>"111111011",
  14921=>"000000000",
  14922=>"000000000",
  14923=>"000111111",
  14924=>"001001000",
  14925=>"110010000",
  14926=>"000000000",
  14927=>"111111111",
  14928=>"000000000",
  14929=>"111111000",
  14930=>"000100100",
  14931=>"000000101",
  14932=>"011000000",
  14933=>"000100110",
  14934=>"001111111",
  14935=>"011000000",
  14936=>"111111111",
  14937=>"000000000",
  14938=>"000011001",
  14939=>"000000100",
  14940=>"000110000",
  14941=>"000000000",
  14942=>"001111000",
  14943=>"100100100",
  14944=>"110111111",
  14945=>"000000111",
  14946=>"100010111",
  14947=>"000000000",
  14948=>"001000000",
  14949=>"101000100",
  14950=>"111001001",
  14951=>"010011000",
  14952=>"111111001",
  14953=>"010011011",
  14954=>"000110110",
  14955=>"111111111",
  14956=>"111011001",
  14957=>"010111110",
  14958=>"000000000",
  14959=>"000000000",
  14960=>"100111111",
  14961=>"100110100",
  14962=>"111010000",
  14963=>"001011111",
  14964=>"000000111",
  14965=>"000001011",
  14966=>"000000001",
  14967=>"000000100",
  14968=>"000000000",
  14969=>"000100100",
  14970=>"111011011",
  14971=>"000000000",
  14972=>"011011011",
  14973=>"111111111",
  14974=>"111111111",
  14975=>"001001000",
  14976=>"000000000",
  14977=>"000001011",
  14978=>"000000000",
  14979=>"000111000",
  14980=>"111101101",
  14981=>"100101000",
  14982=>"101111000",
  14983=>"001001000",
  14984=>"000101111",
  14985=>"010010001",
  14986=>"001000000",
  14987=>"110111110",
  14988=>"111111111",
  14989=>"000000000",
  14990=>"000101111",
  14991=>"000000111",
  14992=>"111111111",
  14993=>"011011000",
  14994=>"111111111",
  14995=>"110110110",
  14996=>"000000000",
  14997=>"000100000",
  14998=>"000000000",
  14999=>"101101101",
  15000=>"100000000",
  15001=>"000000100",
  15002=>"111111111",
  15003=>"111111111",
  15004=>"000000000",
  15005=>"101101000",
  15006=>"000111100",
  15007=>"000110010",
  15008=>"010000100",
  15009=>"000000000",
  15010=>"000001101",
  15011=>"000000000",
  15012=>"011001101",
  15013=>"000001111",
  15014=>"000000111",
  15015=>"111111111",
  15016=>"101111101",
  15017=>"000000000",
  15018=>"000101000",
  15019=>"000011010",
  15020=>"110111111",
  15021=>"111111111",
  15022=>"001111111",
  15023=>"111111111",
  15024=>"000000000",
  15025=>"000111111",
  15026=>"111111111",
  15027=>"000000000",
  15028=>"000000000",
  15029=>"110000000",
  15030=>"011111111",
  15031=>"111111111",
  15032=>"000111100",
  15033=>"111000111",
  15034=>"010000000",
  15035=>"111011001",
  15036=>"111111111",
  15037=>"101111110",
  15038=>"000000000",
  15039=>"111001101",
  15040=>"001000000",
  15041=>"110111111",
  15042=>"000100000",
  15043=>"000001000",
  15044=>"010010011",
  15045=>"000000000",
  15046=>"000000100",
  15047=>"001100100",
  15048=>"110000110",
  15049=>"001001000",
  15050=>"000111111",
  15051=>"111111111",
  15052=>"000000111",
  15053=>"111111111",
  15054=>"100110000",
  15055=>"000000100",
  15056=>"110000011",
  15057=>"111011000",
  15058=>"011000000",
  15059=>"111111111",
  15060=>"011000111",
  15061=>"000001001",
  15062=>"110111001",
  15063=>"000000000",
  15064=>"101101111",
  15065=>"100000000",
  15066=>"000000000",
  15067=>"001100000",
  15068=>"000000000",
  15069=>"001000000",
  15070=>"000011111",
  15071=>"001011011",
  15072=>"111110000",
  15073=>"110111000",
  15074=>"000000000",
  15075=>"100100000",
  15076=>"000000000",
  15077=>"111111001",
  15078=>"000000000",
  15079=>"111100000",
  15080=>"101111000",
  15081=>"111111111",
  15082=>"111000000",
  15083=>"111111111",
  15084=>"111111111",
  15085=>"000000000",
  15086=>"000000001",
  15087=>"101000000",
  15088=>"000000100",
  15089=>"111111111",
  15090=>"000000111",
  15091=>"001101110",
  15092=>"111101000",
  15093=>"011001001",
  15094=>"110100110",
  15095=>"111111100",
  15096=>"101111000",
  15097=>"111000000",
  15098=>"000000000",
  15099=>"111111111",
  15100=>"110111111",
  15101=>"000000000",
  15102=>"110111111",
  15103=>"111111111",
  15104=>"000000000",
  15105=>"011011111",
  15106=>"111111111",
  15107=>"111111111",
  15108=>"000100100",
  15109=>"000000010",
  15110=>"111101111",
  15111=>"000111111",
  15112=>"111111110",
  15113=>"101101111",
  15114=>"001100111",
  15115=>"000000000",
  15116=>"111111111",
  15117=>"111111111",
  15118=>"000000111",
  15119=>"001001111",
  15120=>"111110111",
  15121=>"001001000",
  15122=>"111111001",
  15123=>"000000000",
  15124=>"110111110",
  15125=>"000000001",
  15126=>"110110111",
  15127=>"011111000",
  15128=>"111111011",
  15129=>"111111111",
  15130=>"001011011",
  15131=>"000000000",
  15132=>"110100100",
  15133=>"000000000",
  15134=>"000101000",
  15135=>"111111000",
  15136=>"110111111",
  15137=>"000000000",
  15138=>"110110111",
  15139=>"000100100",
  15140=>"100100111",
  15141=>"001011011",
  15142=>"111001001",
  15143=>"100110111",
  15144=>"110111111",
  15145=>"111111111",
  15146=>"001001011",
  15147=>"111111000",
  15148=>"100110110",
  15149=>"001001001",
  15150=>"101101000",
  15151=>"001000000",
  15152=>"000100000",
  15153=>"010000000",
  15154=>"010000011",
  15155=>"000011000",
  15156=>"000000000",
  15157=>"111111110",
  15158=>"101101100",
  15159=>"100100111",
  15160=>"111111011",
  15161=>"001111001",
  15162=>"011010000",
  15163=>"111000000",
  15164=>"000000000",
  15165=>"000000000",
  15166=>"000000000",
  15167=>"000000000",
  15168=>"000000111",
  15169=>"111111111",
  15170=>"000000000",
  15171=>"000000111",
  15172=>"000001000",
  15173=>"000000001",
  15174=>"000000000",
  15175=>"111111111",
  15176=>"000011001",
  15177=>"110000000",
  15178=>"000000000",
  15179=>"100000001",
  15180=>"000000101",
  15181=>"000000000",
  15182=>"000000000",
  15183=>"100110111",
  15184=>"111011001",
  15185=>"000000000",
  15186=>"000000111",
  15187=>"111111110",
  15188=>"000001001",
  15189=>"000010010",
  15190=>"110111111",
  15191=>"011011100",
  15192=>"001111111",
  15193=>"111111000",
  15194=>"001111011",
  15195=>"111100000",
  15196=>"111111111",
  15197=>"111111100",
  15198=>"101101001",
  15199=>"100110110",
  15200=>"000000000",
  15201=>"111111111",
  15202=>"011101111",
  15203=>"100110100",
  15204=>"011001111",
  15205=>"110101000",
  15206=>"100100000",
  15207=>"111111111",
  15208=>"001011111",
  15209=>"101111111",
  15210=>"000000000",
  15211=>"111111011",
  15212=>"111111111",
  15213=>"110000000",
  15214=>"000000000",
  15215=>"000000000",
  15216=>"000100000",
  15217=>"110110110",
  15218=>"110100000",
  15219=>"111111111",
  15220=>"010111110",
  15221=>"000100110",
  15222=>"100111001",
  15223=>"000001000",
  15224=>"000000000",
  15225=>"111011000",
  15226=>"001001011",
  15227=>"010110111",
  15228=>"000000001",
  15229=>"000001001",
  15230=>"000011001",
  15231=>"000000000",
  15232=>"011001001",
  15233=>"111111111",
  15234=>"000000001",
  15235=>"000111111",
  15236=>"000000000",
  15237=>"100100100",
  15238=>"000000011",
  15239=>"000001000",
  15240=>"101111111",
  15241=>"100100110",
  15242=>"100100101",
  15243=>"000000111",
  15244=>"100110100",
  15245=>"000000001",
  15246=>"000000100",
  15247=>"111111011",
  15248=>"000100100",
  15249=>"111111111",
  15250=>"100000000",
  15251=>"000000001",
  15252=>"011111111",
  15253=>"000000000",
  15254=>"100000001",
  15255=>"101001001",
  15256=>"001111100",
  15257=>"010010011",
  15258=>"111110111",
  15259=>"100100111",
  15260=>"000000000",
  15261=>"000000111",
  15262=>"111111111",
  15263=>"000011011",
  15264=>"000000000",
  15265=>"010000000",
  15266=>"001111011",
  15267=>"000000000",
  15268=>"000000000",
  15269=>"000000000",
  15270=>"000000000",
  15271=>"111011000",
  15272=>"000000000",
  15273=>"101001000",
  15274=>"100100000",
  15275=>"111000000",
  15276=>"111111111",
  15277=>"000001000",
  15278=>"000000000",
  15279=>"000111111",
  15280=>"011111111",
  15281=>"000000000",
  15282=>"000000001",
  15283=>"000000001",
  15284=>"111111010",
  15285=>"111111111",
  15286=>"000100111",
  15287=>"100110010",
  15288=>"000000000",
  15289=>"000100000",
  15290=>"100111001",
  15291=>"000000100",
  15292=>"011011001",
  15293=>"100001001",
  15294=>"111111111",
  15295=>"101101111",
  15296=>"100111110",
  15297=>"000000000",
  15298=>"000000000",
  15299=>"001000000",
  15300=>"111111111",
  15301=>"000000001",
  15302=>"100100110",
  15303=>"111000000",
  15304=>"000000000",
  15305=>"111111001",
  15306=>"000000000",
  15307=>"111111000",
  15308=>"111111111",
  15309=>"101000000",
  15310=>"011100111",
  15311=>"111111111",
  15312=>"000011011",
  15313=>"001001000",
  15314=>"000000000",
  15315=>"100111111",
  15316=>"000001111",
  15317=>"100110000",
  15318=>"011111111",
  15319=>"100000000",
  15320=>"000000111",
  15321=>"011001011",
  15322=>"100101000",
  15323=>"100111111",
  15324=>"000000000",
  15325=>"000100111",
  15326=>"111111100",
  15327=>"001000000",
  15328=>"111111111",
  15329=>"000000000",
  15330=>"100001001",
  15331=>"101100100",
  15332=>"000000011",
  15333=>"100000000",
  15334=>"101111111",
  15335=>"000000000",
  15336=>"000000100",
  15337=>"000111000",
  15338=>"100000000",
  15339=>"101111110",
  15340=>"000000000",
  15341=>"100000000",
  15342=>"100000111",
  15343=>"111011001",
  15344=>"011011111",
  15345=>"111111111",
  15346=>"111001000",
  15347=>"111111111",
  15348=>"111111111",
  15349=>"000000000",
  15350=>"001001000",
  15351=>"110000010",
  15352=>"000100110",
  15353=>"111111111",
  15354=>"000000100",
  15355=>"000000111",
  15356=>"000011111",
  15357=>"011010000",
  15358=>"111111110",
  15359=>"111011111",
  15360=>"010110111",
  15361=>"111111111",
  15362=>"100000000",
  15363=>"101100100",
  15364=>"011101111",
  15365=>"000000010",
  15366=>"000011011",
  15367=>"000000000",
  15368=>"000000000",
  15369=>"000000000",
  15370=>"000000000",
  15371=>"111111101",
  15372=>"110110110",
  15373=>"000000000",
  15374=>"000000000",
  15375=>"000000000",
  15376=>"000101001",
  15377=>"000000111",
  15378=>"111111111",
  15379=>"110111111",
  15380=>"000000101",
  15381=>"111000000",
  15382=>"000000001",
  15383=>"100100111",
  15384=>"110000000",
  15385=>"011111011",
  15386=>"111001001",
  15387=>"111111111",
  15388=>"000000000",
  15389=>"111110000",
  15390=>"111111111",
  15391=>"000000000",
  15392=>"111000000",
  15393=>"000000001",
  15394=>"000001111",
  15395=>"111111111",
  15396=>"000000000",
  15397=>"000000100",
  15398=>"111111111",
  15399=>"111010111",
  15400=>"000000100",
  15401=>"000000000",
  15402=>"000000000",
  15403=>"000000100",
  15404=>"001010010",
  15405=>"100000000",
  15406=>"111100000",
  15407=>"100000111",
  15408=>"011111111",
  15409=>"010111111",
  15410=>"000000011",
  15411=>"100000001",
  15412=>"110010000",
  15413=>"111111110",
  15414=>"001001000",
  15415=>"011001000",
  15416=>"000101111",
  15417=>"000000111",
  15418=>"100100111",
  15419=>"111111100",
  15420=>"111101000",
  15421=>"111101001",
  15422=>"111100111",
  15423=>"111111101",
  15424=>"000000000",
  15425=>"100111111",
  15426=>"000001011",
  15427=>"001011000",
  15428=>"000100000",
  15429=>"110110111",
  15430=>"111010010",
  15431=>"111010000",
  15432=>"011011001",
  15433=>"111111111",
  15434=>"111111111",
  15435=>"111111000",
  15436=>"111111001",
  15437=>"000000000",
  15438=>"000000100",
  15439=>"000100111",
  15440=>"001000000",
  15441=>"000000110",
  15442=>"111111111",
  15443=>"000000000",
  15444=>"000111111",
  15445=>"111111111",
  15446=>"111110110",
  15447=>"111111111",
  15448=>"001001001",
  15449=>"111111001",
  15450=>"111011001",
  15451=>"000000000",
  15452=>"100000001",
  15453=>"000000000",
  15454=>"111111111",
  15455=>"000000010",
  15456=>"111000000",
  15457=>"110111011",
  15458=>"111111111",
  15459=>"010110001",
  15460=>"011111111",
  15461=>"111000000",
  15462=>"000100111",
  15463=>"000000000",
  15464=>"000000000",
  15465=>"111111111",
  15466=>"100001001",
  15467=>"111111111",
  15468=>"001111111",
  15469=>"000000000",
  15470=>"000000000",
  15471=>"000000000",
  15472=>"111111111",
  15473=>"000000000",
  15474=>"010010000",
  15475=>"100100111",
  15476=>"000000000",
  15477=>"001000000",
  15478=>"111110111",
  15479=>"000000000",
  15480=>"000001001",
  15481=>"000111111",
  15482=>"111001011",
  15483=>"100111111",
  15484=>"110110100",
  15485=>"000000000",
  15486=>"000000000",
  15487=>"000000000",
  15488=>"000000000",
  15489=>"000000000",
  15490=>"111000000",
  15491=>"100000000",
  15492=>"000000000",
  15493=>"111111000",
  15494=>"111111111",
  15495=>"011000000",
  15496=>"000000000",
  15497=>"011011010",
  15498=>"000000000",
  15499=>"111111101",
  15500=>"111111111",
  15501=>"000000000",
  15502=>"001001000",
  15503=>"111111111",
  15504=>"000000000",
  15505=>"000000000",
  15506=>"000111111",
  15507=>"111111011",
  15508=>"000000000",
  15509=>"001001111",
  15510=>"100111111",
  15511=>"000000000",
  15512=>"111111111",
  15513=>"111111111",
  15514=>"000000100",
  15515=>"111111011",
  15516=>"100000000",
  15517=>"000000000",
  15518=>"001000100",
  15519=>"000001101",
  15520=>"110000000",
  15521=>"000011000",
  15522=>"000010001",
  15523=>"001001001",
  15524=>"110010110",
  15525=>"110111111",
  15526=>"111111000",
  15527=>"000000001",
  15528=>"111111011",
  15529=>"000000001",
  15530=>"100101111",
  15531=>"000000000",
  15532=>"111011111",
  15533=>"111011111",
  15534=>"111111111",
  15535=>"110001000",
  15536=>"111111111",
  15537=>"001000000",
  15538=>"111111110",
  15539=>"111111000",
  15540=>"000100111",
  15541=>"011110100",
  15542=>"000000000",
  15543=>"111111111",
  15544=>"111111111",
  15545=>"000001000",
  15546=>"011011011",
  15547=>"111011000",
  15548=>"111111111",
  15549=>"000101100",
  15550=>"001001111",
  15551=>"110111111",
  15552=>"111011011",
  15553=>"000000000",
  15554=>"111111101",
  15555=>"000000011",
  15556=>"111111000",
  15557=>"000000111",
  15558=>"001011001",
  15559=>"111011001",
  15560=>"100111000",
  15561=>"000000000",
  15562=>"111111001",
  15563=>"000000111",
  15564=>"111111111",
  15565=>"111111111",
  15566=>"111011000",
  15567=>"100100000",
  15568=>"011000110",
  15569=>"110000000",
  15570=>"111100110",
  15571=>"000000000",
  15572=>"001000111",
  15573=>"110110110",
  15574=>"010110010",
  15575=>"111111111",
  15576=>"111111111",
  15577=>"111111111",
  15578=>"111100000",
  15579=>"111111111",
  15580=>"001001001",
  15581=>"111111111",
  15582=>"000000000",
  15583=>"001001011",
  15584=>"000000111",
  15585=>"110000000",
  15586=>"000000000",
  15587=>"111111111",
  15588=>"000011111",
  15589=>"100000000",
  15590=>"111111111",
  15591=>"000000000",
  15592=>"000000110",
  15593=>"000000000",
  15594=>"000000000",
  15595=>"100110111",
  15596=>"111111000",
  15597=>"110110110",
  15598=>"000110111",
  15599=>"111111111",
  15600=>"000000000",
  15601=>"111111111",
  15602=>"111111111",
  15603=>"000010000",
  15604=>"111001000",
  15605=>"000000000",
  15606=>"011000000",
  15607=>"110110000",
  15608=>"111111111",
  15609=>"111111111",
  15610=>"011011010",
  15611=>"110111110",
  15612=>"000111111",
  15613=>"000000100",
  15614=>"000000001",
  15615=>"000000000",
  15616=>"011001111",
  15617=>"011011111",
  15618=>"000000000",
  15619=>"000000000",
  15620=>"001001000",
  15621=>"000000000",
  15622=>"110111100",
  15623=>"110000101",
  15624=>"000000001",
  15625=>"000100000",
  15626=>"101111111",
  15627=>"111111111",
  15628=>"110000000",
  15629=>"111000000",
  15630=>"000000000",
  15631=>"110111111",
  15632=>"000100111",
  15633=>"101000000",
  15634=>"111111111",
  15635=>"100111101",
  15636=>"001111111",
  15637=>"110111000",
  15638=>"111110110",
  15639=>"000000000",
  15640=>"111111111",
  15641=>"111111111",
  15642=>"111111111",
  15643=>"000110110",
  15644=>"000000000",
  15645=>"111111111",
  15646=>"000000000",
  15647=>"000000000",
  15648=>"000000001",
  15649=>"111111111",
  15650=>"111000000",
  15651=>"111111111",
  15652=>"001000000",
  15653=>"111101101",
  15654=>"011000000",
  15655=>"000000100",
  15656=>"000001000",
  15657=>"000000000",
  15658=>"000000011",
  15659=>"111100000",
  15660=>"111000000",
  15661=>"011000000",
  15662=>"111101000",
  15663=>"111111011",
  15664=>"000000000",
  15665=>"000000000",
  15666=>"011111111",
  15667=>"111111111",
  15668=>"111100000",
  15669=>"000110110",
  15670=>"011101101",
  15671=>"111000000",
  15672=>"000000000",
  15673=>"001000000",
  15674=>"111101100",
  15675=>"100110110",
  15676=>"110111111",
  15677=>"111001000",
  15678=>"010110000",
  15679=>"111011000",
  15680=>"000000000",
  15681=>"001000100",
  15682=>"000000000",
  15683=>"111111111",
  15684=>"011010110",
  15685=>"100100100",
  15686=>"000000110",
  15687=>"000100000",
  15688=>"000000000",
  15689=>"001000000",
  15690=>"000000010",
  15691=>"100100100",
  15692=>"001101111",
  15693=>"001101111",
  15694=>"001001000",
  15695=>"111111111",
  15696=>"000000000",
  15697=>"100100100",
  15698=>"000000000",
  15699=>"000000000",
  15700=>"000000000",
  15701=>"011011001",
  15702=>"111100000",
  15703=>"000000000",
  15704=>"111111000",
  15705=>"101101101",
  15706=>"111111111",
  15707=>"101111100",
  15708=>"100000010",
  15709=>"000000000",
  15710=>"000000100",
  15711=>"011111110",
  15712=>"000000001",
  15713=>"111100111",
  15714=>"001111111",
  15715=>"111111111",
  15716=>"111111001",
  15717=>"000111111",
  15718=>"000000000",
  15719=>"111101100",
  15720=>"011000001",
  15721=>"000000000",
  15722=>"100000110",
  15723=>"000000000",
  15724=>"110010010",
  15725=>"000111111",
  15726=>"000111111",
  15727=>"010010000",
  15728=>"111111111",
  15729=>"111001010",
  15730=>"111111101",
  15731=>"000011011",
  15732=>"111111111",
  15733=>"000000000",
  15734=>"001000110",
  15735=>"000000000",
  15736=>"111111111",
  15737=>"000100111",
  15738=>"000000000",
  15739=>"111111111",
  15740=>"000000000",
  15741=>"111111111",
  15742=>"100111101",
  15743=>"111111111",
  15744=>"000001001",
  15745=>"111001101",
  15746=>"111111001",
  15747=>"110111110",
  15748=>"100111111",
  15749=>"011111111",
  15750=>"100000000",
  15751=>"000111111",
  15752=>"000000000",
  15753=>"000000001",
  15754=>"111111011",
  15755=>"000000000",
  15756=>"001111111",
  15757=>"001001111",
  15758=>"111111110",
  15759=>"110100000",
  15760=>"000000000",
  15761=>"101000000",
  15762=>"110010000",
  15763=>"011011111",
  15764=>"001000000",
  15765=>"000000000",
  15766=>"111111101",
  15767=>"010000000",
  15768=>"000000000",
  15769=>"101111111",
  15770=>"111111111",
  15771=>"100000000",
  15772=>"110110000",
  15773=>"000000000",
  15774=>"001001011",
  15775=>"100000000",
  15776=>"111111111",
  15777=>"110000000",
  15778=>"001001000",
  15779=>"111111111",
  15780=>"000000001",
  15781=>"000010010",
  15782=>"001001000",
  15783=>"000000000",
  15784=>"111111111",
  15785=>"111111111",
  15786=>"111111111",
  15787=>"111111111",
  15788=>"111111111",
  15789=>"111000000",
  15790=>"011000000",
  15791=>"111111011",
  15792=>"101011001",
  15793=>"111111111",
  15794=>"100000000",
  15795=>"111111111",
  15796=>"000000000",
  15797=>"111111111",
  15798=>"111111111",
  15799=>"000101111",
  15800=>"010101111",
  15801=>"000000000",
  15802=>"011111111",
  15803=>"000000000",
  15804=>"111111011",
  15805=>"111111111",
  15806=>"111111111",
  15807=>"111101100",
  15808=>"101111111",
  15809=>"011111111",
  15810=>"000000000",
  15811=>"000000000",
  15812=>"011010001",
  15813=>"000111111",
  15814=>"111011000",
  15815=>"000111111",
  15816=>"000000000",
  15817=>"111011000",
  15818=>"001001111",
  15819=>"111111111",
  15820=>"111111111",
  15821=>"110110000",
  15822=>"111111111",
  15823=>"100110110",
  15824=>"000000000",
  15825=>"111100000",
  15826=>"111111101",
  15827=>"111100000",
  15828=>"111111111",
  15829=>"111111111",
  15830=>"111111000",
  15831=>"000000100",
  15832=>"001001111",
  15833=>"101111110",
  15834=>"111110010",
  15835=>"011001001",
  15836=>"000000000",
  15837=>"111100100",
  15838=>"000000000",
  15839=>"011011111",
  15840=>"000000000",
  15841=>"000011011",
  15842=>"111111001",
  15843=>"111111111",
  15844=>"100111111",
  15845=>"111111111",
  15846=>"110000000",
  15847=>"111111111",
  15848=>"000001000",
  15849=>"000000000",
  15850=>"011000000",
  15851=>"000000001",
  15852=>"111111101",
  15853=>"000000000",
  15854=>"100100101",
  15855=>"000111111",
  15856=>"000000011",
  15857=>"000000000",
  15858=>"001101111",
  15859=>"100111111",
  15860=>"111111111",
  15861=>"000000111",
  15862=>"000001000",
  15863=>"000000000",
  15864=>"000011011",
  15865=>"111111111",
  15866=>"000000000",
  15867=>"111111111",
  15868=>"000000000",
  15869=>"111000000",
  15870=>"100001001",
  15871=>"000000010",
  15872=>"100100100",
  15873=>"100100100",
  15874=>"111111111",
  15875=>"000000011",
  15876=>"000110100",
  15877=>"001011111",
  15878=>"111111111",
  15879=>"001000101",
  15880=>"100111110",
  15881=>"111101111",
  15882=>"000001000",
  15883=>"001001001",
  15884=>"000111111",
  15885=>"000001111",
  15886=>"000111011",
  15887=>"111100000",
  15888=>"000100100",
  15889=>"000110001",
  15890=>"000000000",
  15891=>"000000000",
  15892=>"000000000",
  15893=>"000000110",
  15894=>"111111111",
  15895=>"001011011",
  15896=>"111111101",
  15897=>"111111100",
  15898=>"001001000",
  15899=>"111110110",
  15900=>"000000110",
  15901=>"111111111",
  15902=>"110110111",
  15903=>"000000100",
  15904=>"000000011",
  15905=>"000000000",
  15906=>"100000000",
  15907=>"001000111",
  15908=>"000000000",
  15909=>"111111000",
  15910=>"000110110",
  15911=>"000000010",
  15912=>"001011111",
  15913=>"110111111",
  15914=>"111100111",
  15915=>"111111100",
  15916=>"010110000",
  15917=>"111111001",
  15918=>"000000111",
  15919=>"000000110",
  15920=>"000000001",
  15921=>"111000000",
  15922=>"000000001",
  15923=>"100100000",
  15924=>"111110111",
  15925=>"000001011",
  15926=>"000010000",
  15927=>"101000111",
  15928=>"000000011",
  15929=>"111111111",
  15930=>"101000000",
  15931=>"110101100",
  15932=>"000001111",
  15933=>"100000000",
  15934=>"000000001",
  15935=>"001001111",
  15936=>"111101000",
  15937=>"100000000",
  15938=>"000000111",
  15939=>"111110100",
  15940=>"000000111",
  15941=>"011111111",
  15942=>"111111101",
  15943=>"000000000",
  15944=>"111111001",
  15945=>"111101111",
  15946=>"111110000",
  15947=>"001111111",
  15948=>"111111000",
  15949=>"001011001",
  15950=>"111100000",
  15951=>"000000000",
  15952=>"111111111",
  15953=>"110111111",
  15954=>"111111111",
  15955=>"000000100",
  15956=>"111111111",
  15957=>"000000000",
  15958=>"100101111",
  15959=>"010000011",
  15960=>"011011110",
  15961=>"000000000",
  15962=>"000000000",
  15963=>"111011011",
  15964=>"011001001",
  15965=>"000000000",
  15966=>"111111100",
  15967=>"111110000",
  15968=>"000000000",
  15969=>"111111011",
  15970=>"000000000",
  15971=>"000000111",
  15972=>"011001011",
  15973=>"100000111",
  15974=>"011001111",
  15975=>"000001001",
  15976=>"001000000",
  15977=>"111111011",
  15978=>"001000000",
  15979=>"010000111",
  15980=>"000000000",
  15981=>"000000111",
  15982=>"011000000",
  15983=>"000000000",
  15984=>"010000000",
  15985=>"111111111",
  15986=>"000010010",
  15987=>"000000000",
  15988=>"000000000",
  15989=>"001000001",
  15990=>"000001001",
  15991=>"000000000",
  15992=>"111111111",
  15993=>"111111011",
  15994=>"000010011",
  15995=>"000111011",
  15996=>"111111111",
  15997=>"011011011",
  15998=>"000000000",
  15999=>"000011111",
  16000=>"111111111",
  16001=>"000000000",
  16002=>"000000000",
  16003=>"101101110",
  16004=>"000000000",
  16005=>"010000000",
  16006=>"111110100",
  16007=>"000000100",
  16008=>"111010000",
  16009=>"110111111",
  16010=>"000011111",
  16011=>"111000111",
  16012=>"000000000",
  16013=>"111111110",
  16014=>"111111110",
  16015=>"111111111",
  16016=>"001000000",
  16017=>"000000000",
  16018=>"000110000",
  16019=>"101111110",
  16020=>"111001001",
  16021=>"000000000",
  16022=>"010000000",
  16023=>"000000000",
  16024=>"001000000",
  16025=>"101000111",
  16026=>"010000101",
  16027=>"101111101",
  16028=>"000000000",
  16029=>"111001111",
  16030=>"111011011",
  16031=>"111111000",
  16032=>"000101001",
  16033=>"111100001",
  16034=>"111111000",
  16035=>"101100111",
  16036=>"000000010",
  16037=>"111111101",
  16038=>"000111111",
  16039=>"111111111",
  16040=>"000000000",
  16041=>"111111111",
  16042=>"000000000",
  16043=>"111111111",
  16044=>"000000000",
  16045=>"000001111",
  16046=>"000000000",
  16047=>"000111111",
  16048=>"000000000",
  16049=>"111110000",
  16050=>"010111110",
  16051=>"011011000",
  16052=>"111011010",
  16053=>"000000000",
  16054=>"111011011",
  16055=>"111111111",
  16056=>"111111111",
  16057=>"010000111",
  16058=>"011000000",
  16059=>"001001111",
  16060=>"000000100",
  16061=>"001111000",
  16062=>"111110000",
  16063=>"111111101",
  16064=>"111111111",
  16065=>"001001111",
  16066=>"111111010",
  16067=>"111111000",
  16068=>"011011111",
  16069=>"000000101",
  16070=>"010000011",
  16071=>"000000110",
  16072=>"000110111",
  16073=>"000000011",
  16074=>"000000001",
  16075=>"001110111",
  16076=>"111111101",
  16077=>"111011000",
  16078=>"100000000",
  16079=>"000000011",
  16080=>"000010000",
  16081=>"000011111",
  16082=>"000000101",
  16083=>"000000000",
  16084=>"111000000",
  16085=>"111101001",
  16086=>"011010011",
  16087=>"111111110",
  16088=>"111100000",
  16089=>"111111111",
  16090=>"111000100",
  16091=>"001000001",
  16092=>"110111111",
  16093=>"000000010",
  16094=>"001111000",
  16095=>"001010010",
  16096=>"111111111",
  16097=>"000000000",
  16098=>"000001111",
  16099=>"100100000",
  16100=>"111011000",
  16101=>"110110100",
  16102=>"011111111",
  16103=>"000000101",
  16104=>"111100111",
  16105=>"111000000",
  16106=>"000110111",
  16107=>"000000000",
  16108=>"000000100",
  16109=>"000000001",
  16110=>"000001111",
  16111=>"011111000",
  16112=>"100111111",
  16113=>"111111000",
  16114=>"000000000",
  16115=>"000000001",
  16116=>"111111000",
  16117=>"110100100",
  16118=>"000100000",
  16119=>"111111111",
  16120=>"001000000",
  16121=>"000000001",
  16122=>"101001000",
  16123=>"111001000",
  16124=>"000000111",
  16125=>"001001000",
  16126=>"010010111",
  16127=>"110100101",
  16128=>"011001111",
  16129=>"111110110",
  16130=>"000000100",
  16131=>"111111000",
  16132=>"000000100",
  16133=>"111101001",
  16134=>"000000000",
  16135=>"111000000",
  16136=>"000000110",
  16137=>"000000100",
  16138=>"100100100",
  16139=>"111111111",
  16140=>"110100111",
  16141=>"000000011",
  16142=>"111111111",
  16143=>"000011111",
  16144=>"100001000",
  16145=>"000000000",
  16146=>"000000111",
  16147=>"101000000",
  16148=>"010010111",
  16149=>"100100000",
  16150=>"110110110",
  16151=>"011011111",
  16152=>"111111000",
  16153=>"000000001",
  16154=>"000000000",
  16155=>"000000000",
  16156=>"101011111",
  16157=>"110000000",
  16158=>"001000000",
  16159=>"100110000",
  16160=>"111011001",
  16161=>"111111111",
  16162=>"111111011",
  16163=>"000000111",
  16164=>"111100110",
  16165=>"000011011",
  16166=>"111111111",
  16167=>"000110111",
  16168=>"111111111",
  16169=>"011000000",
  16170=>"001000000",
  16171=>"000010011",
  16172=>"011010010",
  16173=>"100110111",
  16174=>"111111000",
  16175=>"111011000",
  16176=>"001011111",
  16177=>"010111111",
  16178=>"001001011",
  16179=>"000000001",
  16180=>"000000000",
  16181=>"000000111",
  16182=>"000111011",
  16183=>"111111111",
  16184=>"000000000",
  16185=>"000000011",
  16186=>"111010000",
  16187=>"000000101",
  16188=>"111001001",
  16189=>"001000110",
  16190=>"111111000",
  16191=>"111111001",
  16192=>"111111111",
  16193=>"111011000",
  16194=>"111111111",
  16195=>"011111111",
  16196=>"110100110",
  16197=>"100110000",
  16198=>"000110011",
  16199=>"000111111",
  16200=>"000000000",
  16201=>"010000000",
  16202=>"111111000",
  16203=>"011111110",
  16204=>"000000000",
  16205=>"001011111",
  16206=>"111111111",
  16207=>"000000100",
  16208=>"000001111",
  16209=>"001001000",
  16210=>"111111110",
  16211=>"001011011",
  16212=>"000110110",
  16213=>"011000000",
  16214=>"000101111",
  16215=>"000000000",
  16216=>"101001111",
  16217=>"001000000",
  16218=>"101001000",
  16219=>"000100110",
  16220=>"001101101",
  16221=>"111011000",
  16222=>"000000111",
  16223=>"001001000",
  16224=>"111111111",
  16225=>"001001000",
  16226=>"101001011",
  16227=>"111001000",
  16228=>"011111011",
  16229=>"111111111",
  16230=>"000101100",
  16231=>"001001001",
  16232=>"110110111",
  16233=>"101000000",
  16234=>"111111111",
  16235=>"001001101",
  16236=>"110111111",
  16237=>"000000110",
  16238=>"001001000",
  16239=>"100000000",
  16240=>"000000111",
  16241=>"111111011",
  16242=>"000000111",
  16243=>"110110000",
  16244=>"000000100",
  16245=>"000000100",
  16246=>"000000100",
  16247=>"001110100",
  16248=>"000011111",
  16249=>"000000000",
  16250=>"011011111",
  16251=>"011011111",
  16252=>"000000000",
  16253=>"001011111",
  16254=>"000001011",
  16255=>"111000000",
  16256=>"100111111",
  16257=>"000101111",
  16258=>"000110110",
  16259=>"111101000",
  16260=>"000110111",
  16261=>"111100110",
  16262=>"000111111",
  16263=>"001011111",
  16264=>"111111111",
  16265=>"000110110",
  16266=>"111110100",
  16267=>"111111111",
  16268=>"111111111",
  16269=>"100000001",
  16270=>"101000111",
  16271=>"111111010",
  16272=>"000000111",
  16273=>"000111111",
  16274=>"111111111",
  16275=>"011000000",
  16276=>"000000111",
  16277=>"011111111",
  16278=>"000000000",
  16279=>"000011111",
  16280=>"111000101",
  16281=>"111111111",
  16282=>"011001001",
  16283=>"011000000",
  16284=>"111111010",
  16285=>"000000011",
  16286=>"111011011",
  16287=>"110111111",
  16288=>"011111011",
  16289=>"011011011",
  16290=>"100101111",
  16291=>"000000001",
  16292=>"101001001",
  16293=>"111111111",
  16294=>"111000001",
  16295=>"111111110",
  16296=>"100000100",
  16297=>"011111111",
  16298=>"101111000",
  16299=>"101001000",
  16300=>"111111111",
  16301=>"001001000",
  16302=>"111111111",
  16303=>"111000000",
  16304=>"000000000",
  16305=>"111010000",
  16306=>"111111111",
  16307=>"000000000",
  16308=>"101100000",
  16309=>"000000011",
  16310=>"111100000",
  16311=>"000000010",
  16312=>"111111111",
  16313=>"000000000",
  16314=>"000000001",
  16315=>"011011001",
  16316=>"000000111",
  16317=>"110000000",
  16318=>"111111100",
  16319=>"000000001",
  16320=>"111001000",
  16321=>"111111111",
  16322=>"000000000",
  16323=>"000001111",
  16324=>"110010111",
  16325=>"001000001",
  16326=>"001111111",
  16327=>"011001000",
  16328=>"011000100",
  16329=>"111111111",
  16330=>"001011111",
  16331=>"101100010",
  16332=>"111011000",
  16333=>"000100111",
  16334=>"011111100",
  16335=>"111110011",
  16336=>"001000111",
  16337=>"111111000",
  16338=>"111110110",
  16339=>"110000000",
  16340=>"000001001",
  16341=>"111111111",
  16342=>"001001011",
  16343=>"100101111",
  16344=>"111111111",
  16345=>"011111011",
  16346=>"111111000",
  16347=>"000000110",
  16348=>"111010000",
  16349=>"000000000",
  16350=>"111010111",
  16351=>"000000000",
  16352=>"011101111",
  16353=>"110000000",
  16354=>"011110111",
  16355=>"111111101",
  16356=>"000001001",
  16357=>"001001000",
  16358=>"111111111",
  16359=>"000000110",
  16360=>"011111011",
  16361=>"000101101",
  16362=>"000001011",
  16363=>"111111100",
  16364=>"000001001",
  16365=>"000100100",
  16366=>"101101111",
  16367=>"000000100",
  16368=>"011001000",
  16369=>"000011011",
  16370=>"100110111",
  16371=>"111000001",
  16372=>"000000000",
  16373=>"000010000",
  16374=>"110111111",
  16375=>"010010111",
  16376=>"000000111",
  16377=>"001000000",
  16378=>"010110110",
  16379=>"111111110",
  16380=>"001000111",
  16381=>"100101111",
  16382=>"000001111",
  16383=>"011010110",
  16384=>"001001000",
  16385=>"000000011",
  16386=>"000000101",
  16387=>"111001001",
  16388=>"010010001",
  16389=>"000000000",
  16390=>"000000010",
  16391=>"100111110",
  16392=>"111111111",
  16393=>"011001001",
  16394=>"110100101",
  16395=>"110011001",
  16396=>"100000101",
  16397=>"111111111",
  16398=>"111111111",
  16399=>"011000111",
  16400=>"111111111",
  16401=>"111111000",
  16402=>"000000101",
  16403=>"000000000",
  16404=>"000000000",
  16405=>"001100000",
  16406=>"100111101",
  16407=>"110100111",
  16408=>"001000000",
  16409=>"011001000",
  16410=>"111111111",
  16411=>"111101011",
  16412=>"000000111",
  16413=>"111110100",
  16414=>"111111111",
  16415=>"001011111",
  16416=>"000000000",
  16417=>"111101000",
  16418=>"001001001",
  16419=>"111111111",
  16420=>"000000100",
  16421=>"100100110",
  16422=>"000000000",
  16423=>"001111111",
  16424=>"100000111",
  16425=>"000001011",
  16426=>"001000000",
  16427=>"111111111",
  16428=>"000000100",
  16429=>"011110000",
  16430=>"111110111",
  16431=>"001001111",
  16432=>"000000101",
  16433=>"000000100",
  16434=>"000000100",
  16435=>"000000000",
  16436=>"101101101",
  16437=>"110110100",
  16438=>"010000000",
  16439=>"000000000",
  16440=>"111111111",
  16441=>"000001111",
  16442=>"111111111",
  16443=>"111000000",
  16444=>"000000100",
  16445=>"000000000",
  16446=>"101111111",
  16447=>"000000000",
  16448=>"111111111",
  16449=>"001001100",
  16450=>"110110111",
  16451=>"011111111",
  16452=>"000000000",
  16453=>"111110111",
  16454=>"110100111",
  16455=>"110000000",
  16456=>"111111111",
  16457=>"111111111",
  16458=>"000000100",
  16459=>"000110100",
  16460=>"111001000",
  16461=>"011000000",
  16462=>"011001011",
  16463=>"110111111",
  16464=>"000001011",
  16465=>"010000000",
  16466=>"000000000",
  16467=>"111111111",
  16468=>"000000000",
  16469=>"010010000",
  16470=>"000011011",
  16471=>"000000000",
  16472=>"011111111",
  16473=>"111100100",
  16474=>"110111101",
  16475=>"001011101",
  16476=>"000000010",
  16477=>"111111111",
  16478=>"001001111",
  16479=>"111001000",
  16480=>"101000001",
  16481=>"000001000",
  16482=>"110110100",
  16483=>"000000111",
  16484=>"111111110",
  16485=>"000000000",
  16486=>"011111100",
  16487=>"111111111",
  16488=>"111100101",
  16489=>"000001010",
  16490=>"000011000",
  16491=>"111111100",
  16492=>"000110110",
  16493=>"000000011",
  16494=>"000000000",
  16495=>"111111100",
  16496=>"111011001",
  16497=>"111111111",
  16498=>"101101101",
  16499=>"111111111",
  16500=>"111111101",
  16501=>"010110000",
  16502=>"000001000",
  16503=>"011011000",
  16504=>"100111100",
  16505=>"110101000",
  16506=>"111110111",
  16507=>"111011000",
  16508=>"100100100",
  16509=>"111101111",
  16510=>"111111111",
  16511=>"010000000",
  16512=>"000000000",
  16513=>"011101000",
  16514=>"111111101",
  16515=>"111111111",
  16516=>"000001111",
  16517=>"000000100",
  16518=>"111111010",
  16519=>"100100111",
  16520=>"100000000",
  16521=>"111111111",
  16522=>"000101111",
  16523=>"000000000",
  16524=>"000000010",
  16525=>"001011101",
  16526=>"111111110",
  16527=>"111111111",
  16528=>"000000100",
  16529=>"000000000",
  16530=>"001111001",
  16531=>"000000011",
  16532=>"001000000",
  16533=>"111000010",
  16534=>"000000100",
  16535=>"100100100",
  16536=>"001001000",
  16537=>"111011000",
  16538=>"111110010",
  16539=>"111111111",
  16540=>"000000000",
  16541=>"011000000",
  16542=>"001011000",
  16543=>"111000010",
  16544=>"111110110",
  16545=>"000000000",
  16546=>"010000100",
  16547=>"111111111",
  16548=>"110110011",
  16549=>"001001111",
  16550=>"000000101",
  16551=>"011011011",
  16552=>"011111011",
  16553=>"111011111",
  16554=>"000000000",
  16555=>"010010100",
  16556=>"000000000",
  16557=>"000000100",
  16558=>"110111010",
  16559=>"110100100",
  16560=>"000000000",
  16561=>"110010110",
  16562=>"000100000",
  16563=>"000000000",
  16564=>"111111011",
  16565=>"000100000",
  16566=>"100000000",
  16567=>"111011111",
  16568=>"111010000",
  16569=>"101001111",
  16570=>"111110100",
  16571=>"101101101",
  16572=>"000000000",
  16573=>"001001000",
  16574=>"001000000",
  16575=>"111110000",
  16576=>"111000000",
  16577=>"000000000",
  16578=>"111110100",
  16579=>"000000010",
  16580=>"000000101",
  16581=>"000000000",
  16582=>"110000001",
  16583=>"101101001",
  16584=>"000000011",
  16585=>"111010010",
  16586=>"111111000",
  16587=>"110000000",
  16588=>"111011000",
  16589=>"001111110",
  16590=>"111111111",
  16591=>"000000000",
  16592=>"111100101",
  16593=>"111101101",
  16594=>"000100111",
  16595=>"111111111",
  16596=>"111111110",
  16597=>"100110111",
  16598=>"111000000",
  16599=>"011101000",
  16600=>"000000000",
  16601=>"000000000",
  16602=>"000000000",
  16603=>"000001000",
  16604=>"001100000",
  16605=>"100000000",
  16606=>"000000000",
  16607=>"000000000",
  16608=>"001111111",
  16609=>"000000000",
  16610=>"000110110",
  16611=>"000001111",
  16612=>"000000000",
  16613=>"111111100",
  16614=>"111101111",
  16615=>"111110110",
  16616=>"000000010",
  16617=>"000111111",
  16618=>"111011010",
  16619=>"000000000",
  16620=>"000000100",
  16621=>"110111111",
  16622=>"000101111",
  16623=>"000000111",
  16624=>"111110011",
  16625=>"000000000",
  16626=>"110111111",
  16627=>"000100001",
  16628=>"111111111",
  16629=>"111011000",
  16630=>"001000000",
  16631=>"000000000",
  16632=>"111111100",
  16633=>"000000000",
  16634=>"000000101",
  16635=>"111111101",
  16636=>"000100000",
  16637=>"000000111",
  16638=>"000001111",
  16639=>"111110000",
  16640=>"111001111",
  16641=>"110111111",
  16642=>"111111111",
  16643=>"001011011",
  16644=>"000000000",
  16645=>"010010110",
  16646=>"000000000",
  16647=>"001011000",
  16648=>"000010110",
  16649=>"000000000",
  16650=>"111111111",
  16651=>"000000001",
  16652=>"000000000",
  16653=>"101111111",
  16654=>"010000001",
  16655=>"000100110",
  16656=>"000000000",
  16657=>"100110111",
  16658=>"111000000",
  16659=>"000000001",
  16660=>"000000011",
  16661=>"000000000",
  16662=>"001011111",
  16663=>"000000100",
  16664=>"111111111",
  16665=>"111111001",
  16666=>"111110000",
  16667=>"000000000",
  16668=>"111111111",
  16669=>"111101001",
  16670=>"000000000",
  16671=>"111111111",
  16672=>"001101101",
  16673=>"100100101",
  16674=>"111000101",
  16675=>"111111000",
  16676=>"100000000",
  16677=>"000000001",
  16678=>"000000000",
  16679=>"111011000",
  16680=>"000001011",
  16681=>"111111111",
  16682=>"000001001",
  16683=>"101111111",
  16684=>"111001000",
  16685=>"011110111",
  16686=>"000000101",
  16687=>"000000111",
  16688=>"111001000",
  16689=>"000000000",
  16690=>"110100111",
  16691=>"000000000",
  16692=>"111111111",
  16693=>"101001111",
  16694=>"000000110",
  16695=>"101101111",
  16696=>"000000000",
  16697=>"100000100",
  16698=>"111111000",
  16699=>"111011111",
  16700=>"111110110",
  16701=>"111111100",
  16702=>"000000010",
  16703=>"100000000",
  16704=>"001111111",
  16705=>"001000000",
  16706=>"101001001",
  16707=>"111111000",
  16708=>"000001101",
  16709=>"111111111",
  16710=>"000011011",
  16711=>"110111101",
  16712=>"000000000",
  16713=>"000000111",
  16714=>"000000111",
  16715=>"000101101",
  16716=>"100000000",
  16717=>"001001111",
  16718=>"110110111",
  16719=>"000000000",
  16720=>"111100100",
  16721=>"000111010",
  16722=>"111111001",
  16723=>"000000111",
  16724=>"100100111",
  16725=>"011011011",
  16726=>"000000101",
  16727=>"011001000",
  16728=>"111111111",
  16729=>"001001111",
  16730=>"111001111",
  16731=>"100000000",
  16732=>"000000000",
  16733=>"111111111",
  16734=>"000000000",
  16735=>"100100100",
  16736=>"000000000",
  16737=>"111100000",
  16738=>"100111111",
  16739=>"000100111",
  16740=>"100100110",
  16741=>"000001001",
  16742=>"000001010",
  16743=>"000000000",
  16744=>"100111111",
  16745=>"000000101",
  16746=>"000000000",
  16747=>"111111111",
  16748=>"110110000",
  16749=>"110110111",
  16750=>"111101101",
  16751=>"111111111",
  16752=>"000100110",
  16753=>"011011011",
  16754=>"000000001",
  16755=>"001011111",
  16756=>"000000010",
  16757=>"100000100",
  16758=>"001001000",
  16759=>"001001111",
  16760=>"011001100",
  16761=>"001111111",
  16762=>"000111110",
  16763=>"011111111",
  16764=>"000001011",
  16765=>"111111010",
  16766=>"000000000",
  16767=>"011000100",
  16768=>"110110100",
  16769=>"000000000",
  16770=>"111000000",
  16771=>"000000010",
  16772=>"001111111",
  16773=>"000000000",
  16774=>"001011011",
  16775=>"010010011",
  16776=>"111110100",
  16777=>"000000000",
  16778=>"000000000",
  16779=>"000000000",
  16780=>"101001111",
  16781=>"010011111",
  16782=>"110100100",
  16783=>"000000000",
  16784=>"000000000",
  16785=>"100100100",
  16786=>"111110100",
  16787=>"001001000",
  16788=>"111111000",
  16789=>"000000000",
  16790=>"100010000",
  16791=>"000011010",
  16792=>"111111100",
  16793=>"001011011",
  16794=>"111111001",
  16795=>"100100000",
  16796=>"001000110",
  16797=>"110111011",
  16798=>"000000000",
  16799=>"001011111",
  16800=>"000000000",
  16801=>"011010110",
  16802=>"101101110",
  16803=>"000001111",
  16804=>"000111111",
  16805=>"000000000",
  16806=>"111111111",
  16807=>"000111111",
  16808=>"111111111",
  16809=>"100100100",
  16810=>"000111111",
  16811=>"101111101",
  16812=>"000011011",
  16813=>"000001000",
  16814=>"000011011",
  16815=>"001000110",
  16816=>"110110000",
  16817=>"000000000",
  16818=>"001100100",
  16819=>"110111111",
  16820=>"111111111",
  16821=>"000000000",
  16822=>"100011100",
  16823=>"111001011",
  16824=>"001111111",
  16825=>"111111111",
  16826=>"000010111",
  16827=>"000010010",
  16828=>"001001001",
  16829=>"110000000",
  16830=>"100101110",
  16831=>"000101111",
  16832=>"000000111",
  16833=>"111111111",
  16834=>"111000000",
  16835=>"000000000",
  16836=>"011011000",
  16837=>"000000100",
  16838=>"001001100",
  16839=>"000000100",
  16840=>"110101111",
  16841=>"011000000",
  16842=>"011001000",
  16843=>"111111111",
  16844=>"111111111",
  16845=>"000111111",
  16846=>"111001101",
  16847=>"000000000",
  16848=>"000001111",
  16849=>"010100100",
  16850=>"000111111",
  16851=>"100100100",
  16852=>"000000000",
  16853=>"000010000",
  16854=>"000000000",
  16855=>"001000000",
  16856=>"110111110",
  16857=>"000000000",
  16858=>"111111111",
  16859=>"000000001",
  16860=>"000000011",
  16861=>"111110000",
  16862=>"100100100",
  16863=>"010010011",
  16864=>"101111111",
  16865=>"010110011",
  16866=>"111111110",
  16867=>"000001000",
  16868=>"111111111",
  16869=>"111111111",
  16870=>"110000000",
  16871=>"000000000",
  16872=>"111111011",
  16873=>"000000000",
  16874=>"000000000",
  16875=>"011011000",
  16876=>"111111111",
  16877=>"111111011",
  16878=>"111111111",
  16879=>"000000000",
  16880=>"110100110",
  16881=>"000100100",
  16882=>"111011011",
  16883=>"000011001",
  16884=>"111000110",
  16885=>"111111111",
  16886=>"000000000",
  16887=>"001111111",
  16888=>"001000001",
  16889=>"001001001",
  16890=>"000000011",
  16891=>"111111111",
  16892=>"010010110",
  16893=>"000000000",
  16894=>"111111111",
  16895=>"000000110",
  16896=>"111111000",
  16897=>"110000000",
  16898=>"011011111",
  16899=>"110100111",
  16900=>"111101100",
  16901=>"000011111",
  16902=>"111011000",
  16903=>"111011111",
  16904=>"000000111",
  16905=>"000000111",
  16906=>"101111111",
  16907=>"111111001",
  16908=>"111001011",
  16909=>"111111111",
  16910=>"100101111",
  16911=>"111111111",
  16912=>"000110111",
  16913=>"111111111",
  16914=>"001011000",
  16915=>"011111111",
  16916=>"111000000",
  16917=>"000111111",
  16918=>"110111000",
  16919=>"111101100",
  16920=>"000000111",
  16921=>"110100111",
  16922=>"111111011",
  16923=>"110000101",
  16924=>"000100101",
  16925=>"000111111",
  16926=>"111001111",
  16927=>"000000111",
  16928=>"001101101",
  16929=>"000000100",
  16930=>"000000000",
  16931=>"110110111",
  16932=>"000110000",
  16933=>"000000010",
  16934=>"111000000",
  16935=>"000111111",
  16936=>"111000000",
  16937=>"000000111",
  16938=>"011001000",
  16939=>"000000000",
  16940=>"101000000",
  16941=>"011111000",
  16942=>"000010001",
  16943=>"110111100",
  16944=>"011111111",
  16945=>"111000000",
  16946=>"011000000",
  16947=>"000000000",
  16948=>"001000000",
  16949=>"111111110",
  16950=>"000000110",
  16951=>"111110111",
  16952=>"001010111",
  16953=>"000111111",
  16954=>"100000000",
  16955=>"111110100",
  16956=>"111010000",
  16957=>"111111101",
  16958=>"001111011",
  16959=>"000000111",
  16960=>"000111111",
  16961=>"000000001",
  16962=>"111001111",
  16963=>"110000101",
  16964=>"000011101",
  16965=>"111111001",
  16966=>"111001111",
  16967=>"111000000",
  16968=>"011001001",
  16969=>"000000000",
  16970=>"000000000",
  16971=>"000100000",
  16972=>"001001111",
  16973=>"000000001",
  16974=>"000000000",
  16975=>"111111000",
  16976=>"000101111",
  16977=>"100101111",
  16978=>"000000011",
  16979=>"111111000",
  16980=>"000000000",
  16981=>"000000101",
  16982=>"111100000",
  16983=>"111000000",
  16984=>"000111111",
  16985=>"011111011",
  16986=>"000110111",
  16987=>"100000100",
  16988=>"000000101",
  16989=>"000000001",
  16990=>"000010000",
  16991=>"110000000",
  16992=>"000000000",
  16993=>"000000111",
  16994=>"011011000",
  16995=>"111111000",
  16996=>"001001000",
  16997=>"000000001",
  16998=>"100100110",
  16999=>"111111111",
  17000=>"000100000",
  17001=>"011111111",
  17002=>"111111110",
  17003=>"111111100",
  17004=>"110111000",
  17005=>"000000000",
  17006=>"000000000",
  17007=>"011011110",
  17008=>"001110000",
  17009=>"100111111",
  17010=>"000100111",
  17011=>"101100100",
  17012=>"111111000",
  17013=>"100111111",
  17014=>"000001111",
  17015=>"101000000",
  17016=>"000000011",
  17017=>"000101011",
  17018=>"000000000",
  17019=>"000111111",
  17020=>"111010000",
  17021=>"110100110",
  17022=>"000000110",
  17023=>"001000100",
  17024=>"001000000",
  17025=>"000100111",
  17026=>"001001100",
  17027=>"000100000",
  17028=>"000110100",
  17029=>"100000000",
  17030=>"010111111",
  17031=>"000111111",
  17032=>"000000000",
  17033=>"111010000",
  17034=>"001101000",
  17035=>"001100000",
  17036=>"111010111",
  17037=>"111000000",
  17038=>"111000000",
  17039=>"111110001",
  17040=>"000100110",
  17041=>"000111001",
  17042=>"000000000",
  17043=>"111111111",
  17044=>"001111111",
  17045=>"111101111",
  17046=>"000000000",
  17047=>"000000000",
  17048=>"001001111",
  17049=>"111111111",
  17050=>"011000001",
  17051=>"000011000",
  17052=>"111111111",
  17053=>"100001001",
  17054=>"000000111",
  17055=>"111111111",
  17056=>"000000000",
  17057=>"111111101",
  17058=>"011111011",
  17059=>"010111111",
  17060=>"111001000",
  17061=>"010000000",
  17062=>"000111111",
  17063=>"111101011",
  17064=>"000000000",
  17065=>"101000000",
  17066=>"111011000",
  17067=>"000000111",
  17068=>"000000000",
  17069=>"000000111",
  17070=>"011100000",
  17071=>"000000001",
  17072=>"100110110",
  17073=>"001001011",
  17074=>"010111111",
  17075=>"000111111",
  17076=>"111111100",
  17077=>"000000000",
  17078=>"110000000",
  17079=>"000001111",
  17080=>"000000000",
  17081=>"111111000",
  17082=>"110100100",
  17083=>"011101101",
  17084=>"000000111",
  17085=>"111001001",
  17086=>"001111000",
  17087=>"111111111",
  17088=>"111111111",
  17089=>"100111111",
  17090=>"000011111",
  17091=>"000000000",
  17092=>"000000000",
  17093=>"000000111",
  17094=>"101111011",
  17095=>"111111100",
  17096=>"000011011",
  17097=>"001000101",
  17098=>"000000111",
  17099=>"111111100",
  17100=>"111001001",
  17101=>"000111111",
  17102=>"110000100",
  17103=>"111100000",
  17104=>"000000111",
  17105=>"110111111",
  17106=>"111000001",
  17107=>"011111001",
  17108=>"111111000",
  17109=>"111100110",
  17110=>"000000000",
  17111=>"111001000",
  17112=>"000001011",
  17113=>"111100110",
  17114=>"000000110",
  17115=>"000111001",
  17116=>"001101100",
  17117=>"000000000",
  17118=>"000111111",
  17119=>"000000100",
  17120=>"000000000",
  17121=>"000100111",
  17122=>"000000110",
  17123=>"000000000",
  17124=>"110000000",
  17125=>"011000000",
  17126=>"111111101",
  17127=>"110110011",
  17128=>"000000001",
  17129=>"001001001",
  17130=>"111111111",
  17131=>"111001000",
  17132=>"000111111",
  17133=>"010111111",
  17134=>"010110111",
  17135=>"000000111",
  17136=>"000000011",
  17137=>"011001111",
  17138=>"111111001",
  17139=>"000100000",
  17140=>"011010001",
  17141=>"110000011",
  17142=>"000000100",
  17143=>"111111000",
  17144=>"000000111",
  17145=>"111101100",
  17146=>"000000000",
  17147=>"110000000",
  17148=>"100100000",
  17149=>"111111110",
  17150=>"000000111",
  17151=>"111111111",
  17152=>"100000000",
  17153=>"110000000",
  17154=>"111111111",
  17155=>"000000000",
  17156=>"100100100",
  17157=>"010110110",
  17158=>"111111001",
  17159=>"001000000",
  17160=>"001001001",
  17161=>"000000000",
  17162=>"000111111",
  17163=>"000000001",
  17164=>"110110000",
  17165=>"000000000",
  17166=>"000000000",
  17167=>"000110110",
  17168=>"000000000",
  17169=>"111111111",
  17170=>"000100111",
  17171=>"101111000",
  17172=>"010110000",
  17173=>"111000110",
  17174=>"110100100",
  17175=>"111111100",
  17176=>"111111000",
  17177=>"111000111",
  17178=>"001000111",
  17179=>"101000111",
  17180=>"010000000",
  17181=>"001111111",
  17182=>"111111111",
  17183=>"000000111",
  17184=>"110110000",
  17185=>"100101111",
  17186=>"000000111",
  17187=>"001101111",
  17188=>"001000000",
  17189=>"111111111",
  17190=>"111111111",
  17191=>"000111111",
  17192=>"010011111",
  17193=>"001000000",
  17194=>"011110000",
  17195=>"000111111",
  17196=>"001000000",
  17197=>"001111111",
  17198=>"000001101",
  17199=>"110000000",
  17200=>"000010101",
  17201=>"010110111",
  17202=>"111100100",
  17203=>"001000101",
  17204=>"000000000",
  17205=>"001000000",
  17206=>"110000111",
  17207=>"111111111",
  17208=>"000000000",
  17209=>"111111111",
  17210=>"000000001",
  17211=>"110110000",
  17212=>"000001000",
  17213=>"000000000",
  17214=>"111100000",
  17215=>"111000000",
  17216=>"000000110",
  17217=>"100101111",
  17218=>"000000010",
  17219=>"100000000",
  17220=>"010110111",
  17221=>"111011000",
  17222=>"100100000",
  17223=>"101101111",
  17224=>"000000000",
  17225=>"000000101",
  17226=>"101000000",
  17227=>"000000000",
  17228=>"100000111",
  17229=>"000001011",
  17230=>"011111111",
  17231=>"001001000",
  17232=>"010010000",
  17233=>"010110111",
  17234=>"000000000",
  17235=>"111001000",
  17236=>"000001000",
  17237=>"111111011",
  17238=>"000000000",
  17239=>"111111111",
  17240=>"001111100",
  17241=>"000000000",
  17242=>"111111000",
  17243=>"101001000",
  17244=>"000000111",
  17245=>"111101001",
  17246=>"110000111",
  17247=>"111111111",
  17248=>"111000000",
  17249=>"111111000",
  17250=>"100100110",
  17251=>"111000000",
  17252=>"111011000",
  17253=>"000000000",
  17254=>"000110000",
  17255=>"000001111",
  17256=>"000000001",
  17257=>"001011001",
  17258=>"000000000",
  17259=>"001001111",
  17260=>"000000011",
  17261=>"110100100",
  17262=>"000000110",
  17263=>"011011110",
  17264=>"000000111",
  17265=>"010010111",
  17266=>"000000101",
  17267=>"111101100",
  17268=>"111111111",
  17269=>"110110111",
  17270=>"000000001",
  17271=>"000010111",
  17272=>"011000000",
  17273=>"000101101",
  17274=>"111101000",
  17275=>"000000000",
  17276=>"011000000",
  17277=>"000000100",
  17278=>"000100100",
  17279=>"011011111",
  17280=>"110110111",
  17281=>"000000011",
  17282=>"111110100",
  17283=>"111000000",
  17284=>"111000000",
  17285=>"111110100",
  17286=>"000000100",
  17287=>"111000110",
  17288=>"000000000",
  17289=>"011111111",
  17290=>"000001001",
  17291=>"110111111",
  17292=>"110111101",
  17293=>"101001000",
  17294=>"110110111",
  17295=>"111111011",
  17296=>"111111011",
  17297=>"110000000",
  17298=>"100000000",
  17299=>"000110110",
  17300=>"000100000",
  17301=>"001000000",
  17302=>"111111111",
  17303=>"100101000",
  17304=>"110111011",
  17305=>"111011011",
  17306=>"000100001",
  17307=>"001000000",
  17308=>"000001001",
  17309=>"001000111",
  17310=>"001000000",
  17311=>"000000000",
  17312=>"000000000",
  17313=>"101111111",
  17314=>"000000110",
  17315=>"111000011",
  17316=>"000111111",
  17317=>"000000000",
  17318=>"111111000",
  17319=>"000011100",
  17320=>"001001001",
  17321=>"000000111",
  17322=>"000001111",
  17323=>"111111111",
  17324=>"000000000",
  17325=>"000001111",
  17326=>"001111111",
  17327=>"111111110",
  17328=>"011011111",
  17329=>"111100110",
  17330=>"000000101",
  17331=>"000101111",
  17332=>"000000000",
  17333=>"000111111",
  17334=>"000000000",
  17335=>"000111101",
  17336=>"000000000",
  17337=>"011111001",
  17338=>"111001100",
  17339=>"010000010",
  17340=>"111111111",
  17341=>"101100111",
  17342=>"011000111",
  17343=>"100110010",
  17344=>"100111011",
  17345=>"101101111",
  17346=>"111111111",
  17347=>"000000100",
  17348=>"100101111",
  17349=>"000000111",
  17350=>"001001000",
  17351=>"000000000",
  17352=>"111000000",
  17353=>"111111111",
  17354=>"000000000",
  17355=>"001111111",
  17356=>"111000000",
  17357=>"111111111",
  17358=>"111000000",
  17359=>"000011010",
  17360=>"000000010",
  17361=>"000111111",
  17362=>"111111111",
  17363=>"111111001",
  17364=>"000110000",
  17365=>"111000000",
  17366=>"000000000",
  17367=>"111100100",
  17368=>"000001001",
  17369=>"000100101",
  17370=>"110100111",
  17371=>"111001111",
  17372=>"111111111",
  17373=>"111110100",
  17374=>"101101101",
  17375=>"110000001",
  17376=>"111010000",
  17377=>"110111111",
  17378=>"111000000",
  17379=>"000000010",
  17380=>"000110111",
  17381=>"001000101",
  17382=>"111011111",
  17383=>"111000000",
  17384=>"001000000",
  17385=>"111111101",
  17386=>"000101111",
  17387=>"111111000",
  17388=>"000000111",
  17389=>"011111110",
  17390=>"000001011",
  17391=>"011010011",
  17392=>"111000000",
  17393=>"000000000",
  17394=>"111000001",
  17395=>"000000000",
  17396=>"111100000",
  17397=>"111111111",
  17398=>"111111000",
  17399=>"100000001",
  17400=>"111111111",
  17401=>"011011000",
  17402=>"100110111",
  17403=>"111111111",
  17404=>"000000100",
  17405=>"011011011",
  17406=>"000011011",
  17407=>"000000000",
  17408=>"000000000",
  17409=>"000000000",
  17410=>"100101111",
  17411=>"111111111",
  17412=>"000000000",
  17413=>"110110111",
  17414=>"011011011",
  17415=>"111111111",
  17416=>"110111101",
  17417=>"000000001",
  17418=>"111111000",
  17419=>"111111101",
  17420=>"100000100",
  17421=>"000000000",
  17422=>"000110111",
  17423=>"111110000",
  17424=>"111111111",
  17425=>"000011000",
  17426=>"000000000",
  17427=>"000000001",
  17428=>"000111111",
  17429=>"100000000",
  17430=>"100101111",
  17431=>"001001100",
  17432=>"111111111",
  17433=>"101000000",
  17434=>"000000000",
  17435=>"100100011",
  17436=>"111001000",
  17437=>"000000000",
  17438=>"111111111",
  17439=>"111110100",
  17440=>"110111011",
  17441=>"000000000",
  17442=>"001101111",
  17443=>"101000000",
  17444=>"110001000",
  17445=>"000000100",
  17446=>"111011011",
  17447=>"100000000",
  17448=>"000000000",
  17449=>"111111000",
  17450=>"111000000",
  17451=>"111111111",
  17452=>"000000100",
  17453=>"111111111",
  17454=>"111111100",
  17455=>"111111111",
  17456=>"001000001",
  17457=>"111111010",
  17458=>"101110110",
  17459=>"000000000",
  17460=>"111111111",
  17461=>"110111110",
  17462=>"111000110",
  17463=>"000000101",
  17464=>"000001000",
  17465=>"000000111",
  17466=>"101001000",
  17467=>"011000001",
  17468=>"101001000",
  17469=>"111000001",
  17470=>"100000000",
  17471=>"110100000",
  17472=>"101000001",
  17473=>"111011001",
  17474=>"000000001",
  17475=>"000000001",
  17476=>"111100000",
  17477=>"111111111",
  17478=>"011000000",
  17479=>"000000000",
  17480=>"111011111",
  17481=>"111000111",
  17482=>"111111010",
  17483=>"111110111",
  17484=>"000000100",
  17485=>"000000000",
  17486=>"100100111",
  17487=>"101000011",
  17488=>"000000111",
  17489=>"001000000",
  17490=>"111000000",
  17491=>"011111111",
  17492=>"111111111",
  17493=>"111111011",
  17494=>"111111011",
  17495=>"000111010",
  17496=>"111000000",
  17497=>"100000000",
  17498=>"111000000",
  17499=>"110111111",
  17500=>"011111111",
  17501=>"000000010",
  17502=>"111111000",
  17503=>"000000000",
  17504=>"000000000",
  17505=>"000000001",
  17506=>"000100001",
  17507=>"111000001",
  17508=>"101110101",
  17509=>"111100111",
  17510=>"000000000",
  17511=>"111111001",
  17512=>"111111111",
  17513=>"000000000",
  17514=>"000001111",
  17515=>"100000111",
  17516=>"001000000",
  17517=>"001100000",
  17518=>"111001001",
  17519=>"111110001",
  17520=>"001001111",
  17521=>"100110110",
  17522=>"000010111",
  17523=>"111001101",
  17524=>"011011011",
  17525=>"001011111",
  17526=>"111111001",
  17527=>"111011000",
  17528=>"000000000",
  17529=>"000000001",
  17530=>"000000000",
  17531=>"111111001",
  17532=>"100100110",
  17533=>"000000111",
  17534=>"000000000",
  17535=>"111111111",
  17536=>"000000000",
  17537=>"111111111",
  17538=>"111111000",
  17539=>"000000001",
  17540=>"000000011",
  17541=>"000000000",
  17542=>"111111111",
  17543=>"000000110",
  17544=>"000000000",
  17545=>"111011111",
  17546=>"000011111",
  17547=>"100111111",
  17548=>"111110111",
  17549=>"000000000",
  17550=>"111111111",
  17551=>"111111111",
  17552=>"000000000",
  17553=>"111111111",
  17554=>"011110110",
  17555=>"011011001",
  17556=>"011011101",
  17557=>"010011011",
  17558=>"001000000",
  17559=>"000000000",
  17560=>"001000000",
  17561=>"100110010",
  17562=>"111111111",
  17563=>"001000000",
  17564=>"100000000",
  17565=>"010111111",
  17566=>"000000000",
  17567=>"111000000",
  17568=>"111111101",
  17569=>"000000000",
  17570=>"011000000",
  17571=>"000000011",
  17572=>"111000000",
  17573=>"011011111",
  17574=>"111001111",
  17575=>"001111111",
  17576=>"000000000",
  17577=>"011011001",
  17578=>"000000000",
  17579=>"111111011",
  17580=>"000110110",
  17581=>"000000000",
  17582=>"111111110",
  17583=>"000000111",
  17584=>"011111000",
  17585=>"011010010",
  17586=>"111111010",
  17587=>"000000111",
  17588=>"011100000",
  17589=>"110111111",
  17590=>"110111011",
  17591=>"111111000",
  17592=>"000100111",
  17593=>"011011111",
  17594=>"011001001",
  17595=>"000000000",
  17596=>"000000111",
  17597=>"111111111",
  17598=>"000000000",
  17599=>"111000000",
  17600=>"110011000",
  17601=>"111100111",
  17602=>"110000000",
  17603=>"000000000",
  17604=>"110111111",
  17605=>"000000000",
  17606=>"000000001",
  17607=>"001000000",
  17608=>"000111111",
  17609=>"100100110",
  17610=>"001000010",
  17611=>"001000000",
  17612=>"111001111",
  17613=>"000000000",
  17614=>"111010000",
  17615=>"000000000",
  17616=>"111000000",
  17617=>"000100000",
  17618=>"111011001",
  17619=>"000110110",
  17620=>"111111111",
  17621=>"111111111",
  17622=>"000001000",
  17623=>"000111000",
  17624=>"111111000",
  17625=>"111111111",
  17626=>"100100110",
  17627=>"001011111",
  17628=>"100000000",
  17629=>"001001000",
  17630=>"110111000",
  17631=>"000011011",
  17632=>"100101001",
  17633=>"110010001",
  17634=>"110111111",
  17635=>"000000000",
  17636=>"000000000",
  17637=>"000111100",
  17638=>"100100110",
  17639=>"010110000",
  17640=>"101000000",
  17641=>"110111111",
  17642=>"111111000",
  17643=>"111111111",
  17644=>"000000000",
  17645=>"111111100",
  17646=>"000100000",
  17647=>"101000000",
  17648=>"100000100",
  17649=>"000111111",
  17650=>"001111111",
  17651=>"000000011",
  17652=>"111111010",
  17653=>"001000100",
  17654=>"011101001",
  17655=>"000000000",
  17656=>"000000000",
  17657=>"000000000",
  17658=>"111111010",
  17659=>"000100111",
  17660=>"111110000",
  17661=>"001001111",
  17662=>"011111111",
  17663=>"000000000",
  17664=>"111100101",
  17665=>"110111011",
  17666=>"000111000",
  17667=>"111111011",
  17668=>"100111011",
  17669=>"000111011",
  17670=>"000000000",
  17671=>"111111011",
  17672=>"000001000",
  17673=>"000000000",
  17674=>"011000001",
  17675=>"111111011",
  17676=>"001000000",
  17677=>"111110100",
  17678=>"111111000",
  17679=>"111111000",
  17680=>"111111111",
  17681=>"000000001",
  17682=>"001000000",
  17683=>"000000010",
  17684=>"000000011",
  17685=>"111111111",
  17686=>"101111111",
  17687=>"001001000",
  17688=>"011111111",
  17689=>"111111111",
  17690=>"101101101",
  17691=>"000000000",
  17692=>"000000000",
  17693=>"111011111",
  17694=>"000000000",
  17695=>"111101000",
  17696=>"110010000",
  17697=>"011000000",
  17698=>"111111110",
  17699=>"101111000",
  17700=>"000000000",
  17701=>"000000000",
  17702=>"000000000",
  17703=>"110110001",
  17704=>"100000000",
  17705=>"000000000",
  17706=>"111111111",
  17707=>"111111111",
  17708=>"000000111",
  17709=>"111101101",
  17710=>"000000011",
  17711=>"111111010",
  17712=>"111010110",
  17713=>"010000000",
  17714=>"000000000",
  17715=>"101001101",
  17716=>"000000011",
  17717=>"000000000",
  17718=>"000000000",
  17719=>"100000000",
  17720=>"110110100",
  17721=>"110000000",
  17722=>"000000001",
  17723=>"001000000",
  17724=>"000000000",
  17725=>"010011100",
  17726=>"111011111",
  17727=>"011011001",
  17728=>"000101111",
  17729=>"111111110",
  17730=>"000000000",
  17731=>"000000111",
  17732=>"000000111",
  17733=>"000000000",
  17734=>"111111111",
  17735=>"000000000",
  17736=>"000000000",
  17737=>"000000000",
  17738=>"000111111",
  17739=>"100001000",
  17740=>"000000111",
  17741=>"100000000",
  17742=>"100000000",
  17743=>"000001110",
  17744=>"000000001",
  17745=>"000000000",
  17746=>"001000011",
  17747=>"111110000",
  17748=>"000111110",
  17749=>"011000000",
  17750=>"111111111",
  17751=>"000000000",
  17752=>"111001000",
  17753=>"000000000",
  17754=>"000001111",
  17755=>"000111100",
  17756=>"000000000",
  17757=>"000000110",
  17758=>"001111111",
  17759=>"000110000",
  17760=>"000000000",
  17761=>"111000101",
  17762=>"011010110",
  17763=>"111111111",
  17764=>"100001011",
  17765=>"000000000",
  17766=>"010000000",
  17767=>"001111111",
  17768=>"111111100",
  17769=>"110100000",
  17770=>"000010000",
  17771=>"001100100",
  17772=>"011111111",
  17773=>"001000101",
  17774=>"111111111",
  17775=>"001000000",
  17776=>"001011010",
  17777=>"111110111",
  17778=>"000000000",
  17779=>"110111111",
  17780=>"000000000",
  17781=>"000000111",
  17782=>"011011000",
  17783=>"000000000",
  17784=>"000000000",
  17785=>"111011111",
  17786=>"000000111",
  17787=>"001101111",
  17788=>"000111111",
  17789=>"111001001",
  17790=>"111011000",
  17791=>"001001000",
  17792=>"111111011",
  17793=>"111111000",
  17794=>"111111000",
  17795=>"000000000",
  17796=>"011000001",
  17797=>"010011011",
  17798=>"110111111",
  17799=>"111111011",
  17800=>"001000101",
  17801=>"111111011",
  17802=>"100000110",
  17803=>"111111000",
  17804=>"000101111",
  17805=>"000000000",
  17806=>"111111100",
  17807=>"000000000",
  17808=>"000000001",
  17809=>"000100111",
  17810=>"111111000",
  17811=>"001001000",
  17812=>"000000000",
  17813=>"000010000",
  17814=>"011000011",
  17815=>"000111111",
  17816=>"111111111",
  17817=>"011001000",
  17818=>"000000001",
  17819=>"100000000",
  17820=>"001010111",
  17821=>"111111111",
  17822=>"100111111",
  17823=>"011111111",
  17824=>"110110011",
  17825=>"011000001",
  17826=>"111111111",
  17827=>"011000100",
  17828=>"111111010",
  17829=>"111111111",
  17830=>"001000000",
  17831=>"111110100",
  17832=>"100000111",
  17833=>"000000000",
  17834=>"000000110",
  17835=>"000000100",
  17836=>"000000000",
  17837=>"000000000",
  17838=>"011011000",
  17839=>"111011001",
  17840=>"111110110",
  17841=>"111111000",
  17842=>"001001000",
  17843=>"000000000",
  17844=>"010011000",
  17845=>"000000011",
  17846=>"001011111",
  17847=>"000000000",
  17848=>"111111101",
  17849=>"111111011",
  17850=>"011000000",
  17851=>"110111111",
  17852=>"111111000",
  17853=>"000001111",
  17854=>"111000000",
  17855=>"100010111",
  17856=>"000000000",
  17857=>"101111100",
  17858=>"000000000",
  17859=>"111111111",
  17860=>"111110000",
  17861=>"001011111",
  17862=>"000110111",
  17863=>"100100101",
  17864=>"000000000",
  17865=>"101111111",
  17866=>"000000000",
  17867=>"000000101",
  17868=>"111100100",
  17869=>"100100001",
  17870=>"001000000",
  17871=>"000000100",
  17872=>"110111111",
  17873=>"111111111",
  17874=>"001101111",
  17875=>"111111111",
  17876=>"111110010",
  17877=>"001000000",
  17878=>"111100000",
  17879=>"011111001",
  17880=>"100100101",
  17881=>"111111110",
  17882=>"111110000",
  17883=>"001101000",
  17884=>"111000101",
  17885=>"111111110",
  17886=>"000000000",
  17887=>"000001101",
  17888=>"111000100",
  17889=>"111111111",
  17890=>"111111110",
  17891=>"111100000",
  17892=>"101101111",
  17893=>"111111110",
  17894=>"110111111",
  17895=>"111111111",
  17896=>"001001011",
  17897=>"111111111",
  17898=>"111100000",
  17899=>"111111111",
  17900=>"000100000",
  17901=>"000000100",
  17902=>"000000000",
  17903=>"000101111",
  17904=>"000000000",
  17905=>"000111110",
  17906=>"000110110",
  17907=>"011000000",
  17908=>"000000000",
  17909=>"111111111",
  17910=>"111000000",
  17911=>"011001000",
  17912=>"000100000",
  17913=>"011001001",
  17914=>"100000000",
  17915=>"111111100",
  17916=>"000000001",
  17917=>"000000000",
  17918=>"101000000",
  17919=>"111111111",
  17920=>"011101000",
  17921=>"111111111",
  17922=>"111111111",
  17923=>"000000111",
  17924=>"000000000",
  17925=>"111110010",
  17926=>"000000000",
  17927=>"111111111",
  17928=>"001001111",
  17929=>"001000000",
  17930=>"111111111",
  17931=>"000010010",
  17932=>"111000000",
  17933=>"111111000",
  17934=>"111110100",
  17935=>"001000000",
  17936=>"001111001",
  17937=>"011111111",
  17938=>"011111111",
  17939=>"000000000",
  17940=>"001000000",
  17941=>"111111010",
  17942=>"010000000",
  17943=>"011111111",
  17944=>"111111111",
  17945=>"111011001",
  17946=>"001001001",
  17947=>"111111111",
  17948=>"111100101",
  17949=>"010111111",
  17950=>"110110110",
  17951=>"000000111",
  17952=>"001000000",
  17953=>"010010000",
  17954=>"000000011",
  17955=>"111111111",
  17956=>"001000000",
  17957=>"010110010",
  17958=>"000011011",
  17959=>"000001111",
  17960=>"000111001",
  17961=>"000000000",
  17962=>"111011111",
  17963=>"111110110",
  17964=>"110111111",
  17965=>"111111001",
  17966=>"111000000",
  17967=>"011000000",
  17968=>"011110110",
  17969=>"001001000",
  17970=>"100011000",
  17971=>"000010110",
  17972=>"000000000",
  17973=>"111011011",
  17974=>"111111000",
  17975=>"000110111",
  17976=>"111000110",
  17977=>"011001000",
  17978=>"000000000",
  17979=>"100101111",
  17980=>"111000000",
  17981=>"000000000",
  17982=>"000010000",
  17983=>"011000000",
  17984=>"110001001",
  17985=>"111000011",
  17986=>"001111001",
  17987=>"000000011",
  17988=>"001001000",
  17989=>"110100000",
  17990=>"001000000",
  17991=>"111000000",
  17992=>"110000000",
  17993=>"000000000",
  17994=>"110101111",
  17995=>"111001001",
  17996=>"111111001",
  17997=>"000000001",
  17998=>"000111111",
  17999=>"111100000",
  18000=>"011001001",
  18001=>"111100000",
  18002=>"000100111",
  18003=>"101111111",
  18004=>"001000000",
  18005=>"000000000",
  18006=>"110000111",
  18007=>"010010111",
  18008=>"000000000",
  18009=>"111000000",
  18010=>"111011011",
  18011=>"011001001",
  18012=>"011011111",
  18013=>"001111111",
  18014=>"111011111",
  18015=>"111000000",
  18016=>"000000111",
  18017=>"110111111",
  18018=>"101110100",
  18019=>"000000000",
  18020=>"000000000",
  18021=>"111000000",
  18022=>"111111110",
  18023=>"000000000",
  18024=>"110000000",
  18025=>"000000100",
  18026=>"111001001",
  18027=>"011101111",
  18028=>"000000001",
  18029=>"111110000",
  18030=>"111100000",
  18031=>"101001111",
  18032=>"010110100",
  18033=>"111111111",
  18034=>"111111100",
  18035=>"111000000",
  18036=>"111010000",
  18037=>"111111111",
  18038=>"001000000",
  18039=>"000000101",
  18040=>"111000000",
  18041=>"111110000",
  18042=>"000000000",
  18043=>"010011010",
  18044=>"111111100",
  18045=>"011111111",
  18046=>"010100000",
  18047=>"011010000",
  18048=>"001111111",
  18049=>"110110010",
  18050=>"000000111",
  18051=>"000000110",
  18052=>"000000110",
  18053=>"111100111",
  18054=>"000000000",
  18055=>"010010010",
  18056=>"001011111",
  18057=>"101101101",
  18058=>"000000000",
  18059=>"111100100",
  18060=>"011011111",
  18061=>"011010000",
  18062=>"111110100",
  18063=>"100000000",
  18064=>"111111001",
  18065=>"000011011",
  18066=>"001000000",
  18067=>"000000000",
  18068=>"010010000",
  18069=>"000010010",
  18070=>"111100001",
  18071=>"111001111",
  18072=>"111111110",
  18073=>"001100100",
  18074=>"000000110",
  18075=>"000111011",
  18076=>"000000001",
  18077=>"001000000",
  18078=>"111001000",
  18079=>"111111111",
  18080=>"000000000",
  18081=>"010010000",
  18082=>"111000000",
  18083=>"111111000",
  18084=>"011001011",
  18085=>"000110110",
  18086=>"111011011",
  18087=>"111111001",
  18088=>"001000100",
  18089=>"111000101",
  18090=>"001111000",
  18091=>"010111111",
  18092=>"011001111",
  18093=>"010111110",
  18094=>"100000000",
  18095=>"111111111",
  18096=>"011000000",
  18097=>"111110010",
  18098=>"111111111",
  18099=>"010000000",
  18100=>"110100000",
  18101=>"000001011",
  18102=>"000011111",
  18103=>"001111011",
  18104=>"000000111",
  18105=>"000000001",
  18106=>"101000001",
  18107=>"111111001",
  18108=>"000000000",
  18109=>"000000011",
  18110=>"000000000",
  18111=>"001000111",
  18112=>"100111111",
  18113=>"110000100",
  18114=>"111111111",
  18115=>"111110111",
  18116=>"111000100",
  18117=>"110111000",
  18118=>"000000000",
  18119=>"000000000",
  18120=>"000101111",
  18121=>"111000000",
  18122=>"000110100",
  18123=>"101000000",
  18124=>"111111111",
  18125=>"000111011",
  18126=>"000000011",
  18127=>"011111111",
  18128=>"000000000",
  18129=>"001101111",
  18130=>"000111111",
  18131=>"111000000",
  18132=>"011000000",
  18133=>"111001000",
  18134=>"111001000",
  18135=>"000000000",
  18136=>"000111000",
  18137=>"111011001",
  18138=>"000000000",
  18139=>"001001111",
  18140=>"000001011",
  18141=>"111010110",
  18142=>"010111111",
  18143=>"000000000",
  18144=>"111111111",
  18145=>"000000111",
  18146=>"111111000",
  18147=>"000000000",
  18148=>"011000000",
  18149=>"100100000",
  18150=>"000000011",
  18151=>"111111110",
  18152=>"100110111",
  18153=>"011000100",
  18154=>"111100000",
  18155=>"110000000",
  18156=>"000100100",
  18157=>"001001001",
  18158=>"000000001",
  18159=>"101001001",
  18160=>"100111111",
  18161=>"100111011",
  18162=>"011111111",
  18163=>"110111001",
  18164=>"000010000",
  18165=>"111101001",
  18166=>"000111111",
  18167=>"110100000",
  18168=>"000111001",
  18169=>"000000011",
  18170=>"000001111",
  18171=>"000111111",
  18172=>"110100000",
  18173=>"000000000",
  18174=>"000000110",
  18175=>"111111110",
  18176=>"111111011",
  18177=>"111110100",
  18178=>"111111110",
  18179=>"111111000",
  18180=>"000000111",
  18181=>"000000111",
  18182=>"111111111",
  18183=>"110111111",
  18184=>"110111110",
  18185=>"001001001",
  18186=>"111000000",
  18187=>"111111111",
  18188=>"000000001",
  18189=>"110010001",
  18190=>"111000111",
  18191=>"000011000",
  18192=>"000000110",
  18193=>"010000000",
  18194=>"011000000",
  18195=>"111010111",
  18196=>"001001000",
  18197=>"111111111",
  18198=>"001000000",
  18199=>"010010111",
  18200=>"011111111",
  18201=>"101111000",
  18202=>"000110111",
  18203=>"000001011",
  18204=>"011111000",
  18205=>"000000000",
  18206=>"100111111",
  18207=>"000100000",
  18208=>"000000010",
  18209=>"111101001",
  18210=>"000111111",
  18211=>"111111111",
  18212=>"100100111",
  18213=>"100000000",
  18214=>"100000000",
  18215=>"000110111",
  18216=>"000010000",
  18217=>"100000000",
  18218=>"000010011",
  18219=>"000000010",
  18220=>"000000000",
  18221=>"000110110",
  18222=>"111111111",
  18223=>"001001000",
  18224=>"111111111",
  18225=>"000000000",
  18226=>"110111011",
  18227=>"000000011",
  18228=>"010001011",
  18229=>"011010110",
  18230=>"000000111",
  18231=>"111111111",
  18232=>"000011000",
  18233=>"111000000",
  18234=>"011000111",
  18235=>"001001100",
  18236=>"110110010",
  18237=>"010000101",
  18238=>"010010000",
  18239=>"000000001",
  18240=>"011000000",
  18241=>"111111101",
  18242=>"111011110",
  18243=>"110100000",
  18244=>"000000011",
  18245=>"001111101",
  18246=>"001011110",
  18247=>"111111000",
  18248=>"011001110",
  18249=>"000001111",
  18250=>"111111110",
  18251=>"111000000",
  18252=>"000111011",
  18253=>"000000000",
  18254=>"000100111",
  18255=>"100001011",
  18256=>"100001000",
  18257=>"000000000",
  18258=>"111100000",
  18259=>"011000000",
  18260=>"000100110",
  18261=>"111110010",
  18262=>"111111000",
  18263=>"110111111",
  18264=>"111111111",
  18265=>"000000101",
  18266=>"110010000",
  18267=>"111111111",
  18268=>"000001001",
  18269=>"110110111",
  18270=>"011011011",
  18271=>"111101101",
  18272=>"000000001",
  18273=>"110111111",
  18274=>"111111011",
  18275=>"101100100",
  18276=>"100100000",
  18277=>"000100000",
  18278=>"000101111",
  18279=>"001101111",
  18280=>"111100000",
  18281=>"000000111",
  18282=>"000111101",
  18283=>"000000000",
  18284=>"000100111",
  18285=>"001011111",
  18286=>"000110111",
  18287=>"100000000",
  18288=>"000010111",
  18289=>"000000010",
  18290=>"000010111",
  18291=>"000000000",
  18292=>"111101001",
  18293=>"110100000",
  18294=>"101000000",
  18295=>"000000010",
  18296=>"101000110",
  18297=>"111001111",
  18298=>"011111111",
  18299=>"000000110",
  18300=>"111010010",
  18301=>"000100111",
  18302=>"000000111",
  18303=>"111101000",
  18304=>"111001001",
  18305=>"000110110",
  18306=>"111000000",
  18307=>"111001000",
  18308=>"000000111",
  18309=>"000100110",
  18310=>"111111110",
  18311=>"000000000",
  18312=>"000111110",
  18313=>"111101111",
  18314=>"111000000",
  18315=>"111101101",
  18316=>"111111111",
  18317=>"111111100",
  18318=>"000000111",
  18319=>"100000111",
  18320=>"011011011",
  18321=>"000110000",
  18322=>"000111111",
  18323=>"011011010",
  18324=>"000111111",
  18325=>"000000000",
  18326=>"001100111",
  18327=>"110000000",
  18328=>"000000000",
  18329=>"001110110",
  18330=>"111111000",
  18331=>"001001001",
  18332=>"000000111",
  18333=>"000110010",
  18334=>"001000000",
  18335=>"000000000",
  18336=>"000000000",
  18337=>"000111011",
  18338=>"111111100",
  18339=>"000011011",
  18340=>"110110000",
  18341=>"011001000",
  18342=>"000000000",
  18343=>"100111110",
  18344=>"000000000",
  18345=>"000000000",
  18346=>"111111111",
  18347=>"011000000",
  18348=>"101000000",
  18349=>"000001001",
  18350=>"100001101",
  18351=>"111000000",
  18352=>"001000100",
  18353=>"000000001",
  18354=>"101100000",
  18355=>"111000000",
  18356=>"111111001",
  18357=>"111111111",
  18358=>"111111100",
  18359=>"000000000",
  18360=>"000000000",
  18361=>"001011111",
  18362=>"111111000",
  18363=>"111110110",
  18364=>"000100111",
  18365=>"111000000",
  18366=>"111111111",
  18367=>"111110101",
  18368=>"111111001",
  18369=>"111001000",
  18370=>"111111111",
  18371=>"000111111",
  18372=>"000000000",
  18373=>"011011011",
  18374=>"000000001",
  18375=>"111000000",
  18376=>"000000001",
  18377=>"000010111",
  18378=>"000000001",
  18379=>"000010010",
  18380=>"111111111",
  18381=>"000110110",
  18382=>"001000000",
  18383=>"111010111",
  18384=>"111000010",
  18385=>"111111000",
  18386=>"011011111",
  18387=>"000000010",
  18388=>"100110100",
  18389=>"000000111",
  18390=>"000000000",
  18391=>"000000000",
  18392=>"001000100",
  18393=>"000000000",
  18394=>"111000000",
  18395=>"000000001",
  18396=>"111111110",
  18397=>"000000001",
  18398=>"101000011",
  18399=>"001000000",
  18400=>"011111000",
  18401=>"111111000",
  18402=>"111001000",
  18403=>"110000000",
  18404=>"011010000",
  18405=>"011000110",
  18406=>"000000001",
  18407=>"001000000",
  18408=>"111110111",
  18409=>"001001001",
  18410=>"110111011",
  18411=>"000000000",
  18412=>"001000000",
  18413=>"000011011",
  18414=>"001000000",
  18415=>"000110111",
  18416=>"111100000",
  18417=>"001001111",
  18418=>"000000111",
  18419=>"111001000",
  18420=>"000001111",
  18421=>"000000000",
  18422=>"111111111",
  18423=>"001111110",
  18424=>"000001001",
  18425=>"100111011",
  18426=>"100000000",
  18427=>"010000000",
  18428=>"100000100",
  18429=>"110111100",
  18430=>"111000000",
  18431=>"000000000",
  18432=>"111111000",
  18433=>"110110111",
  18434=>"111011000",
  18435=>"111110101",
  18436=>"001001001",
  18437=>"000001111",
  18438=>"111111111",
  18439=>"110000111",
  18440=>"101000000",
  18441=>"100000000",
  18442=>"001000000",
  18443=>"111101001",
  18444=>"111011111",
  18445=>"111101111",
  18446=>"100100000",
  18447=>"000000101",
  18448=>"100000000",
  18449=>"111001001",
  18450=>"001111111",
  18451=>"111111111",
  18452=>"110110000",
  18453=>"001000111",
  18454=>"010011111",
  18455=>"001000000",
  18456=>"000001000",
  18457=>"110001111",
  18458=>"001111110",
  18459=>"100100111",
  18460=>"100111110",
  18461=>"111111111",
  18462=>"001111100",
  18463=>"100111111",
  18464=>"111111111",
  18465=>"000001001",
  18466=>"000000000",
  18467=>"011111111",
  18468=>"000011111",
  18469=>"000000110",
  18470=>"001000111",
  18471=>"101100000",
  18472=>"001001111",
  18473=>"011011000",
  18474=>"111111111",
  18475=>"111111000",
  18476=>"001010000",
  18477=>"011111111",
  18478=>"111000000",
  18479=>"100000000",
  18480=>"011111111",
  18481=>"000111111",
  18482=>"111101000",
  18483=>"111111000",
  18484=>"000000000",
  18485=>"111100000",
  18486=>"001000111",
  18487=>"000011111",
  18488=>"000110000",
  18489=>"111110111",
  18490=>"110110000",
  18491=>"111000100",
  18492=>"000000000",
  18493=>"101100111",
  18494=>"110111111",
  18495=>"111111111",
  18496=>"000111011",
  18497=>"000000000",
  18498=>"111101100",
  18499=>"101000101",
  18500=>"000111111",
  18501=>"011111000",
  18502=>"111111110",
  18503=>"111110111",
  18504=>"101111111",
  18505=>"111000000",
  18506=>"000000111",
  18507=>"000000000",
  18508=>"111111111",
  18509=>"110110111",
  18510=>"000000100",
  18511=>"001000100",
  18512=>"000000111",
  18513=>"011000000",
  18514=>"111001000",
  18515=>"100001000",
  18516=>"111101101",
  18517=>"000000000",
  18518=>"011111111",
  18519=>"000111000",
  18520=>"001000000",
  18521=>"101000001",
  18522=>"111110010",
  18523=>"101111111",
  18524=>"000000000",
  18525=>"111101111",
  18526=>"100001001",
  18527=>"000000000",
  18528=>"000000000",
  18529=>"111000011",
  18530=>"000000110",
  18531=>"000000111",
  18532=>"111111010",
  18533=>"111111111",
  18534=>"111010000",
  18535=>"011001000",
  18536=>"111111010",
  18537=>"111111011",
  18538=>"111100111",
  18539=>"111111010",
  18540=>"111111111",
  18541=>"101111000",
  18542=>"000000000",
  18543=>"111110010",
  18544=>"011011011",
  18545=>"110100111",
  18546=>"100100000",
  18547=>"001010000",
  18548=>"101000000",
  18549=>"001001001",
  18550=>"101000000",
  18551=>"111111100",
  18552=>"000111111",
  18553=>"110110111",
  18554=>"111111111",
  18555=>"111111111",
  18556=>"000001000",
  18557=>"000000100",
  18558=>"111111111",
  18559=>"111111111",
  18560=>"010011010",
  18561=>"001001011",
  18562=>"011000111",
  18563=>"111110000",
  18564=>"110110011",
  18565=>"000000111",
  18566=>"111111111",
  18567=>"111001001",
  18568=>"111111011",
  18569=>"000000111",
  18570=>"000000001",
  18571=>"111111111",
  18572=>"111000001",
  18573=>"000000001",
  18574=>"100100100",
  18575=>"111111100",
  18576=>"001000000",
  18577=>"111111111",
  18578=>"110111001",
  18579=>"110000000",
  18580=>"100110111",
  18581=>"000000100",
  18582=>"010010110",
  18583=>"010000000",
  18584=>"001001001",
  18585=>"000000000",
  18586=>"001000000",
  18587=>"100100101",
  18588=>"110111111",
  18589=>"111111101",
  18590=>"111111111",
  18591=>"000000000",
  18592=>"111111100",
  18593=>"110000000",
  18594=>"101111110",
  18595=>"000110111",
  18596=>"111111101",
  18597=>"110100001",
  18598=>"111101111",
  18599=>"001100111",
  18600=>"001000000",
  18601=>"001001101",
  18602=>"011000000",
  18603=>"110111000",
  18604=>"011011001",
  18605=>"000101011",
  18606=>"111011010",
  18607=>"000000111",
  18608=>"100100111",
  18609=>"111100101",
  18610=>"111111111",
  18611=>"111111111",
  18612=>"111101111",
  18613=>"000000000",
  18614=>"111111111",
  18615=>"000000000",
  18616=>"111111111",
  18617=>"110111111",
  18618=>"000000100",
  18619=>"101001011",
  18620=>"001000000",
  18621=>"000000000",
  18622=>"110100000",
  18623=>"111101111",
  18624=>"000000010",
  18625=>"111111111",
  18626=>"111111111",
  18627=>"001001111",
  18628=>"000000000",
  18629=>"000011011",
  18630=>"000100000",
  18631=>"111100101",
  18632=>"000111111",
  18633=>"111111111",
  18634=>"000000000",
  18635=>"000000000",
  18636=>"100110000",
  18637=>"101011000",
  18638=>"111110111",
  18639=>"111110111",
  18640=>"011111111",
  18641=>"000000111",
  18642=>"000000111",
  18643=>"011001000",
  18644=>"100100000",
  18645=>"111000001",
  18646=>"000000000",
  18647=>"000110010",
  18648=>"111111111",
  18649=>"111000001",
  18650=>"111111111",
  18651=>"100000011",
  18652=>"011111111",
  18653=>"000010110",
  18654=>"111001001",
  18655=>"001101000",
  18656=>"101100101",
  18657=>"011011001",
  18658=>"011011010",
  18659=>"111111111",
  18660=>"100101001",
  18661=>"000011001",
  18662=>"011011000",
  18663=>"001000000",
  18664=>"111111100",
  18665=>"000000111",
  18666=>"111111111",
  18667=>"000010011",
  18668=>"000110111",
  18669=>"111011010",
  18670=>"111000100",
  18671=>"111111111",
  18672=>"000000000",
  18673=>"111110100",
  18674=>"000000010",
  18675=>"111011111",
  18676=>"011000101",
  18677=>"111111100",
  18678=>"100100100",
  18679=>"111111011",
  18680=>"001000000",
  18681=>"000111111",
  18682=>"111111111",
  18683=>"000011111",
  18684=>"000000010",
  18685=>"011110100",
  18686=>"011011001",
  18687=>"111111000",
  18688=>"001000101",
  18689=>"000000101",
  18690=>"111111000",
  18691=>"101111111",
  18692=>"111101001",
  18693=>"010010111",
  18694=>"000110110",
  18695=>"000110111",
  18696=>"001000001",
  18697=>"000000001",
  18698=>"001000000",
  18699=>"111111011",
  18700=>"011000000",
  18701=>"001001001",
  18702=>"111111111",
  18703=>"111011000",
  18704=>"111000000",
  18705=>"000110100",
  18706=>"000000011",
  18707=>"000111111",
  18708=>"111111111",
  18709=>"101001001",
  18710=>"110111111",
  18711=>"100000001",
  18712=>"001001101",
  18713=>"000000011",
  18714=>"000000110",
  18715=>"000000111",
  18716=>"111111001",
  18717=>"111111100",
  18718=>"011111000",
  18719=>"011000111",
  18720=>"101101111",
  18721=>"000001000",
  18722=>"000110001",
  18723=>"000111111",
  18724=>"000000011",
  18725=>"000000000",
  18726=>"000100000",
  18727=>"111110100",
  18728=>"000000000",
  18729=>"000100100",
  18730=>"001111111",
  18731=>"011011000",
  18732=>"000001111",
  18733=>"111110100",
  18734=>"111111111",
  18735=>"001000000",
  18736=>"111111101",
  18737=>"111000111",
  18738=>"011111000",
  18739=>"000000000",
  18740=>"111001000",
  18741=>"000000011",
  18742=>"111111000",
  18743=>"000000000",
  18744=>"011011111",
  18745=>"001000011",
  18746=>"111100000",
  18747=>"111110000",
  18748=>"111111000",
  18749=>"111111111",
  18750=>"000100110",
  18751=>"111000111",
  18752=>"100000111",
  18753=>"111111101",
  18754=>"000101111",
  18755=>"000000000",
  18756=>"000111111",
  18757=>"100001011",
  18758=>"110111111",
  18759=>"000001111",
  18760=>"111111101",
  18761=>"011001111",
  18762=>"000000000",
  18763=>"000000000",
  18764=>"111000000",
  18765=>"000001011",
  18766=>"111111111",
  18767=>"000010111",
  18768=>"011011100",
  18769=>"000000001",
  18770=>"111111001",
  18771=>"001010111",
  18772=>"111111111",
  18773=>"000000000",
  18774=>"010000000",
  18775=>"000101100",
  18776=>"110111111",
  18777=>"111101111",
  18778=>"111111111",
  18779=>"001000100",
  18780=>"110100100",
  18781=>"111010000",
  18782=>"110000101",
  18783=>"000000100",
  18784=>"000000001",
  18785=>"101011001",
  18786=>"000100001",
  18787=>"011000000",
  18788=>"000001011",
  18789=>"111111011",
  18790=>"111011000",
  18791=>"001000000",
  18792=>"000010000",
  18793=>"000000000",
  18794=>"111110111",
  18795=>"011011111",
  18796=>"111001001",
  18797=>"010010000",
  18798=>"011111011",
  18799=>"111001100",
  18800=>"011101111",
  18801=>"000010010",
  18802=>"111011011",
  18803=>"000000111",
  18804=>"111111111",
  18805=>"111001001",
  18806=>"111111111",
  18807=>"000000011",
  18808=>"001001000",
  18809=>"100001111",
  18810=>"000011111",
  18811=>"000000000",
  18812=>"111111000",
  18813=>"000000000",
  18814=>"000111010",
  18815=>"000000110",
  18816=>"001000000",
  18817=>"000001011",
  18818=>"100111111",
  18819=>"011111111",
  18820=>"111000000",
  18821=>"011111111",
  18822=>"010111110",
  18823=>"111000000",
  18824=>"000000111",
  18825=>"000000000",
  18826=>"101101111",
  18827=>"000000000",
  18828=>"011010000",
  18829=>"100100100",
  18830=>"111000000",
  18831=>"001000000",
  18832=>"111111111",
  18833=>"000000000",
  18834=>"001001000",
  18835=>"111010110",
  18836=>"000011001",
  18837=>"110000010",
  18838=>"111111000",
  18839=>"111101001",
  18840=>"101001000",
  18841=>"000000111",
  18842=>"000001111",
  18843=>"111100000",
  18844=>"000101001",
  18845=>"111110000",
  18846=>"111100000",
  18847=>"000000011",
  18848=>"111111101",
  18849=>"111000000",
  18850=>"011011000",
  18851=>"111001111",
  18852=>"111111000",
  18853=>"000000000",
  18854=>"111111111",
  18855=>"000000000",
  18856=>"011011001",
  18857=>"011011011",
  18858=>"111111010",
  18859=>"100001111",
  18860=>"111111111",
  18861=>"000000110",
  18862=>"111111001",
  18863=>"101111111",
  18864=>"111100000",
  18865=>"001000000",
  18866=>"000110110",
  18867=>"111000000",
  18868=>"111111000",
  18869=>"000000000",
  18870=>"001000111",
  18871=>"111111000",
  18872=>"000100011",
  18873=>"111111111",
  18874=>"111000000",
  18875=>"000000000",
  18876=>"011111000",
  18877=>"000000111",
  18878=>"011011000",
  18879=>"100100101",
  18880=>"111111111",
  18881=>"100101111",
  18882=>"111111101",
  18883=>"110000111",
  18884=>"111111000",
  18885=>"111000000",
  18886=>"111111111",
  18887=>"011011011",
  18888=>"111000001",
  18889=>"110100100",
  18890=>"111111111",
  18891=>"000001111",
  18892=>"100100111",
  18893=>"000000100",
  18894=>"000000011",
  18895=>"010011001",
  18896=>"111110000",
  18897=>"000000101",
  18898=>"000000001",
  18899=>"000000111",
  18900=>"000100111",
  18901=>"101000000",
  18902=>"111111111",
  18903=>"111111010",
  18904=>"000000100",
  18905=>"111111111",
  18906=>"111111000",
  18907=>"000000000",
  18908=>"000001001",
  18909=>"110000001",
  18910=>"111000111",
  18911=>"100100111",
  18912=>"000000111",
  18913=>"011000000",
  18914=>"000000111",
  18915=>"010111110",
  18916=>"011110111",
  18917=>"001111101",
  18918=>"000000000",
  18919=>"111110010",
  18920=>"011000000",
  18921=>"000011000",
  18922=>"000000011",
  18923=>"100100111",
  18924=>"111001000",
  18925=>"111101111",
  18926=>"111111000",
  18927=>"011000111",
  18928=>"100000100",
  18929=>"000000000",
  18930=>"000111111",
  18931=>"001101100",
  18932=>"000111111",
  18933=>"000000000",
  18934=>"111111001",
  18935=>"100111111",
  18936=>"000010111",
  18937=>"011011001",
  18938=>"111111000",
  18939=>"000011110",
  18940=>"111111111",
  18941=>"001000001",
  18942=>"111111100",
  18943=>"100101001",
  18944=>"001001110",
  18945=>"001001001",
  18946=>"001001111",
  18947=>"001111101",
  18948=>"010110010",
  18949=>"100000101",
  18950=>"110111111",
  18951=>"111111111",
  18952=>"011001011",
  18953=>"000001100",
  18954=>"110110000",
  18955=>"110010011",
  18956=>"000100111",
  18957=>"111111010",
  18958=>"000100100",
  18959=>"110110000",
  18960=>"110000000",
  18961=>"000110100",
  18962=>"000111110",
  18963=>"000000010",
  18964=>"001000001",
  18965=>"000000101",
  18966=>"000010111",
  18967=>"000000101",
  18968=>"111110100",
  18969=>"111110100",
  18970=>"101001111",
  18971=>"001000000",
  18972=>"111000111",
  18973=>"011011001",
  18974=>"011011001",
  18975=>"001001011",
  18976=>"010111111",
  18977=>"111111000",
  18978=>"100110111",
  18979=>"111110000",
  18980=>"101011001",
  18981=>"111111111",
  18982=>"011111011",
  18983=>"101101111",
  18984=>"000000101",
  18985=>"101001000",
  18986=>"000000000",
  18987=>"001000101",
  18988=>"000000011",
  18989=>"010111111",
  18990=>"111000001",
  18991=>"011101000",
  18992=>"010000001",
  18993=>"010000000",
  18994=>"000000000",
  18995=>"000000000",
  18996=>"000000000",
  18997=>"111110000",
  18998=>"000000000",
  18999=>"000000111",
  19000=>"000000000",
  19001=>"000000000",
  19002=>"110110010",
  19003=>"000000011",
  19004=>"001000100",
  19005=>"111110000",
  19006=>"100100000",
  19007=>"110000000",
  19008=>"000110111",
  19009=>"000000001",
  19010=>"110000000",
  19011=>"111100110",
  19012=>"010000000",
  19013=>"111111111",
  19014=>"000000000",
  19015=>"111111111",
  19016=>"011011001",
  19017=>"000000010",
  19018=>"000000100",
  19019=>"000000000",
  19020=>"100000110",
  19021=>"000000111",
  19022=>"000000011",
  19023=>"111111110",
  19024=>"110110110",
  19025=>"111110000",
  19026=>"000000001",
  19027=>"000000000",
  19028=>"000000000",
  19029=>"000001111",
  19030=>"000000000",
  19031=>"000111001",
  19032=>"110110011",
  19033=>"101000111",
  19034=>"000011111",
  19035=>"000000100",
  19036=>"111111111",
  19037=>"111000001",
  19038=>"000000001",
  19039=>"100100100",
  19040=>"001111010",
  19041=>"100000000",
  19042=>"000000111",
  19043=>"000111111",
  19044=>"100000000",
  19045=>"111000000",
  19046=>"000000000",
  19047=>"000000000",
  19048=>"000111111",
  19049=>"001001111",
  19050=>"101001000",
  19051=>"000111011",
  19052=>"111111111",
  19053=>"000000111",
  19054=>"001001111",
  19055=>"110111111",
  19056=>"000000111",
  19057=>"110110111",
  19058=>"000000000",
  19059=>"111100000",
  19060=>"000000000",
  19061=>"000000000",
  19062=>"001001101",
  19063=>"001001001",
  19064=>"111001001",
  19065=>"111011011",
  19066=>"001001000",
  19067=>"011010000",
  19068=>"110110100",
  19069=>"111110110",
  19070=>"111101111",
  19071=>"100111111",
  19072=>"000101111",
  19073=>"011000111",
  19074=>"000100110",
  19075=>"011001100",
  19076=>"001001111",
  19077=>"101000000",
  19078=>"001001110",
  19079=>"001001111",
  19080=>"000001111",
  19081=>"010000010",
  19082=>"010000000",
  19083=>"111010011",
  19084=>"111111111",
  19085=>"100100011",
  19086=>"110110000",
  19087=>"000000100",
  19088=>"001001111",
  19089=>"000000001",
  19090=>"000000000",
  19091=>"111111101",
  19092=>"000000000",
  19093=>"110000000",
  19094=>"000100000",
  19095=>"000000001",
  19096=>"111001001",
  19097=>"111111111",
  19098=>"110110110",
  19099=>"000000000",
  19100=>"100110111",
  19101=>"001000000",
  19102=>"100000000",
  19103=>"001001111",
  19104=>"000001111",
  19105=>"110000000",
  19106=>"001001101",
  19107=>"110111110",
  19108=>"001001001",
  19109=>"101011111",
  19110=>"111001111",
  19111=>"111110000",
  19112=>"101001001",
  19113=>"001000111",
  19114=>"110110101",
  19115=>"000111111",
  19116=>"101000000",
  19117=>"001001001",
  19118=>"101101101",
  19119=>"110110000",
  19120=>"000000000",
  19121=>"100100100",
  19122=>"111111111",
  19123=>"000101001",
  19124=>"111111000",
  19125=>"001000101",
  19126=>"000001101",
  19127=>"000110110",
  19128=>"000000000",
  19129=>"010010111",
  19130=>"001001101",
  19131=>"100100111",
  19132=>"001101111",
  19133=>"111111101",
  19134=>"000000000",
  19135=>"110011001",
  19136=>"110010010",
  19137=>"001000000",
  19138=>"000111010",
  19139=>"111111111",
  19140=>"100001010",
  19141=>"001001101",
  19142=>"111111011",
  19143=>"000000101",
  19144=>"011000000",
  19145=>"111111111",
  19146=>"110000000",
  19147=>"011011111",
  19148=>"101100000",
  19149=>"000001000",
  19150=>"101111111",
  19151=>"001000100",
  19152=>"000010110",
  19153=>"001000000",
  19154=>"111011111",
  19155=>"000000111",
  19156=>"000000000",
  19157=>"000000000",
  19158=>"011000111",
  19159=>"001111111",
  19160=>"000100100",
  19161=>"000000001",
  19162=>"111000000",
  19163=>"101111001",
  19164=>"110110000",
  19165=>"111111000",
  19166=>"111111110",
  19167=>"001001001",
  19168=>"000000000",
  19169=>"011001001",
  19170=>"000110111",
  19171=>"000000101",
  19172=>"010110110",
  19173=>"000000011",
  19174=>"111111111",
  19175=>"110110111",
  19176=>"010111111",
  19177=>"111001000",
  19178=>"100110111",
  19179=>"111101111",
  19180=>"110111111",
  19181=>"000000011",
  19182=>"110110011",
  19183=>"100000101",
  19184=>"010111111",
  19185=>"111111111",
  19186=>"010110111",
  19187=>"000000001",
  19188=>"100000111",
  19189=>"001001011",
  19190=>"111111011",
  19191=>"110000000",
  19192=>"000001111",
  19193=>"110111111",
  19194=>"100010110",
  19195=>"011111011",
  19196=>"100111111",
  19197=>"110110110",
  19198=>"111001001",
  19199=>"000000000",
  19200=>"101000001",
  19201=>"100101101",
  19202=>"110110111",
  19203=>"111111110",
  19204=>"110101000",
  19205=>"000000000",
  19206=>"111111011",
  19207=>"110010000",
  19208=>"000000100",
  19209=>"001111111",
  19210=>"000000101",
  19211=>"000101111",
  19212=>"101000111",
  19213=>"110000000",
  19214=>"000000000",
  19215=>"000000000",
  19216=>"000000110",
  19217=>"000000101",
  19218=>"000000000",
  19219=>"110110010",
  19220=>"010010110",
  19221=>"110010000",
  19222=>"001100111",
  19223=>"010000000",
  19224=>"111001001",
  19225=>"001111111",
  19226=>"111111110",
  19227=>"000111110",
  19228=>"000000000",
  19229=>"011000000",
  19230=>"010000010",
  19231=>"111111110",
  19232=>"110111000",
  19233=>"111111001",
  19234=>"110010000",
  19235=>"110110111",
  19236=>"101001000",
  19237=>"000000000",
  19238=>"101111100",
  19239=>"110110010",
  19240=>"001000000",
  19241=>"110111111",
  19242=>"110110010",
  19243=>"010010011",
  19244=>"111111011",
  19245=>"111111111",
  19246=>"000000010",
  19247=>"000001110",
  19248=>"100110010",
  19249=>"000000000",
  19250=>"001001001",
  19251=>"011000000",
  19252=>"000100000",
  19253=>"001000011",
  19254=>"110110111",
  19255=>"110111111",
  19256=>"000111011",
  19257=>"111001111",
  19258=>"010001000",
  19259=>"111111111",
  19260=>"000000000",
  19261=>"001101001",
  19262=>"000000000",
  19263=>"000000101",
  19264=>"010011011",
  19265=>"111101000",
  19266=>"100000000",
  19267=>"000000000",
  19268=>"000000000",
  19269=>"111111111",
  19270=>"111111111",
  19271=>"000110110",
  19272=>"111000000",
  19273=>"000001000",
  19274=>"001111111",
  19275=>"110110100",
  19276=>"000000000",
  19277=>"000001111",
  19278=>"000000000",
  19279=>"111111000",
  19280=>"000000000",
  19281=>"000000001",
  19282=>"111000100",
  19283=>"101101001",
  19284=>"000000000",
  19285=>"011011011",
  19286=>"111001000",
  19287=>"111110111",
  19288=>"000001011",
  19289=>"000110111",
  19290=>"110110110",
  19291=>"000000111",
  19292=>"010001111",
  19293=>"000000000",
  19294=>"000001101",
  19295=>"110110110",
  19296=>"100101001",
  19297=>"000000111",
  19298=>"110100100",
  19299=>"101100101",
  19300=>"000100110",
  19301=>"111111000",
  19302=>"111010010",
  19303=>"000000001",
  19304=>"011111111",
  19305=>"011010011",
  19306=>"111111111",
  19307=>"000000111",
  19308=>"000110111",
  19309=>"001100110",
  19310=>"000000110",
  19311=>"110111111",
  19312=>"110100110",
  19313=>"010111000",
  19314=>"110000000",
  19315=>"110110110",
  19316=>"010011011",
  19317=>"000000000",
  19318=>"000000000",
  19319=>"001001001",
  19320=>"000000000",
  19321=>"111001101",
  19322=>"011111001",
  19323=>"001001000",
  19324=>"110110110",
  19325=>"000000111",
  19326=>"000000101",
  19327=>"000100000",
  19328=>"000110110",
  19329=>"110110111",
  19330=>"111101100",
  19331=>"000000000",
  19332=>"110001001",
  19333=>"011111011",
  19334=>"000000001",
  19335=>"001001111",
  19336=>"000001001",
  19337=>"000000110",
  19338=>"000000000",
  19339=>"000011011",
  19340=>"111001111",
  19341=>"111111111",
  19342=>"000110111",
  19343=>"111010000",
  19344=>"000000001",
  19345=>"100100111",
  19346=>"110110111",
  19347=>"000000000",
  19348=>"001001011",
  19349=>"000000000",
  19350=>"010100110",
  19351=>"001001011",
  19352=>"001111111",
  19353=>"000000000",
  19354=>"000001111",
  19355=>"000000001",
  19356=>"111111111",
  19357=>"111001111",
  19358=>"001001001",
  19359=>"111111111",
  19360=>"111111111",
  19361=>"111111111",
  19362=>"000000010",
  19363=>"111001111",
  19364=>"100100001",
  19365=>"111011000",
  19366=>"111000001",
  19367=>"010010010",
  19368=>"111111111",
  19369=>"110000000",
  19370=>"010000111",
  19371=>"000000001",
  19372=>"100110110",
  19373=>"000000100",
  19374=>"100000000",
  19375=>"111111111",
  19376=>"100000100",
  19377=>"000000000",
  19378=>"111111111",
  19379=>"110111100",
  19380=>"111111010",
  19381=>"111000000",
  19382=>"111111111",
  19383=>"100000000",
  19384=>"001001111",
  19385=>"110111110",
  19386=>"111100100",
  19387=>"001001000",
  19388=>"111001001",
  19389=>"000000111",
  19390=>"000110101",
  19391=>"000000110",
  19392=>"000000011",
  19393=>"011001111",
  19394=>"000010011",
  19395=>"011111111",
  19396=>"110110010",
  19397=>"101001000",
  19398=>"001001001",
  19399=>"001011111",
  19400=>"000000000",
  19401=>"001001111",
  19402=>"001101101",
  19403=>"100100000",
  19404=>"111111011",
  19405=>"111111111",
  19406=>"000000000",
  19407=>"001001001",
  19408=>"000000001",
  19409=>"011011000",
  19410=>"111111111",
  19411=>"011001100",
  19412=>"000000100",
  19413=>"111111110",
  19414=>"000010001",
  19415=>"010111111",
  19416=>"000000000",
  19417=>"110110110",
  19418=>"111111100",
  19419=>"000000101",
  19420=>"100111101",
  19421=>"111101101",
  19422=>"111111001",
  19423=>"100111111",
  19424=>"001001111",
  19425=>"111011110",
  19426=>"000001011",
  19427=>"100000011",
  19428=>"111101001",
  19429=>"111111001",
  19430=>"110110010",
  19431=>"111001000",
  19432=>"000000000",
  19433=>"110110111",
  19434=>"001000000",
  19435=>"111110000",
  19436=>"111111111",
  19437=>"000000100",
  19438=>"001111000",
  19439=>"111111010",
  19440=>"001001001",
  19441=>"100110110",
  19442=>"110110010",
  19443=>"111100000",
  19444=>"111111111",
  19445=>"111111011",
  19446=>"000010011",
  19447=>"011001011",
  19448=>"111001011",
  19449=>"000000100",
  19450=>"000000111",
  19451=>"101111111",
  19452=>"000001011",
  19453=>"001011111",
  19454=>"000110000",
  19455=>"000000001",
  19456=>"000010110",
  19457=>"000110111",
  19458=>"111000011",
  19459=>"000111000",
  19460=>"111111110",
  19461=>"000000101",
  19462=>"000000111",
  19463=>"111111111",
  19464=>"111111111",
  19465=>"110100000",
  19466=>"000111111",
  19467=>"000010000",
  19468=>"111110100",
  19469=>"000000000",
  19470=>"010011111",
  19471=>"000110111",
  19472=>"111111110",
  19473=>"000000011",
  19474=>"111000000",
  19475=>"011000000",
  19476=>"000000000",
  19477=>"111101111",
  19478=>"011111111",
  19479=>"001001000",
  19480=>"000000000",
  19481=>"001000000",
  19482=>"111100100",
  19483=>"110111111",
  19484=>"011010111",
  19485=>"111000000",
  19486=>"110001001",
  19487=>"000000000",
  19488=>"001000000",
  19489=>"111000111",
  19490=>"111111011",
  19491=>"000000000",
  19492=>"111001001",
  19493=>"110100000",
  19494=>"100100000",
  19495=>"111101001",
  19496=>"000001011",
  19497=>"111100111",
  19498=>"011011001",
  19499=>"111111011",
  19500=>"000000011",
  19501=>"111111111",
  19502=>"110010000",
  19503=>"010000011",
  19504=>"111111110",
  19505=>"000111101",
  19506=>"000111111",
  19507=>"000000000",
  19508=>"110100000",
  19509=>"110111111",
  19510=>"000000000",
  19511=>"110000001",
  19512=>"111011111",
  19513=>"111111000",
  19514=>"111001000",
  19515=>"000100000",
  19516=>"000000011",
  19517=>"000010000",
  19518=>"000110000",
  19519=>"111000111",
  19520=>"111011000",
  19521=>"111111110",
  19522=>"010111111",
  19523=>"001001000",
  19524=>"110111011",
  19525=>"000000111",
  19526=>"111000000",
  19527=>"111111000",
  19528=>"011011011",
  19529=>"000000000",
  19530=>"111111111",
  19531=>"000000001",
  19532=>"000001011",
  19533=>"000000000",
  19534=>"100000000",
  19535=>"110000000",
  19536=>"000000110",
  19537=>"100000001",
  19538=>"111111111",
  19539=>"010110111",
  19540=>"000111000",
  19541=>"111111111",
  19542=>"111001001",
  19543=>"000000011",
  19544=>"010111110",
  19545=>"111001111",
  19546=>"100111111",
  19547=>"001000000",
  19548=>"101101100",
  19549=>"111111111",
  19550=>"001000000",
  19551=>"110110000",
  19552=>"000000000",
  19553=>"000000000",
  19554=>"111111000",
  19555=>"111000001",
  19556=>"111111010",
  19557=>"001000111",
  19558=>"000100000",
  19559=>"111111110",
  19560=>"000000000",
  19561=>"000000000",
  19562=>"001000110",
  19563=>"111110010",
  19564=>"000001000",
  19565=>"111000001",
  19566=>"000000111",
  19567=>"000000000",
  19568=>"000000000",
  19569=>"001001000",
  19570=>"100110000",
  19571=>"101111111",
  19572=>"000001001",
  19573=>"111111000",
  19574=>"010001111",
  19575=>"000100000",
  19576=>"001000000",
  19577=>"000000000",
  19578=>"111111000",
  19579=>"111000000",
  19580=>"000011111",
  19581=>"100100110",
  19582=>"000000001",
  19583=>"000001001",
  19584=>"100000000",
  19585=>"000000111",
  19586=>"100100000",
  19587=>"110111111",
  19588=>"111111111",
  19589=>"000000111",
  19590=>"110011010",
  19591=>"000000111",
  19592=>"000111111",
  19593=>"001100110",
  19594=>"000000111",
  19595=>"111111111",
  19596=>"110111111",
  19597=>"000110111",
  19598=>"100000000",
  19599=>"111000110",
  19600=>"000001000",
  19601=>"000111111",
  19602=>"000000001",
  19603=>"011111111",
  19604=>"000000000",
  19605=>"111110000",
  19606=>"000000110",
  19607=>"111000000",
  19608=>"000000000",
  19609=>"110100111",
  19610=>"111111000",
  19611=>"110100111",
  19612=>"000000000",
  19613=>"001111100",
  19614=>"111111110",
  19615=>"010000111",
  19616=>"100000000",
  19617=>"111111111",
  19618=>"000011111",
  19619=>"111111111",
  19620=>"011001000",
  19621=>"000000111",
  19622=>"110111111",
  19623=>"011010000",
  19624=>"011111111",
  19625=>"111111101",
  19626=>"000000000",
  19627=>"000110110",
  19628=>"110111000",
  19629=>"111010000",
  19630=>"101111001",
  19631=>"111111001",
  19632=>"000100011",
  19633=>"000000000",
  19634=>"011111001",
  19635=>"000000001",
  19636=>"110110110",
  19637=>"001111111",
  19638=>"000100110",
  19639=>"010010110",
  19640=>"111111111",
  19641=>"000000000",
  19642=>"000000010",
  19643=>"111111111",
  19644=>"000000111",
  19645=>"001111111",
  19646=>"110111101",
  19647=>"000000111",
  19648=>"100000000",
  19649=>"111000110",
  19650=>"001001011",
  19651=>"000111111",
  19652=>"000000000",
  19653=>"111111000",
  19654=>"011111111",
  19655=>"111110110",
  19656=>"101001011",
  19657=>"011111000",
  19658=>"000000001",
  19659=>"000000111",
  19660=>"000000000",
  19661=>"000000000",
  19662=>"111111111",
  19663=>"000000000",
  19664=>"001001101",
  19665=>"000000000",
  19666=>"000000111",
  19667=>"111000011",
  19668=>"000000100",
  19669=>"110011001",
  19670=>"110000000",
  19671=>"000000000",
  19672=>"011001111",
  19673=>"010000111",
  19674=>"000000000",
  19675=>"000000010",
  19676=>"100000000",
  19677=>"000000000",
  19678=>"111000001",
  19679=>"000000110",
  19680=>"111101111",
  19681=>"001000000",
  19682=>"110000110",
  19683=>"101111111",
  19684=>"011101111",
  19685=>"100000001",
  19686=>"110000000",
  19687=>"010111111",
  19688=>"011011011",
  19689=>"000000100",
  19690=>"000111111",
  19691=>"101000000",
  19692=>"111111111",
  19693=>"000000110",
  19694=>"001000000",
  19695=>"000111110",
  19696=>"111000000",
  19697=>"000111000",
  19698=>"001011111",
  19699=>"000000110",
  19700=>"000000000",
  19701=>"011011000",
  19702=>"001000001",
  19703=>"110000000",
  19704=>"101001111",
  19705=>"000000000",
  19706=>"100000000",
  19707=>"111100000",
  19708=>"111111000",
  19709=>"111011011",
  19710=>"100000000",
  19711=>"111010000",
  19712=>"101110111",
  19713=>"111010010",
  19714=>"111100100",
  19715=>"111100000",
  19716=>"111011111",
  19717=>"111101101",
  19718=>"000000000",
  19719=>"111111111",
  19720=>"111110110",
  19721=>"000111001",
  19722=>"000000011",
  19723=>"110110100",
  19724=>"001000111",
  19725=>"000000000",
  19726=>"000000000",
  19727=>"000111001",
  19728=>"010000000",
  19729=>"100111111",
  19730=>"001000000",
  19731=>"111111111",
  19732=>"010000111",
  19733=>"111111100",
  19734=>"011001011",
  19735=>"111110000",
  19736=>"111111111",
  19737=>"000001111",
  19738=>"000000000",
  19739=>"000000000",
  19740=>"110110010",
  19741=>"111111111",
  19742=>"000110111",
  19743=>"100100111",
  19744=>"011111111",
  19745=>"110110000",
  19746=>"000000011",
  19747=>"001011000",
  19748=>"000000000",
  19749=>"000000000",
  19750=>"000111111",
  19751=>"000000000",
  19752=>"111111011",
  19753=>"010111100",
  19754=>"111001000",
  19755=>"000000101",
  19756=>"001000000",
  19757=>"000001000",
  19758=>"111111111",
  19759=>"000111000",
  19760=>"000000000",
  19761=>"111100000",
  19762=>"111010000",
  19763=>"000000001",
  19764=>"111111111",
  19765=>"000001101",
  19766=>"101100110",
  19767=>"000000000",
  19768=>"111111111",
  19769=>"000000000",
  19770=>"000000111",
  19771=>"110110111",
  19772=>"000000000",
  19773=>"000000100",
  19774=>"111111111",
  19775=>"000111111",
  19776=>"111111111",
  19777=>"101111000",
  19778=>"111001000",
  19779=>"101111000",
  19780=>"100110001",
  19781=>"100110111",
  19782=>"010111110",
  19783=>"111111111",
  19784=>"000100000",
  19785=>"111000001",
  19786=>"110111111",
  19787=>"111001001",
  19788=>"111001000",
  19789=>"000000000",
  19790=>"000101111",
  19791=>"000000000",
  19792=>"000000001",
  19793=>"100111111",
  19794=>"111111111",
  19795=>"110111100",
  19796=>"000000000",
  19797=>"001010001",
  19798=>"000111111",
  19799=>"111110100",
  19800=>"000101111",
  19801=>"111111111",
  19802=>"000111001",
  19803=>"100010010",
  19804=>"001001000",
  19805=>"000101001",
  19806=>"111000000",
  19807=>"000110111",
  19808=>"111111111",
  19809=>"000000000",
  19810=>"111100000",
  19811=>"000000000",
  19812=>"010011110",
  19813=>"000111000",
  19814=>"000000000",
  19815=>"011011000",
  19816=>"111000000",
  19817=>"000000111",
  19818=>"111111000",
  19819=>"000011111",
  19820=>"111100100",
  19821=>"010111110",
  19822=>"111010000",
  19823=>"001001001",
  19824=>"111111000",
  19825=>"000110000",
  19826=>"001001001",
  19827=>"110100001",
  19828=>"000000000",
  19829=>"111111001",
  19830=>"000010111",
  19831=>"111001000",
  19832=>"110110110",
  19833=>"000000111",
  19834=>"000000000",
  19835=>"100000110",
  19836=>"111111111",
  19837=>"110110111",
  19838=>"111000000",
  19839=>"111000000",
  19840=>"001011000",
  19841=>"111111000",
  19842=>"100100110",
  19843=>"000000000",
  19844=>"111011000",
  19845=>"000000000",
  19846=>"111000001",
  19847=>"000111111",
  19848=>"101000000",
  19849=>"000100111",
  19850=>"000000100",
  19851=>"110000100",
  19852=>"111111111",
  19853=>"111110110",
  19854=>"111000000",
  19855=>"011011000",
  19856=>"000111101",
  19857=>"011000011",
  19858=>"100000001",
  19859=>"000000001",
  19860=>"111111111",
  19861=>"000011000",
  19862=>"111010010",
  19863=>"010111110",
  19864=>"110111110",
  19865=>"011000000",
  19866=>"111110111",
  19867=>"000011000",
  19868=>"011011001",
  19869=>"000001001",
  19870=>"000000000",
  19871=>"000000000",
  19872=>"000000000",
  19873=>"010000100",
  19874=>"000000111",
  19875=>"001111101",
  19876=>"111000000",
  19877=>"111111111",
  19878=>"000001111",
  19879=>"000111001",
  19880=>"100100111",
  19881=>"110001001",
  19882=>"111111111",
  19883=>"000000000",
  19884=>"000000000",
  19885=>"000000100",
  19886=>"101000000",
  19887=>"000111111",
  19888=>"111111111",
  19889=>"001000000",
  19890=>"110111111",
  19891=>"000000000",
  19892=>"000101111",
  19893=>"111100111",
  19894=>"011011011",
  19895=>"000000100",
  19896=>"001001001",
  19897=>"001000001",
  19898=>"011110110",
  19899=>"111001000",
  19900=>"111111111",
  19901=>"111111111",
  19902=>"011001000",
  19903=>"011000000",
  19904=>"111111111",
  19905=>"000111001",
  19906=>"000000000",
  19907=>"011010010",
  19908=>"000000001",
  19909=>"011111111",
  19910=>"100010000",
  19911=>"111111000",
  19912=>"111010000",
  19913=>"001000000",
  19914=>"101101000",
  19915=>"000101111",
  19916=>"000000110",
  19917=>"111000111",
  19918=>"000000010",
  19919=>"111000000",
  19920=>"111101000",
  19921=>"111111111",
  19922=>"000000000",
  19923=>"011010000",
  19924=>"000000000",
  19925=>"111010000",
  19926=>"000000000",
  19927=>"110110000",
  19928=>"000100111",
  19929=>"101111111",
  19930=>"111111111",
  19931=>"000111101",
  19932=>"111111011",
  19933=>"000000111",
  19934=>"111101000",
  19935=>"001000000",
  19936=>"110111111",
  19937=>"010000000",
  19938=>"000111111",
  19939=>"111100000",
  19940=>"001001111",
  19941=>"101000010",
  19942=>"000000100",
  19943=>"111110000",
  19944=>"100000000",
  19945=>"000100111",
  19946=>"111000100",
  19947=>"111111111",
  19948=>"111111011",
  19949=>"110110111",
  19950=>"111111111",
  19951=>"111000010",
  19952=>"000111010",
  19953=>"000000000",
  19954=>"001000000",
  19955=>"110111000",
  19956=>"011000001",
  19957=>"000000000",
  19958=>"110111111",
  19959=>"110110110",
  19960=>"001011111",
  19961=>"100001001",
  19962=>"111000000",
  19963=>"111111101",
  19964=>"101000110",
  19965=>"111110000",
  19966=>"000101111",
  19967=>"111011011",
  19968=>"111001000",
  19969=>"111101001",
  19970=>"111011000",
  19971=>"111111111",
  19972=>"111110110",
  19973=>"110111111",
  19974=>"111000001",
  19975=>"111000000",
  19976=>"000000000",
  19977=>"010111111",
  19978=>"000000000",
  19979=>"000000000",
  19980=>"011001011",
  19981=>"001011111",
  19982=>"101101101",
  19983=>"100111111",
  19984=>"000111111",
  19985=>"100110111",
  19986=>"000000111",
  19987=>"000000000",
  19988=>"000000000",
  19989=>"001001111",
  19990=>"000011011",
  19991=>"001001011",
  19992=>"110110111",
  19993=>"000010111",
  19994=>"000000000",
  19995=>"000000011",
  19996=>"000000000",
  19997=>"111111111",
  19998=>"011001001",
  19999=>"100100000",
  20000=>"111111110",
  20001=>"110111111",
  20002=>"111100000",
  20003=>"111111001",
  20004=>"000000000",
  20005=>"111011001",
  20006=>"000000000",
  20007=>"000000000",
  20008=>"000000000",
  20009=>"111111111",
  20010=>"000000000",
  20011=>"101111111",
  20012=>"111101111",
  20013=>"001000000",
  20014=>"000000000",
  20015=>"001000000",
  20016=>"111111011",
  20017=>"011011111",
  20018=>"000000011",
  20019=>"000000000",
  20020=>"111111111",
  20021=>"010111111",
  20022=>"111011011",
  20023=>"000000000",
  20024=>"001111111",
  20025=>"000001000",
  20026=>"001000110",
  20027=>"000000000",
  20028=>"000000000",
  20029=>"111101001",
  20030=>"101110110",
  20031=>"100100110",
  20032=>"110101011",
  20033=>"000101101",
  20034=>"001111010",
  20035=>"100110111",
  20036=>"001001001",
  20037=>"111111110",
  20038=>"111111000",
  20039=>"000000000",
  20040=>"111111011",
  20041=>"000111000",
  20042=>"110111111",
  20043=>"000001000",
  20044=>"000100110",
  20045=>"000000001",
  20046=>"111010000",
  20047=>"011000000",
  20048=>"000011010",
  20049=>"100101101",
  20050=>"111111011",
  20051=>"111111111",
  20052=>"111111100",
  20053=>"010010000",
  20054=>"111001111",
  20055=>"111111111",
  20056=>"000000110",
  20057=>"000110111",
  20058=>"100111111",
  20059=>"100100110",
  20060=>"000000000",
  20061=>"000001111",
  20062=>"100110111",
  20063=>"000000000",
  20064=>"000000101",
  20065=>"000000110",
  20066=>"111010111",
  20067=>"000000000",
  20068=>"000010110",
  20069=>"100100101",
  20070=>"111111111",
  20071=>"111111110",
  20072=>"111111111",
  20073=>"111111111",
  20074=>"111011111",
  20075=>"000001000",
  20076=>"111111100",
  20077=>"100110110",
  20078=>"111111000",
  20079=>"000001001",
  20080=>"110111001",
  20081=>"011011000",
  20082=>"011111111",
  20083=>"000000000",
  20084=>"000000000",
  20085=>"111111000",
  20086=>"000111111",
  20087=>"111100100",
  20088=>"000000000",
  20089=>"000000000",
  20090=>"111111111",
  20091=>"000000000",
  20092=>"111110110",
  20093=>"111111010",
  20094=>"000000001",
  20095=>"000000000",
  20096=>"000000000",
  20097=>"011000000",
  20098=>"000000000",
  20099=>"010000010",
  20100=>"111111011",
  20101=>"111000000",
  20102=>"110110000",
  20103=>"011111000",
  20104=>"000101111",
  20105=>"000000000",
  20106=>"000100111",
  20107=>"000001111",
  20108=>"110011000",
  20109=>"111110111",
  20110=>"000000100",
  20111=>"100001000",
  20112=>"110111111",
  20113=>"111111110",
  20114=>"000000000",
  20115=>"101100111",
  20116=>"100111111",
  20117=>"001001000",
  20118=>"111111011",
  20119=>"110111111",
  20120=>"110111110",
  20121=>"000000000",
  20122=>"100000000",
  20123=>"110110110",
  20124=>"111111111",
  20125=>"110110010",
  20126=>"000000000",
  20127=>"111001001",
  20128=>"111111001",
  20129=>"001000000",
  20130=>"111111110",
  20131=>"111111111",
  20132=>"110001001",
  20133=>"000000110",
  20134=>"111111111",
  20135=>"111011000",
  20136=>"000001001",
  20137=>"000000000",
  20138=>"000000000",
  20139=>"000000111",
  20140=>"010111010",
  20141=>"111111111",
  20142=>"111001011",
  20143=>"000000000",
  20144=>"110110111",
  20145=>"110110100",
  20146=>"111111111",
  20147=>"000111111",
  20148=>"111111000",
  20149=>"111111111",
  20150=>"000111011",
  20151=>"001000000",
  20152=>"111110010",
  20153=>"101001000",
  20154=>"111000111",
  20155=>"110111011",
  20156=>"111111101",
  20157=>"111111111",
  20158=>"111000000",
  20159=>"000001000",
  20160=>"011011011",
  20161=>"111010110",
  20162=>"001000000",
  20163=>"000000000",
  20164=>"000000000",
  20165=>"100111110",
  20166=>"010111111",
  20167=>"000000000",
  20168=>"000011000",
  20169=>"001011111",
  20170=>"010010000",
  20171=>"011001111",
  20172=>"000000000",
  20173=>"111111011",
  20174=>"111011001",
  20175=>"011111011",
  20176=>"111111110",
  20177=>"001001001",
  20178=>"111111111",
  20179=>"000000000",
  20180=>"111000000",
  20181=>"111110111",
  20182=>"000001000",
  20183=>"111111111",
  20184=>"011111000",
  20185=>"000000010",
  20186=>"111110000",
  20187=>"111111111",
  20188=>"001000001",
  20189=>"000010010",
  20190=>"011111111",
  20191=>"000001101",
  20192=>"000000000",
  20193=>"000100111",
  20194=>"101001001",
  20195=>"110000001",
  20196=>"100100110",
  20197=>"000000010",
  20198=>"011011000",
  20199=>"111011011",
  20200=>"011111011",
  20201=>"110110000",
  20202=>"111111111",
  20203=>"111111101",
  20204=>"000000000",
  20205=>"111111111",
  20206=>"000000110",
  20207=>"111111000",
  20208=>"000000010",
  20209=>"100111001",
  20210=>"100100111",
  20211=>"111100110",
  20212=>"111111111",
  20213=>"001001000",
  20214=>"001011011",
  20215=>"111111111",
  20216=>"001001000",
  20217=>"000000000",
  20218=>"000000010",
  20219=>"000000000",
  20220=>"000000110",
  20221=>"000111011",
  20222=>"111111111",
  20223=>"110010111",
  20224=>"000000111",
  20225=>"011011111",
  20226=>"101111111",
  20227=>"011111111",
  20228=>"000000000",
  20229=>"100000000",
  20230=>"111000000",
  20231=>"010010111",
  20232=>"101111111",
  20233=>"000101111",
  20234=>"000000000",
  20235=>"110000000",
  20236=>"001001001",
  20237=>"000000000",
  20238=>"111111111",
  20239=>"000000000",
  20240=>"100000001",
  20241=>"011000011",
  20242=>"000000000",
  20243=>"111011011",
  20244=>"000001011",
  20245=>"111111001",
  20246=>"111111111",
  20247=>"111111111",
  20248=>"111111111",
  20249=>"100000000",
  20250=>"011111111",
  20251=>"100000000",
  20252=>"111111110",
  20253=>"101111101",
  20254=>"001000000",
  20255=>"100000011",
  20256=>"011011011",
  20257=>"110110110",
  20258=>"000011011",
  20259=>"011000111",
  20260=>"000000001",
  20261=>"000000110",
  20262=>"000000000",
  20263=>"110111111",
  20264=>"111111111",
  20265=>"111111111",
  20266=>"000001011",
  20267=>"000000000",
  20268=>"111111111",
  20269=>"011011111",
  20270=>"111111111",
  20271=>"000000101",
  20272=>"000000000",
  20273=>"111000000",
  20274=>"011100111",
  20275=>"001111111",
  20276=>"111000000",
  20277=>"111010000",
  20278=>"111111101",
  20279=>"111111111",
  20280=>"000000000",
  20281=>"111111000",
  20282=>"000111111",
  20283=>"000001000",
  20284=>"000000000",
  20285=>"111000100",
  20286=>"111001001",
  20287=>"000000110",
  20288=>"000000110",
  20289=>"111001001",
  20290=>"100000000",
  20291=>"111000000",
  20292=>"000000000",
  20293=>"101111111",
  20294=>"111111111",
  20295=>"000000000",
  20296=>"000000001",
  20297=>"000000000",
  20298=>"110000000",
  20299=>"000000000",
  20300=>"011000000",
  20301=>"011001000",
  20302=>"111111111",
  20303=>"101000000",
  20304=>"110100110",
  20305=>"110110111",
  20306=>"100000100",
  20307=>"000110110",
  20308=>"000000010",
  20309=>"100100100",
  20310=>"000000000",
  20311=>"000000001",
  20312=>"000000000",
  20313=>"110000000",
  20314=>"000001111",
  20315=>"100110111",
  20316=>"010000000",
  20317=>"000000000",
  20318=>"000000000",
  20319=>"111111111",
  20320=>"000000000",
  20321=>"111111111",
  20322=>"000110110",
  20323=>"110000000",
  20324=>"001001011",
  20325=>"111111111",
  20326=>"001000000",
  20327=>"000000000",
  20328=>"001001001",
  20329=>"000000000",
  20330=>"000000000",
  20331=>"000000000",
  20332=>"110000000",
  20333=>"111100100",
  20334=>"111111000",
  20335=>"000000000",
  20336=>"010111111",
  20337=>"111001000",
  20338=>"111111110",
  20339=>"100100110",
  20340=>"111111111",
  20341=>"101101100",
  20342=>"100110000",
  20343=>"000000101",
  20344=>"110000000",
  20345=>"000000000",
  20346=>"000000000",
  20347=>"111101111",
  20348=>"111111100",
  20349=>"001000000",
  20350=>"000000000",
  20351=>"111111111",
  20352=>"111011011",
  20353=>"111011001",
  20354=>"111101100",
  20355=>"111111111",
  20356=>"000111111",
  20357=>"111111100",
  20358=>"011011110",
  20359=>"000000101",
  20360=>"111111111",
  20361=>"000000001",
  20362=>"000000000",
  20363=>"000110111",
  20364=>"111111111",
  20365=>"001000000",
  20366=>"000000010",
  20367=>"000000001",
  20368=>"000000111",
  20369=>"111100100",
  20370=>"010000000",
  20371=>"000000000",
  20372=>"000000111",
  20373=>"100100000",
  20374=>"011111011",
  20375=>"111111110",
  20376=>"111111111",
  20377=>"100100111",
  20378=>"000000100",
  20379=>"000110001",
  20380=>"111111111",
  20381=>"111011111",
  20382=>"111111111",
  20383=>"000000000",
  20384=>"111111101",
  20385=>"011111111",
  20386=>"111111111",
  20387=>"110111111",
  20388=>"111011001",
  20389=>"000000000",
  20390=>"000000000",
  20391=>"000111111",
  20392=>"000000001",
  20393=>"111111111",
  20394=>"111000000",
  20395=>"000000000",
  20396=>"011000000",
  20397=>"001100111",
  20398=>"000001111",
  20399=>"100000111",
  20400=>"010111111",
  20401=>"000000000",
  20402=>"111000000",
  20403=>"100000111",
  20404=>"000000000",
  20405=>"100111111",
  20406=>"100000000",
  20407=>"000010111",
  20408=>"000000100",
  20409=>"000001011",
  20410=>"011000111",
  20411=>"111111111",
  20412=>"000000000",
  20413=>"111011111",
  20414=>"000000000",
  20415=>"111011111",
  20416=>"000000000",
  20417=>"001000000",
  20418=>"000000000",
  20419=>"111111111",
  20420=>"111110110",
  20421=>"111111111",
  20422=>"111001001",
  20423=>"100100011",
  20424=>"000000000",
  20425=>"000101110",
  20426=>"100010000",
  20427=>"111111011",
  20428=>"000000011",
  20429=>"101011111",
  20430=>"001000000",
  20431=>"000000000",
  20432=>"000000000",
  20433=>"101101001",
  20434=>"001111100",
  20435=>"111111101",
  20436=>"111100110",
  20437=>"011011111",
  20438=>"110000111",
  20439=>"100100110",
  20440=>"110111111",
  20441=>"011001011",
  20442=>"001001011",
  20443=>"111111111",
  20444=>"011001001",
  20445=>"000001011",
  20446=>"111011001",
  20447=>"001000111",
  20448=>"000100000",
  20449=>"110110111",
  20450=>"000110111",
  20451=>"111000000",
  20452=>"000000111",
  20453=>"000001001",
  20454=>"000000010",
  20455=>"000000000",
  20456=>"000000011",
  20457=>"111111111",
  20458=>"111111101",
  20459=>"000001000",
  20460=>"011001011",
  20461=>"111111111",
  20462=>"000000000",
  20463=>"111111111",
  20464=>"111101011",
  20465=>"000101111",
  20466=>"111111111",
  20467=>"111111110",
  20468=>"011011111",
  20469=>"000000000",
  20470=>"011111101",
  20471=>"000011011",
  20472=>"000000000",
  20473=>"001000111",
  20474=>"111111000",
  20475=>"111111111",
  20476=>"000000000",
  20477=>"000000000",
  20478=>"001011000",
  20479=>"000000000",
  20480=>"101111111",
  20481=>"100111100",
  20482=>"000000111",
  20483=>"101000000",
  20484=>"111111111",
  20485=>"010010000",
  20486=>"000000000",
  20487=>"100100101",
  20488=>"000100111",
  20489=>"111111111",
  20490=>"111111111",
  20491=>"011011001",
  20492=>"000000001",
  20493=>"111000100",
  20494=>"000111101",
  20495=>"000111100",
  20496=>"111000000",
  20497=>"011111111",
  20498=>"011001111",
  20499=>"001011000",
  20500=>"111111000",
  20501=>"000000000",
  20502=>"111000000",
  20503=>"001011111",
  20504=>"111111110",
  20505=>"110011001",
  20506=>"111111110",
  20507=>"000000001",
  20508=>"010111011",
  20509=>"000000000",
  20510=>"111001001",
  20511=>"110110111",
  20512=>"000100000",
  20513=>"000000001",
  20514=>"100100111",
  20515=>"110111111",
  20516=>"111111111",
  20517=>"000000000",
  20518=>"011011000",
  20519=>"011001000",
  20520=>"000000000",
  20521=>"000000000",
  20522=>"111111111",
  20523=>"111111111",
  20524=>"000000100",
  20525=>"111000000",
  20526=>"111001001",
  20527=>"010000100",
  20528=>"101000011",
  20529=>"110111111",
  20530=>"111111111",
  20531=>"001000000",
  20532=>"101100110",
  20533=>"000000001",
  20534=>"111000000",
  20535=>"111010011",
  20536=>"111111001",
  20537=>"000000000",
  20538=>"000000000",
  20539=>"001000000",
  20540=>"000100111",
  20541=>"111111111",
  20542=>"010010111",
  20543=>"000111111",
  20544=>"000100100",
  20545=>"110110110",
  20546=>"001010000",
  20547=>"000000000",
  20548=>"110110110",
  20549=>"001111111",
  20550=>"000000000",
  20551=>"000000000",
  20552=>"011011111",
  20553=>"000000000",
  20554=>"000100110",
  20555=>"101000000",
  20556=>"000000001",
  20557=>"000000000",
  20558=>"110111000",
  20559=>"000000110",
  20560=>"111000000",
  20561=>"000000000",
  20562=>"000000110",
  20563=>"101001111",
  20564=>"001001111",
  20565=>"111111111",
  20566=>"111111111",
  20567=>"111111111",
  20568=>"000110111",
  20569=>"000000000",
  20570=>"010111111",
  20571=>"001001111",
  20572=>"011111111",
  20573=>"010000111",
  20574=>"111111111",
  20575=>"100110110",
  20576=>"110100000",
  20577=>"111111111",
  20578=>"001111001",
  20579=>"110100000",
  20580=>"000001000",
  20581=>"000000000",
  20582=>"111111111",
  20583=>"111111100",
  20584=>"000111111",
  20585=>"000000111",
  20586=>"111111001",
  20587=>"010110111",
  20588=>"011011111",
  20589=>"000000010",
  20590=>"111111111",
  20591=>"010111111",
  20592=>"000000000",
  20593=>"111110100",
  20594=>"111100110",
  20595=>"100101100",
  20596=>"000000000",
  20597=>"011010010",
  20598=>"000000110",
  20599=>"011011011",
  20600=>"000000000",
  20601=>"001001001",
  20602=>"011011011",
  20603=>"000000000",
  20604=>"000001011",
  20605=>"111010111",
  20606=>"111111000",
  20607=>"111111100",
  20608=>"111111000",
  20609=>"000000111",
  20610=>"111111111",
  20611=>"110110111",
  20612=>"000000000",
  20613=>"000000000",
  20614=>"000100000",
  20615=>"110011010",
  20616=>"000011011",
  20617=>"000100110",
  20618=>"110111111",
  20619=>"100000000",
  20620=>"000000000",
  20621=>"111010110",
  20622=>"111001001",
  20623=>"001001111",
  20624=>"001111111",
  20625=>"111111101",
  20626=>"111110110",
  20627=>"111100110",
  20628=>"001001001",
  20629=>"110110000",
  20630=>"001001100",
  20631=>"111111000",
  20632=>"111111101",
  20633=>"111111111",
  20634=>"000000111",
  20635=>"111101100",
  20636=>"000000000",
  20637=>"101111010",
  20638=>"110000000",
  20639=>"001001000",
  20640=>"000110000",
  20641=>"000000010",
  20642=>"000000000",
  20643=>"111111111",
  20644=>"010011111",
  20645=>"000000000",
  20646=>"111111111",
  20647=>"111110110",
  20648=>"111111101",
  20649=>"111111111",
  20650=>"000011111",
  20651=>"000000100",
  20652=>"110110110",
  20653=>"001001001",
  20654=>"100000001",
  20655=>"111111111",
  20656=>"000001000",
  20657=>"100100100",
  20658=>"110110110",
  20659=>"000000000",
  20660=>"111111011",
  20661=>"011011000",
  20662=>"111110111",
  20663=>"111110000",
  20664=>"111111111",
  20665=>"111111000",
  20666=>"111111111",
  20667=>"000000001",
  20668=>"000000000",
  20669=>"011000000",
  20670=>"000001000",
  20671=>"000000001",
  20672=>"000000111",
  20673=>"000110110",
  20674=>"000000000",
  20675=>"111111001",
  20676=>"000000000",
  20677=>"111111111",
  20678=>"000000001",
  20679=>"111110111",
  20680=>"111111111",
  20681=>"000000100",
  20682=>"011000000",
  20683=>"111111110",
  20684=>"111111111",
  20685=>"111111111",
  20686=>"110111000",
  20687=>"001111111",
  20688=>"100011111",
  20689=>"001001000",
  20690=>"011000000",
  20691=>"000001111",
  20692=>"111000101",
  20693=>"000000001",
  20694=>"000000000",
  20695=>"111110100",
  20696=>"001000000",
  20697=>"110110100",
  20698=>"000000000",
  20699=>"000000110",
  20700=>"011000000",
  20701=>"111111111",
  20702=>"111111101",
  20703=>"011100111",
  20704=>"100001001",
  20705=>"000111111",
  20706=>"000101111",
  20707=>"111000000",
  20708=>"110000111",
  20709=>"110110100",
  20710=>"011111111",
  20711=>"101111111",
  20712=>"111010000",
  20713=>"100000001",
  20714=>"100110110",
  20715=>"000000000",
  20716=>"000000000",
  20717=>"111111111",
  20718=>"111011000",
  20719=>"000001000",
  20720=>"011000000",
  20721=>"110000100",
  20722=>"000010000",
  20723=>"000000000",
  20724=>"000000100",
  20725=>"001011011",
  20726=>"000100110",
  20727=>"000001011",
  20728=>"000001111",
  20729=>"001111111",
  20730=>"000001111",
  20731=>"000000000",
  20732=>"111111111",
  20733=>"000000000",
  20734=>"011111111",
  20735=>"011011111",
  20736=>"000000000",
  20737=>"111111111",
  20738=>"111111011",
  20739=>"010111010",
  20740=>"000100100",
  20741=>"111011000",
  20742=>"111111111",
  20743=>"001001011",
  20744=>"000110110",
  20745=>"110111111",
  20746=>"000000000",
  20747=>"111111111",
  20748=>"111111110",
  20749=>"011011111",
  20750=>"110110110",
  20751=>"001001001",
  20752=>"000000010",
  20753=>"111011001",
  20754=>"001000011",
  20755=>"011000111",
  20756=>"011011000",
  20757=>"101111001",
  20758=>"111011011",
  20759=>"000000110",
  20760=>"111111111",
  20761=>"000110111",
  20762=>"000000000",
  20763=>"011011011",
  20764=>"111111110",
  20765=>"110000001",
  20766=>"111111111",
  20767=>"000100010",
  20768=>"011011001",
  20769=>"000000111",
  20770=>"011111111",
  20771=>"000011011",
  20772=>"000000000",
  20773=>"011011000",
  20774=>"110000001",
  20775=>"110110111",
  20776=>"111101100",
  20777=>"111001000",
  20778=>"100100100",
  20779=>"110111111",
  20780=>"011100000",
  20781=>"110000000",
  20782=>"000000000",
  20783=>"000100100",
  20784=>"111111001",
  20785=>"001000100",
  20786=>"111111111",
  20787=>"111000000",
  20788=>"000000000",
  20789=>"000000000",
  20790=>"001111100",
  20791=>"110100000",
  20792=>"011101111",
  20793=>"001111111",
  20794=>"000000011",
  20795=>"000000000",
  20796=>"101111111",
  20797=>"000000000",
  20798=>"000111111",
  20799=>"000000100",
  20800=>"100001001",
  20801=>"000000100",
  20802=>"110111101",
  20803=>"100000111",
  20804=>"111001000",
  20805=>"000000000",
  20806=>"100101101",
  20807=>"011010000",
  20808=>"010010110",
  20809=>"111111000",
  20810=>"000000000",
  20811=>"100110100",
  20812=>"111010000",
  20813=>"011001000",
  20814=>"010110110",
  20815=>"001101100",
  20816=>"000010011",
  20817=>"010000011",
  20818=>"100110110",
  20819=>"000000000",
  20820=>"111111111",
  20821=>"111111111",
  20822=>"111111111",
  20823=>"111111101",
  20824=>"001000000",
  20825=>"111111010",
  20826=>"111111111",
  20827=>"000000100",
  20828=>"000000001",
  20829=>"000000000",
  20830=>"001011010",
  20831=>"111111111",
  20832=>"001001011",
  20833=>"000000000",
  20834=>"110000000",
  20835=>"110111001",
  20836=>"110110111",
  20837=>"001001001",
  20838=>"110000000",
  20839=>"000000000",
  20840=>"000111001",
  20841=>"000000001",
  20842=>"000000000",
  20843=>"101001001",
  20844=>"000000000",
  20845=>"010010000",
  20846=>"010111011",
  20847=>"111111111",
  20848=>"111101100",
  20849=>"111010000",
  20850=>"111111110",
  20851=>"010000001",
  20852=>"011111011",
  20853=>"100100111",
  20854=>"000000001",
  20855=>"111111111",
  20856=>"111111001",
  20857=>"111111001",
  20858=>"010000100",
  20859=>"100100100",
  20860=>"100111101",
  20861=>"110110111",
  20862=>"011001011",
  20863=>"111111000",
  20864=>"010110111",
  20865=>"111111111",
  20866=>"010111111",
  20867=>"000000000",
  20868=>"010011011",
  20869=>"000000000",
  20870=>"111011000",
  20871=>"000001001",
  20872=>"000000000",
  20873=>"100110110",
  20874=>"111111000",
  20875=>"111111111",
  20876=>"111111111",
  20877=>"001001001",
  20878=>"100000000",
  20879=>"000000000",
  20880=>"111111111",
  20881=>"110111111",
  20882=>"000000111",
  20883=>"001001001",
  20884=>"111111111",
  20885=>"001001000",
  20886=>"011111111",
  20887=>"001001011",
  20888=>"111111111",
  20889=>"111000110",
  20890=>"000111111",
  20891=>"111101011",
  20892=>"111111111",
  20893=>"000000000",
  20894=>"001000000",
  20895=>"111111111",
  20896=>"011001000",
  20897=>"111011011",
  20898=>"110111100",
  20899=>"000000000",
  20900=>"000000100",
  20901=>"111111011",
  20902=>"110010010",
  20903=>"000000000",
  20904=>"100100000",
  20905=>"000000100",
  20906=>"011000111",
  20907=>"101001000",
  20908=>"001000000",
  20909=>"011111111",
  20910=>"000100110",
  20911=>"011111111",
  20912=>"001000000",
  20913=>"111111111",
  20914=>"101000000",
  20915=>"000000100",
  20916=>"000100000",
  20917=>"000000110",
  20918=>"110110111",
  20919=>"101000000",
  20920=>"000000011",
  20921=>"111001100",
  20922=>"100111100",
  20923=>"111111110",
  20924=>"000000000",
  20925=>"111001101",
  20926=>"000101101",
  20927=>"011011011",
  20928=>"100011000",
  20929=>"000000000",
  20930=>"000000000",
  20931=>"111111111",
  20932=>"111111111",
  20933=>"000000000",
  20934=>"000000000",
  20935=>"111111111",
  20936=>"111110110",
  20937=>"001100110",
  20938=>"111100100",
  20939=>"000111111",
  20940=>"000000000",
  20941=>"111001000",
  20942=>"011111110",
  20943=>"001000000",
  20944=>"000000111",
  20945=>"110111111",
  20946=>"000000000",
  20947=>"111111111",
  20948=>"000000011",
  20949=>"111111111",
  20950=>"010000000",
  20951=>"001001111",
  20952=>"000111011",
  20953=>"001101111",
  20954=>"111111001",
  20955=>"011011000",
  20956=>"000001000",
  20957=>"001011000",
  20958=>"111111000",
  20959=>"111111011",
  20960=>"000000110",
  20961=>"111111111",
  20962=>"111111111",
  20963=>"000000000",
  20964=>"111111111",
  20965=>"011011111",
  20966=>"101100100",
  20967=>"010000000",
  20968=>"000000000",
  20969=>"000101101",
  20970=>"110110000",
  20971=>"000001011",
  20972=>"000000000",
  20973=>"000000100",
  20974=>"100100111",
  20975=>"010000000",
  20976=>"001111111",
  20977=>"000000000",
  20978=>"011011011",
  20979=>"000001000",
  20980=>"000000110",
  20981=>"111111001",
  20982=>"000000000",
  20983=>"111100100",
  20984=>"111111110",
  20985=>"000100100",
  20986=>"001011111",
  20987=>"100000000",
  20988=>"000000100",
  20989=>"111011011",
  20990=>"001000000",
  20991=>"100001001",
  20992=>"110101111",
  20993=>"010111011",
  20994=>"111011000",
  20995=>"111010000",
  20996=>"001001111",
  20997=>"100111111",
  20998=>"111111010",
  20999=>"111111111",
  21000=>"111011011",
  21001=>"001001011",
  21002=>"000000000",
  21003=>"111111111",
  21004=>"110110111",
  21005=>"000001001",
  21006=>"101111111",
  21007=>"000111111",
  21008=>"111101000",
  21009=>"111110100",
  21010=>"011011111",
  21011=>"001000001",
  21012=>"111011011",
  21013=>"000111111",
  21014=>"010111111",
  21015=>"100111011",
  21016=>"000100100",
  21017=>"110110111",
  21018=>"111111001",
  21019=>"100110100",
  21020=>"111101111",
  21021=>"010000000",
  21022=>"001011011",
  21023=>"000000001",
  21024=>"010000111",
  21025=>"000000110",
  21026=>"100110110",
  21027=>"101111111",
  21028=>"111000000",
  21029=>"000000000",
  21030=>"000000000",
  21031=>"000000110",
  21032=>"111111111",
  21033=>"010111110",
  21034=>"000001111",
  21035=>"111111110",
  21036=>"110111111",
  21037=>"000000000",
  21038=>"001000010",
  21039=>"000001111",
  21040=>"111111111",
  21041=>"000000111",
  21042=>"100100100",
  21043=>"111100000",
  21044=>"110110111",
  21045=>"100100110",
  21046=>"110110111",
  21047=>"000000000",
  21048=>"111111111",
  21049=>"001111101",
  21050=>"111111111",
  21051=>"111000000",
  21052=>"111111111",
  21053=>"111110111",
  21054=>"000011111",
  21055=>"000000000",
  21056=>"000100111",
  21057=>"000000001",
  21058=>"000000000",
  21059=>"001000111",
  21060=>"000001001",
  21061=>"111111111",
  21062=>"000000000",
  21063=>"111111110",
  21064=>"011111000",
  21065=>"000011000",
  21066=>"010000000",
  21067=>"111111111",
  21068=>"111101010",
  21069=>"000000001",
  21070=>"001000000",
  21071=>"111001001",
  21072=>"000000000",
  21073=>"000001111",
  21074=>"000000000",
  21075=>"001001101",
  21076=>"110110000",
  21077=>"000000110",
  21078=>"111000000",
  21079=>"111111111",
  21080=>"111000100",
  21081=>"101000000",
  21082=>"111111111",
  21083=>"110110010",
  21084=>"000110111",
  21085=>"011000000",
  21086=>"111111111",
  21087=>"000000000",
  21088=>"000110110",
  21089=>"001011011",
  21090=>"111101000",
  21091=>"001011111",
  21092=>"111111000",
  21093=>"000000001",
  21094=>"000000010",
  21095=>"010011010",
  21096=>"111011001",
  21097=>"111011011",
  21098=>"011111111",
  21099=>"111111110",
  21100=>"101001011",
  21101=>"110000000",
  21102=>"111000011",
  21103=>"000000100",
  21104=>"111111101",
  21105=>"000001111",
  21106=>"011011111",
  21107=>"000100110",
  21108=>"000000000",
  21109=>"000100000",
  21110=>"000111111",
  21111=>"000111111",
  21112=>"001111001",
  21113=>"000000000",
  21114=>"000000000",
  21115=>"000111111",
  21116=>"111011011",
  21117=>"000000000",
  21118=>"000000000",
  21119=>"100101111",
  21120=>"000000111",
  21121=>"011000010",
  21122=>"101001000",
  21123=>"101101001",
  21124=>"000101000",
  21125=>"000100000",
  21126=>"001001001",
  21127=>"001001010",
  21128=>"100000000",
  21129=>"111000111",
  21130=>"111111111",
  21131=>"000000100",
  21132=>"000000000",
  21133=>"111111111",
  21134=>"111111111",
  21135=>"111111111",
  21136=>"011101111",
  21137=>"000000000",
  21138=>"100110111",
  21139=>"001000000",
  21140=>"000000000",
  21141=>"111000000",
  21142=>"000111111",
  21143=>"111001001",
  21144=>"000000100",
  21145=>"111111111",
  21146=>"111100110",
  21147=>"001001001",
  21148=>"111000000",
  21149=>"100101111",
  21150=>"111111001",
  21151=>"010000010",
  21152=>"111111111",
  21153=>"000011001",
  21154=>"001111111",
  21155=>"111111111",
  21156=>"011011001",
  21157=>"000000001",
  21158=>"111111111",
  21159=>"000011001",
  21160=>"111111111",
  21161=>"000000000",
  21162=>"111111110",
  21163=>"000000000",
  21164=>"001111111",
  21165=>"111100000",
  21166=>"000000101",
  21167=>"000111111",
  21168=>"000111111",
  21169=>"011111110",
  21170=>"111111111",
  21171=>"111111111",
  21172=>"110010001",
  21173=>"001010000",
  21174=>"000000000",
  21175=>"111001000",
  21176=>"000000100",
  21177=>"111111111",
  21178=>"000000000",
  21179=>"110110100",
  21180=>"001000000",
  21181=>"010000100",
  21182=>"000010110",
  21183=>"000000000",
  21184=>"111000111",
  21185=>"000000000",
  21186=>"000000000",
  21187=>"101101111",
  21188=>"000000000",
  21189=>"000000011",
  21190=>"100000000",
  21191=>"111111010",
  21192=>"011111000",
  21193=>"111111111",
  21194=>"111101111",
  21195=>"000000000",
  21196=>"101000000",
  21197=>"100100000",
  21198=>"111111001",
  21199=>"100000111",
  21200=>"000000111",
  21201=>"000001111",
  21202=>"111000000",
  21203=>"111111110",
  21204=>"111111100",
  21205=>"111111110",
  21206=>"001000000",
  21207=>"000000110",
  21208=>"111111110",
  21209=>"110111111",
  21210=>"111111111",
  21211=>"000000001",
  21212=>"110110010",
  21213=>"000000000",
  21214=>"000111111",
  21215=>"000000111",
  21216=>"100000111",
  21217=>"000000111",
  21218=>"000001111",
  21219=>"111111000",
  21220=>"111111111",
  21221=>"011011111",
  21222=>"000000000",
  21223=>"000000000",
  21224=>"000000000",
  21225=>"111111100",
  21226=>"101001000",
  21227=>"000000100",
  21228=>"001000101",
  21229=>"000101111",
  21230=>"000000000",
  21231=>"000000000",
  21232=>"000000000",
  21233=>"111111110",
  21234=>"111111111",
  21235=>"000100100",
  21236=>"111000100",
  21237=>"000000101",
  21238=>"111111111",
  21239=>"111111111",
  21240=>"000000011",
  21241=>"110111110",
  21242=>"000000000",
  21243=>"111000000",
  21244=>"011001001",
  21245=>"001001001",
  21246=>"001000000",
  21247=>"000000000",
  21248=>"000000000",
  21249=>"101100100",
  21250=>"111111000",
  21251=>"000011000",
  21252=>"100110110",
  21253=>"010111110",
  21254=>"111111101",
  21255=>"111111111",
  21256=>"111111010",
  21257=>"010000000",
  21258=>"011000100",
  21259=>"111111111",
  21260=>"111110110",
  21261=>"000000000",
  21262=>"000000000",
  21263=>"000000000",
  21264=>"001001100",
  21265=>"000000100",
  21266=>"111111111",
  21267=>"111111011",
  21268=>"111111000",
  21269=>"001000000",
  21270=>"111100100",
  21271=>"000000000",
  21272=>"000000000",
  21273=>"110100000",
  21274=>"111111111",
  21275=>"011000000",
  21276=>"000001011",
  21277=>"000000001",
  21278=>"000101111",
  21279=>"001011111",
  21280=>"111110000",
  21281=>"010111111",
  21282=>"111111110",
  21283=>"001001111",
  21284=>"000000000",
  21285=>"000000111",
  21286=>"111111111",
  21287=>"100111010",
  21288=>"001011010",
  21289=>"111001001",
  21290=>"101000000",
  21291=>"100100101",
  21292=>"111111000",
  21293=>"001001100",
  21294=>"101001000",
  21295=>"011111111",
  21296=>"111111000",
  21297=>"001110111",
  21298=>"001000110",
  21299=>"111011000",
  21300=>"111111111",
  21301=>"000000000",
  21302=>"001111110",
  21303=>"111101101",
  21304=>"110010000",
  21305=>"100000000",
  21306=>"011010000",
  21307=>"100000100",
  21308=>"000000100",
  21309=>"000110110",
  21310=>"111101000",
  21311=>"110100000",
  21312=>"100111111",
  21313=>"000000000",
  21314=>"111110010",
  21315=>"000111111",
  21316=>"000001111",
  21317=>"000000000",
  21318=>"111111000",
  21319=>"000000100",
  21320=>"000000000",
  21321=>"000000000",
  21322=>"101111111",
  21323=>"111001101",
  21324=>"000000000",
  21325=>"001001111",
  21326=>"101000000",
  21327=>"000001101",
  21328=>"001000100",
  21329=>"111111000",
  21330=>"111000000",
  21331=>"000000001",
  21332=>"011000000",
  21333=>"011001000",
  21334=>"011010111",
  21335=>"000000000",
  21336=>"111111111",
  21337=>"100000000",
  21338=>"101111000",
  21339=>"000000000",
  21340=>"111110110",
  21341=>"000110111",
  21342=>"111111010",
  21343=>"000000000",
  21344=>"000001111",
  21345=>"000000000",
  21346=>"000100111",
  21347=>"011001001",
  21348=>"111111111",
  21349=>"000000000",
  21350=>"000000111",
  21351=>"111111111",
  21352=>"001001111",
  21353=>"000111111",
  21354=>"101101111",
  21355=>"100100101",
  21356=>"110011111",
  21357=>"000000111",
  21358=>"000000000",
  21359=>"000111111",
  21360=>"000000010",
  21361=>"111111111",
  21362=>"000000110",
  21363=>"001001000",
  21364=>"111111000",
  21365=>"000000000",
  21366=>"000000000",
  21367=>"110110100",
  21368=>"111111000",
  21369=>"111111000",
  21370=>"000000110",
  21371=>"011111111",
  21372=>"101111000",
  21373=>"110100111",
  21374=>"000000000",
  21375=>"000111111",
  21376=>"111111111",
  21377=>"000000100",
  21378=>"110111111",
  21379=>"000000000",
  21380=>"000000101",
  21381=>"000000000",
  21382=>"000000110",
  21383=>"000000000",
  21384=>"111000000",
  21385=>"000000000",
  21386=>"100000000",
  21387=>"010110111",
  21388=>"111100111",
  21389=>"100100101",
  21390=>"000000000",
  21391=>"000001111",
  21392=>"000100100",
  21393=>"111111111",
  21394=>"000000000",
  21395=>"111000000",
  21396=>"111111111",
  21397=>"000000000",
  21398=>"111111010",
  21399=>"111111110",
  21400=>"100101111",
  21401=>"101111001",
  21402=>"000110111",
  21403=>"000000111",
  21404=>"011000000",
  21405=>"111001001",
  21406=>"110110111",
  21407=>"111111111",
  21408=>"110110110",
  21409=>"111111110",
  21410=>"111111111",
  21411=>"000000000",
  21412=>"100100101",
  21413=>"111000000",
  21414=>"111001100",
  21415=>"000000000",
  21416=>"111001001",
  21417=>"111100000",
  21418=>"001000101",
  21419=>"000000000",
  21420=>"001101001",
  21421=>"000000000",
  21422=>"000000001",
  21423=>"000100100",
  21424=>"111111111",
  21425=>"111001000",
  21426=>"111110111",
  21427=>"001000000",
  21428=>"111111111",
  21429=>"000001111",
  21430=>"000000111",
  21431=>"111111111",
  21432=>"101111000",
  21433=>"111101100",
  21434=>"101000000",
  21435=>"111011011",
  21436=>"111111111",
  21437=>"001001000",
  21438=>"011111000",
  21439=>"111100110",
  21440=>"111111111",
  21441=>"001001001",
  21442=>"111111000",
  21443=>"100111111",
  21444=>"111111111",
  21445=>"001001101",
  21446=>"010000000",
  21447=>"000000101",
  21448=>"111000000",
  21449=>"000010111",
  21450=>"000000001",
  21451=>"010000001",
  21452=>"000001000",
  21453=>"000000000",
  21454=>"101101111",
  21455=>"000111111",
  21456=>"111100100",
  21457=>"101001000",
  21458=>"000000000",
  21459=>"011000000",
  21460=>"001000100",
  21461=>"001000001",
  21462=>"111111000",
  21463=>"011001001",
  21464=>"000100101",
  21465=>"000000101",
  21466=>"111111111",
  21467=>"000000000",
  21468=>"111111111",
  21469=>"111000000",
  21470=>"110100000",
  21471=>"000101111",
  21472=>"000101111",
  21473=>"000111111",
  21474=>"011111111",
  21475=>"010000000",
  21476=>"111001111",
  21477=>"111110000",
  21478=>"000101111",
  21479=>"110110110",
  21480=>"000000001",
  21481=>"111111111",
  21482=>"000000000",
  21483=>"111111111",
  21484=>"101111111",
  21485=>"000110000",
  21486=>"111001111",
  21487=>"111111111",
  21488=>"000000000",
  21489=>"000000000",
  21490=>"100100101",
  21491=>"000111111",
  21492=>"111001000",
  21493=>"111111111",
  21494=>"101100100",
  21495=>"001001000",
  21496=>"001011011",
  21497=>"111010010",
  21498=>"000000101",
  21499=>"111111100",
  21500=>"100111001",
  21501=>"001000000",
  21502=>"111000101",
  21503=>"101000000",
  21504=>"000000011",
  21505=>"000000110",
  21506=>"000100111",
  21507=>"111111111",
  21508=>"000001011",
  21509=>"111110111",
  21510=>"110100000",
  21511=>"000000000",
  21512=>"011111111",
  21513=>"000111111",
  21514=>"110111111",
  21515=>"000000000",
  21516=>"100000000",
  21517=>"111001111",
  21518=>"000100111",
  21519=>"000100111",
  21520=>"001000110",
  21521=>"000010110",
  21522=>"111111111",
  21523=>"000011001",
  21524=>"000000000",
  21525=>"111101111",
  21526=>"111111111",
  21527=>"011111001",
  21528=>"011011000",
  21529=>"000000001",
  21530=>"000000111",
  21531=>"000000000",
  21532=>"000000000",
  21533=>"000001111",
  21534=>"111111110",
  21535=>"011001111",
  21536=>"000110110",
  21537=>"100111001",
  21538=>"110000100",
  21539=>"000000000",
  21540=>"000000000",
  21541=>"000111111",
  21542=>"000100000",
  21543=>"000000000",
  21544=>"100001101",
  21545=>"010111110",
  21546=>"000000000",
  21547=>"110000101",
  21548=>"011000010",
  21549=>"100111111",
  21550=>"000000001",
  21551=>"000000000",
  21552=>"111111001",
  21553=>"000000001",
  21554=>"111111111",
  21555=>"000111111",
  21556=>"111011000",
  21557=>"000110111",
  21558=>"000000001",
  21559=>"100100000",
  21560=>"111111111",
  21561=>"000000101",
  21562=>"101000000",
  21563=>"001000000",
  21564=>"000001001",
  21565=>"111000000",
  21566=>"100110011",
  21567=>"111000000",
  21568=>"011000000",
  21569=>"000001000",
  21570=>"111011011",
  21571=>"111111111",
  21572=>"000000000",
  21573=>"111111111",
  21574=>"111110111",
  21575=>"111111111",
  21576=>"100111111",
  21577=>"000000101",
  21578=>"110000000",
  21579=>"111010000",
  21580=>"111111111",
  21581=>"000000000",
  21582=>"000000000",
  21583=>"011000101",
  21584=>"011001000",
  21585=>"011111100",
  21586=>"111111111",
  21587=>"110111111",
  21588=>"000000000",
  21589=>"000000000",
  21590=>"011001001",
  21591=>"001001001",
  21592=>"010011111",
  21593=>"111111101",
  21594=>"000000001",
  21595=>"000000000",
  21596=>"000000011",
  21597=>"000010111",
  21598=>"111111111",
  21599=>"111110111",
  21600=>"010110111",
  21601=>"000000000",
  21602=>"000000000",
  21603=>"000000000",
  21604=>"001001001",
  21605=>"111100000",
  21606=>"111111111",
  21607=>"111111111",
  21608=>"000101111",
  21609=>"011011001",
  21610=>"000000111",
  21611=>"000000000",
  21612=>"000000000",
  21613=>"000000000",
  21614=>"001011011",
  21615=>"000000010",
  21616=>"111000000",
  21617=>"011000011",
  21618=>"111110010",
  21619=>"000000001",
  21620=>"111000000",
  21621=>"000110000",
  21622=>"111111111",
  21623=>"111111111",
  21624=>"000100000",
  21625=>"000000000",
  21626=>"011111101",
  21627=>"000000000",
  21628=>"110110000",
  21629=>"000000000",
  21630=>"000000000",
  21631=>"000000000",
  21632=>"000000000",
  21633=>"111111111",
  21634=>"111000000",
  21635=>"011011101",
  21636=>"111111111",
  21637=>"100000000",
  21638=>"111001111",
  21639=>"000000110",
  21640=>"110110110",
  21641=>"111101000",
  21642=>"000000011",
  21643=>"011000000",
  21644=>"111111111",
  21645=>"110100100",
  21646=>"011001001",
  21647=>"110111111",
  21648=>"011010000",
  21649=>"000000111",
  21650=>"111111110",
  21651=>"111111111",
  21652=>"111111110",
  21653=>"000000000",
  21654=>"000000111",
  21655=>"000000000",
  21656=>"000000000",
  21657=>"000000000",
  21658=>"000000000",
  21659=>"110111111",
  21660=>"111101000",
  21661=>"111110000",
  21662=>"011111111",
  21663=>"000000000",
  21664=>"011000100",
  21665=>"110100000",
  21666=>"111000110",
  21667=>"000000011",
  21668=>"000000000",
  21669=>"110110111",
  21670=>"011001000",
  21671=>"011111100",
  21672=>"100000000",
  21673=>"111100000",
  21674=>"000000000",
  21675=>"000111111",
  21676=>"111111001",
  21677=>"000000100",
  21678=>"111111111",
  21679=>"111110011",
  21680=>"010000000",
  21681=>"000100111",
  21682=>"111111111",
  21683=>"000101111",
  21684=>"000000001",
  21685=>"000000101",
  21686=>"000000001",
  21687=>"000000111",
  21688=>"001001011",
  21689=>"111111111",
  21690=>"000000000",
  21691=>"000000001",
  21692=>"000000000",
  21693=>"111000111",
  21694=>"111111110",
  21695=>"111111111",
  21696=>"111111111",
  21697=>"000011011",
  21698=>"110011000",
  21699=>"111111111",
  21700=>"001001111",
  21701=>"011110000",
  21702=>"011101100",
  21703=>"000101011",
  21704=>"000011000",
  21705=>"000000000",
  21706=>"001001111",
  21707=>"000010000",
  21708=>"111011111",
  21709=>"000110000",
  21710=>"111111111",
  21711=>"000000000",
  21712=>"110110000",
  21713=>"000100111",
  21714=>"100000000",
  21715=>"000000000",
  21716=>"111111100",
  21717=>"011011111",
  21718=>"000110000",
  21719=>"000001101",
  21720=>"101111111",
  21721=>"000000001",
  21722=>"111000000",
  21723=>"000000111",
  21724=>"000111111",
  21725=>"001011111",
  21726=>"111111111",
  21727=>"111111101",
  21728=>"000100110",
  21729=>"000000110",
  21730=>"111111000",
  21731=>"111000000",
  21732=>"000000000",
  21733=>"000101111",
  21734=>"110111111",
  21735=>"111111111",
  21736=>"111011000",
  21737=>"111000010",
  21738=>"111110111",
  21739=>"111111111",
  21740=>"111011000",
  21741=>"111010000",
  21742=>"111111111",
  21743=>"000000000",
  21744=>"110100111",
  21745=>"000000001",
  21746=>"000000000",
  21747=>"000000101",
  21748=>"111111111",
  21749=>"011001001",
  21750=>"000110111",
  21751=>"111111111",
  21752=>"000111111",
  21753=>"000000000",
  21754=>"000001001",
  21755=>"111111111",
  21756=>"100111111",
  21757=>"011011111",
  21758=>"111111110",
  21759=>"111100101",
  21760=>"011001101",
  21761=>"100100100",
  21762=>"000000000",
  21763=>"000111111",
  21764=>"111111111",
  21765=>"111001101",
  21766=>"111110000",
  21767=>"000011001",
  21768=>"111111111",
  21769=>"001001000",
  21770=>"000000111",
  21771=>"011011111",
  21772=>"000000011",
  21773=>"111111100",
  21774=>"000001111",
  21775=>"110000000",
  21776=>"000000000",
  21777=>"000000000",
  21778=>"111000101",
  21779=>"011111111",
  21780=>"000100110",
  21781=>"000010111",
  21782=>"110111100",
  21783=>"001000000",
  21784=>"010000111",
  21785=>"111111111",
  21786=>"110011011",
  21787=>"000000000",
  21788=>"001011011",
  21789=>"000001111",
  21790=>"111000000",
  21791=>"110111111",
  21792=>"100100111",
  21793=>"011111111",
  21794=>"111111110",
  21795=>"111111111",
  21796=>"100100111",
  21797=>"011000000",
  21798=>"001001001",
  21799=>"111111000",
  21800=>"111111111",
  21801=>"111000001",
  21802=>"111100101",
  21803=>"001000100",
  21804=>"000000000",
  21805=>"000000000",
  21806=>"000000000",
  21807=>"000001010",
  21808=>"110111111",
  21809=>"001000000",
  21810=>"110001000",
  21811=>"000000000",
  21812=>"000000000",
  21813=>"011000000",
  21814=>"000000001",
  21815=>"111111100",
  21816=>"000000000",
  21817=>"111001000",
  21818=>"111111001",
  21819=>"000000010",
  21820=>"000010010",
  21821=>"101101110",
  21822=>"000000000",
  21823=>"000000000",
  21824=>"000000111",
  21825=>"111111010",
  21826=>"000011011",
  21827=>"111000000",
  21828=>"000001111",
  21829=>"011001000",
  21830=>"000000000",
  21831=>"110111111",
  21832=>"000000000",
  21833=>"000000000",
  21834=>"111000000",
  21835=>"110110000",
  21836=>"000000000",
  21837=>"000000000",
  21838=>"111111011",
  21839=>"010000000",
  21840=>"110111111",
  21841=>"000000000",
  21842=>"110111001",
  21843=>"000000000",
  21844=>"011000000",
  21845=>"011011011",
  21846=>"111111000",
  21847=>"000001000",
  21848=>"000000000",
  21849=>"000100001",
  21850=>"000000000",
  21851=>"111111111",
  21852=>"000110010",
  21853=>"000000111",
  21854=>"110010000",
  21855=>"111111011",
  21856=>"000000000",
  21857=>"110000000",
  21858=>"111111011",
  21859=>"000000000",
  21860=>"000001000",
  21861=>"110111100",
  21862=>"111100000",
  21863=>"000000111",
  21864=>"011011010",
  21865=>"111111100",
  21866=>"001111011",
  21867=>"111000110",
  21868=>"100010111",
  21869=>"111110000",
  21870=>"000000000",
  21871=>"111111111",
  21872=>"000010001",
  21873=>"000010111",
  21874=>"010100000",
  21875=>"111101111",
  21876=>"111100000",
  21877=>"011111111",
  21878=>"111000000",
  21879=>"010000000",
  21880=>"000000000",
  21881=>"000000000",
  21882=>"000000000",
  21883=>"000000000",
  21884=>"000000000",
  21885=>"111111100",
  21886=>"000111111",
  21887=>"000000110",
  21888=>"000001111",
  21889=>"110100000",
  21890=>"101111001",
  21891=>"001000000",
  21892=>"000000000",
  21893=>"111111000",
  21894=>"111000000",
  21895=>"110110111",
  21896=>"000000000",
  21897=>"111110000",
  21898=>"000000000",
  21899=>"001000000",
  21900=>"111111111",
  21901=>"000000000",
  21902=>"000000111",
  21903=>"000000000",
  21904=>"000000000",
  21905=>"111100000",
  21906=>"000000111",
  21907=>"000000000",
  21908=>"001000000",
  21909=>"000100000",
  21910=>"001000000",
  21911=>"111111111",
  21912=>"001111111",
  21913=>"011001110",
  21914=>"100100000",
  21915=>"000010111",
  21916=>"111001001",
  21917=>"000000010",
  21918=>"000000000",
  21919=>"101000000",
  21920=>"100100000",
  21921=>"111111100",
  21922=>"111100101",
  21923=>"001111111",
  21924=>"001111001",
  21925=>"111111000",
  21926=>"011000000",
  21927=>"000000000",
  21928=>"000000000",
  21929=>"110000000",
  21930=>"111110110",
  21931=>"010111101",
  21932=>"000000000",
  21933=>"111111110",
  21934=>"111011101",
  21935=>"011011001",
  21936=>"011000000",
  21937=>"010000000",
  21938=>"000000000",
  21939=>"111111111",
  21940=>"111111111",
  21941=>"111100100",
  21942=>"001001000",
  21943=>"000110101",
  21944=>"000000000",
  21945=>"111011000",
  21946=>"100000000",
  21947=>"100111111",
  21948=>"000111111",
  21949=>"000000000",
  21950=>"011110111",
  21951=>"100100100",
  21952=>"000000110",
  21953=>"010000000",
  21954=>"011001111",
  21955=>"111110111",
  21956=>"000000111",
  21957=>"000001001",
  21958=>"000000100",
  21959=>"000101111",
  21960=>"000000000",
  21961=>"000000000",
  21962=>"111000001",
  21963=>"111111111",
  21964=>"101101111",
  21965=>"111111111",
  21966=>"000000000",
  21967=>"111111100",
  21968=>"110110000",
  21969=>"111111001",
  21970=>"000000000",
  21971=>"001111111",
  21972=>"100000001",
  21973=>"111111100",
  21974=>"000000111",
  21975=>"011000110",
  21976=>"000000000",
  21977=>"011001000",
  21978=>"000011111",
  21979=>"111111110",
  21980=>"110111111",
  21981=>"100001011",
  21982=>"111111001",
  21983=>"111110000",
  21984=>"111111110",
  21985=>"111111111",
  21986=>"000011010",
  21987=>"111110000",
  21988=>"011000000",
  21989=>"111111111",
  21990=>"000000000",
  21991=>"101100001",
  21992=>"110000001",
  21993=>"111111111",
  21994=>"000000000",
  21995=>"011111011",
  21996=>"000000000",
  21997=>"000000000",
  21998=>"000000000",
  21999=>"111111111",
  22000=>"000000000",
  22001=>"111011000",
  22002=>"000001111",
  22003=>"111111000",
  22004=>"001000101",
  22005=>"000000000",
  22006=>"110110100",
  22007=>"110111110",
  22008=>"001000111",
  22009=>"111111011",
  22010=>"000110110",
  22011=>"111111011",
  22012=>"101111111",
  22013=>"000000000",
  22014=>"111111110",
  22015=>"000001111",
  22016=>"110110000",
  22017=>"111000010",
  22018=>"111000000",
  22019=>"000000000",
  22020=>"000100111",
  22021=>"000000011",
  22022=>"000000000",
  22023=>"111101100",
  22024=>"000000000",
  22025=>"011111000",
  22026=>"000000000",
  22027=>"010010001",
  22028=>"011011011",
  22029=>"110111111",
  22030=>"110110110",
  22031=>"000000000",
  22032=>"001001111",
  22033=>"000000000",
  22034=>"000000011",
  22035=>"111111111",
  22036=>"111111000",
  22037=>"111111001",
  22038=>"000000001",
  22039=>"100101100",
  22040=>"111011011",
  22041=>"000100111",
  22042=>"000000111",
  22043=>"011011001",
  22044=>"011011001",
  22045=>"000111111",
  22046=>"100000000",
  22047=>"111111000",
  22048=>"001011111",
  22049=>"110111111",
  22050=>"000000111",
  22051=>"010000100",
  22052=>"000000110",
  22053=>"100100111",
  22054=>"111110000",
  22055=>"000000111",
  22056=>"111111000",
  22057=>"000000000",
  22058=>"111000111",
  22059=>"111001010",
  22060=>"000000000",
  22061=>"111111111",
  22062=>"000000111",
  22063=>"000000000",
  22064=>"000000100",
  22065=>"111111111",
  22066=>"111011011",
  22067=>"111111000",
  22068=>"000000000",
  22069=>"010110000",
  22070=>"000000011",
  22071=>"111111111",
  22072=>"000000111",
  22073=>"000000111",
  22074=>"000000000",
  22075=>"110000000",
  22076=>"000100000",
  22077=>"001101000",
  22078=>"011111110",
  22079=>"000000110",
  22080=>"000000000",
  22081=>"100111111",
  22082=>"111111110",
  22083=>"111111000",
  22084=>"000000001",
  22085=>"000000000",
  22086=>"101000001",
  22087=>"111111000",
  22088=>"000000100",
  22089=>"001000000",
  22090=>"001000000",
  22091=>"111111111",
  22092=>"011010000",
  22093=>"000000001",
  22094=>"000000001",
  22095=>"111000000",
  22096=>"101001000",
  22097=>"000000111",
  22098=>"000000111",
  22099=>"011000001",
  22100=>"000000001",
  22101=>"001111111",
  22102=>"100000000",
  22103=>"000000000",
  22104=>"000000111",
  22105=>"101000000",
  22106=>"111111001",
  22107=>"111111100",
  22108=>"000000011",
  22109=>"111111001",
  22110=>"000111111",
  22111=>"111111110",
  22112=>"000000000",
  22113=>"000001011",
  22114=>"000000000",
  22115=>"001001000",
  22116=>"000100111",
  22117=>"000000000",
  22118=>"011011000",
  22119=>"000000000",
  22120=>"111111111",
  22121=>"000100101",
  22122=>"000000111",
  22123=>"110011000",
  22124=>"110111000",
  22125=>"000000000",
  22126=>"000000001",
  22127=>"111111111",
  22128=>"000001101",
  22129=>"111111111",
  22130=>"100000101",
  22131=>"000010110",
  22132=>"000000000",
  22133=>"110111101",
  22134=>"000000000",
  22135=>"000000000",
  22136=>"000111111",
  22137=>"000000000",
  22138=>"000000111",
  22139=>"000001000",
  22140=>"110111011",
  22141=>"110011010",
  22142=>"000101111",
  22143=>"000000000",
  22144=>"000110110",
  22145=>"000000000",
  22146=>"111010010",
  22147=>"001000111",
  22148=>"011010000",
  22149=>"000000111",
  22150=>"000100000",
  22151=>"000111111",
  22152=>"111001011",
  22153=>"001011011",
  22154=>"000000111",
  22155=>"000000110",
  22156=>"111111000",
  22157=>"000100111",
  22158=>"111111000",
  22159=>"111111000",
  22160=>"100000111",
  22161=>"000000000",
  22162=>"000000000",
  22163=>"000100111",
  22164=>"000000110",
  22165=>"000111111",
  22166=>"000000001",
  22167=>"000000111",
  22168=>"000100111",
  22169=>"111111000",
  22170=>"000001111",
  22171=>"000111111",
  22172=>"111111110",
  22173=>"000000000",
  22174=>"111111011",
  22175=>"000000111",
  22176=>"000000000",
  22177=>"001000000",
  22178=>"000000000",
  22179=>"000000000",
  22180=>"011111111",
  22181=>"000000100",
  22182=>"111000000",
  22183=>"000100100",
  22184=>"111011000",
  22185=>"000000000",
  22186=>"101100000",
  22187=>"011001001",
  22188=>"111111111",
  22189=>"111111000",
  22190=>"011111111",
  22191=>"111001001",
  22192=>"011000010",
  22193=>"000110110",
  22194=>"111111111",
  22195=>"000000001",
  22196=>"011011011",
  22197=>"001000011",
  22198=>"111111000",
  22199=>"110111111",
  22200=>"111111111",
  22201=>"111111000",
  22202=>"001000000",
  22203=>"000010000",
  22204=>"000000000",
  22205=>"111001000",
  22206=>"000001001",
  22207=>"000100111",
  22208=>"111111111",
  22209=>"000001111",
  22210=>"000001111",
  22211=>"111110000",
  22212=>"111111011",
  22213=>"000000011",
  22214=>"111111000",
  22215=>"000000000",
  22216=>"000000010",
  22217=>"011001001",
  22218=>"111011111",
  22219=>"000000000",
  22220=>"111111000",
  22221=>"110111111",
  22222=>"111111101",
  22223=>"000001111",
  22224=>"000000001",
  22225=>"000000111",
  22226=>"010011111",
  22227=>"000000111",
  22228=>"010111001",
  22229=>"111111011",
  22230=>"111111111",
  22231=>"111111000",
  22232=>"111111000",
  22233=>"100111110",
  22234=>"111001001",
  22235=>"000000000",
  22236=>"111111111",
  22237=>"111111000",
  22238=>"011011111",
  22239=>"000000111",
  22240=>"111111000",
  22241=>"010010000",
  22242=>"000000000",
  22243=>"111011111",
  22244=>"110110110",
  22245=>"111111001",
  22246=>"111111111",
  22247=>"111100000",
  22248=>"001000000",
  22249=>"110000000",
  22250=>"001111111",
  22251=>"011011011",
  22252=>"011111000",
  22253=>"000000111",
  22254=>"110111000",
  22255=>"000111001",
  22256=>"000100100",
  22257=>"111111111",
  22258=>"000000111",
  22259=>"001000111",
  22260=>"000000111",
  22261=>"110110100",
  22262=>"001011011",
  22263=>"111111000",
  22264=>"000000000",
  22265=>"000000000",
  22266=>"111011000",
  22267=>"111110010",
  22268=>"001000000",
  22269=>"001001111",
  22270=>"000000011",
  22271=>"111111000",
  22272=>"000000000",
  22273=>"101001001",
  22274=>"000000111",
  22275=>"001000000",
  22276=>"110000101",
  22277=>"011000000",
  22278=>"000000000",
  22279=>"000000000",
  22280=>"000001111",
  22281=>"000000100",
  22282=>"111111011",
  22283=>"000000111",
  22284=>"111000000",
  22285=>"000000111",
  22286=>"101111010",
  22287=>"111000000",
  22288=>"011000000",
  22289=>"001000001",
  22290=>"000000111",
  22291=>"011011000",
  22292=>"000110000",
  22293=>"000000011",
  22294=>"111111001",
  22295=>"000111101",
  22296=>"000000111",
  22297=>"111111111",
  22298=>"000000111",
  22299=>"110110010",
  22300=>"000000000",
  22301=>"111111111",
  22302=>"111111011",
  22303=>"111100100",
  22304=>"000100111",
  22305=>"111111000",
  22306=>"110000000",
  22307=>"100100100",
  22308=>"100000001",
  22309=>"111001000",
  22310=>"000000111",
  22311=>"010011111",
  22312=>"000101011",
  22313=>"000000010",
  22314=>"001001011",
  22315=>"110111111",
  22316=>"111010000",
  22317=>"001111011",
  22318=>"000010000",
  22319=>"111111000",
  22320=>"111110011",
  22321=>"100000111",
  22322=>"111111000",
  22323=>"000000001",
  22324=>"000000000",
  22325=>"111100100",
  22326=>"000000110",
  22327=>"000000100",
  22328=>"101000111",
  22329=>"101000111",
  22330=>"000000010",
  22331=>"110110111",
  22332=>"001001011",
  22333=>"111111001",
  22334=>"000000111",
  22335=>"000000000",
  22336=>"100100101",
  22337=>"001111111",
  22338=>"111111111",
  22339=>"000000000",
  22340=>"000000111",
  22341=>"111010000",
  22342=>"111111111",
  22343=>"001001000",
  22344=>"000000111",
  22345=>"011000000",
  22346=>"101111000",
  22347=>"010011011",
  22348=>"111111111",
  22349=>"111101101",
  22350=>"000000000",
  22351=>"011000000",
  22352=>"011011010",
  22353=>"000000111",
  22354=>"110111111",
  22355=>"111011000",
  22356=>"000000000",
  22357=>"011011001",
  22358=>"000000000",
  22359=>"111111111",
  22360=>"100110000",
  22361=>"000000000",
  22362=>"000010110",
  22363=>"000000111",
  22364=>"001111111",
  22365=>"111000000",
  22366=>"000000000",
  22367=>"111110000",
  22368=>"111110111",
  22369=>"111111111",
  22370=>"010100000",
  22371=>"010000100",
  22372=>"000000001",
  22373=>"000000111",
  22374=>"111010111",
  22375=>"000000111",
  22376=>"111111111",
  22377=>"000000010",
  22378=>"000000000",
  22379=>"110111000",
  22380=>"010001001",
  22381=>"000000000",
  22382=>"011001000",
  22383=>"110000011",
  22384=>"111100000",
  22385=>"000000111",
  22386=>"111111011",
  22387=>"111111111",
  22388=>"000000000",
  22389=>"100100100",
  22390=>"000000110",
  22391=>"110111111",
  22392=>"111010110",
  22393=>"111111001",
  22394=>"111111111",
  22395=>"000000110",
  22396=>"000000111",
  22397=>"000000000",
  22398=>"000000101",
  22399=>"111111010",
  22400=>"111111000",
  22401=>"111111010",
  22402=>"010000000",
  22403=>"001011111",
  22404=>"010010111",
  22405=>"000010110",
  22406=>"000000000",
  22407=>"111111110",
  22408=>"000001011",
  22409=>"000000111",
  22410=>"000000001",
  22411=>"010000111",
  22412=>"110010000",
  22413=>"100000000",
  22414=>"000000111",
  22415=>"100100000",
  22416=>"000000111",
  22417=>"111111110",
  22418=>"000011111",
  22419=>"110100110",
  22420=>"111010000",
  22421=>"000011000",
  22422=>"101101000",
  22423=>"010001011",
  22424=>"110111010",
  22425=>"110111000",
  22426=>"011000000",
  22427=>"000000111",
  22428=>"110111000",
  22429=>"000001000",
  22430=>"001000111",
  22431=>"000000000",
  22432=>"111100010",
  22433=>"110110111",
  22434=>"111111100",
  22435=>"111000000",
  22436=>"000110110",
  22437=>"000111011",
  22438=>"111001000",
  22439=>"000000111",
  22440=>"110000000",
  22441=>"000000000",
  22442=>"011001100",
  22443=>"001000011",
  22444=>"100000000",
  22445=>"000000111",
  22446=>"000000100",
  22447=>"000000111",
  22448=>"000011000",
  22449=>"111111111",
  22450=>"000111000",
  22451=>"000000001",
  22452=>"111111111",
  22453=>"011001000",
  22454=>"100001111",
  22455=>"111001000",
  22456=>"000000000",
  22457=>"000010011",
  22458=>"001000001",
  22459=>"000000111",
  22460=>"110110000",
  22461=>"000000000",
  22462=>"000011111",
  22463=>"001000111",
  22464=>"111111111",
  22465=>"111111111",
  22466=>"111111111",
  22467=>"000000001",
  22468=>"110100100",
  22469=>"000100111",
  22470=>"000000000",
  22471=>"100110100",
  22472=>"001101111",
  22473=>"111110100",
  22474=>"111111000",
  22475=>"111111111",
  22476=>"111000000",
  22477=>"111010000",
  22478=>"111001000",
  22479=>"000011111",
  22480=>"000000000",
  22481=>"111111001",
  22482=>"000000000",
  22483=>"111111100",
  22484=>"011111000",
  22485=>"100100100",
  22486=>"000111111",
  22487=>"010011111",
  22488=>"101011111",
  22489=>"000000011",
  22490=>"110110111",
  22491=>"100000000",
  22492=>"010000001",
  22493=>"111111000",
  22494=>"000000000",
  22495=>"000000000",
  22496=>"111111111",
  22497=>"011000000",
  22498=>"000001111",
  22499=>"000000000",
  22500=>"000000010",
  22501=>"000000000",
  22502=>"000001111",
  22503=>"111111011",
  22504=>"111111110",
  22505=>"111111110",
  22506=>"000000111",
  22507=>"111011100",
  22508=>"000000000",
  22509=>"100110000",
  22510=>"000000000",
  22511=>"000110111",
  22512=>"000000111",
  22513=>"011011111",
  22514=>"000000000",
  22515=>"111000000",
  22516=>"101000000",
  22517=>"111110000",
  22518=>"111100111",
  22519=>"001111111",
  22520=>"000000111",
  22521=>"110000000",
  22522=>"100001000",
  22523=>"001000111",
  22524=>"111111000",
  22525=>"110111100",
  22526=>"100000000",
  22527=>"000000001",
  22528=>"011000000",
  22529=>"111111111",
  22530=>"111111111",
  22531=>"111111111",
  22532=>"001001011",
  22533=>"100110110",
  22534=>"001111111",
  22535=>"111111111",
  22536=>"111111111",
  22537=>"000000111",
  22538=>"110111111",
  22539=>"111111100",
  22540=>"111111111",
  22541=>"001001001",
  22542=>"000000100",
  22543=>"111111111",
  22544=>"000000000",
  22545=>"001000000",
  22546=>"001101000",
  22547=>"111111111",
  22548=>"100110110",
  22549=>"000000000",
  22550=>"001000000",
  22551=>"000000001",
  22552=>"000000110",
  22553=>"001001010",
  22554=>"011111111",
  22555=>"100111110",
  22556=>"000000000",
  22557=>"111111110",
  22558=>"111111110",
  22559=>"111111111",
  22560=>"111101000",
  22561=>"000000001",
  22562=>"111111101",
  22563=>"100000101",
  22564=>"111000000",
  22565=>"000000000",
  22566=>"100000000",
  22567=>"111111000",
  22568=>"001001001",
  22569=>"111111111",
  22570=>"000000000",
  22571=>"111001001",
  22572=>"000000100",
  22573=>"011011111",
  22574=>"111111111",
  22575=>"000000000",
  22576=>"001001111",
  22577=>"000000000",
  22578=>"111111100",
  22579=>"000111100",
  22580=>"110010010",
  22581=>"101111100",
  22582=>"110111011",
  22583=>"000000101",
  22584=>"000001011",
  22585=>"100001101",
  22586=>"000000000",
  22587=>"000000000",
  22588=>"111111111",
  22589=>"111110000",
  22590=>"111011011",
  22591=>"111111110",
  22592=>"111111100",
  22593=>"000000110",
  22594=>"000000000",
  22595=>"001001001",
  22596=>"000110110",
  22597=>"111111011",
  22598=>"000100110",
  22599=>"000000000",
  22600=>"111111011",
  22601=>"000000111",
  22602=>"111111111",
  22603=>"000000000",
  22604=>"000000000",
  22605=>"001000001",
  22606=>"000000000",
  22607=>"000000000",
  22608=>"110010111",
  22609=>"011111111",
  22610=>"100000000",
  22611=>"111110111",
  22612=>"000000000",
  22613=>"000000000",
  22614=>"111100000",
  22615=>"110100111",
  22616=>"111000000",
  22617=>"000000000",
  22618=>"111001000",
  22619=>"000000011",
  22620=>"011111111",
  22621=>"100110110",
  22622=>"111101001",
  22623=>"111111111",
  22624=>"010010000",
  22625=>"000000000",
  22626=>"000000000",
  22627=>"011111111",
  22628=>"101011011",
  22629=>"000000111",
  22630=>"111110010",
  22631=>"000000000",
  22632=>"011010000",
  22633=>"111111010",
  22634=>"111111111",
  22635=>"000000000",
  22636=>"011000000",
  22637=>"000000000",
  22638=>"110100000",
  22639=>"111000111",
  22640=>"000110111",
  22641=>"110100111",
  22642=>"000000000",
  22643=>"000100111",
  22644=>"111111111",
  22645=>"000000111",
  22646=>"000000000",
  22647=>"111111110",
  22648=>"000111111",
  22649=>"000000000",
  22650=>"000001101",
  22651=>"000000000",
  22652=>"001000000",
  22653=>"011011001",
  22654=>"000000101",
  22655=>"111111111",
  22656=>"000000000",
  22657=>"011000000",
  22658=>"011011011",
  22659=>"000111011",
  22660=>"111000001",
  22661=>"111000000",
  22662=>"100111111",
  22663=>"111001011",
  22664=>"111111101",
  22665=>"111100000",
  22666=>"000000000",
  22667=>"101010000",
  22668=>"100111111",
  22669=>"000000000",
  22670=>"000000000",
  22671=>"000000000",
  22672=>"000010000",
  22673=>"110110111",
  22674=>"001000000",
  22675=>"011111000",
  22676=>"111111111",
  22677=>"000000100",
  22678=>"111000000",
  22679=>"000000000",
  22680=>"001111111",
  22681=>"011001000",
  22682=>"111111111",
  22683=>"000100110",
  22684=>"000000000",
  22685=>"000100111",
  22686=>"000000001",
  22687=>"000000000",
  22688=>"000111111",
  22689=>"011000000",
  22690=>"000000111",
  22691=>"000000000",
  22692=>"111001111",
  22693=>"000000000",
  22694=>"000000000",
  22695=>"010000111",
  22696=>"111111111",
  22697=>"000000000",
  22698=>"001000000",
  22699=>"001111111",
  22700=>"110000000",
  22701=>"111111001",
  22702=>"111111001",
  22703=>"000000000",
  22704=>"111000000",
  22705=>"000000000",
  22706=>"010111010",
  22707=>"111111000",
  22708=>"100100000",
  22709=>"000000000",
  22710=>"110110110",
  22711=>"111111111",
  22712=>"000000000",
  22713=>"000001011",
  22714=>"111000000",
  22715=>"001001000",
  22716=>"111111111",
  22717=>"111111111",
  22718=>"011010110",
  22719=>"000001101",
  22720=>"111001000",
  22721=>"000000000",
  22722=>"111111111",
  22723=>"111111111",
  22724=>"000000000",
  22725=>"111111111",
  22726=>"000001001",
  22727=>"000000000",
  22728=>"000101111",
  22729=>"111010000",
  22730=>"100111111",
  22731=>"111111000",
  22732=>"000000100",
  22733=>"000000000",
  22734=>"111001010",
  22735=>"111111110",
  22736=>"000000100",
  22737=>"111000000",
  22738=>"111011110",
  22739=>"000000000",
  22740=>"111011010",
  22741=>"111000000",
  22742=>"111001000",
  22743=>"111111111",
  22744=>"001000111",
  22745=>"111111111",
  22746=>"111111111",
  22747=>"110011001",
  22748=>"000000000",
  22749=>"000010000",
  22750=>"000100111",
  22751=>"111111111",
  22752=>"011010111",
  22753=>"010010111",
  22754=>"000111111",
  22755=>"000000000",
  22756=>"000000000",
  22757=>"000000100",
  22758=>"000001000",
  22759=>"001001000",
  22760=>"001000000",
  22761=>"111111111",
  22762=>"111100100",
  22763=>"111010000",
  22764=>"000000000",
  22765=>"111111111",
  22766=>"000000001",
  22767=>"111100111",
  22768=>"110111111",
  22769=>"000000111",
  22770=>"010000010",
  22771=>"111111001",
  22772=>"000000000",
  22773=>"001001001",
  22774=>"100100110",
  22775=>"001000000",
  22776=>"111011000",
  22777=>"111111111",
  22778=>"110110110",
  22779=>"000000000",
  22780=>"000000011",
  22781=>"001100101",
  22782=>"111001001",
  22783=>"000000000",
  22784=>"000001001",
  22785=>"100100100",
  22786=>"111111111",
  22787=>"000000111",
  22788=>"000000000",
  22789=>"000010111",
  22790=>"001000000",
  22791=>"100111111",
  22792=>"010111011",
  22793=>"111111111",
  22794=>"000000000",
  22795=>"100100001",
  22796=>"111111100",
  22797=>"111111001",
  22798=>"100000000",
  22799=>"111111101",
  22800=>"100101001",
  22801=>"011111111",
  22802=>"110111111",
  22803=>"000000000",
  22804=>"000000000",
  22805=>"000111111",
  22806=>"100000000",
  22807=>"001000000",
  22808=>"110110111",
  22809=>"000000110",
  22810=>"000000000",
  22811=>"100110110",
  22812=>"111111111",
  22813=>"111110100",
  22814=>"111000000",
  22815=>"110111111",
  22816=>"111000000",
  22817=>"001111000",
  22818=>"000111000",
  22819=>"100100110",
  22820=>"000000000",
  22821=>"111111111",
  22822=>"001000000",
  22823=>"111111111",
  22824=>"111011011",
  22825=>"000000000",
  22826=>"101000011",
  22827=>"111111111",
  22828=>"000000000",
  22829=>"110001001",
  22830=>"111110011",
  22831=>"100001000",
  22832=>"000000100",
  22833=>"111111111",
  22834=>"100111111",
  22835=>"001000011",
  22836=>"000000000",
  22837=>"001111101",
  22838=>"001001001",
  22839=>"000101111",
  22840=>"000000000",
  22841=>"000000000",
  22842=>"000000000",
  22843=>"011000000",
  22844=>"011001001",
  22845=>"111111111",
  22846=>"111000000",
  22847=>"001000000",
  22848=>"000000100",
  22849=>"111111100",
  22850=>"100100111",
  22851=>"000001111",
  22852=>"100101111",
  22853=>"000001111",
  22854=>"000000000",
  22855=>"111111111",
  22856=>"111111111",
  22857=>"110110110",
  22858=>"101000001",
  22859=>"100101000",
  22860=>"000001011",
  22861=>"001111111",
  22862=>"111111111",
  22863=>"000000001",
  22864=>"101101101",
  22865=>"111111110",
  22866=>"110111111",
  22867=>"000001001",
  22868=>"000000000",
  22869=>"000000010",
  22870=>"100111111",
  22871=>"000011111",
  22872=>"111111111",
  22873=>"111110000",
  22874=>"000110111",
  22875=>"100100000",
  22876=>"001111111",
  22877=>"111011111",
  22878=>"000100110",
  22879=>"011001001",
  22880=>"000000001",
  22881=>"000000000",
  22882=>"110111111",
  22883=>"000000011",
  22884=>"000000000",
  22885=>"111111111",
  22886=>"000000000",
  22887=>"000001000",
  22888=>"101101001",
  22889=>"111111111",
  22890=>"111111000",
  22891=>"000011111",
  22892=>"001001001",
  22893=>"111111000",
  22894=>"000000000",
  22895=>"110000000",
  22896=>"111100000",
  22897=>"111000011",
  22898=>"111101100",
  22899=>"001001000",
  22900=>"000000000",
  22901=>"000000101",
  22902=>"111111111",
  22903=>"100100100",
  22904=>"001000011",
  22905=>"111101000",
  22906=>"000000100",
  22907=>"000000000",
  22908=>"000000111",
  22909=>"011111101",
  22910=>"000100100",
  22911=>"000000000",
  22912=>"100010110",
  22913=>"001001001",
  22914=>"111111110",
  22915=>"000000100",
  22916=>"000000000",
  22917=>"111111110",
  22918=>"000000000",
  22919=>"111011111",
  22920=>"111111110",
  22921=>"000000000",
  22922=>"100100100",
  22923=>"000000111",
  22924=>"000000000",
  22925=>"101000000",
  22926=>"100101101",
  22927=>"100111110",
  22928=>"000001101",
  22929=>"100100100",
  22930=>"000000000",
  22931=>"111111000",
  22932=>"000000010",
  22933=>"110000000",
  22934=>"111111011",
  22935=>"000111111",
  22936=>"011101000",
  22937=>"010000000",
  22938=>"111111111",
  22939=>"000000111",
  22940=>"000000000",
  22941=>"000000001",
  22942=>"011000000",
  22943=>"110110111",
  22944=>"111000000",
  22945=>"100100101",
  22946=>"111001000",
  22947=>"111000000",
  22948=>"001001001",
  22949=>"000000000",
  22950=>"111111111",
  22951=>"011111111",
  22952=>"000000000",
  22953=>"111111111",
  22954=>"111111111",
  22955=>"110110000",
  22956=>"000000000",
  22957=>"100111111",
  22958=>"011011010",
  22959=>"111111100",
  22960=>"110010000",
  22961=>"111111111",
  22962=>"101101111",
  22963=>"111111111",
  22964=>"000000111",
  22965=>"110100000",
  22966=>"000001011",
  22967=>"000000111",
  22968=>"011011000",
  22969=>"011111000",
  22970=>"111110010",
  22971=>"111101111",
  22972=>"011111000",
  22973=>"111111011",
  22974=>"001000000",
  22975=>"111011111",
  22976=>"000000001",
  22977=>"110111111",
  22978=>"111111111",
  22979=>"111111111",
  22980=>"111100111",
  22981=>"011111111",
  22982=>"000000000",
  22983=>"111001001",
  22984=>"101111111",
  22985=>"000111111",
  22986=>"000000000",
  22987=>"001000000",
  22988=>"000000111",
  22989=>"000000000",
  22990=>"000001000",
  22991=>"111111111",
  22992=>"100110111",
  22993=>"001000001",
  22994=>"011001001",
  22995=>"000000111",
  22996=>"111111000",
  22997=>"111111001",
  22998=>"100110111",
  22999=>"101111111",
  23000=>"000000100",
  23001=>"000000000",
  23002=>"010001111",
  23003=>"100000000",
  23004=>"000000001",
  23005=>"001001000",
  23006=>"001000000",
  23007=>"001001011",
  23008=>"010000111",
  23009=>"111111101",
  23010=>"111110110",
  23011=>"000000011",
  23012=>"011111111",
  23013=>"000000000",
  23014=>"010110110",
  23015=>"011000000",
  23016=>"001001111",
  23017=>"111110000",
  23018=>"111110000",
  23019=>"111111111",
  23020=>"000000101",
  23021=>"000100101",
  23022=>"111111111",
  23023=>"001000000",
  23024=>"111001011",
  23025=>"111000111",
  23026=>"000000000",
  23027=>"111111000",
  23028=>"100100111",
  23029=>"111111111",
  23030=>"100000000",
  23031=>"000111111",
  23032=>"111111001",
  23033=>"000000000",
  23034=>"111000000",
  23035=>"000001001",
  23036=>"111110000",
  23037=>"100110111",
  23038=>"010110110",
  23039=>"000000000",
  23040=>"111111000",
  23041=>"000011000",
  23042=>"000000000",
  23043=>"111111000",
  23044=>"011111111",
  23045=>"000100000",
  23046=>"011111111",
  23047=>"111000000",
  23048=>"111111000",
  23049=>"111111001",
  23050=>"111111000",
  23051=>"000110110",
  23052=>"001111111",
  23053=>"101001100",
  23054=>"110001111",
  23055=>"101101000",
  23056=>"101111111",
  23057=>"000000100",
  23058=>"000000100",
  23059=>"000111110",
  23060=>"011000000",
  23061=>"111111111",
  23062=>"101001001",
  23063=>"000011111",
  23064=>"111111011",
  23065=>"000011011",
  23066=>"000000111",
  23067=>"000000000",
  23068=>"111110000",
  23069=>"100111111",
  23070=>"000011001",
  23071=>"000010100",
  23072=>"111111000",
  23073=>"111111111",
  23074=>"000010011",
  23075=>"000000000",
  23076=>"111111011",
  23077=>"110100111",
  23078=>"100011011",
  23079=>"111111101",
  23080=>"110100100",
  23081=>"000000000",
  23082=>"001001101",
  23083=>"000000100",
  23084=>"110111111",
  23085=>"101101111",
  23086=>"111111000",
  23087=>"000000001",
  23088=>"100011000",
  23089=>"001000000",
  23090=>"000000100",
  23091=>"011000000",
  23092=>"000000000",
  23093=>"001001001",
  23094=>"000000000",
  23095=>"001000010",
  23096=>"000000100",
  23097=>"110110111",
  23098=>"000100111",
  23099=>"110111111",
  23100=>"111111111",
  23101=>"000000110",
  23102=>"000011011",
  23103=>"111111111",
  23104=>"000001111",
  23105=>"111011010",
  23106=>"111001000",
  23107=>"111011001",
  23108=>"001001011",
  23109=>"100100000",
  23110=>"000000001",
  23111=>"000000000",
  23112=>"100100000",
  23113=>"000000111",
  23114=>"111000001",
  23115=>"111111110",
  23116=>"110011011",
  23117=>"000000000",
  23118=>"000000000",
  23119=>"000000111",
  23120=>"111111111",
  23121=>"111011011",
  23122=>"000000000",
  23123=>"111111000",
  23124=>"000000000",
  23125=>"010111111",
  23126=>"111111111",
  23127=>"101111111",
  23128=>"001111111",
  23129=>"000000000",
  23130=>"000011111",
  23131=>"001000111",
  23132=>"001111111",
  23133=>"111111111",
  23134=>"000000111",
  23135=>"011111111",
  23136=>"000000000",
  23137=>"000000111",
  23138=>"000000000",
  23139=>"000000000",
  23140=>"111111101",
  23141=>"000000000",
  23142=>"000000000",
  23143=>"111001001",
  23144=>"111111111",
  23145=>"000000101",
  23146=>"111111111",
  23147=>"110010110",
  23148=>"100100110",
  23149=>"111111111",
  23150=>"000000000",
  23151=>"100000000",
  23152=>"000000000",
  23153=>"110000001",
  23154=>"011111001",
  23155=>"111111111",
  23156=>"000000000",
  23157=>"111111111",
  23158=>"000000000",
  23159=>"000000000",
  23160=>"111111000",
  23161=>"000111000",
  23162=>"000100100",
  23163=>"111111000",
  23164=>"011000011",
  23165=>"000000000",
  23166=>"000000000",
  23167=>"111000000",
  23168=>"111111111",
  23169=>"110110000",
  23170=>"000001001",
  23171=>"110110111",
  23172=>"000000101",
  23173=>"000000111",
  23174=>"001001000",
  23175=>"111111111",
  23176=>"111100100",
  23177=>"111101001",
  23178=>"111000000",
  23179=>"000000000",
  23180=>"000011000",
  23181=>"110110110",
  23182=>"111111111",
  23183=>"000000000",
  23184=>"111111111",
  23185=>"000100000",
  23186=>"000000000",
  23187=>"000111111",
  23188=>"111101111",
  23189=>"000000000",
  23190=>"111111111",
  23191=>"011100111",
  23192=>"000001111",
  23193=>"000000000",
  23194=>"011011111",
  23195=>"111011001",
  23196=>"001000000",
  23197=>"111111000",
  23198=>"001000100",
  23199=>"111111111",
  23200=>"100100111",
  23201=>"000100000",
  23202=>"111111011",
  23203=>"000000000",
  23204=>"001001111",
  23205=>"000111011",
  23206=>"000000000",
  23207=>"011011111",
  23208=>"011000000",
  23209=>"000000100",
  23210=>"000000000",
  23211=>"000000000",
  23212=>"111010111",
  23213=>"111011000",
  23214=>"111111111",
  23215=>"111111111",
  23216=>"000000000",
  23217=>"000001000",
  23218=>"111011011",
  23219=>"000100110",
  23220=>"111111000",
  23221=>"100101111",
  23222=>"101000000",
  23223=>"111000000",
  23224=>"000000000",
  23225=>"111111111",
  23226=>"101101111",
  23227=>"011011000",
  23228=>"111001000",
  23229=>"111011000",
  23230=>"000000000",
  23231=>"111111111",
  23232=>"111000111",
  23233=>"000111111",
  23234=>"111101100",
  23235=>"000000000",
  23236=>"111111011",
  23237=>"000000000",
  23238=>"111111111",
  23239=>"001000000",
  23240=>"111001001",
  23241=>"011000000",
  23242=>"110111010",
  23243=>"101101101",
  23244=>"110111111",
  23245=>"111111111",
  23246=>"111001000",
  23247=>"011111111",
  23248=>"000000000",
  23249=>"111111000",
  23250=>"000000000",
  23251=>"111011111",
  23252=>"100110001",
  23253=>"110111111",
  23254=>"000000000",
  23255=>"000000000",
  23256=>"111100100",
  23257=>"000001000",
  23258=>"111111111",
  23259=>"111111011",
  23260=>"111111111",
  23261=>"111111111",
  23262=>"111111111",
  23263=>"000000000",
  23264=>"000000000",
  23265=>"110111111",
  23266=>"000000000",
  23267=>"110111111",
  23268=>"011111000",
  23269=>"100000000",
  23270=>"111111011",
  23271=>"000011101",
  23272=>"111000000",
  23273=>"011111111",
  23274=>"000000101",
  23275=>"011111111",
  23276=>"101111111",
  23277=>"000000111",
  23278=>"000000100",
  23279=>"000000000",
  23280=>"111101100",
  23281=>"000000100",
  23282=>"110110000",
  23283=>"111111111",
  23284=>"110111111",
  23285=>"100000001",
  23286=>"011100000",
  23287=>"000000000",
  23288=>"000111110",
  23289=>"111111011",
  23290=>"001001001",
  23291=>"111111111",
  23292=>"111111100",
  23293=>"000111010",
  23294=>"001000101",
  23295=>"111001101",
  23296=>"001111111",
  23297=>"011111010",
  23298=>"111001000",
  23299=>"000000100",
  23300=>"111111000",
  23301=>"110000000",
  23302=>"100111111",
  23303=>"011011111",
  23304=>"111110111",
  23305=>"111000000",
  23306=>"101000000",
  23307=>"111110100",
  23308=>"000000000",
  23309=>"100110111",
  23310=>"001000000",
  23311=>"000000011",
  23312=>"110100000",
  23313=>"110110000",
  23314=>"000000000",
  23315=>"000111100",
  23316=>"100100000",
  23317=>"100111100",
  23318=>"001001111",
  23319=>"000000000",
  23320=>"110110110",
  23321=>"000000001",
  23322=>"000000000",
  23323=>"111100111",
  23324=>"011001001",
  23325=>"110111100",
  23326=>"111101100",
  23327=>"000000000",
  23328=>"111111110",
  23329=>"000110111",
  23330=>"000000000",
  23331=>"110000000",
  23332=>"000111111",
  23333=>"000000000",
  23334=>"110000000",
  23335=>"000110111",
  23336=>"000000100",
  23337=>"101111111",
  23338=>"000000000",
  23339=>"111111111",
  23340=>"011111111",
  23341=>"110100000",
  23342=>"000000000",
  23343=>"011011001",
  23344=>"111111110",
  23345=>"101100111",
  23346=>"111111000",
  23347=>"000000111",
  23348=>"000000000",
  23349=>"000100110",
  23350=>"011111111",
  23351=>"000000000",
  23352=>"000000000",
  23353=>"000000000",
  23354=>"101000000",
  23355=>"000000000",
  23356=>"100100100",
  23357=>"001000110",
  23358=>"111111101",
  23359=>"111101001",
  23360=>"101111110",
  23361=>"111111111",
  23362=>"001000111",
  23363=>"000101100",
  23364=>"111111001",
  23365=>"000000001",
  23366=>"111111111",
  23367=>"000000111",
  23368=>"000000000",
  23369=>"111000000",
  23370=>"111111000",
  23371=>"111111111",
  23372=>"111111111",
  23373=>"111011111",
  23374=>"000000000",
  23375=>"110100110",
  23376=>"000000100",
  23377=>"111111000",
  23378=>"111110000",
  23379=>"111111011",
  23380=>"000000000",
  23381=>"111111111",
  23382=>"000000100",
  23383=>"010100110",
  23384=>"111110100",
  23385=>"000000000",
  23386=>"111000110",
  23387=>"111111110",
  23388=>"000111101",
  23389=>"111111111",
  23390=>"000000000",
  23391=>"000001000",
  23392=>"111110111",
  23393=>"000000000",
  23394=>"000100111",
  23395=>"111111111",
  23396=>"111111111",
  23397=>"000000000",
  23398=>"110111101",
  23399=>"000000000",
  23400=>"111100111",
  23401=>"011011000",
  23402=>"001000000",
  23403=>"000000000",
  23404=>"000000000",
  23405=>"011011110",
  23406=>"111111000",
  23407=>"011011011",
  23408=>"000000001",
  23409=>"101101111",
  23410=>"011110111",
  23411=>"000000100",
  23412=>"000000000",
  23413=>"000000000",
  23414=>"111111110",
  23415=>"010010000",
  23416=>"000000000",
  23417=>"000000000",
  23418=>"000000000",
  23419=>"000000010",
  23420=>"000000000",
  23421=>"001111111",
  23422=>"100110110",
  23423=>"111111110",
  23424=>"000000001",
  23425=>"110111111",
  23426=>"011011001",
  23427=>"000100111",
  23428=>"111111111",
  23429=>"101000000",
  23430=>"101100111",
  23431=>"000001000",
  23432=>"000000111",
  23433=>"111111111",
  23434=>"000000000",
  23435=>"000111111",
  23436=>"111111010",
  23437=>"000000000",
  23438=>"111111111",
  23439=>"111101001",
  23440=>"111000000",
  23441=>"000000000",
  23442=>"101100000",
  23443=>"001001001",
  23444=>"111111111",
  23445=>"000000011",
  23446=>"000100000",
  23447=>"001000000",
  23448=>"111110100",
  23449=>"000000000",
  23450=>"101001011",
  23451=>"011001000",
  23452=>"100000000",
  23453=>"000000000",
  23454=>"000100101",
  23455=>"001001001",
  23456=>"101101111",
  23457=>"100101001",
  23458=>"100000000",
  23459=>"000000000",
  23460=>"011111111",
  23461=>"101001000",
  23462=>"111111000",
  23463=>"111110100",
  23464=>"111111000",
  23465=>"000000000",
  23466=>"000000000",
  23467=>"111110111",
  23468=>"111111111",
  23469=>"111011011",
  23470=>"111001000",
  23471=>"000000000",
  23472=>"111111111",
  23473=>"000000000",
  23474=>"111100111",
  23475=>"000000000",
  23476=>"111111001",
  23477=>"000010111",
  23478=>"000000000",
  23479=>"000000000",
  23480=>"000111111",
  23481=>"111111011",
  23482=>"000000000",
  23483=>"100100000",
  23484=>"001001000",
  23485=>"111111111",
  23486=>"111111110",
  23487=>"001011011",
  23488=>"000000000",
  23489=>"111111111",
  23490=>"000000000",
  23491=>"000000111",
  23492=>"000100100",
  23493=>"001001011",
  23494=>"000000001",
  23495=>"000000000",
  23496=>"111111111",
  23497=>"111111001",
  23498=>"000000000",
  23499=>"111111000",
  23500=>"111000000",
  23501=>"111110111",
  23502=>"000000000",
  23503=>"000111111",
  23504=>"000000110",
  23505=>"110110000",
  23506=>"001111111",
  23507=>"111111000",
  23508=>"011011011",
  23509=>"111111111",
  23510=>"111011000",
  23511=>"110110110",
  23512=>"110110000",
  23513=>"111100000",
  23514=>"000000000",
  23515=>"001000000",
  23516=>"111111111",
  23517=>"000000000",
  23518=>"011000111",
  23519=>"001111111",
  23520=>"111101111",
  23521=>"010010000",
  23522=>"111111111",
  23523=>"000000000",
  23524=>"111111011",
  23525=>"111011000",
  23526=>"000000111",
  23527=>"111111111",
  23528=>"111111000",
  23529=>"000000010",
  23530=>"100000000",
  23531=>"100000000",
  23532=>"000000000",
  23533=>"101100111",
  23534=>"111110111",
  23535=>"100000000",
  23536=>"000000000",
  23537=>"111101000",
  23538=>"000000000",
  23539=>"000000000",
  23540=>"111111111",
  23541=>"000010000",
  23542=>"111111111",
  23543=>"001000000",
  23544=>"000000000",
  23545=>"100100100",
  23546=>"000000000",
  23547=>"000000000",
  23548=>"011011111",
  23549=>"111111011",
  23550=>"111111111",
  23551=>"000000000",
  23552=>"001000001",
  23553=>"111111000",
  23554=>"000000101",
  23555=>"000000000",
  23556=>"001001111",
  23557=>"011010010",
  23558=>"000000000",
  23559=>"111000100",
  23560=>"000000000",
  23561=>"000100000",
  23562=>"000000000",
  23563=>"000000000",
  23564=>"100111111",
  23565=>"110100110",
  23566=>"110110111",
  23567=>"111111111",
  23568=>"110000001",
  23569=>"000111111",
  23570=>"001011011",
  23571=>"011111111",
  23572=>"001001000",
  23573=>"100000000",
  23574=>"111111111",
  23575=>"001000000",
  23576=>"010110110",
  23577=>"111111100",
  23578=>"111001010",
  23579=>"111001001",
  23580=>"111111000",
  23581=>"000000001",
  23582=>"111110110",
  23583=>"000100110",
  23584=>"001111111",
  23585=>"000000110",
  23586=>"000000000",
  23587=>"111111111",
  23588=>"011111111",
  23589=>"110111111",
  23590=>"001000011",
  23591=>"000000000",
  23592=>"000000000",
  23593=>"111000110",
  23594=>"000000010",
  23595=>"001000001",
  23596=>"111111111",
  23597=>"011011000",
  23598=>"001100111",
  23599=>"001000000",
  23600=>"001000110",
  23601=>"000000000",
  23602=>"000000000",
  23603=>"100110111",
  23604=>"100111111",
  23605=>"001001010",
  23606=>"000000000",
  23607=>"000000000",
  23608=>"000000000",
  23609=>"111000100",
  23610=>"111111110",
  23611=>"001111010",
  23612=>"001000011",
  23613=>"111111111",
  23614=>"000111000",
  23615=>"111111111",
  23616=>"000000111",
  23617=>"110000001",
  23618=>"000110111",
  23619=>"001000011",
  23620=>"110010010",
  23621=>"000000110",
  23622=>"010010000",
  23623=>"111100100",
  23624=>"110110110",
  23625=>"000000000",
  23626=>"110010000",
  23627=>"100000001",
  23628=>"011010000",
  23629=>"011111111",
  23630=>"110110000",
  23631=>"000000000",
  23632=>"110000000",
  23633=>"010001000",
  23634=>"000000000",
  23635=>"000000000",
  23636=>"111111111",
  23637=>"110100100",
  23638=>"100000111",
  23639=>"011011011",
  23640=>"111111111",
  23641=>"001001001",
  23642=>"111111111",
  23643=>"111011111",
  23644=>"011100000",
  23645=>"011111010",
  23646=>"000000000",
  23647=>"000100001",
  23648=>"001001101",
  23649=>"111000000",
  23650=>"000011011",
  23651=>"111111111",
  23652=>"000000000",
  23653=>"000000111",
  23654=>"011111111",
  23655=>"000000011",
  23656=>"000000000",
  23657=>"101111110",
  23658=>"000000001",
  23659=>"011011000",
  23660=>"000000000",
  23661=>"000000001",
  23662=>"000000000",
  23663=>"000000001",
  23664=>"001000000",
  23665=>"111111111",
  23666=>"100100100",
  23667=>"111111111",
  23668=>"011001001",
  23669=>"111111111",
  23670=>"010010010",
  23671=>"000000000",
  23672=>"000000000",
  23673=>"000001000",
  23674=>"000000000",
  23675=>"110110111",
  23676=>"010110110",
  23677=>"110110110",
  23678=>"000000000",
  23679=>"000000000",
  23680=>"000100110",
  23681=>"111111111",
  23682=>"110110110",
  23683=>"110110100",
  23684=>"001111111",
  23685=>"000000000",
  23686=>"111111000",
  23687=>"000010111",
  23688=>"111111111",
  23689=>"111111001",
  23690=>"110110110",
  23691=>"001000000",
  23692=>"100000000",
  23693=>"111111011",
  23694=>"111111111",
  23695=>"011011011",
  23696=>"000000000",
  23697=>"000000000",
  23698=>"111111111",
  23699=>"000000000",
  23700=>"000111111",
  23701=>"000000110",
  23702=>"111111111",
  23703=>"000000000",
  23704=>"000000011",
  23705=>"000000001",
  23706=>"011010000",
  23707=>"010111110",
  23708=>"011000111",
  23709=>"111011001",
  23710=>"111111000",
  23711=>"000000001",
  23712=>"111110011",
  23713=>"111001000",
  23714=>"111111111",
  23715=>"001001000",
  23716=>"000000000",
  23717=>"111100110",
  23718=>"000111111",
  23719=>"011001001",
  23720=>"101000111",
  23721=>"000000000",
  23722=>"010111111",
  23723=>"111111111",
  23724=>"001000010",
  23725=>"000010000",
  23726=>"000000000",
  23727=>"111110001",
  23728=>"011000111",
  23729=>"111101000",
  23730=>"000111111",
  23731=>"000000110",
  23732=>"000110011",
  23733=>"000000001",
  23734=>"111111110",
  23735=>"110100111",
  23736=>"111111001",
  23737=>"001001001",
  23738=>"000110111",
  23739=>"011011111",
  23740=>"001000001",
  23741=>"100111100",
  23742=>"110110101",
  23743=>"000000000",
  23744=>"111100100",
  23745=>"111011111",
  23746=>"111011011",
  23747=>"010000000",
  23748=>"111111111",
  23749=>"010110001",
  23750=>"000000010",
  23751=>"001010111",
  23752=>"010000000",
  23753=>"000000001",
  23754=>"110010011",
  23755=>"111111111",
  23756=>"110111111",
  23757=>"111111000",
  23758=>"111110110",
  23759=>"011011010",
  23760=>"111000000",
  23761=>"110100110",
  23762=>"111100001",
  23763=>"000000000",
  23764=>"101101001",
  23765=>"000000100",
  23766=>"111111111",
  23767=>"001000001",
  23768=>"000000111",
  23769=>"000000000",
  23770=>"100100000",
  23771=>"001011111",
  23772=>"000000000",
  23773=>"001000000",
  23774=>"111011111",
  23775=>"011000000",
  23776=>"101000000",
  23777=>"001000000",
  23778=>"111111111",
  23779=>"011001111",
  23780=>"111111111",
  23781=>"000011011",
  23782=>"110111110",
  23783=>"000000000",
  23784=>"001001001",
  23785=>"001001000",
  23786=>"101000001",
  23787=>"111111111",
  23788=>"000000000",
  23789=>"111111101",
  23790=>"001000110",
  23791=>"111111110",
  23792=>"110110011",
  23793=>"001001011",
  23794=>"000000000",
  23795=>"000000001",
  23796=>"011111111",
  23797=>"000100111",
  23798=>"000001011",
  23799=>"111111111",
  23800=>"111011011",
  23801=>"000000000",
  23802=>"111100110",
  23803=>"001000000",
  23804=>"000000100",
  23805=>"111011001",
  23806=>"111111111",
  23807=>"111001011",
  23808=>"100000000",
  23809=>"000011011",
  23810=>"000100110",
  23811=>"000000000",
  23812=>"000000000",
  23813=>"100000000",
  23814=>"011000000",
  23815=>"101111111",
  23816=>"111110111",
  23817=>"100110110",
  23818=>"010011011",
  23819=>"111111000",
  23820=>"111111111",
  23821=>"000001011",
  23822=>"000000111",
  23823=>"011011011",
  23824=>"111111111",
  23825=>"111110111",
  23826=>"000000000",
  23827=>"111111111",
  23828=>"000000000",
  23829=>"000000000",
  23830=>"110111111",
  23831=>"111011011",
  23832=>"101001000",
  23833=>"111111111",
  23834=>"111011011",
  23835=>"000000000",
  23836=>"000011110",
  23837=>"101111111",
  23838=>"111000000",
  23839=>"111111101",
  23840=>"000011001",
  23841=>"100100100",
  23842=>"000000000",
  23843=>"111001101",
  23844=>"110110010",
  23845=>"111111111",
  23846=>"000000001",
  23847=>"111111111",
  23848=>"000000000",
  23849=>"001001011",
  23850=>"111111111",
  23851=>"100100110",
  23852=>"111111111",
  23853=>"000000000",
  23854=>"000000000",
  23855=>"000000000",
  23856=>"010010110",
  23857=>"001001000",
  23858=>"111111110",
  23859=>"100111111",
  23860=>"001001111",
  23861=>"000000000",
  23862=>"001000000",
  23863=>"000000000",
  23864=>"110111111",
  23865=>"000001111",
  23866=>"000101101",
  23867=>"000000100",
  23868=>"111110011",
  23869=>"111010000",
  23870=>"011111111",
  23871=>"110111111",
  23872=>"111110110",
  23873=>"111111000",
  23874=>"000000110",
  23875=>"111111111",
  23876=>"111110010",
  23877=>"001001001",
  23878=>"110100100",
  23879=>"000000000",
  23880=>"111111111",
  23881=>"111111111",
  23882=>"000000000",
  23883=>"011111111",
  23884=>"111001000",
  23885=>"000000000",
  23886=>"111111111",
  23887=>"000000000",
  23888=>"001000010",
  23889=>"001111111",
  23890=>"101000001",
  23891=>"000000001",
  23892=>"000000000",
  23893=>"001001011",
  23894=>"000000000",
  23895=>"111111111",
  23896=>"111111111",
  23897=>"111111111",
  23898=>"000000000",
  23899=>"111111111",
  23900=>"000000000",
  23901=>"000000000",
  23902=>"111000011",
  23903=>"111011111",
  23904=>"000000111",
  23905=>"111001000",
  23906=>"111111001",
  23907=>"011000000",
  23908=>"000000000",
  23909=>"000000001",
  23910=>"000000000",
  23911=>"010010000",
  23912=>"111110100",
  23913=>"100100100",
  23914=>"000000000",
  23915=>"111110000",
  23916=>"001000000",
  23917=>"000100100",
  23918=>"000010000",
  23919=>"101000101",
  23920=>"000000001",
  23921=>"000000100",
  23922=>"000111000",
  23923=>"000110111",
  23924=>"110000100",
  23925=>"000000000",
  23926=>"111001000",
  23927=>"110110110",
  23928=>"111101111",
  23929=>"111111111",
  23930=>"111000000",
  23931=>"111000011",
  23932=>"111000000",
  23933=>"001000000",
  23934=>"001000000",
  23935=>"111111111",
  23936=>"000000000",
  23937=>"100000000",
  23938=>"000111111",
  23939=>"111111000",
  23940=>"000000000",
  23941=>"000000000",
  23942=>"000000000",
  23943=>"100000000",
  23944=>"111000100",
  23945=>"111111111",
  23946=>"010010010",
  23947=>"101111001",
  23948=>"111111111",
  23949=>"001011111",
  23950=>"000001111",
  23951=>"000000000",
  23952=>"000010011",
  23953=>"000000001",
  23954=>"000000111",
  23955=>"111001111",
  23956=>"000000000",
  23957=>"000101000",
  23958=>"000000010",
  23959=>"000010000",
  23960=>"011011111",
  23961=>"110000000",
  23962=>"111111011",
  23963=>"100111111",
  23964=>"000000011",
  23965=>"111111110",
  23966=>"000000011",
  23967=>"111111011",
  23968=>"001001001",
  23969=>"010011000",
  23970=>"111100101",
  23971=>"000100110",
  23972=>"111111111",
  23973=>"000000000",
  23974=>"000000000",
  23975=>"000000000",
  23976=>"000000000",
  23977=>"010000110",
  23978=>"000000000",
  23979=>"111110000",
  23980=>"000000000",
  23981=>"011000111",
  23982=>"000000100",
  23983=>"111111010",
  23984=>"000000000",
  23985=>"111111111",
  23986=>"000000110",
  23987=>"111111111",
  23988=>"111111000",
  23989=>"111111111",
  23990=>"111111111",
  23991=>"111111111",
  23992=>"011111000",
  23993=>"111111111",
  23994=>"011110110",
  23995=>"000000000",
  23996=>"000000000",
  23997=>"111111111",
  23998=>"111001000",
  23999=>"000010010",
  24000=>"011111011",
  24001=>"000000000",
  24002=>"000000000",
  24003=>"111111111",
  24004=>"111111111",
  24005=>"001010110",
  24006=>"011011011",
  24007=>"101100100",
  24008=>"111011011",
  24009=>"000000000",
  24010=>"000000000",
  24011=>"100110111",
  24012=>"000000000",
  24013=>"000001000",
  24014=>"000000000",
  24015=>"000000000",
  24016=>"101000000",
  24017=>"001000000",
  24018=>"000000001",
  24019=>"110111110",
  24020=>"110000000",
  24021=>"111011110",
  24022=>"001011011",
  24023=>"110110110",
  24024=>"000000001",
  24025=>"111111011",
  24026=>"111000000",
  24027=>"110100000",
  24028=>"000000000",
  24029=>"111111111",
  24030=>"000000000",
  24031=>"010010000",
  24032=>"001001001",
  24033=>"111111111",
  24034=>"000100000",
  24035=>"000000000",
  24036=>"000111111",
  24037=>"111111111",
  24038=>"111100111",
  24039=>"000001111",
  24040=>"111111111",
  24041=>"000000110",
  24042=>"000100100",
  24043=>"001011111",
  24044=>"111000000",
  24045=>"111111111",
  24046=>"101111111",
  24047=>"100000001",
  24048=>"000000000",
  24049=>"111111001",
  24050=>"001111111",
  24051=>"111000000",
  24052=>"000000000",
  24053=>"000000000",
  24054=>"000000010",
  24055=>"001000011",
  24056=>"010111010",
  24057=>"001000010",
  24058=>"111111000",
  24059=>"101000101",
  24060=>"000000000",
  24061=>"000000001",
  24062=>"000100011",
  24063=>"100111111",
  24064=>"000001111",
  24065=>"101000000",
  24066=>"101000000",
  24067=>"000000000",
  24068=>"111111111",
  24069=>"110100100",
  24070=>"110111110",
  24071=>"001001001",
  24072=>"111111111",
  24073=>"100111111",
  24074=>"111101100",
  24075=>"110100000",
  24076=>"110110110",
  24077=>"111111111",
  24078=>"000100111",
  24079=>"101000001",
  24080=>"111111001",
  24081=>"000010000",
  24082=>"000000001",
  24083=>"010000010",
  24084=>"100000100",
  24085=>"000001001",
  24086=>"111111111",
  24087=>"011111010",
  24088=>"110000000",
  24089=>"110110110",
  24090=>"111111001",
  24091=>"111000100",
  24092=>"111111111",
  24093=>"000000001",
  24094=>"001001011",
  24095=>"000000001",
  24096=>"000000100",
  24097=>"000000110",
  24098=>"011001001",
  24099=>"111111111",
  24100=>"111111111",
  24101=>"000001011",
  24102=>"110111010",
  24103=>"000000111",
  24104=>"110110111",
  24105=>"000000000",
  24106=>"100100100",
  24107=>"000011001",
  24108=>"111111111",
  24109=>"010011001",
  24110=>"111001001",
  24111=>"000000101",
  24112=>"000000000",
  24113=>"111111110",
  24114=>"110110110",
  24115=>"000000000",
  24116=>"001001001",
  24117=>"000000000",
  24118=>"111110111",
  24119=>"000000001",
  24120=>"000000000",
  24121=>"111101111",
  24122=>"111111111",
  24123=>"111000001",
  24124=>"100101111",
  24125=>"001000101",
  24126=>"110100100",
  24127=>"001001101",
  24128=>"110111111",
  24129=>"001001011",
  24130=>"110110110",
  24131=>"111111111",
  24132=>"001001011",
  24133=>"000000000",
  24134=>"100100111",
  24135=>"000000000",
  24136=>"000000100",
  24137=>"000000000",
  24138=>"111000000",
  24139=>"100100100",
  24140=>"000011111",
  24141=>"000001000",
  24142=>"100000111",
  24143=>"001011101",
  24144=>"000000001",
  24145=>"001100000",
  24146=>"000000110",
  24147=>"111101011",
  24148=>"111111000",
  24149=>"110000110",
  24150=>"111100100",
  24151=>"111110010",
  24152=>"111110010",
  24153=>"100000000",
  24154=>"111111011",
  24155=>"111111110",
  24156=>"001001001",
  24157=>"000001001",
  24158=>"110110110",
  24159=>"111111111",
  24160=>"011111111",
  24161=>"000000101",
  24162=>"000000110",
  24163=>"001001111",
  24164=>"110001000",
  24165=>"111111111",
  24166=>"000000010",
  24167=>"000000000",
  24168=>"100000100",
  24169=>"000000000",
  24170=>"000000000",
  24171=>"111110000",
  24172=>"001001000",
  24173=>"011001001",
  24174=>"111111000",
  24175=>"110111111",
  24176=>"011000000",
  24177=>"110110110",
  24178=>"100000000",
  24179=>"100100100",
  24180=>"000000000",
  24181=>"000000000",
  24182=>"111111111",
  24183=>"000001101",
  24184=>"000000110",
  24185=>"000000000",
  24186=>"111111111",
  24187=>"000000000",
  24188=>"101111011",
  24189=>"000000000",
  24190=>"000000001",
  24191=>"000000000",
  24192=>"000000111",
  24193=>"110010000",
  24194=>"111111000",
  24195=>"111111010",
  24196=>"111111110",
  24197=>"001000010",
  24198=>"001111111",
  24199=>"000000000",
  24200=>"000000000",
  24201=>"111111111",
  24202=>"111111111",
  24203=>"111101000",
  24204=>"110110000",
  24205=>"001001000",
  24206=>"111110110",
  24207=>"011101111",
  24208=>"101000001",
  24209=>"001000000",
  24210=>"000100111",
  24211=>"011010110",
  24212=>"110000010",
  24213=>"011011000",
  24214=>"001000001",
  24215=>"101001001",
  24216=>"000000000",
  24217=>"111111011",
  24218=>"000000000",
  24219=>"000000000",
  24220=>"110110110",
  24221=>"000101101",
  24222=>"111111010",
  24223=>"111111111",
  24224=>"111111111",
  24225=>"000111001",
  24226=>"100000111",
  24227=>"000010000",
  24228=>"110111111",
  24229=>"111110111",
  24230=>"001001101",
  24231=>"100101101",
  24232=>"000111111",
  24233=>"000100110",
  24234=>"111110110",
  24235=>"101111111",
  24236=>"000000110",
  24237=>"110111111",
  24238=>"110100000",
  24239=>"000000101",
  24240=>"000001011",
  24241=>"111111100",
  24242=>"011111111",
  24243=>"111000000",
  24244=>"000000100",
  24245=>"000001011",
  24246=>"000000000",
  24247=>"111111111",
  24248=>"000000101",
  24249=>"111111111",
  24250=>"111000000",
  24251=>"110110000",
  24252=>"000000000",
  24253=>"110100110",
  24254=>"111111111",
  24255=>"101000000",
  24256=>"000000000",
  24257=>"000000000",
  24258=>"000001001",
  24259=>"001000001",
  24260=>"111111111",
  24261=>"000000000",
  24262=>"000001000",
  24263=>"000000000",
  24264=>"001001010",
  24265=>"111111111",
  24266=>"111111110",
  24267=>"000000000",
  24268=>"000000010",
  24269=>"111111001",
  24270=>"000000011",
  24271=>"110111000",
  24272=>"110110100",
  24273=>"000110111",
  24274=>"000000001",
  24275=>"100000000",
  24276=>"111111111",
  24277=>"000000000",
  24278=>"100100100",
  24279=>"111111111",
  24280=>"000000110",
  24281=>"000000101",
  24282=>"111111111",
  24283=>"011000111",
  24284=>"000000000",
  24285=>"110001000",
  24286=>"110100000",
  24287=>"110000000",
  24288=>"100000111",
  24289=>"000110111",
  24290=>"100111011",
  24291=>"111110110",
  24292=>"000010000",
  24293=>"011001011",
  24294=>"110000000",
  24295=>"111111111",
  24296=>"000110010",
  24297=>"111111111",
  24298=>"000001111",
  24299=>"011111111",
  24300=>"111111111",
  24301=>"011111111",
  24302=>"111000000",
  24303=>"111001001",
  24304=>"111111000",
  24305=>"111111111",
  24306=>"111111111",
  24307=>"000000001",
  24308=>"001011111",
  24309=>"110110111",
  24310=>"011111011",
  24311=>"101101000",
  24312=>"001001000",
  24313=>"001001001",
  24314=>"000000000",
  24315=>"101111111",
  24316=>"111111101",
  24317=>"001001010",
  24318=>"110000000",
  24319=>"000000111",
  24320=>"000000101",
  24321=>"100000000",
  24322=>"000000000",
  24323=>"100100100",
  24324=>"100100111",
  24325=>"010000110",
  24326=>"001000000",
  24327=>"111010010",
  24328=>"000000000",
  24329=>"101101000",
  24330=>"011111111",
  24331=>"111100100",
  24332=>"111001001",
  24333=>"111111111",
  24334=>"000000000",
  24335=>"111111111",
  24336=>"010111101",
  24337=>"111110010",
  24338=>"100101100",
  24339=>"100100000",
  24340=>"111111110",
  24341=>"111111111",
  24342=>"001000000",
  24343=>"001000001",
  24344=>"001001001",
  24345=>"111000000",
  24346=>"100101000",
  24347=>"011011001",
  24348=>"000000001",
  24349=>"000000000",
  24350=>"000000000",
  24351=>"111111111",
  24352=>"110100000",
  24353=>"110110110",
  24354=>"000000000",
  24355=>"000000000",
  24356=>"100000101",
  24357=>"111111111",
  24358=>"001000101",
  24359=>"111101100",
  24360=>"001100000",
  24361=>"001000001",
  24362=>"111111010",
  24363=>"111100100",
  24364=>"111011011",
  24365=>"001011111",
  24366=>"101000111",
  24367=>"111111010",
  24368=>"111110110",
  24369=>"000000000",
  24370=>"000000000",
  24371=>"000000100",
  24372=>"000000000",
  24373=>"000000000",
  24374=>"111011010",
  24375=>"111111010",
  24376=>"100010010",
  24377=>"111111111",
  24378=>"111111101",
  24379=>"111111111",
  24380=>"000000100",
  24381=>"110000000",
  24382=>"111100100",
  24383=>"000000000",
  24384=>"111100111",
  24385=>"000000001",
  24386=>"100000000",
  24387=>"111111111",
  24388=>"000110111",
  24389=>"000000000",
  24390=>"011111111",
  24391=>"111111110",
  24392=>"101111111",
  24393=>"000110110",
  24394=>"111111111",
  24395=>"001001011",
  24396=>"000000001",
  24397=>"110100001",
  24398=>"010011011",
  24399=>"000000100",
  24400=>"000000010",
  24401=>"000001111",
  24402=>"110100111",
  24403=>"000001000",
  24404=>"010000100",
  24405=>"000000000",
  24406=>"000000000",
  24407=>"100000000",
  24408=>"000000010",
  24409=>"000000000",
  24410=>"111111101",
  24411=>"111111111",
  24412=>"111000000",
  24413=>"000000000",
  24414=>"001000000",
  24415=>"111111110",
  24416=>"000100111",
  24417=>"101100100",
  24418=>"110000100",
  24419=>"100110000",
  24420=>"110110010",
  24421=>"101000000",
  24422=>"000000111",
  24423=>"000000111",
  24424=>"111001000",
  24425=>"000000000",
  24426=>"001001110",
  24427=>"111111111",
  24428=>"000000000",
  24429=>"000000000",
  24430=>"111100000",
  24431=>"111100100",
  24432=>"000000101",
  24433=>"000100111",
  24434=>"001101001",
  24435=>"000000110",
  24436=>"100000100",
  24437=>"110110111",
  24438=>"000000000",
  24439=>"111111110",
  24440=>"111111111",
  24441=>"001001101",
  24442=>"010001000",
  24443=>"000000001",
  24444=>"001000110",
  24445=>"000001001",
  24446=>"110111111",
  24447=>"101000100",
  24448=>"110110110",
  24449=>"111111111",
  24450=>"110110111",
  24451=>"110110100",
  24452=>"001111111",
  24453=>"001101100",
  24454=>"000000000",
  24455=>"111111110",
  24456=>"100000000",
  24457=>"011010010",
  24458=>"000000000",
  24459=>"101001101",
  24460=>"101101111",
  24461=>"111111111",
  24462=>"000010010",
  24463=>"111111001",
  24464=>"111101001",
  24465=>"111111011",
  24466=>"100000001",
  24467=>"000000101",
  24468=>"110000111",
  24469=>"000010000",
  24470=>"111000000",
  24471=>"111101101",
  24472=>"111000000",
  24473=>"111111111",
  24474=>"001001001",
  24475=>"110110000",
  24476=>"000000000",
  24477=>"011110111",
  24478=>"001001001",
  24479=>"111111000",
  24480=>"000110111",
  24481=>"110100000",
  24482=>"111110000",
  24483=>"111111001",
  24484=>"001000000",
  24485=>"000001111",
  24486=>"111101111",
  24487=>"001011001",
  24488=>"001000000",
  24489=>"000000111",
  24490=>"110110111",
  24491=>"001000000",
  24492=>"111111110",
  24493=>"011111111",
  24494=>"110100100",
  24495=>"000000000",
  24496=>"000000100",
  24497=>"000000000",
  24498=>"110110110",
  24499=>"010000010",
  24500=>"001000001",
  24501=>"001000000",
  24502=>"100000000",
  24503=>"001000000",
  24504=>"000000100",
  24505=>"111110000",
  24506=>"100000000",
  24507=>"000001001",
  24508=>"001011001",
  24509=>"000000000",
  24510=>"111101111",
  24511=>"100000000",
  24512=>"000100100",
  24513=>"111111111",
  24514=>"111111111",
  24515=>"111011000",
  24516=>"111001001",
  24517=>"111010000",
  24518=>"101100001",
  24519=>"101000001",
  24520=>"010000000",
  24521=>"111010000",
  24522=>"001000111",
  24523=>"111001000",
  24524=>"001000000",
  24525=>"011011111",
  24526=>"101000000",
  24527=>"100000000",
  24528=>"001001001",
  24529=>"111111011",
  24530=>"000000000",
  24531=>"000000011",
  24532=>"100100100",
  24533=>"001001001",
  24534=>"000100110",
  24535=>"011111010",
  24536=>"000000000",
  24537=>"111111111",
  24538=>"000000110",
  24539=>"111110010",
  24540=>"111111111",
  24541=>"001000001",
  24542=>"011011011",
  24543=>"010000001",
  24544=>"000000001",
  24545=>"000000001",
  24546=>"110111111",
  24547=>"000000000",
  24548=>"011001000",
  24549=>"000000000",
  24550=>"100101101",
  24551=>"100100111",
  24552=>"000000000",
  24553=>"111111000",
  24554=>"000011000",
  24555=>"000000000",
  24556=>"111001111",
  24557=>"000111110",
  24558=>"001101111",
  24559=>"001111001",
  24560=>"011011011",
  24561=>"000000000",
  24562=>"110000100",
  24563=>"001000000",
  24564=>"000000000",
  24565=>"010000000",
  24566=>"010000000",
  24567=>"000000000",
  24568=>"000000111",
  24569=>"011000001",
  24570=>"110110100",
  24571=>"101000100",
  24572=>"001000110",
  24573=>"111111111",
  24574=>"111011011",
  24575=>"000000011",
  24576=>"111100000",
  24577=>"111111001",
  24578=>"111000000",
  24579=>"110111011",
  24580=>"000100110",
  24581=>"000000111",
  24582=>"000000000",
  24583=>"111111101",
  24584=>"111111000",
  24585=>"001011011",
  24586=>"000000000",
  24587=>"001000000",
  24588=>"101111111",
  24589=>"110100001",
  24590=>"111111101",
  24591=>"111111111",
  24592=>"111111111",
  24593=>"000101101",
  24594=>"011011111",
  24595=>"100100000",
  24596=>"000100000",
  24597=>"111000000",
  24598=>"111111111",
  24599=>"000100100",
  24600=>"000100000",
  24601=>"000011111",
  24602=>"000001111",
  24603=>"001001001",
  24604=>"000000000",
  24605=>"000000000",
  24606=>"011111111",
  24607=>"111111111",
  24608=>"111111110",
  24609=>"100000000",
  24610=>"001111110",
  24611=>"000000000",
  24612=>"000000000",
  24613=>"000000001",
  24614=>"111111000",
  24615=>"100111000",
  24616=>"000001000",
  24617=>"111001000",
  24618=>"110111011",
  24619=>"000000011",
  24620=>"111101110",
  24621=>"000111111",
  24622=>"111110100",
  24623=>"111111111",
  24624=>"110111111",
  24625=>"000011111",
  24626=>"000000110",
  24627=>"111101000",
  24628=>"110111000",
  24629=>"111111100",
  24630=>"111111110",
  24631=>"111010000",
  24632=>"000000000",
  24633=>"011001011",
  24634=>"000000000",
  24635=>"010111111",
  24636=>"111000000",
  24637=>"111101101",
  24638=>"111100000",
  24639=>"000000000",
  24640=>"111111101",
  24641=>"111111111",
  24642=>"000111110",
  24643=>"011111111",
  24644=>"111110110",
  24645=>"010001001",
  24646=>"000000000",
  24647=>"000000000",
  24648=>"001001101",
  24649=>"111111111",
  24650=>"111100000",
  24651=>"111001011",
  24652=>"111111100",
  24653=>"111111111",
  24654=>"100000001",
  24655=>"000111111",
  24656=>"111111000",
  24657=>"001011111",
  24658=>"000000000",
  24659=>"111101000",
  24660=>"000111111",
  24661=>"000001011",
  24662=>"000000000",
  24663=>"111111111",
  24664=>"111000000",
  24665=>"000100111",
  24666=>"110111111",
  24667=>"100100000",
  24668=>"001001101",
  24669=>"111111001",
  24670=>"000000000",
  24671=>"001111111",
  24672=>"111000000",
  24673=>"000000000",
  24674=>"111111001",
  24675=>"000111111",
  24676=>"111000000",
  24677=>"110010000",
  24678=>"111011001",
  24679=>"000000000",
  24680=>"000111010",
  24681=>"110000000",
  24682=>"111000110",
  24683=>"000000000",
  24684=>"001111111",
  24685=>"000000000",
  24686=>"011111111",
  24687=>"111111111",
  24688=>"001000000",
  24689=>"111101000",
  24690=>"111111101",
  24691=>"111111000",
  24692=>"000000000",
  24693=>"100111111",
  24694=>"000000000",
  24695=>"011111111",
  24696=>"100111101",
  24697=>"011111111",
  24698=>"011011011",
  24699=>"000000000",
  24700=>"101111000",
  24701=>"111111111",
  24702=>"000001000",
  24703=>"001111111",
  24704=>"111000010",
  24705=>"101111111",
  24706=>"110110110",
  24707=>"000000000",
  24708=>"111111011",
  24709=>"111101000",
  24710=>"111111000",
  24711=>"111001000",
  24712=>"001000000",
  24713=>"110001001",
  24714=>"000000000",
  24715=>"111111111",
  24716=>"111111001",
  24717=>"111011000",
  24718=>"111111111",
  24719=>"111111011",
  24720=>"000000000",
  24721=>"000101100",
  24722=>"000000000",
  24723=>"000110111",
  24724=>"000001000",
  24725=>"001000000",
  24726=>"110111111",
  24727=>"111111110",
  24728=>"000000000",
  24729=>"011001110",
  24730=>"111111110",
  24731=>"000000000",
  24732=>"110111000",
  24733=>"110110000",
  24734=>"111000000",
  24735=>"111000000",
  24736=>"111111001",
  24737=>"111111000",
  24738=>"000100111",
  24739=>"111111111",
  24740=>"010001001",
  24741=>"000000101",
  24742=>"111111100",
  24743=>"101111100",
  24744=>"000000000",
  24745=>"111111111",
  24746=>"111111111",
  24747=>"001000000",
  24748=>"000110111",
  24749=>"111111110",
  24750=>"111011000",
  24751=>"000000000",
  24752=>"000000000",
  24753=>"000111100",
  24754=>"000111111",
  24755=>"000000000",
  24756=>"111111111",
  24757=>"111100101",
  24758=>"000000001",
  24759=>"111000000",
  24760=>"110011001",
  24761=>"000110111",
  24762=>"000000000",
  24763=>"111011000",
  24764=>"001111111",
  24765=>"110111000",
  24766=>"000100110",
  24767=>"000000001",
  24768=>"000110111",
  24769=>"000000000",
  24770=>"111111111",
  24771=>"111111111",
  24772=>"001110000",
  24773=>"010000000",
  24774=>"000010111",
  24775=>"001000000",
  24776=>"100001000",
  24777=>"111111111",
  24778=>"100101000",
  24779=>"000001001",
  24780=>"011111111",
  24781=>"000000111",
  24782=>"000111111",
  24783=>"000000000",
  24784=>"000000111",
  24785=>"100110011",
  24786=>"111111111",
  24787=>"000000010",
  24788=>"000000000",
  24789=>"110111111",
  24790=>"011000000",
  24791=>"000000100",
  24792=>"000000000",
  24793=>"111111110",
  24794=>"000000000",
  24795=>"000011011",
  24796=>"111001000",
  24797=>"000000000",
  24798=>"000000000",
  24799=>"110111000",
  24800=>"100000000",
  24801=>"000000001",
  24802=>"111111001",
  24803=>"111011000",
  24804=>"100111111",
  24805=>"111111101",
  24806=>"011111111",
  24807=>"111000000",
  24808=>"000000111",
  24809=>"111101001",
  24810=>"110111111",
  24811=>"111101111",
  24812=>"110111111",
  24813=>"001011010",
  24814=>"111111100",
  24815=>"000000000",
  24816=>"000111111",
  24817=>"011000000",
  24818=>"000111001",
  24819=>"111111000",
  24820=>"111111111",
  24821=>"000110111",
  24822=>"000100100",
  24823=>"111111111",
  24824=>"001000000",
  24825=>"000000000",
  24826=>"100000000",
  24827=>"011110111",
  24828=>"000000000",
  24829=>"001001100",
  24830=>"111011111",
  24831=>"001000000",
  24832=>"110111111",
  24833=>"010000000",
  24834=>"111111111",
  24835=>"111000000",
  24836=>"000000000",
  24837=>"000100000",
  24838=>"111111000",
  24839=>"111110101",
  24840=>"111111011",
  24841=>"000000111",
  24842=>"100001111",
  24843=>"110100100",
  24844=>"111101000",
  24845=>"000001100",
  24846=>"110101000",
  24847=>"111010000",
  24848=>"111111111",
  24849=>"011111001",
  24850=>"000000000",
  24851=>"011111000",
  24852=>"111111001",
  24853=>"011111000",
  24854=>"001111100",
  24855=>"000000011",
  24856=>"001111111",
  24857=>"000000000",
  24858=>"011011000",
  24859=>"111111111",
  24860=>"001000000",
  24861=>"000000000",
  24862=>"000111111",
  24863=>"000000000",
  24864=>"101000000",
  24865=>"000000110",
  24866=>"000000000",
  24867=>"111111111",
  24868=>"111011011",
  24869=>"110111101",
  24870=>"010111000",
  24871=>"111111001",
  24872=>"000000000",
  24873=>"111111011",
  24874=>"111111001",
  24875=>"111111000",
  24876=>"000000000",
  24877=>"001111011",
  24878=>"111111010",
  24879=>"000000000",
  24880=>"000111000",
  24881=>"100111111",
  24882=>"000000001",
  24883=>"001000000",
  24884=>"000000000",
  24885=>"010001101",
  24886=>"111011111",
  24887=>"110000000",
  24888=>"000000000",
  24889=>"111000000",
  24890=>"111111111",
  24891=>"000111111",
  24892=>"111000000",
  24893=>"011111100",
  24894=>"100111000",
  24895=>"110100000",
  24896=>"111111001",
  24897=>"111111000",
  24898=>"111111111",
  24899=>"000111111",
  24900=>"000000100",
  24901=>"111111111",
  24902=>"000011111",
  24903=>"111000000",
  24904=>"100111001",
  24905=>"001010010",
  24906=>"111111011",
  24907=>"000100100",
  24908=>"111000000",
  24909=>"111111110",
  24910=>"001000000",
  24911=>"100100000",
  24912=>"111111011",
  24913=>"000001101",
  24914=>"000111110",
  24915=>"011001000",
  24916=>"011000000",
  24917=>"000000000",
  24918=>"111111111",
  24919=>"001010000",
  24920=>"001000000",
  24921=>"000000000",
  24922=>"011000000",
  24923=>"000000000",
  24924=>"110110000",
  24925=>"000111111",
  24926=>"111000001",
  24927=>"001111000",
  24928=>"000100111",
  24929=>"000000001",
  24930=>"101101001",
  24931=>"000100111",
  24932=>"000001111",
  24933=>"110110000",
  24934=>"101000000",
  24935=>"111111111",
  24936=>"011011001",
  24937=>"111111111",
  24938=>"000000000",
  24939=>"101100000",
  24940=>"111111110",
  24941=>"000000001",
  24942=>"110110110",
  24943=>"000000000",
  24944=>"111111111",
  24945=>"111111111",
  24946=>"111111110",
  24947=>"111111000",
  24948=>"100000000",
  24949=>"111111110",
  24950=>"001111000",
  24951=>"110110111",
  24952=>"111111111",
  24953=>"000111000",
  24954=>"001001000",
  24955=>"111000000",
  24956=>"000000110",
  24957=>"111111101",
  24958=>"111111111",
  24959=>"110111111",
  24960=>"111101100",
  24961=>"111001001",
  24962=>"100110110",
  24963=>"000100000",
  24964=>"000000111",
  24965=>"000100110",
  24966=>"100000001",
  24967=>"011011001",
  24968=>"000000000",
  24969=>"000001000",
  24970=>"111111000",
  24971=>"010111000",
  24972=>"000111111",
  24973=>"000101110",
  24974=>"111110100",
  24975=>"010110111",
  24976=>"001000000",
  24977=>"000000000",
  24978=>"000000000",
  24979=>"001001000",
  24980=>"111111110",
  24981=>"000000010",
  24982=>"000001000",
  24983=>"111110000",
  24984=>"111100000",
  24985=>"101101000",
  24986=>"111000000",
  24987=>"000101001",
  24988=>"111111111",
  24989=>"000000000",
  24990=>"111011011",
  24991=>"000000000",
  24992=>"110011000",
  24993=>"111110000",
  24994=>"111000111",
  24995=>"111111111",
  24996=>"111111111",
  24997=>"000111111",
  24998=>"000000000",
  24999=>"000000110",
  25000=>"000000000",
  25001=>"000000111",
  25002=>"111111111",
  25003=>"111111000",
  25004=>"010010000",
  25005=>"100000000",
  25006=>"111000000",
  25007=>"000111111",
  25008=>"000000000",
  25009=>"000000000",
  25010=>"011111111",
  25011=>"100000100",
  25012=>"111111011",
  25013=>"001000000",
  25014=>"000101111",
  25015=>"110000000",
  25016=>"000000000",
  25017=>"111111111",
  25018=>"101000000",
  25019=>"111111100",
  25020=>"111011000",
  25021=>"001001000",
  25022=>"111111101",
  25023=>"000001101",
  25024=>"000000000",
  25025=>"000111111",
  25026=>"111110010",
  25027=>"000000000",
  25028=>"111111111",
  25029=>"100000010",
  25030=>"111001111",
  25031=>"110110111",
  25032=>"011000000",
  25033=>"000100111",
  25034=>"011000000",
  25035=>"000000000",
  25036=>"000000000",
  25037=>"111111111",
  25038=>"000000001",
  25039=>"010111111",
  25040=>"110100000",
  25041=>"011000000",
  25042=>"001001001",
  25043=>"000000001",
  25044=>"111111111",
  25045=>"000101101",
  25046=>"000100111",
  25047=>"011001001",
  25048=>"000000000",
  25049=>"001001001",
  25050=>"000000000",
  25051=>"111101000",
  25052=>"000000001",
  25053=>"110111000",
  25054=>"111011000",
  25055=>"000001011",
  25056=>"011111111",
  25057=>"111000000",
  25058=>"000000000",
  25059=>"111101001",
  25060=>"111111000",
  25061=>"000000110",
  25062=>"111111000",
  25063=>"000000000",
  25064=>"111111000",
  25065=>"000000000",
  25066=>"111111011",
  25067=>"000000111",
  25068=>"000000111",
  25069=>"001001101",
  25070=>"001001001",
  25071=>"110010000",
  25072=>"000000000",
  25073=>"000000000",
  25074=>"000100000",
  25075=>"111110000",
  25076=>"000000000",
  25077=>"000000111",
  25078=>"000000111",
  25079=>"000001000",
  25080=>"100000011",
  25081=>"000100101",
  25082=>"001111111",
  25083=>"000000000",
  25084=>"000000000",
  25085=>"111111011",
  25086=>"001000000",
  25087=>"000000000",
  25088=>"000111111",
  25089=>"111000100",
  25090=>"000011111",
  25091=>"000000100",
  25092=>"100111111",
  25093=>"001101001",
  25094=>"000100110",
  25095=>"111111111",
  25096=>"011011111",
  25097=>"000000000",
  25098=>"111111111",
  25099=>"000000000",
  25100=>"110111100",
  25101=>"100100000",
  25102=>"000000111",
  25103=>"110111110",
  25104=>"111100100",
  25105=>"000110111",
  25106=>"000000101",
  25107=>"111010000",
  25108=>"111000000",
  25109=>"111111111",
  25110=>"000000000",
  25111=>"111011011",
  25112=>"001111111",
  25113=>"100100100",
  25114=>"111000000",
  25115=>"000000111",
  25116=>"100000000",
  25117=>"111110000",
  25118=>"111101001",
  25119=>"000000010",
  25120=>"000001001",
  25121=>"111110101",
  25122=>"000001101",
  25123=>"000000000",
  25124=>"111111111",
  25125=>"000111111",
  25126=>"000001110",
  25127=>"000000111",
  25128=>"001001000",
  25129=>"100000000",
  25130=>"100001001",
  25131=>"100000001",
  25132=>"111111001",
  25133=>"000000111",
  25134=>"111011000",
  25135=>"010100100",
  25136=>"000011111",
  25137=>"000000100",
  25138=>"011111111",
  25139=>"100000001",
  25140=>"110101101",
  25141=>"011011000",
  25142=>"011111111",
  25143=>"000000000",
  25144=>"000000111",
  25145=>"000000111",
  25146=>"110111000",
  25147=>"110010000",
  25148=>"000000110",
  25149=>"011110110",
  25150=>"110111110",
  25151=>"111011001",
  25152=>"110000011",
  25153=>"111111000",
  25154=>"010111111",
  25155=>"110100111",
  25156=>"111001001",
  25157=>"111110100",
  25158=>"111000000",
  25159=>"000000100",
  25160=>"111111011",
  25161=>"000000000",
  25162=>"000110000",
  25163=>"000000001",
  25164=>"000000111",
  25165=>"001011101",
  25166=>"000000000",
  25167=>"111000001",
  25168=>"011000000",
  25169=>"001100000",
  25170=>"000000111",
  25171=>"001011111",
  25172=>"000000000",
  25173=>"100000111",
  25174=>"000000001",
  25175=>"000000111",
  25176=>"000000000",
  25177=>"000000000",
  25178=>"111111000",
  25179=>"011011011",
  25180=>"110111111",
  25181=>"111000000",
  25182=>"000111001",
  25183=>"111110000",
  25184=>"000000000",
  25185=>"000000111",
  25186=>"000000101",
  25187=>"111000111",
  25188=>"000000000",
  25189=>"000000000",
  25190=>"110100000",
  25191=>"000000000",
  25192=>"111111111",
  25193=>"010000000",
  25194=>"000011111",
  25195=>"000000000",
  25196=>"001001011",
  25197=>"000000011",
  25198=>"000000000",
  25199=>"000000111",
  25200=>"111000001",
  25201=>"000111111",
  25202=>"111111111",
  25203=>"000001000",
  25204=>"000000000",
  25205=>"110110111",
  25206=>"011000000",
  25207=>"000000000",
  25208=>"111111111",
  25209=>"000000100",
  25210=>"000000000",
  25211=>"111000000",
  25212=>"000011111",
  25213=>"001001111",
  25214=>"000000000",
  25215=>"111111111",
  25216=>"110000000",
  25217=>"110000000",
  25218=>"111111000",
  25219=>"111101100",
  25220=>"111011010",
  25221=>"101000000",
  25222=>"000000111",
  25223=>"000000000",
  25224=>"101011001",
  25225=>"100000000",
  25226=>"000000000",
  25227=>"000000000",
  25228=>"111001010",
  25229=>"010000000",
  25230=>"000100101",
  25231=>"000000000",
  25232=>"000000111",
  25233=>"000001011",
  25234=>"110110000",
  25235=>"000000111",
  25236=>"000000111",
  25237=>"000010111",
  25238=>"111000000",
  25239=>"111000111",
  25240=>"000000000",
  25241=>"111111110",
  25242=>"101000000",
  25243=>"011000000",
  25244=>"000000000",
  25245=>"111000000",
  25246=>"111111000",
  25247=>"000000000",
  25248=>"000000000",
  25249=>"000000111",
  25250=>"111101000",
  25251=>"000000000",
  25252=>"000000111",
  25253=>"000111111",
  25254=>"101000111",
  25255=>"000111110",
  25256=>"011001000",
  25257=>"000000110",
  25258=>"111000110",
  25259=>"111111111",
  25260=>"000000000",
  25261=>"100001111",
  25262=>"101111111",
  25263=>"000000000",
  25264=>"111000000",
  25265=>"111111001",
  25266=>"111111111",
  25267=>"000100111",
  25268=>"111000000",
  25269=>"000001101",
  25270=>"000000011",
  25271=>"000000011",
  25272=>"111000000",
  25273=>"011000000",
  25274=>"000001000",
  25275=>"000000111",
  25276=>"100000000",
  25277=>"111111000",
  25278=>"101111111",
  25279=>"000000000",
  25280=>"011111011",
  25281=>"000000111",
  25282=>"000000111",
  25283=>"111111101",
  25284=>"111111111",
  25285=>"000000011",
  25286=>"001000000",
  25287=>"000000111",
  25288=>"111000000",
  25289=>"110111111",
  25290=>"000000100",
  25291=>"001111111",
  25292=>"111110110",
  25293=>"000110111",
  25294=>"000000100",
  25295=>"000111000",
  25296=>"000111111",
  25297=>"000000000",
  25298=>"000111111",
  25299=>"000000000",
  25300=>"111111000",
  25301=>"001111111",
  25302=>"111111101",
  25303=>"000100101",
  25304=>"101111101",
  25305=>"000111111",
  25306=>"001111000",
  25307=>"111110000",
  25308=>"000111111",
  25309=>"001000000",
  25310=>"110110111",
  25311=>"111100111",
  25312=>"111001000",
  25313=>"001000000",
  25314=>"000111111",
  25315=>"111111100",
  25316=>"000000000",
  25317=>"111111100",
  25318=>"001000111",
  25319=>"000000000",
  25320=>"111111110",
  25321=>"111110110",
  25322=>"000000101",
  25323=>"111111111",
  25324=>"011000111",
  25325=>"011000011",
  25326=>"000000111",
  25327=>"000000000",
  25328=>"000000000",
  25329=>"111110011",
  25330=>"000000000",
  25331=>"001001111",
  25332=>"110111111",
  25333=>"111001001",
  25334=>"000110110",
  25335=>"011000000",
  25336=>"110100111",
  25337=>"000000000",
  25338=>"000000111",
  25339=>"000000111",
  25340=>"111011000",
  25341=>"111000110",
  25342=>"111111000",
  25343=>"000001111",
  25344=>"111111111",
  25345=>"110110110",
  25346=>"011111000",
  25347=>"111000100",
  25348=>"100110100",
  25349=>"000000100",
  25350=>"110100000",
  25351=>"011000000",
  25352=>"101000000",
  25353=>"000000000",
  25354=>"000000000",
  25355=>"000011111",
  25356=>"000000111",
  25357=>"111111111",
  25358=>"111101100",
  25359=>"000000011",
  25360=>"111111110",
  25361=>"000000000",
  25362=>"111000000",
  25363=>"000100111",
  25364=>"111111111",
  25365=>"000000111",
  25366=>"011011001",
  25367=>"000000111",
  25368=>"000111111",
  25369=>"100000110",
  25370=>"100111111",
  25371=>"000111111",
  25372=>"100100100",
  25373=>"011011000",
  25374=>"000000000",
  25375=>"000101111",
  25376=>"000001011",
  25377=>"001011111",
  25378=>"000000110",
  25379=>"101111000",
  25380=>"111000000",
  25381=>"111101100",
  25382=>"000000001",
  25383=>"011011010",
  25384=>"111111110",
  25385=>"000010111",
  25386=>"000001111",
  25387=>"111101111",
  25388=>"000000100",
  25389=>"000100110",
  25390=>"000101001",
  25391=>"000000110",
  25392=>"111111001",
  25393=>"000010111",
  25394=>"111111000",
  25395=>"111100111",
  25396=>"100000000",
  25397=>"000000011",
  25398=>"001000000",
  25399=>"111000000",
  25400=>"010110000",
  25401=>"111111000",
  25402=>"111111111",
  25403=>"000000100",
  25404=>"011001111",
  25405=>"101111100",
  25406=>"110111111",
  25407=>"000111000",
  25408=>"000000111",
  25409=>"000100110",
  25410=>"000000101",
  25411=>"111111010",
  25412=>"000000100",
  25413=>"001000000",
  25414=>"111000000",
  25415=>"000000000",
  25416=>"000100010",
  25417=>"000000000",
  25418=>"100011111",
  25419=>"000100110",
  25420=>"000000000",
  25421=>"000000000",
  25422=>"000110111",
  25423=>"110001001",
  25424=>"000000010",
  25425=>"000000111",
  25426=>"101111010",
  25427=>"000000000",
  25428=>"000000111",
  25429=>"011111110",
  25430=>"101111000",
  25431=>"111111111",
  25432=>"111111000",
  25433=>"000000000",
  25434=>"000101111",
  25435=>"111101000",
  25436=>"101111111",
  25437=>"010111111",
  25438=>"111000000",
  25439=>"111111111",
  25440=>"000000111",
  25441=>"000000111",
  25442=>"011110000",
  25443=>"100000000",
  25444=>"110111111",
  25445=>"000000000",
  25446=>"000000000",
  25447=>"000000111",
  25448=>"001101111",
  25449=>"111000000",
  25450=>"110000101",
  25451=>"111110000",
  25452=>"111111111",
  25453=>"001000000",
  25454=>"000000110",
  25455=>"000111111",
  25456=>"000000010",
  25457=>"000000111",
  25458=>"000000000",
  25459=>"111110110",
  25460=>"000000100",
  25461=>"000000000",
  25462=>"000000000",
  25463=>"100000111",
  25464=>"111110000",
  25465=>"110011001",
  25466=>"000100100",
  25467=>"011111000",
  25468=>"000000101",
  25469=>"000000100",
  25470=>"000000000",
  25471=>"111111000",
  25472=>"000110011",
  25473=>"000100110",
  25474=>"111001001",
  25475=>"000111111",
  25476=>"001001111",
  25477=>"000000111",
  25478=>"000000000",
  25479=>"001000000",
  25480=>"111000000",
  25481=>"100111111",
  25482=>"010000000",
  25483=>"111111111",
  25484=>"000000011",
  25485=>"001001111",
  25486=>"000000001",
  25487=>"000111111",
  25488=>"000000111",
  25489=>"000000000",
  25490=>"011001000",
  25491=>"110100000",
  25492=>"111111000",
  25493=>"000001000",
  25494=>"000111111",
  25495=>"000000000",
  25496=>"000110111",
  25497=>"111000000",
  25498=>"000111111",
  25499=>"001111111",
  25500=>"011001000",
  25501=>"010000000",
  25502=>"111001111",
  25503=>"111111110",
  25504=>"111111111",
  25505=>"000110111",
  25506=>"001001011",
  25507=>"001000000",
  25508=>"101111111",
  25509=>"000111111",
  25510=>"000000000",
  25511=>"000000000",
  25512=>"000000000",
  25513=>"011000101",
  25514=>"001001101",
  25515=>"001011011",
  25516=>"000000000",
  25517=>"111111110",
  25518=>"110000000",
  25519=>"001001010",
  25520=>"110111111",
  25521=>"111010000",
  25522=>"000000000",
  25523=>"111000111",
  25524=>"000001111",
  25525=>"001000000",
  25526=>"001111111",
  25527=>"111000000",
  25528=>"111111000",
  25529=>"111111111",
  25530=>"111110000",
  25531=>"111111111",
  25532=>"111111111",
  25533=>"110111111",
  25534=>"010111111",
  25535=>"110110000",
  25536=>"111111010",
  25537=>"111100111",
  25538=>"111000111",
  25539=>"000100000",
  25540=>"000111101",
  25541=>"001111111",
  25542=>"000000100",
  25543=>"110110000",
  25544=>"000000000",
  25545=>"000000000",
  25546=>"101000000",
  25547=>"000000000",
  25548=>"111000000",
  25549=>"111001000",
  25550=>"000000100",
  25551=>"000000000",
  25552=>"000011111",
  25553=>"000000011",
  25554=>"100110101",
  25555=>"101101111",
  25556=>"011111110",
  25557=>"111111000",
  25558=>"001001100",
  25559=>"111110110",
  25560=>"000010011",
  25561=>"011000000",
  25562=>"000000110",
  25563=>"000000001",
  25564=>"000111111",
  25565=>"001111111",
  25566=>"100111101",
  25567=>"000000000",
  25568=>"111100111",
  25569=>"110111111",
  25570=>"000000000",
  25571=>"000111110",
  25572=>"001001000",
  25573=>"100000000",
  25574=>"000000011",
  25575=>"111000000",
  25576=>"000011111",
  25577=>"010111111",
  25578=>"000000000",
  25579=>"000000111",
  25580=>"000111111",
  25581=>"001000100",
  25582=>"111111011",
  25583=>"001000000",
  25584=>"110111111",
  25585=>"000111111",
  25586=>"000000000",
  25587=>"011111111",
  25588=>"101111000",
  25589=>"111000000",
  25590=>"000000110",
  25591=>"100000101",
  25592=>"000111111",
  25593=>"100111110",
  25594=>"100111111",
  25595=>"111111111",
  25596=>"000111111",
  25597=>"000000000",
  25598=>"111001000",
  25599=>"100000000",
  25600=>"000000000",
  25601=>"111000000",
  25602=>"111101111",
  25603=>"000000001",
  25604=>"100000000",
  25605=>"111101101",
  25606=>"000000000",
  25607=>"100110000",
  25608=>"000000000",
  25609=>"111110111",
  25610=>"000000000",
  25611=>"000111111",
  25612=>"000100000",
  25613=>"100100100",
  25614=>"111001111",
  25615=>"110111111",
  25616=>"000100100",
  25617=>"000110000",
  25618=>"000111001",
  25619=>"111100100",
  25620=>"110111110",
  25621=>"000000000",
  25622=>"000000100",
  25623=>"110110000",
  25624=>"100000000",
  25625=>"010011001",
  25626=>"111000000",
  25627=>"110010000",
  25628=>"111001001",
  25629=>"000000000",
  25630=>"111001001",
  25631=>"000011111",
  25632=>"111111111",
  25633=>"111111111",
  25634=>"000001010",
  25635=>"111110010",
  25636=>"111011001",
  25637=>"000000100",
  25638=>"111000111",
  25639=>"111111111",
  25640=>"110000000",
  25641=>"000000000",
  25642=>"000000000",
  25643=>"000000000",
  25644=>"111111111",
  25645=>"000000000",
  25646=>"001010000",
  25647=>"000000000",
  25648=>"100000000",
  25649=>"000000111",
  25650=>"000111011",
  25651=>"001001011",
  25652=>"000010000",
  25653=>"000101001",
  25654=>"011001001",
  25655=>"000100100",
  25656=>"000000111",
  25657=>"100100100",
  25658=>"000000000",
  25659=>"001000000",
  25660=>"111001111",
  25661=>"100000000",
  25662=>"000100100",
  25663=>"000000000",
  25664=>"000101111",
  25665=>"010111010",
  25666=>"000110000",
  25667=>"111101000",
  25668=>"100000000",
  25669=>"011001000",
  25670=>"111111010",
  25671=>"000000000",
  25672=>"111111110",
  25673=>"111100000",
  25674=>"000000110",
  25675=>"111011111",
  25676=>"110110000",
  25677=>"000000110",
  25678=>"110111000",
  25679=>"111101111",
  25680=>"100000100",
  25681=>"110111011",
  25682=>"000110000",
  25683=>"111101110",
  25684=>"110110111",
  25685=>"110110000",
  25686=>"100100110",
  25687=>"000000000",
  25688=>"000000000",
  25689=>"111101001",
  25690=>"000000000",
  25691=>"111111111",
  25692=>"111111111",
  25693=>"111111111",
  25694=>"111000000",
  25695=>"110110110",
  25696=>"000000001",
  25697=>"011001000",
  25698=>"000000011",
  25699=>"111111111",
  25700=>"001000000",
  25701=>"111111111",
  25702=>"001011011",
  25703=>"010000000",
  25704=>"110111111",
  25705=>"000000000",
  25706=>"111111111",
  25707=>"110111111",
  25708=>"111111111",
  25709=>"111111111",
  25710=>"111111101",
  25711=>"111111111",
  25712=>"000000000",
  25713=>"111111110",
  25714=>"000000000",
  25715=>"001011111",
  25716=>"111001000",
  25717=>"111111111",
  25718=>"111111110",
  25719=>"011111000",
  25720=>"111111111",
  25721=>"110000101",
  25722=>"000000000",
  25723=>"111000000",
  25724=>"101111111",
  25725=>"000101111",
  25726=>"000000000",
  25727=>"111111100",
  25728=>"000000110",
  25729=>"111111101",
  25730=>"111111111",
  25731=>"111111111",
  25732=>"111111001",
  25733=>"100111111",
  25734=>"111111000",
  25735=>"111111010",
  25736=>"111111000",
  25737=>"111111001",
  25738=>"000000000",
  25739=>"000000111",
  25740=>"110111111",
  25741=>"011011011",
  25742=>"010011111",
  25743=>"000011011",
  25744=>"111111011",
  25745=>"101111111",
  25746=>"100000110",
  25747=>"000100100",
  25748=>"000000111",
  25749=>"000101011",
  25750=>"111111111",
  25751=>"111111000",
  25752=>"111111111",
  25753=>"111111000",
  25754=>"111111001",
  25755=>"000010000",
  25756=>"110100111",
  25757=>"111111110",
  25758=>"111111111",
  25759=>"000000000",
  25760=>"000000000",
  25761=>"000000000",
  25762=>"000000000",
  25763=>"000000000",
  25764=>"100111111",
  25765=>"111111111",
  25766=>"000000000",
  25767=>"011111111",
  25768=>"111111111",
  25769=>"111111100",
  25770=>"000000000",
  25771=>"000000000",
  25772=>"111001000",
  25773=>"001111110",
  25774=>"111111111",
  25775=>"000111111",
  25776=>"000000000",
  25777=>"000000100",
  25778=>"111111111",
  25779=>"000000000",
  25780=>"111111011",
  25781=>"100000000",
  25782=>"000000001",
  25783=>"000000000",
  25784=>"000000000",
  25785=>"111111111",
  25786=>"101111111",
  25787=>"100000000",
  25788=>"111001001",
  25789=>"010000000",
  25790=>"111111010",
  25791=>"110110100",
  25792=>"101100101",
  25793=>"000000100",
  25794=>"000100000",
  25795=>"000000000",
  25796=>"111111111",
  25797=>"111111111",
  25798=>"011111110",
  25799=>"110111111",
  25800=>"000001000",
  25801=>"000000000",
  25802=>"100000000",
  25803=>"000000000",
  25804=>"000111111",
  25805=>"111111111",
  25806=>"110000000",
  25807=>"111100001",
  25808=>"011001000",
  25809=>"001011000",
  25810=>"111011011",
  25811=>"000110111",
  25812=>"000011111",
  25813=>"110110111",
  25814=>"000000000",
  25815=>"010010111",
  25816=>"110100000",
  25817=>"011010000",
  25818=>"000111000",
  25819=>"000111011",
  25820=>"000000000",
  25821=>"000100110",
  25822=>"000000110",
  25823=>"110000000",
  25824=>"000000111",
  25825=>"111111111",
  25826=>"000010111",
  25827=>"000000000",
  25828=>"000000111",
  25829=>"111111111",
  25830=>"000000000",
  25831=>"110111111",
  25832=>"111111000",
  25833=>"010010001",
  25834=>"111000000",
  25835=>"111111111",
  25836=>"111111111",
  25837=>"011000100",
  25838=>"110100111",
  25839=>"000000000",
  25840=>"100110111",
  25841=>"111111110",
  25842=>"111111111",
  25843=>"111111111",
  25844=>"111111111",
  25845=>"111001000",
  25846=>"000011010",
  25847=>"111100000",
  25848=>"111000000",
  25849=>"110000000",
  25850=>"100000000",
  25851=>"111111000",
  25852=>"111111101",
  25853=>"010000001",
  25854=>"111101111",
  25855=>"000000000",
  25856=>"010010000",
  25857=>"001001000",
  25858=>"100111111",
  25859=>"010000000",
  25860=>"111111000",
  25861=>"000000000",
  25862=>"111111100",
  25863=>"000010110",
  25864=>"000000100",
  25865=>"000110111",
  25866=>"100100000",
  25867=>"111111111",
  25868=>"000001101",
  25869=>"111111111",
  25870=>"111111111",
  25871=>"000001001",
  25872=>"100110100",
  25873=>"000100000",
  25874=>"000000011",
  25875=>"000111111",
  25876=>"000111111",
  25877=>"111111111",
  25878=>"001011010",
  25879=>"100000111",
  25880=>"000000001",
  25881=>"000000000",
  25882=>"000000000",
  25883=>"100111100",
  25884=>"110111111",
  25885=>"000000000",
  25886=>"111111111",
  25887=>"000000111",
  25888=>"001011011",
  25889=>"110111111",
  25890=>"111111111",
  25891=>"111111010",
  25892=>"111100100",
  25893=>"110111000",
  25894=>"100110100",
  25895=>"111111111",
  25896=>"110100000",
  25897=>"000110110",
  25898=>"111111001",
  25899=>"110001001",
  25900=>"000000110",
  25901=>"001000000",
  25902=>"001000011",
  25903=>"111111111",
  25904=>"110111110",
  25905=>"101000011",
  25906=>"000000000",
  25907=>"001101101",
  25908=>"000000000",
  25909=>"110000000",
  25910=>"110000000",
  25911=>"110111010",
  25912=>"001000000",
  25913=>"000001111",
  25914=>"111111110",
  25915=>"000000000",
  25916=>"011111111",
  25917=>"000000001",
  25918=>"000111111",
  25919=>"000111111",
  25920=>"000000000",
  25921=>"111111000",
  25922=>"000000000",
  25923=>"111111111",
  25924=>"111111111",
  25925=>"000111111",
  25926=>"000000001",
  25927=>"111111111",
  25928=>"111100111",
  25929=>"000000000",
  25930=>"111010000",
  25931=>"100100000",
  25932=>"110111100",
  25933=>"111000000",
  25934=>"110111111",
  25935=>"111011001",
  25936=>"110110111",
  25937=>"000000000",
  25938=>"111100110",
  25939=>"100000000",
  25940=>"000000000",
  25941=>"011011111",
  25942=>"111101111",
  25943=>"000000000",
  25944=>"111001011",
  25945=>"100000000",
  25946=>"100101000",
  25947=>"111111000",
  25948=>"000000000",
  25949=>"110111111",
  25950=>"010010110",
  25951=>"111000000",
  25952=>"111110000",
  25953=>"000000000",
  25954=>"111000000",
  25955=>"101101101",
  25956=>"110111000",
  25957=>"101001111",
  25958=>"110111111",
  25959=>"100000000",
  25960=>"011000000",
  25961=>"111111100",
  25962=>"000000000",
  25963=>"011111110",
  25964=>"100111110",
  25965=>"100000010",
  25966=>"000100111",
  25967=>"000000000",
  25968=>"011101000",
  25969=>"111111111",
  25970=>"110111111",
  25971=>"000100100",
  25972=>"000000001",
  25973=>"111111110",
  25974=>"111000000",
  25975=>"100100000",
  25976=>"110111000",
  25977=>"011111110",
  25978=>"101111111",
  25979=>"010010000",
  25980=>"100110100",
  25981=>"111111111",
  25982=>"000000000",
  25983=>"110110110",
  25984=>"111111000",
  25985=>"111111111",
  25986=>"111111010",
  25987=>"111111111",
  25988=>"110111111",
  25989=>"111010000",
  25990=>"111000000",
  25991=>"001000000",
  25992=>"000001001",
  25993=>"110111111",
  25994=>"111111111",
  25995=>"000000000",
  25996=>"111111111",
  25997=>"001000000",
  25998=>"000000000",
  25999=>"000000000",
  26000=>"101101000",
  26001=>"001111011",
  26002=>"000100000",
  26003=>"110110110",
  26004=>"000000111",
  26005=>"011010011",
  26006=>"000000000",
  26007=>"100000111",
  26008=>"001111001",
  26009=>"001001001",
  26010=>"000000000",
  26011=>"000001001",
  26012=>"111111111",
  26013=>"000000000",
  26014=>"000110111",
  26015=>"000000000",
  26016=>"111101000",
  26017=>"111111001",
  26018=>"111110110",
  26019=>"111111000",
  26020=>"111011011",
  26021=>"000000000",
  26022=>"111111111",
  26023=>"010100111",
  26024=>"000000000",
  26025=>"000000000",
  26026=>"001001111",
  26027=>"000000001",
  26028=>"000010010",
  26029=>"111111111",
  26030=>"111110000",
  26031=>"000001111",
  26032=>"000000000",
  26033=>"100000000",
  26034=>"000001001",
  26035=>"000000111",
  26036=>"100000000",
  26037=>"100110000",
  26038=>"111000111",
  26039=>"000000000",
  26040=>"011000100",
  26041=>"000000100",
  26042=>"000000000",
  26043=>"110100000",
  26044=>"011111111",
  26045=>"111111111",
  26046=>"000000110",
  26047=>"011001000",
  26048=>"111001000",
  26049=>"010111111",
  26050=>"000000000",
  26051=>"111111111",
  26052=>"000010110",
  26053=>"001001011",
  26054=>"001110110",
  26055=>"000110111",
  26056=>"000010010",
  26057=>"111111000",
  26058=>"110111111",
  26059=>"111000000",
  26060=>"111110111",
  26061=>"000000000",
  26062=>"000000000",
  26063=>"000100101",
  26064=>"111111111",
  26065=>"000000000",
  26066=>"000000000",
  26067=>"111111111",
  26068=>"000000000",
  26069=>"100111111",
  26070=>"000111111",
  26071=>"001001011",
  26072=>"001001000",
  26073=>"100000000",
  26074=>"000111111",
  26075=>"000000000",
  26076=>"000000100",
  26077=>"110110110",
  26078=>"000000000",
  26079=>"101111100",
  26080=>"111111011",
  26081=>"001111100",
  26082=>"000000111",
  26083=>"000011000",
  26084=>"111111111",
  26085=>"111111000",
  26086=>"000000001",
  26087=>"111111100",
  26088=>"111111100",
  26089=>"000000000",
  26090=>"111001001",
  26091=>"000000000",
  26092=>"111111011",
  26093=>"010111111",
  26094=>"010001001",
  26095=>"110000000",
  26096=>"100100000",
  26097=>"111100000",
  26098=>"111000000",
  26099=>"000011010",
  26100=>"000010000",
  26101=>"000111111",
  26102=>"100111111",
  26103=>"111011111",
  26104=>"000000000",
  26105=>"000000001",
  26106=>"111111011",
  26107=>"111111111",
  26108=>"111111111",
  26109=>"111111111",
  26110=>"111111111",
  26111=>"111111110",
  26112=>"111111100",
  26113=>"001000000",
  26114=>"111111111",
  26115=>"000111111",
  26116=>"111111111",
  26117=>"110011111",
  26118=>"001011011",
  26119=>"001001111",
  26120=>"011000000",
  26121=>"000000000",
  26122=>"111111111",
  26123=>"001011101",
  26124=>"100110000",
  26125=>"110111111",
  26126=>"011001000",
  26127=>"000000000",
  26128=>"000000100",
  26129=>"000000000",
  26130=>"001000000",
  26131=>"000000001",
  26132=>"000100111",
  26133=>"111001001",
  26134=>"000000000",
  26135=>"011010110",
  26136=>"000000000",
  26137=>"000010110",
  26138=>"000001101",
  26139=>"111000000",
  26140=>"000000000",
  26141=>"101101001",
  26142=>"000110100",
  26143=>"011010000",
  26144=>"111100000",
  26145=>"000000000",
  26146=>"110110110",
  26147=>"011001011",
  26148=>"000000000",
  26149=>"000001001",
  26150=>"100000000",
  26151=>"000000000",
  26152=>"011111111",
  26153=>"111111111",
  26154=>"000000000",
  26155=>"111111100",
  26156=>"111000000",
  26157=>"111111111",
  26158=>"100000101",
  26159=>"111111111",
  26160=>"111111111",
  26161=>"100110110",
  26162=>"000000000",
  26163=>"000000001",
  26164=>"100101001",
  26165=>"111111110",
  26166=>"001000000",
  26167=>"110111111",
  26168=>"000110000",
  26169=>"111111101",
  26170=>"111111111",
  26171=>"111111001",
  26172=>"111111001",
  26173=>"011010000",
  26174=>"000100111",
  26175=>"000000000",
  26176=>"001001000",
  26177=>"111101000",
  26178=>"000000000",
  26179=>"000000000",
  26180=>"100110110",
  26181=>"000011011",
  26182=>"111111101",
  26183=>"000111111",
  26184=>"000000000",
  26185=>"111111000",
  26186=>"000000000",
  26187=>"000000000",
  26188=>"000000111",
  26189=>"111111110",
  26190=>"000000000",
  26191=>"000000000",
  26192=>"111111111",
  26193=>"100100001",
  26194=>"111111111",
  26195=>"111111111",
  26196=>"000000000",
  26197=>"000000000",
  26198=>"000000000",
  26199=>"111111000",
  26200=>"111111111",
  26201=>"111101111",
  26202=>"001000000",
  26203=>"111111100",
  26204=>"000000000",
  26205=>"000000000",
  26206=>"000000000",
  26207=>"111011011",
  26208=>"000000000",
  26209=>"000000000",
  26210=>"110111011",
  26211=>"000000100",
  26212=>"000000000",
  26213=>"011000001",
  26214=>"101000000",
  26215=>"100100111",
  26216=>"000000000",
  26217=>"000000000",
  26218=>"000001000",
  26219=>"000000000",
  26220=>"000100111",
  26221=>"001111111",
  26222=>"000000101",
  26223=>"011110100",
  26224=>"101000001",
  26225=>"111101001",
  26226=>"111010000",
  26227=>"011001001",
  26228=>"000000000",
  26229=>"000100110",
  26230=>"001000000",
  26231=>"000000000",
  26232=>"111010110",
  26233=>"000111111",
  26234=>"100100111",
  26235=>"111111111",
  26236=>"110110110",
  26237=>"111111111",
  26238=>"010111111",
  26239=>"000000000",
  26240=>"000000000",
  26241=>"111111111",
  26242=>"000000000",
  26243=>"011000000",
  26244=>"000000000",
  26245=>"111000111",
  26246=>"000000000",
  26247=>"111111001",
  26248=>"100100110",
  26249=>"000000000",
  26250=>"001000000",
  26251=>"000000001",
  26252=>"000100011",
  26253=>"111001001",
  26254=>"011000000",
  26255=>"111111001",
  26256=>"001000111",
  26257=>"000000000",
  26258=>"010110111",
  26259=>"010000000",
  26260=>"000000000",
  26261=>"000000000",
  26262=>"111111111",
  26263=>"000000111",
  26264=>"000000000",
  26265=>"000000000",
  26266=>"111111000",
  26267=>"000000000",
  26268=>"000000000",
  26269=>"001000110",
  26270=>"011001000",
  26271=>"000001111",
  26272=>"100000000",
  26273=>"111111111",
  26274=>"111111111",
  26275=>"111111111",
  26276=>"000001001",
  26277=>"011011000",
  26278=>"111111110",
  26279=>"111111001",
  26280=>"111001000",
  26281=>"000000001",
  26282=>"111111111",
  26283=>"000000000",
  26284=>"001001011",
  26285=>"110110000",
  26286=>"000000000",
  26287=>"111001111",
  26288=>"000000000",
  26289=>"000000000",
  26290=>"111111010",
  26291=>"111111000",
  26292=>"111101111",
  26293=>"011111000",
  26294=>"011000011",
  26295=>"000001011",
  26296=>"101000001",
  26297=>"111111011",
  26298=>"110001100",
  26299=>"110010000",
  26300=>"000001001",
  26301=>"000100000",
  26302=>"000001001",
  26303=>"111111111",
  26304=>"111111111",
  26305=>"000011011",
  26306=>"000000111",
  26307=>"111000000",
  26308=>"001000000",
  26309=>"000000111",
  26310=>"000000000",
  26311=>"111111111",
  26312=>"000000000",
  26313=>"000000000",
  26314=>"011111111",
  26315=>"000000000",
  26316=>"111111111",
  26317=>"111111111",
  26318=>"110011111",
  26319=>"001101100",
  26320=>"000000000",
  26321=>"100000000",
  26322=>"011001001",
  26323=>"000000000",
  26324=>"111111111",
  26325=>"111111111",
  26326=>"000000001",
  26327=>"111111111",
  26328=>"111111111",
  26329=>"111111111",
  26330=>"000000000",
  26331=>"111111111",
  26332=>"100100111",
  26333=>"111111111",
  26334=>"001001111",
  26335=>"010000000",
  26336=>"000000000",
  26337=>"000000000",
  26338=>"000000000",
  26339=>"111001000",
  26340=>"111010111",
  26341=>"110100010",
  26342=>"000000111",
  26343=>"100000101",
  26344=>"000111010",
  26345=>"111111111",
  26346=>"001000000",
  26347=>"111111101",
  26348=>"111111111",
  26349=>"000000111",
  26350=>"000011111",
  26351=>"111111111",
  26352=>"000010000",
  26353=>"111111110",
  26354=>"111111000",
  26355=>"110100001",
  26356=>"000000000",
  26357=>"111110010",
  26358=>"111110100",
  26359=>"111111000",
  26360=>"000000000",
  26361=>"110111000",
  26362=>"100111000",
  26363=>"001000000",
  26364=>"000001001",
  26365=>"000000000",
  26366=>"111111111",
  26367=>"110000000",
  26368=>"111111000",
  26369=>"011011000",
  26370=>"111111111",
  26371=>"111111111",
  26372=>"000000000",
  26373=>"000000000",
  26374=>"111111111",
  26375=>"111111111",
  26376=>"000000000",
  26377=>"000000100",
  26378=>"111111111",
  26379=>"000000000",
  26380=>"000000000",
  26381=>"111011001",
  26382=>"000001000",
  26383=>"000111111",
  26384=>"011000100",
  26385=>"000000000",
  26386=>"000000000",
  26387=>"011111111",
  26388=>"000000000",
  26389=>"000000000",
  26390=>"000100100",
  26391=>"000000000",
  26392=>"111111000",
  26393=>"111111111",
  26394=>"111111111",
  26395=>"000010110",
  26396=>"010010100",
  26397=>"111101000",
  26398=>"000000000",
  26399=>"000001001",
  26400=>"011111000",
  26401=>"110000000",
  26402=>"111111111",
  26403=>"000000000",
  26404=>"111001111",
  26405=>"110011111",
  26406=>"010011111",
  26407=>"000000000",
  26408=>"111111111",
  26409=>"011001001",
  26410=>"111111101",
  26411=>"101000100",
  26412=>"111111110",
  26413=>"000000000",
  26414=>"000010000",
  26415=>"000000110",
  26416=>"111001001",
  26417=>"000000000",
  26418=>"111110111",
  26419=>"000010111",
  26420=>"111111010",
  26421=>"011001001",
  26422=>"111011110",
  26423=>"001000000",
  26424=>"111111000",
  26425=>"111001111",
  26426=>"111111111",
  26427=>"001111011",
  26428=>"001011111",
  26429=>"111111001",
  26430=>"010110110",
  26431=>"011010000",
  26432=>"001000000",
  26433=>"000000000",
  26434=>"111111111",
  26435=>"000000000",
  26436=>"000000000",
  26437=>"111111111",
  26438=>"000000000",
  26439=>"000000000",
  26440=>"100100110",
  26441=>"111011000",
  26442=>"000011111",
  26443=>"111111100",
  26444=>"000000000",
  26445=>"111111111",
  26446=>"111111111",
  26447=>"010000100",
  26448=>"011111111",
  26449=>"111111111",
  26450=>"000000000",
  26451=>"111111110",
  26452=>"001111001",
  26453=>"011011011",
  26454=>"010000000",
  26455=>"111111111",
  26456=>"111111101",
  26457=>"101000000",
  26458=>"000000000",
  26459=>"111111111",
  26460=>"110100000",
  26461=>"010010000",
  26462=>"111110000",
  26463=>"001001011",
  26464=>"000000000",
  26465=>"111111111",
  26466=>"011011111",
  26467=>"001111111",
  26468=>"110111111",
  26469=>"000000100",
  26470=>"100000000",
  26471=>"110111111",
  26472=>"001100110",
  26473=>"011001001",
  26474=>"001011000",
  26475=>"000000000",
  26476=>"000000000",
  26477=>"111111111",
  26478=>"000001001",
  26479=>"000000000",
  26480=>"000000000",
  26481=>"011111010",
  26482=>"000000000",
  26483=>"111111011",
  26484=>"111111111",
  26485=>"111111111",
  26486=>"001001010",
  26487=>"000000100",
  26488=>"000000000",
  26489=>"000000000",
  26490=>"000000000",
  26491=>"111110110",
  26492=>"111111111",
  26493=>"111100000",
  26494=>"000000000",
  26495=>"111000000",
  26496=>"111111111",
  26497=>"000000000",
  26498=>"111111111",
  26499=>"111111111",
  26500=>"000010111",
  26501=>"100000111",
  26502=>"001000000",
  26503=>"111111111",
  26504=>"001000100",
  26505=>"000000111",
  26506=>"000000011",
  26507=>"000111110",
  26508=>"001001001",
  26509=>"011111001",
  26510=>"011000000",
  26511=>"001000000",
  26512=>"000000000",
  26513=>"001000000",
  26514=>"110111001",
  26515=>"100111111",
  26516=>"111111111",
  26517=>"000000000",
  26518=>"011011011",
  26519=>"000100000",
  26520=>"111111111",
  26521=>"111110110",
  26522=>"100000000",
  26523=>"011011100",
  26524=>"100100000",
  26525=>"111111110",
  26526=>"110111111",
  26527=>"000000000",
  26528=>"111111111",
  26529=>"000000000",
  26530=>"000000000",
  26531=>"001111111",
  26532=>"101001111",
  26533=>"111111111",
  26534=>"111001001",
  26535=>"000010010",
  26536=>"000000000",
  26537=>"111111111",
  26538=>"101100100",
  26539=>"111111011",
  26540=>"000000000",
  26541=>"001001000",
  26542=>"000101000",
  26543=>"000010001",
  26544=>"000000000",
  26545=>"010001001",
  26546=>"111000001",
  26547=>"000000111",
  26548=>"111101111",
  26549=>"111111111",
  26550=>"111111111",
  26551=>"000000000",
  26552=>"000000000",
  26553=>"011011000",
  26554=>"000000010",
  26555=>"000000101",
  26556=>"111111111",
  26557=>"001000000",
  26558=>"001000000",
  26559=>"000000100",
  26560=>"111110011",
  26561=>"000000000",
  26562=>"111111011",
  26563=>"001111111",
  26564=>"101000000",
  26565=>"011011000",
  26566=>"001001000",
  26567=>"111111111",
  26568=>"000000111",
  26569=>"000000000",
  26570=>"000000000",
  26571=>"111111111",
  26572=>"101111001",
  26573=>"000000000",
  26574=>"111000000",
  26575=>"100111111",
  26576=>"001000110",
  26577=>"011011001",
  26578=>"111111111",
  26579=>"111111111",
  26580=>"000001001",
  26581=>"111111111",
  26582=>"100111100",
  26583=>"000100000",
  26584=>"000011001",
  26585=>"000000000",
  26586=>"111111000",
  26587=>"000000000",
  26588=>"000101001",
  26589=>"111111111",
  26590=>"111111111",
  26591=>"010111011",
  26592=>"001000000",
  26593=>"100111111",
  26594=>"000000111",
  26595=>"000111111",
  26596=>"111011001",
  26597=>"111110100",
  26598=>"001000001",
  26599=>"110110110",
  26600=>"010111011",
  26601=>"000000000",
  26602=>"111111110",
  26603=>"000000000",
  26604=>"001101100",
  26605=>"001001001",
  26606=>"000000000",
  26607=>"000000000",
  26608=>"011111111",
  26609=>"000000000",
  26610=>"001000000",
  26611=>"000100000",
  26612=>"000000101",
  26613=>"110110111",
  26614=>"111111100",
  26615=>"000000100",
  26616=>"000000000",
  26617=>"000001001",
  26618=>"000000000",
  26619=>"111111000",
  26620=>"111111111",
  26621=>"111111100",
  26622=>"000000000",
  26623=>"011000000",
  26624=>"000000001",
  26625=>"010111111",
  26626=>"001000000",
  26627=>"111111010",
  26628=>"111101111",
  26629=>"111111111",
  26630=>"111111111",
  26631=>"111001000",
  26632=>"000000000",
  26633=>"111110110",
  26634=>"101101001",
  26635=>"111000000",
  26636=>"101111000",
  26637=>"110111111",
  26638=>"000000000",
  26639=>"111111111",
  26640=>"000000000",
  26641=>"011111110",
  26642=>"000000000",
  26643=>"000000000",
  26644=>"000000000",
  26645=>"001001101",
  26646=>"011111101",
  26647=>"111110000",
  26648=>"000000000",
  26649=>"011011001",
  26650=>"111111111",
  26651=>"111111111",
  26652=>"111111111",
  26653=>"000000000",
  26654=>"000000000",
  26655=>"000000101",
  26656=>"111101001",
  26657=>"111110111",
  26658=>"111001001",
  26659=>"110111111",
  26660=>"101000000",
  26661=>"000000000",
  26662=>"111101011",
  26663=>"110100111",
  26664=>"000110011",
  26665=>"011000100",
  26666=>"111111111",
  26667=>"000011111",
  26668=>"111111000",
  26669=>"110000000",
  26670=>"111111111",
  26671=>"000111111",
  26672=>"001001000",
  26673=>"000000000",
  26674=>"110100000",
  26675=>"000000000",
  26676=>"111111111",
  26677=>"110111111",
  26678=>"111111111",
  26679=>"000000000",
  26680=>"100111000",
  26681=>"000000000",
  26682=>"110110110",
  26683=>"000000000",
  26684=>"000000000",
  26685=>"100100000",
  26686=>"111111000",
  26687=>"111111010",
  26688=>"011011111",
  26689=>"011011011",
  26690=>"000000000",
  26691=>"111000000",
  26692=>"000000000",
  26693=>"111111110",
  26694=>"001000000",
  26695=>"001101111",
  26696=>"000111111",
  26697=>"111000111",
  26698=>"100000000",
  26699=>"110100001",
  26700=>"111111110",
  26701=>"000001000",
  26702=>"000000000",
  26703=>"000000001",
  26704=>"000000100",
  26705=>"000000000",
  26706=>"011111111",
  26707=>"001000000",
  26708=>"100101111",
  26709=>"000000000",
  26710=>"100100111",
  26711=>"111111001",
  26712=>"100000000",
  26713=>"101001111",
  26714=>"111111011",
  26715=>"100110010",
  26716=>"111110000",
  26717=>"000000001",
  26718=>"000000000",
  26719=>"111111111",
  26720=>"011111111",
  26721=>"000000000",
  26722=>"000000111",
  26723=>"001001000",
  26724=>"110110000",
  26725=>"101101000",
  26726=>"000000111",
  26727=>"011001111",
  26728=>"001001111",
  26729=>"111011011",
  26730=>"101111111",
  26731=>"101000111",
  26732=>"001001001",
  26733=>"111111000",
  26734=>"000000011",
  26735=>"111111111",
  26736=>"000010000",
  26737=>"000000111",
  26738=>"010110111",
  26739=>"001010000",
  26740=>"000010010",
  26741=>"000000001",
  26742=>"000000000",
  26743=>"100000001",
  26744=>"001000000",
  26745=>"111111111",
  26746=>"001000001",
  26747=>"000011000",
  26748=>"110110100",
  26749=>"000000000",
  26750=>"101001001",
  26751=>"000000011",
  26752=>"000000111",
  26753=>"101100111",
  26754=>"111111111",
  26755=>"000000000",
  26756=>"001001101",
  26757=>"000000000",
  26758=>"110111000",
  26759=>"111111111",
  26760=>"000000000",
  26761=>"000000111",
  26762=>"111111110",
  26763=>"000000011",
  26764=>"000000000",
  26765=>"100000000",
  26766=>"000000000",
  26767=>"000000000",
  26768=>"001000000",
  26769=>"111010010",
  26770=>"010000000",
  26771=>"000000000",
  26772=>"111011111",
  26773=>"110101000",
  26774=>"000111111",
  26775=>"001001000",
  26776=>"000000000",
  26777=>"111111010",
  26778=>"110110000",
  26779=>"000000000",
  26780=>"111111111",
  26781=>"000000000",
  26782=>"111101000",
  26783=>"000001000",
  26784=>"110000000",
  26785=>"110111111",
  26786=>"110000000",
  26787=>"000111111",
  26788=>"101001001",
  26789=>"000101111",
  26790=>"000000001",
  26791=>"011010000",
  26792=>"001001000",
  26793=>"001011111",
  26794=>"101001001",
  26795=>"111001111",
  26796=>"100111111",
  26797=>"110000000",
  26798=>"111111101",
  26799=>"111101111",
  26800=>"010111000",
  26801=>"111011011",
  26802=>"010011011",
  26803=>"100101000",
  26804=>"011011111",
  26805=>"000001011",
  26806=>"100000000",
  26807=>"000000000",
  26808=>"000101111",
  26809=>"011111111",
  26810=>"100000000",
  26811=>"100000001",
  26812=>"000000001",
  26813=>"000101111",
  26814=>"000000111",
  26815=>"001001000",
  26816=>"111111111",
  26817=>"101111111",
  26818=>"000111111",
  26819=>"111011111",
  26820=>"111111111",
  26821=>"000000000",
  26822=>"001001001",
  26823=>"000000000",
  26824=>"000110111",
  26825=>"111111111",
  26826=>"101000001",
  26827=>"011111111",
  26828=>"000000000",
  26829=>"110110111",
  26830=>"111000000",
  26831=>"111110100",
  26832=>"011111001",
  26833=>"000111111",
  26834=>"101101111",
  26835=>"000000000",
  26836=>"000000000",
  26837=>"011000100",
  26838=>"000000011",
  26839=>"100000111",
  26840=>"111110010",
  26841=>"111000000",
  26842=>"111111111",
  26843=>"111111110",
  26844=>"000100000",
  26845=>"000000000",
  26846=>"000011011",
  26847=>"000000000",
  26848=>"111000000",
  26849=>"000000000",
  26850=>"110110111",
  26851=>"100000000",
  26852=>"001000000",
  26853=>"000001101",
  26854=>"000000000",
  26855=>"000000001",
  26856=>"000000000",
  26857=>"100110010",
  26858=>"000000000",
  26859=>"001001111",
  26860=>"000000000",
  26861=>"011010011",
  26862=>"000110111",
  26863=>"000000000",
  26864=>"000000000",
  26865=>"000011011",
  26866=>"111111011",
  26867=>"000000001",
  26868=>"101001000",
  26869=>"111100100",
  26870=>"111111000",
  26871=>"011000000",
  26872=>"000000000",
  26873=>"000000110",
  26874=>"000000010",
  26875=>"011111000",
  26876=>"000000000",
  26877=>"001001001",
  26878=>"111111111",
  26879=>"000001000",
  26880=>"000000000",
  26881=>"001001001",
  26882=>"101101000",
  26883=>"000000100",
  26884=>"000000000",
  26885=>"111111111",
  26886=>"111111101",
  26887=>"100000010",
  26888=>"100000000",
  26889=>"000000111",
  26890=>"100111001",
  26891=>"111101111",
  26892=>"100000000",
  26893=>"100000000",
  26894=>"000000000",
  26895=>"000000101",
  26896=>"000000001",
  26897=>"111111100",
  26898=>"000000000",
  26899=>"111111001",
  26900=>"001000000",
  26901=>"110110111",
  26902=>"011001001",
  26903=>"001000111",
  26904=>"111111111",
  26905=>"111010000",
  26906=>"111111000",
  26907=>"000000000",
  26908=>"111111111",
  26909=>"110000000",
  26910=>"000000000",
  26911=>"111100000",
  26912=>"011011011",
  26913=>"000000100",
  26914=>"111111111",
  26915=>"001111111",
  26916=>"000100111",
  26917=>"000000001",
  26918=>"111111000",
  26919=>"000000000",
  26920=>"000000000",
  26921=>"111111000",
  26922=>"100100001",
  26923=>"011000001",
  26924=>"000000111",
  26925=>"100101001",
  26926=>"101110000",
  26927=>"000000001",
  26928=>"011010000",
  26929=>"110001000",
  26930=>"000000000",
  26931=>"011011010",
  26932=>"000001000",
  26933=>"010000110",
  26934=>"000000001",
  26935=>"101000000",
  26936=>"000000000",
  26937=>"000101111",
  26938=>"000000001",
  26939=>"111111110",
  26940=>"001000000",
  26941=>"000000000",
  26942=>"111111111",
  26943=>"100000000",
  26944=>"001000000",
  26945=>"111111000",
  26946=>"111100110",
  26947=>"101000000",
  26948=>"000000000",
  26949=>"000000000",
  26950=>"000000000",
  26951=>"000000000",
  26952=>"000000111",
  26953=>"000000100",
  26954=>"100000000",
  26955=>"001011011",
  26956=>"011111000",
  26957=>"111111000",
  26958=>"111111001",
  26959=>"000000000",
  26960=>"001101001",
  26961=>"111111111",
  26962=>"111111110",
  26963=>"000000101",
  26964=>"000000001",
  26965=>"011011011",
  26966=>"100000111",
  26967=>"000000010",
  26968=>"001001000",
  26969=>"111110111",
  26970=>"101000110",
  26971=>"000000001",
  26972=>"000010110",
  26973=>"000000010",
  26974=>"000000110",
  26975=>"111111010",
  26976=>"000000010",
  26977=>"011011011",
  26978=>"001000000",
  26979=>"001000001",
  26980=>"000000000",
  26981=>"000000000",
  26982=>"000000000",
  26983=>"000001010",
  26984=>"100110111",
  26985=>"000000001",
  26986=>"000000010",
  26987=>"000110100",
  26988=>"111111110",
  26989=>"001000000",
  26990=>"000000001",
  26991=>"111111001",
  26992=>"001000011",
  26993=>"000000100",
  26994=>"001000000",
  26995=>"100100100",
  26996=>"010111000",
  26997=>"110111100",
  26998=>"111000000",
  26999=>"110110110",
  27000=>"000000101",
  27001=>"111111111",
  27002=>"111111111",
  27003=>"000000001",
  27004=>"100110110",
  27005=>"001001011",
  27006=>"000000000",
  27007=>"000000000",
  27008=>"000101011",
  27009=>"001011011",
  27010=>"111111010",
  27011=>"000110100",
  27012=>"000000000",
  27013=>"011111111",
  27014=>"011011010",
  27015=>"111111111",
  27016=>"000000000",
  27017=>"111111111",
  27018=>"000001011",
  27019=>"011001000",
  27020=>"101001111",
  27021=>"111111110",
  27022=>"110000000",
  27023=>"111111111",
  27024=>"001000000",
  27025=>"000000000",
  27026=>"000100000",
  27027=>"100000000",
  27028=>"000001111",
  27029=>"000000000",
  27030=>"111111111",
  27031=>"101101000",
  27032=>"111000000",
  27033=>"000000111",
  27034=>"111111111",
  27035=>"111111100",
  27036=>"000000000",
  27037=>"111111110",
  27038=>"001001011",
  27039=>"011000000",
  27040=>"100011001",
  27041=>"011011001",
  27042=>"101101001",
  27043=>"000000000",
  27044=>"000000000",
  27045=>"011011000",
  27046=>"001111111",
  27047=>"010010000",
  27048=>"000000101",
  27049=>"011010110",
  27050=>"000000001",
  27051=>"000000000",
  27052=>"000000101",
  27053=>"111111111",
  27054=>"111111110",
  27055=>"111111001",
  27056=>"000011011",
  27057=>"000000000",
  27058=>"100110100",
  27059=>"000000000",
  27060=>"111111111",
  27061=>"011011001",
  27062=>"000101111",
  27063=>"111111011",
  27064=>"111011000",
  27065=>"111111111",
  27066=>"000010110",
  27067=>"000000000",
  27068=>"011111011",
  27069=>"111111000",
  27070=>"000000000",
  27071=>"001111111",
  27072=>"011011000",
  27073=>"110110010",
  27074=>"000010111",
  27075=>"111111110",
  27076=>"111111111",
  27077=>"110110110",
  27078=>"111111111",
  27079=>"111111111",
  27080=>"100000000",
  27081=>"101001000",
  27082=>"000000101",
  27083=>"000000000",
  27084=>"000000000",
  27085=>"000110000",
  27086=>"111100111",
  27087=>"110111111",
  27088=>"000000000",
  27089=>"101000100",
  27090=>"111010011",
  27091=>"111000000",
  27092=>"001011011",
  27093=>"000000000",
  27094=>"000001111",
  27095=>"111110110",
  27096=>"111111111",
  27097=>"000000001",
  27098=>"000000000",
  27099=>"111101111",
  27100=>"111111000",
  27101=>"110100000",
  27102=>"111111011",
  27103=>"000000100",
  27104=>"000000000",
  27105=>"001001111",
  27106=>"110110111",
  27107=>"000000000",
  27108=>"011000011",
  27109=>"000001111",
  27110=>"000000110",
  27111=>"110110000",
  27112=>"001101000",
  27113=>"111111100",
  27114=>"011011001",
  27115=>"111111110",
  27116=>"000001111",
  27117=>"000110110",
  27118=>"001001000",
  27119=>"000000000",
  27120=>"000000000",
  27121=>"111111111",
  27122=>"111111110",
  27123=>"000000111",
  27124=>"111000000",
  27125=>"000000000",
  27126=>"111111111",
  27127=>"000000000",
  27128=>"111111000",
  27129=>"000001001",
  27130=>"111000000",
  27131=>"111111111",
  27132=>"101111100",
  27133=>"000111111",
  27134=>"001111111",
  27135=>"111111111",
  27136=>"110110100",
  27137=>"000000100",
  27138=>"000000111",
  27139=>"111000111",
  27140=>"000000000",
  27141=>"000001111",
  27142=>"000001111",
  27143=>"100000100",
  27144=>"000000111",
  27145=>"111111000",
  27146=>"000000000",
  27147=>"000000010",
  27148=>"000000000",
  27149=>"111111111",
  27150=>"010000111",
  27151=>"111111111",
  27152=>"000000000",
  27153=>"000000000",
  27154=>"000000001",
  27155=>"000000000",
  27156=>"111111110",
  27157=>"001000100",
  27158=>"011111111",
  27159=>"011011000",
  27160=>"111111111",
  27161=>"101000000",
  27162=>"111110111",
  27163=>"000000111",
  27164=>"000000000",
  27165=>"000000000",
  27166=>"001000000",
  27167=>"111111111",
  27168=>"001000000",
  27169=>"111111011",
  27170=>"111101111",
  27171=>"011001111",
  27172=>"001000000",
  27173=>"000000000",
  27174=>"111111000",
  27175=>"000000100",
  27176=>"000000001",
  27177=>"000000000",
  27178=>"111111111",
  27179=>"000000000",
  27180=>"000101111",
  27181=>"111111001",
  27182=>"111011000",
  27183=>"111110100",
  27184=>"111111111",
  27185=>"000000000",
  27186=>"111001111",
  27187=>"001000000",
  27188=>"000010000",
  27189=>"111011011",
  27190=>"100000000",
  27191=>"000000000",
  27192=>"000000100",
  27193=>"101101000",
  27194=>"000000000",
  27195=>"000000000",
  27196=>"110000000",
  27197=>"001000001",
  27198=>"000000000",
  27199=>"111111001",
  27200=>"111111111",
  27201=>"000000000",
  27202=>"010111011",
  27203=>"110000000",
  27204=>"111111011",
  27205=>"111111111",
  27206=>"001000011",
  27207=>"111111111",
  27208=>"111111111",
  27209=>"000000111",
  27210=>"000000000",
  27211=>"111111111",
  27212=>"111011100",
  27213=>"000011111",
  27214=>"011000000",
  27215=>"000000000",
  27216=>"000000111",
  27217=>"110100000",
  27218=>"111111111",
  27219=>"001000000",
  27220=>"000000000",
  27221=>"000000001",
  27222=>"111111000",
  27223=>"111111100",
  27224=>"110000000",
  27225=>"110000000",
  27226=>"111010000",
  27227=>"010111111",
  27228=>"111111111",
  27229=>"111111111",
  27230=>"010000000",
  27231=>"111011001",
  27232=>"001001111",
  27233=>"000000000",
  27234=>"000000000",
  27235=>"001000100",
  27236=>"011001001",
  27237=>"111001111",
  27238=>"000011000",
  27239=>"110010000",
  27240=>"011111111",
  27241=>"100111111",
  27242=>"111011000",
  27243=>"001000000",
  27244=>"100000000",
  27245=>"000000000",
  27246=>"000110100",
  27247=>"000000000",
  27248=>"000001111",
  27249=>"111111111",
  27250=>"111000000",
  27251=>"111010000",
  27252=>"000000000",
  27253=>"111011111",
  27254=>"000000000",
  27255=>"011011111",
  27256=>"000001111",
  27257=>"100000000",
  27258=>"000000000",
  27259=>"111111111",
  27260=>"111111100",
  27261=>"010000000",
  27262=>"000000000",
  27263=>"000000000",
  27264=>"000000000",
  27265=>"110110110",
  27266=>"111010111",
  27267=>"000000000",
  27268=>"111111110",
  27269=>"000000000",
  27270=>"100110110",
  27271=>"011111111",
  27272=>"111110100",
  27273=>"111100001",
  27274=>"001000000",
  27275=>"000000000",
  27276=>"110000000",
  27277=>"011001000",
  27278=>"111111111",
  27279=>"111000000",
  27280=>"111111111",
  27281=>"111011111",
  27282=>"000000000",
  27283=>"111110111",
  27284=>"000000100",
  27285=>"000000001",
  27286=>"111111111",
  27287=>"111110100",
  27288=>"101111111",
  27289=>"111111111",
  27290=>"011001000",
  27291=>"000000000",
  27292=>"111111111",
  27293=>"100000001",
  27294=>"110000000",
  27295=>"000000010",
  27296=>"001000000",
  27297=>"111011101",
  27298=>"000000000",
  27299=>"111111111",
  27300=>"000000000",
  27301=>"110100101",
  27302=>"111111100",
  27303=>"000100100",
  27304=>"000111111",
  27305=>"000000100",
  27306=>"011000000",
  27307=>"000000000",
  27308=>"011011001",
  27309=>"111111111",
  27310=>"000000000",
  27311=>"000000111",
  27312=>"110111111",
  27313=>"111111001",
  27314=>"111111111",
  27315=>"111111001",
  27316=>"111111000",
  27317=>"111111000",
  27318=>"111101000",
  27319=>"000111111",
  27320=>"111111111",
  27321=>"111111111",
  27322=>"001000000",
  27323=>"100100000",
  27324=>"011111111",
  27325=>"111111100",
  27326=>"000000000",
  27327=>"000000000",
  27328=>"000000000",
  27329=>"000111111",
  27330=>"111111111",
  27331=>"000001000",
  27332=>"111111111",
  27333=>"111111111",
  27334=>"000000000",
  27335=>"000010111",
  27336=>"000000000",
  27337=>"111111111",
  27338=>"100110000",
  27339=>"110110000",
  27340=>"001111111",
  27341=>"111100001",
  27342=>"111011001",
  27343=>"011000000",
  27344=>"000000001",
  27345=>"000010000",
  27346=>"000000001",
  27347=>"000000000",
  27348=>"111111001",
  27349=>"110100100",
  27350=>"000001111",
  27351=>"001000001",
  27352=>"101111111",
  27353=>"111111111",
  27354=>"111000000",
  27355=>"000000000",
  27356=>"100000001",
  27357=>"110110111",
  27358=>"100111111",
  27359=>"000000000",
  27360=>"000000000",
  27361=>"000010111",
  27362=>"011111111",
  27363=>"111001111",
  27364=>"000000000",
  27365=>"111110100",
  27366=>"000000000",
  27367=>"111111111",
  27368=>"000000000",
  27369=>"100000101",
  27370=>"000000101",
  27371=>"110100000",
  27372=>"000011111",
  27373=>"000001001",
  27374=>"111110111",
  27375=>"000111111",
  27376=>"010000000",
  27377=>"111111111",
  27378=>"000000000",
  27379=>"000000000",
  27380=>"110111111",
  27381=>"101100100",
  27382=>"000000000",
  27383=>"000000000",
  27384=>"111111111",
  27385=>"000000000",
  27386=>"000000000",
  27387=>"000000001",
  27388=>"110110111",
  27389=>"000000000",
  27390=>"111110100",
  27391=>"000011011",
  27392=>"000000000",
  27393=>"111111111",
  27394=>"000000000",
  27395=>"000000001",
  27396=>"100000110",
  27397=>"000000000",
  27398=>"100100111",
  27399=>"100000001",
  27400=>"111111111",
  27401=>"000000010",
  27402=>"000111111",
  27403=>"111111111",
  27404=>"101101000",
  27405=>"000001111",
  27406=>"000000000",
  27407=>"010010000",
  27408=>"000000000",
  27409=>"000000001",
  27410=>"111000000",
  27411=>"101000001",
  27412=>"000000000",
  27413=>"111111111",
  27414=>"000101111",
  27415=>"100101111",
  27416=>"111111111",
  27417=>"000000111",
  27418=>"001001000",
  27419=>"000000000",
  27420=>"001111111",
  27421=>"000000000",
  27422=>"000010000",
  27423=>"111111111",
  27424=>"111000000",
  27425=>"001001111",
  27426=>"000000000",
  27427=>"111111111",
  27428=>"111111111",
  27429=>"000000000",
  27430=>"110110000",
  27431=>"000000110",
  27432=>"000000000",
  27433=>"011011011",
  27434=>"111100000",
  27435=>"111111100",
  27436=>"111111111",
  27437=>"101111001",
  27438=>"101110011",
  27439=>"001000000",
  27440=>"000000000",
  27441=>"000000000",
  27442=>"101000100",
  27443=>"111001111",
  27444=>"000000110",
  27445=>"111011010",
  27446=>"111111111",
  27447=>"111110100",
  27448=>"000000000",
  27449=>"111101100",
  27450=>"000100111",
  27451=>"000000000",
  27452=>"111111111",
  27453=>"000010110",
  27454=>"111111111",
  27455=>"010000110",
  27456=>"000000100",
  27457=>"000000000",
  27458=>"000000000",
  27459=>"000101111",
  27460=>"110100111",
  27461=>"011111111",
  27462=>"000001001",
  27463=>"000000000",
  27464=>"111000000",
  27465=>"000000111",
  27466=>"001000000",
  27467=>"111111111",
  27468=>"000000100",
  27469=>"111111010",
  27470=>"100100111",
  27471=>"101111111",
  27472=>"100101111",
  27473=>"000000000",
  27474=>"111110111",
  27475=>"000000100",
  27476=>"000010010",
  27477=>"001001001",
  27478=>"111111111",
  27479=>"110000000",
  27480=>"000000000",
  27481=>"000101111",
  27482=>"000000110",
  27483=>"111100100",
  27484=>"000000100",
  27485=>"111011111",
  27486=>"111111111",
  27487=>"111111111",
  27488=>"111110111",
  27489=>"000000000",
  27490=>"100100001",
  27491=>"000000000",
  27492=>"011111111",
  27493=>"000000000",
  27494=>"000000000",
  27495=>"001101111",
  27496=>"111111111",
  27497=>"111111111",
  27498=>"111111111",
  27499=>"111111111",
  27500=>"000001101",
  27501=>"000000011",
  27502=>"010011010",
  27503=>"111111111",
  27504=>"111111111",
  27505=>"000000010",
  27506=>"000000000",
  27507=>"111111111",
  27508=>"010000000",
  27509=>"111111111",
  27510=>"000001111",
  27511=>"100100000",
  27512=>"111000001",
  27513=>"111111111",
  27514=>"111111111",
  27515=>"110110111",
  27516=>"001001011",
  27517=>"111100111",
  27518=>"111011001",
  27519=>"000000000",
  27520=>"101100100",
  27521=>"000111111",
  27522=>"111111111",
  27523=>"111111000",
  27524=>"010011111",
  27525=>"010000000",
  27526=>"001000000",
  27527=>"111111111",
  27528=>"001001111",
  27529=>"111110010",
  27530=>"111111111",
  27531=>"111111100",
  27532=>"111111111",
  27533=>"111111110",
  27534=>"000000000",
  27535=>"000000100",
  27536=>"000000001",
  27537=>"000101111",
  27538=>"000000011",
  27539=>"111111111",
  27540=>"000000100",
  27541=>"000000000",
  27542=>"111111111",
  27543=>"001000000",
  27544=>"010111111",
  27545=>"000000001",
  27546=>"111111111",
  27547=>"000000000",
  27548=>"111110110",
  27549=>"111000000",
  27550=>"000000001",
  27551=>"000000000",
  27552=>"001001111",
  27553=>"111000100",
  27554=>"110111100",
  27555=>"000000011",
  27556=>"100100100",
  27557=>"000010010",
  27558=>"110111010",
  27559=>"000000000",
  27560=>"000000010",
  27561=>"111111111",
  27562=>"111110110",
  27563=>"111101111",
  27564=>"000000000",
  27565=>"101100000",
  27566=>"111111111",
  27567=>"000000000",
  27568=>"111111111",
  27569=>"000000000",
  27570=>"000000001",
  27571=>"011101111",
  27572=>"000000000",
  27573=>"000000000",
  27574=>"111111111",
  27575=>"111111111",
  27576=>"000000110",
  27577=>"000000000",
  27578=>"000000000",
  27579=>"111000100",
  27580=>"100111111",
  27581=>"101111111",
  27582=>"000000100",
  27583=>"101111111",
  27584=>"111111110",
  27585=>"011011011",
  27586=>"000000001",
  27587=>"111111111",
  27588=>"000000000",
  27589=>"111001001",
  27590=>"100000000",
  27591=>"000110110",
  27592=>"001001001",
  27593=>"000000000",
  27594=>"101000000",
  27595=>"010110100",
  27596=>"000000000",
  27597=>"111111111",
  27598=>"101000100",
  27599=>"110111111",
  27600=>"111111111",
  27601=>"111111111",
  27602=>"000000000",
  27603=>"000000100",
  27604=>"110100110",
  27605=>"000001001",
  27606=>"111111111",
  27607=>"001001000",
  27608=>"001001000",
  27609=>"000001000",
  27610=>"011110011",
  27611=>"111111000",
  27612=>"010011111",
  27613=>"111000001",
  27614=>"111111100",
  27615=>"100000001",
  27616=>"000000000",
  27617=>"000000110",
  27618=>"111111111",
  27619=>"011111101",
  27620=>"111111111",
  27621=>"000000000",
  27622=>"011001000",
  27623=>"111011011",
  27624=>"100000000",
  27625=>"001111111",
  27626=>"100001110",
  27627=>"111111111",
  27628=>"111010111",
  27629=>"000100000",
  27630=>"111111111",
  27631=>"000000010",
  27632=>"000000000",
  27633=>"000100110",
  27634=>"000000000",
  27635=>"111000000",
  27636=>"001000000",
  27637=>"111111101",
  27638=>"000000100",
  27639=>"000000000",
  27640=>"111110100",
  27641=>"001100000",
  27642=>"000111111",
  27643=>"000110110",
  27644=>"011111111",
  27645=>"000000111",
  27646=>"000000000",
  27647=>"111111111",
  27648=>"111111111",
  27649=>"110110000",
  27650=>"111111111",
  27651=>"000100111",
  27652=>"110100111",
  27653=>"111000101",
  27654=>"010000000",
  27655=>"000000111",
  27656=>"000111111",
  27657=>"010111110",
  27658=>"111111111",
  27659=>"111111000",
  27660=>"100110110",
  27661=>"110100111",
  27662=>"000100000",
  27663=>"000000000",
  27664=>"000100000",
  27665=>"000000100",
  27666=>"000010111",
  27667=>"111110000",
  27668=>"000000111",
  27669=>"000111111",
  27670=>"111111111",
  27671=>"011100100",
  27672=>"001001111",
  27673=>"000000011",
  27674=>"001000001",
  27675=>"000000110",
  27676=>"100000110",
  27677=>"110000000",
  27678=>"111111111",
  27679=>"111111000",
  27680=>"101101000",
  27681=>"111111101",
  27682=>"111011111",
  27683=>"010111100",
  27684=>"111111110",
  27685=>"111111111",
  27686=>"000000000",
  27687=>"000101111",
  27688=>"000001101",
  27689=>"000000000",
  27690=>"111111111",
  27691=>"000000001",
  27692=>"000000111",
  27693=>"001111111",
  27694=>"001001001",
  27695=>"000000000",
  27696=>"000000000",
  27697=>"000000000",
  27698=>"000000000",
  27699=>"000000111",
  27700=>"111100000",
  27701=>"001000000",
  27702=>"101000111",
  27703=>"100001111",
  27704=>"111000000",
  27705=>"010010111",
  27706=>"111111111",
  27707=>"111111111",
  27708=>"111100000",
  27709=>"100111111",
  27710=>"110111100",
  27711=>"000000111",
  27712=>"001000000",
  27713=>"000110111",
  27714=>"111111111",
  27715=>"000001000",
  27716=>"000100110",
  27717=>"111111100",
  27718=>"000000111",
  27719=>"000000000",
  27720=>"111111111",
  27721=>"111000010",
  27722=>"111110111",
  27723=>"000000000",
  27724=>"111111111",
  27725=>"000001000",
  27726=>"111000001",
  27727=>"000000000",
  27728=>"000000000",
  27729=>"010000110",
  27730=>"000111111",
  27731=>"011111110",
  27732=>"101000000",
  27733=>"000000100",
  27734=>"000001100",
  27735=>"000001001",
  27736=>"000000000",
  27737=>"001000111",
  27738=>"001000110",
  27739=>"001001001",
  27740=>"000000000",
  27741=>"000000111",
  27742=>"000101100",
  27743=>"110110000",
  27744=>"111111111",
  27745=>"011111011",
  27746=>"000011111",
  27747=>"000000000",
  27748=>"000000000",
  27749=>"000000001",
  27750=>"001000000",
  27751=>"000000000",
  27752=>"001011000",
  27753=>"111011011",
  27754=>"000000111",
  27755=>"000000000",
  27756=>"111111100",
  27757=>"000000000",
  27758=>"111000110",
  27759=>"111010000",
  27760=>"111111011",
  27761=>"000000001",
  27762=>"000000011",
  27763=>"111011101",
  27764=>"101000000",
  27765=>"011111111",
  27766=>"011111111",
  27767=>"111111000",
  27768=>"000000000",
  27769=>"101100100",
  27770=>"001011000",
  27771=>"000000000",
  27772=>"100111100",
  27773=>"111000000",
  27774=>"110111101",
  27775=>"000000000",
  27776=>"000000000",
  27777=>"001001111",
  27778=>"111000000",
  27779=>"000001000",
  27780=>"000000111",
  27781=>"111100111",
  27782=>"111111111",
  27783=>"111111111",
  27784=>"110111111",
  27785=>"000000111",
  27786=>"111111000",
  27787=>"000001000",
  27788=>"100000100",
  27789=>"001000000",
  27790=>"101001110",
  27791=>"010111011",
  27792=>"101111011",
  27793=>"000000000",
  27794=>"000111111",
  27795=>"000000101",
  27796=>"000000011",
  27797=>"110111111",
  27798=>"110111111",
  27799=>"000000000",
  27800=>"000000000",
  27801=>"000000100",
  27802=>"011000000",
  27803=>"100000011",
  27804=>"000000000",
  27805=>"010100100",
  27806=>"100000000",
  27807=>"000111111",
  27808=>"001000000",
  27809=>"101001001",
  27810=>"111111101",
  27811=>"111111111",
  27812=>"000100000",
  27813=>"100000000",
  27814=>"100000000",
  27815=>"111111110",
  27816=>"111111111",
  27817=>"111000000",
  27818=>"111000000",
  27819=>"111011001",
  27820=>"111111000",
  27821=>"000000001",
  27822=>"100101100",
  27823=>"000000000",
  27824=>"111111000",
  27825=>"111111000",
  27826=>"111111111",
  27827=>"000000100",
  27828=>"111111100",
  27829=>"111111111",
  27830=>"000000000",
  27831=>"000111111",
  27832=>"100000110",
  27833=>"010000000",
  27834=>"001000110",
  27835=>"111111001",
  27836=>"001001000",
  27837=>"100101111",
  27838=>"010111110",
  27839=>"000111111",
  27840=>"000000111",
  27841=>"111110111",
  27842=>"011001101",
  27843=>"000111111",
  27844=>"111111111",
  27845=>"000000101",
  27846=>"000000000",
  27847=>"111111111",
  27848=>"000000000",
  27849=>"000000000",
  27850=>"000000000",
  27851=>"000000011",
  27852=>"111111111",
  27853=>"000001101",
  27854=>"100110100",
  27855=>"000111111",
  27856=>"111000001",
  27857=>"000000000",
  27858=>"000000100",
  27859=>"000000000",
  27860=>"111000111",
  27861=>"111111111",
  27862=>"000000111",
  27863=>"000100111",
  27864=>"000000111",
  27865=>"100111111",
  27866=>"111100000",
  27867=>"000110111",
  27868=>"111111111",
  27869=>"111110000",
  27870=>"000000000",
  27871=>"000000111",
  27872=>"111011111",
  27873=>"000010000",
  27874=>"000000000",
  27875=>"111001111",
  27876=>"000000000",
  27877=>"100100000",
  27878=>"000000000",
  27879=>"111111111",
  27880=>"000111111",
  27881=>"111111111",
  27882=>"000000101",
  27883=>"000111111",
  27884=>"101111111",
  27885=>"000111111",
  27886=>"110110000",
  27887=>"110000000",
  27888=>"000001001",
  27889=>"000000000",
  27890=>"000111011",
  27891=>"000000001",
  27892=>"111111111",
  27893=>"111111111",
  27894=>"000000100",
  27895=>"111111111",
  27896=>"000001000",
  27897=>"111111111",
  27898=>"100000100",
  27899=>"111111111",
  27900=>"011011000",
  27901=>"111001101",
  27902=>"111000000",
  27903=>"111111111",
  27904=>"111111111",
  27905=>"100000000",
  27906=>"101101001",
  27907=>"000000000",
  27908=>"111111111",
  27909=>"111111111",
  27910=>"111111101",
  27911=>"100110111",
  27912=>"110110000",
  27913=>"111000000",
  27914=>"111111111",
  27915=>"000100100",
  27916=>"001000000",
  27917=>"111001000",
  27918=>"111111101",
  27919=>"000000111",
  27920=>"000000000",
  27921=>"101000000",
  27922=>"111100111",
  27923=>"111111111",
  27924=>"111111011",
  27925=>"000000111",
  27926=>"111111111",
  27927=>"101100000",
  27928=>"001000000",
  27929=>"000000000",
  27930=>"111111000",
  27931=>"111111111",
  27932=>"000100001",
  27933=>"000000111",
  27934=>"000000000",
  27935=>"111111111",
  27936=>"100100000",
  27937=>"100111101",
  27938=>"000000001",
  27939=>"111111111",
  27940=>"101111111",
  27941=>"000000011",
  27942=>"111111111",
  27943=>"000000111",
  27944=>"011110110",
  27945=>"000000000",
  27946=>"001101101",
  27947=>"011011111",
  27948=>"000000000",
  27949=>"111111011",
  27950=>"000111100",
  27951=>"000100000",
  27952=>"000000000",
  27953=>"111111111",
  27954=>"111000001",
  27955=>"000111111",
  27956=>"001000111",
  27957=>"000101111",
  27958=>"000000011",
  27959=>"000111111",
  27960=>"000000110",
  27961=>"001001111",
  27962=>"011111111",
  27963=>"000111111",
  27964=>"000000000",
  27965=>"111111000",
  27966=>"010000000",
  27967=>"000000000",
  27968=>"000000000",
  27969=>"101000000",
  27970=>"000001101",
  27971=>"011000000",
  27972=>"000001100",
  27973=>"100010110",
  27974=>"000000000",
  27975=>"000000000",
  27976=>"000000000",
  27977=>"000000000",
  27978=>"111101000",
  27979=>"100100000",
  27980=>"000000101",
  27981=>"001001000",
  27982=>"110111111",
  27983=>"001000000",
  27984=>"011011000",
  27985=>"000000000",
  27986=>"111111011",
  27987=>"000000000",
  27988=>"110111111",
  27989=>"011011011",
  27990=>"111111000",
  27991=>"111000000",
  27992=>"000000001",
  27993=>"111111111",
  27994=>"001000000",
  27995=>"000000000",
  27996=>"000100111",
  27997=>"111111111",
  27998=>"000000000",
  27999=>"000000000",
  28000=>"000000101",
  28001=>"111111111",
  28002=>"111110111",
  28003=>"000000100",
  28004=>"110110111",
  28005=>"001000000",
  28006=>"000110111",
  28007=>"110101111",
  28008=>"010111001",
  28009=>"111111111",
  28010=>"000000000",
  28011=>"110100110",
  28012=>"000000000",
  28013=>"000111111",
  28014=>"000000000",
  28015=>"011000000",
  28016=>"111110000",
  28017=>"110000000",
  28018=>"001000000",
  28019=>"011000000",
  28020=>"000111111",
  28021=>"100100100",
  28022=>"110000100",
  28023=>"100111000",
  28024=>"001000000",
  28025=>"000000111",
  28026=>"110000001",
  28027=>"000000000",
  28028=>"111001000",
  28029=>"000000000",
  28030=>"111111000",
  28031=>"000000000",
  28032=>"000000000",
  28033=>"000000110",
  28034=>"111111000",
  28035=>"111111111",
  28036=>"111010111",
  28037=>"000001000",
  28038=>"000000101",
  28039=>"000000100",
  28040=>"010000111",
  28041=>"111111111",
  28042=>"000000000",
  28043=>"111111000",
  28044=>"101111111",
  28045=>"001101001",
  28046=>"000000000",
  28047=>"000001000",
  28048=>"000000000",
  28049=>"100000000",
  28050=>"000100111",
  28051=>"000000000",
  28052=>"011001011",
  28053=>"010111000",
  28054=>"000000001",
  28055=>"000000000",
  28056=>"001111111",
  28057=>"110111000",
  28058=>"100111110",
  28059=>"000000111",
  28060=>"111111111",
  28061=>"000000111",
  28062=>"000000000",
  28063=>"001001000",
  28064=>"000111111",
  28065=>"100000000",
  28066=>"111111111",
  28067=>"010111111",
  28068=>"110111101",
  28069=>"001011010",
  28070=>"111111111",
  28071=>"111111111",
  28072=>"110110100",
  28073=>"101000000",
  28074=>"000001011",
  28075=>"100000000",
  28076=>"001000000",
  28077=>"000000000",
  28078=>"000110111",
  28079=>"000000000",
  28080=>"100111111",
  28081=>"111111111",
  28082=>"000000001",
  28083=>"111111111",
  28084=>"011001001",
  28085=>"011001001",
  28086=>"111111011",
  28087=>"111111001",
  28088=>"000000111",
  28089=>"011001000",
  28090=>"111111111",
  28091=>"001000101",
  28092=>"100111111",
  28093=>"000000000",
  28094=>"000000000",
  28095=>"100111110",
  28096=>"111111000",
  28097=>"111011111",
  28098=>"111111111",
  28099=>"000000111",
  28100=>"000101111",
  28101=>"000100110",
  28102=>"011111000",
  28103=>"011011001",
  28104=>"111111110",
  28105=>"000000000",
  28106=>"100000000",
  28107=>"000000000",
  28108=>"000000111",
  28109=>"000001000",
  28110=>"111000000",
  28111=>"111111111",
  28112=>"011000000",
  28113=>"111111111",
  28114=>"000000011",
  28115=>"111001010",
  28116=>"010111111",
  28117=>"111111111",
  28118=>"000000000",
  28119=>"011011011",
  28120=>"000101111",
  28121=>"100000000",
  28122=>"111111111",
  28123=>"001000000",
  28124=>"100111111",
  28125=>"111001001",
  28126=>"000000100",
  28127=>"001001000",
  28128=>"000000000",
  28129=>"000000000",
  28130=>"001111000",
  28131=>"000000010",
  28132=>"000011111",
  28133=>"101111011",
  28134=>"000000000",
  28135=>"000000111",
  28136=>"000000000",
  28137=>"000000000",
  28138=>"000000111",
  28139=>"110110100",
  28140=>"111111011",
  28141=>"001000100",
  28142=>"000000001",
  28143=>"000000101",
  28144=>"000000000",
  28145=>"000000000",
  28146=>"111100000",
  28147=>"000000000",
  28148=>"001101111",
  28149=>"000000000",
  28150=>"111111111",
  28151=>"110111111",
  28152=>"111111111",
  28153=>"000100100",
  28154=>"110100101",
  28155=>"011011111",
  28156=>"000000000",
  28157=>"100101111",
  28158=>"111000000",
  28159=>"000100000",
  28160=>"100010111",
  28161=>"000000000",
  28162=>"011111111",
  28163=>"000101011",
  28164=>"111111111",
  28165=>"001001110",
  28166=>"000000010",
  28167=>"000101001",
  28168=>"111110000",
  28169=>"000100100",
  28170=>"111111111",
  28171=>"100100100",
  28172=>"100110000",
  28173=>"000000100",
  28174=>"000001001",
  28175=>"111111111",
  28176=>"111101111",
  28177=>"100000000",
  28178=>"111101111",
  28179=>"000011011",
  28180=>"001101111",
  28181=>"111111111",
  28182=>"110111111",
  28183=>"111111001",
  28184=>"111101100",
  28185=>"000110011",
  28186=>"000011111",
  28187=>"000000001",
  28188=>"000000000",
  28189=>"111111000",
  28190=>"111011011",
  28191=>"100000000",
  28192=>"000000000",
  28193=>"001001001",
  28194=>"001001111",
  28195=>"000000000",
  28196=>"000000000",
  28197=>"111111111",
  28198=>"000100110",
  28199=>"110110111",
  28200=>"100110111",
  28201=>"011111111",
  28202=>"000000011",
  28203=>"111111111",
  28204=>"111111111",
  28205=>"111001000",
  28206=>"100000111",
  28207=>"000000011",
  28208=>"000011011",
  28209=>"010011000",
  28210=>"110110110",
  28211=>"100100011",
  28212=>"011011011",
  28213=>"000000110",
  28214=>"000001111",
  28215=>"111111111",
  28216=>"000000111",
  28217=>"111101001",
  28218=>"110111111",
  28219=>"111111111",
  28220=>"100000000",
  28221=>"111111111",
  28222=>"000000000",
  28223=>"000000000",
  28224=>"111001000",
  28225=>"000110000",
  28226=>"011000000",
  28227=>"100111111",
  28228=>"111111111",
  28229=>"111111111",
  28230=>"001000000",
  28231=>"000000000",
  28232=>"111000000",
  28233=>"000000111",
  28234=>"111111111",
  28235=>"000000000",
  28236=>"111111111",
  28237=>"101000000",
  28238=>"101001110",
  28239=>"100000001",
  28240=>"100111011",
  28241=>"001101111",
  28242=>"000000000",
  28243=>"000000100",
  28244=>"000000000",
  28245=>"011111111",
  28246=>"111111110",
  28247=>"001000101",
  28248=>"000011111",
  28249=>"001001000",
  28250=>"101111111",
  28251=>"000000000",
  28252=>"000000000",
  28253=>"111111111",
  28254=>"101100100",
  28255=>"011001001",
  28256=>"000000010",
  28257=>"101111111",
  28258=>"110110101",
  28259=>"000000000",
  28260=>"011111111",
  28261=>"110100110",
  28262=>"000000000",
  28263=>"000000000",
  28264=>"000111000",
  28265=>"011000000",
  28266=>"000010110",
  28267=>"000110111",
  28268=>"000000000",
  28269=>"001111111",
  28270=>"111110100",
  28271=>"000000100",
  28272=>"101101111",
  28273=>"000011111",
  28274=>"000011111",
  28275=>"000000101",
  28276=>"000000000",
  28277=>"111111000",
  28278=>"001011000",
  28279=>"000000000",
  28280=>"000000000",
  28281=>"000111111",
  28282=>"011110100",
  28283=>"000000100",
  28284=>"110111111",
  28285=>"111111111",
  28286=>"110111100",
  28287=>"111111111",
  28288=>"111111111",
  28289=>"101000000",
  28290=>"111110110",
  28291=>"000001000",
  28292=>"111111011",
  28293=>"000000000",
  28294=>"000011011",
  28295=>"000000100",
  28296=>"100000110",
  28297=>"111111111",
  28298=>"000010000",
  28299=>"100100000",
  28300=>"000111111",
  28301=>"000010000",
  28302=>"000100111",
  28303=>"000000000",
  28304=>"001001001",
  28305=>"111111000",
  28306=>"111111101",
  28307=>"000010000",
  28308=>"111011000",
  28309=>"111000000",
  28310=>"000000111",
  28311=>"000000000",
  28312=>"000000000",
  28313=>"111111111",
  28314=>"000000101",
  28315=>"111111110",
  28316=>"001111111",
  28317=>"111111110",
  28318=>"000011111",
  28319=>"000000000",
  28320=>"110110111",
  28321=>"100000000",
  28322=>"000011000",
  28323=>"111111111",
  28324=>"000100110",
  28325=>"000000000",
  28326=>"111101111",
  28327=>"110110111",
  28328=>"000101111",
  28329=>"000000000",
  28330=>"001111111",
  28331=>"101000000",
  28332=>"111011111",
  28333=>"100001000",
  28334=>"000001011",
  28335=>"111111111",
  28336=>"000000000",
  28337=>"100111000",
  28338=>"101001010",
  28339=>"010000000",
  28340=>"111000001",
  28341=>"001000100",
  28342=>"111001001",
  28343=>"000000000",
  28344=>"001011110",
  28345=>"000001111",
  28346=>"011111000",
  28347=>"101100000",
  28348=>"001001101",
  28349=>"111111110",
  28350=>"111111000",
  28351=>"110010000",
  28352=>"000000000",
  28353=>"000000000",
  28354=>"111011011",
  28355=>"000000000",
  28356=>"001100111",
  28357=>"111111001",
  28358=>"011010111",
  28359=>"100001111",
  28360=>"110110111",
  28361=>"000111011",
  28362=>"000000000",
  28363=>"011000000",
  28364=>"111110110",
  28365=>"100111111",
  28366=>"101111111",
  28367=>"110000000",
  28368=>"111110000",
  28369=>"111011011",
  28370=>"111000000",
  28371=>"011111111",
  28372=>"111001101",
  28373=>"000000000",
  28374=>"111001000",
  28375=>"000111111",
  28376=>"011111110",
  28377=>"010111111",
  28378=>"111111111",
  28379=>"111001001",
  28380=>"111111111",
  28381=>"100100100",
  28382=>"000000100",
  28383=>"000000101",
  28384=>"000111011",
  28385=>"011011011",
  28386=>"111111111",
  28387=>"111000000",
  28388=>"111111101",
  28389=>"000010011",
  28390=>"000000000",
  28391=>"111111000",
  28392=>"000000000",
  28393=>"000000000",
  28394=>"111111111",
  28395=>"100101111",
  28396=>"000000000",
  28397=>"111011101",
  28398=>"000000101",
  28399=>"111011000",
  28400=>"011010110",
  28401=>"111000100",
  28402=>"111111111",
  28403=>"000000111",
  28404=>"111111001",
  28405=>"110001001",
  28406=>"110100000",
  28407=>"111011010",
  28408=>"000010000",
  28409=>"000000000",
  28410=>"001111010",
  28411=>"111011000",
  28412=>"101101011",
  28413=>"001001001",
  28414=>"101101100",
  28415=>"100100100",
  28416=>"101100000",
  28417=>"001011011",
  28418=>"111111111",
  28419=>"001000000",
  28420=>"111111111",
  28421=>"000010000",
  28422=>"000000111",
  28423=>"000011100",
  28424=>"111111110",
  28425=>"000000000",
  28426=>"000000000",
  28427=>"100110110",
  28428=>"000001111",
  28429=>"000000000",
  28430=>"000000000",
  28431=>"111111100",
  28432=>"001000000",
  28433=>"100000111",
  28434=>"101111111",
  28435=>"000111001",
  28436=>"000001001",
  28437=>"000000000",
  28438=>"111011111",
  28439=>"100100000",
  28440=>"111111111",
  28441=>"000000100",
  28442=>"111111111",
  28443=>"111100101",
  28444=>"100111111",
  28445=>"001011011",
  28446=>"000000100",
  28447=>"111000101",
  28448=>"100100101",
  28449=>"111000000",
  28450=>"000000001",
  28451=>"000000000",
  28452=>"011000000",
  28453=>"111111110",
  28454=>"001001001",
  28455=>"011011111",
  28456=>"110101111",
  28457=>"001000001",
  28458=>"101000010",
  28459=>"000000101",
  28460=>"101100100",
  28461=>"001011011",
  28462=>"000001000",
  28463=>"000110010",
  28464=>"000011000",
  28465=>"111111111",
  28466=>"111101101",
  28467=>"011010000",
  28468=>"000000000",
  28469=>"111100111",
  28470=>"110000000",
  28471=>"000000000",
  28472=>"111111011",
  28473=>"000000000",
  28474=>"011011100",
  28475=>"110111111",
  28476=>"001001011",
  28477=>"000001011",
  28478=>"000000000",
  28479=>"000000000",
  28480=>"001111001",
  28481=>"000001001",
  28482=>"101111000",
  28483=>"000110111",
  28484=>"000000000",
  28485=>"000111111",
  28486=>"100111111",
  28487=>"110110111",
  28488=>"000000000",
  28489=>"110000000",
  28490=>"000000000",
  28491=>"011000001",
  28492=>"001100101",
  28493=>"100110010",
  28494=>"101110100",
  28495=>"010110110",
  28496=>"000000110",
  28497=>"111111110",
  28498=>"010110111",
  28499=>"000011011",
  28500=>"000000000",
  28501=>"011011001",
  28502=>"111001011",
  28503=>"100000011",
  28504=>"000000000",
  28505=>"001001011",
  28506=>"101111011",
  28507=>"110110111",
  28508=>"000000000",
  28509=>"111101100",
  28510=>"111111111",
  28511=>"000000000",
  28512=>"000000000",
  28513=>"111111111",
  28514=>"111110110",
  28515=>"000000000",
  28516=>"011111111",
  28517=>"000000100",
  28518=>"111111111",
  28519=>"000101001",
  28520=>"110110111",
  28521=>"011110101",
  28522=>"000011000",
  28523=>"111100111",
  28524=>"100110110",
  28525=>"000011001",
  28526=>"000000000",
  28527=>"000000000",
  28528=>"111111111",
  28529=>"011000001",
  28530=>"000000000",
  28531=>"111000001",
  28532=>"000000110",
  28533=>"111110111",
  28534=>"101100000",
  28535=>"000100000",
  28536=>"000000000",
  28537=>"000000110",
  28538=>"111101111",
  28539=>"110000000",
  28540=>"001011000",
  28541=>"000000000",
  28542=>"111100000",
  28543=>"100100110",
  28544=>"000110111",
  28545=>"101101111",
  28546=>"111111111",
  28547=>"000000000",
  28548=>"000111111",
  28549=>"010010111",
  28550=>"111011001",
  28551=>"111000001",
  28552=>"101101101",
  28553=>"000110011",
  28554=>"000000000",
  28555=>"111111111",
  28556=>"000101111",
  28557=>"100100100",
  28558=>"100101111",
  28559=>"000000000",
  28560=>"000010000",
  28561=>"110100110",
  28562=>"110111011",
  28563=>"110110111",
  28564=>"011000000",
  28565=>"000000000",
  28566=>"111111000",
  28567=>"001011111",
  28568=>"111111111",
  28569=>"111100100",
  28570=>"100100000",
  28571=>"000000100",
  28572=>"100111111",
  28573=>"000001001",
  28574=>"111011010",
  28575=>"100111111",
  28576=>"111000000",
  28577=>"000000000",
  28578=>"111011111",
  28579=>"000000000",
  28580=>"000001101",
  28581=>"000000000",
  28582=>"001000000",
  28583=>"111001111",
  28584=>"000000110",
  28585=>"111111111",
  28586=>"111111000",
  28587=>"000000011",
  28588=>"000000100",
  28589=>"000000000",
  28590=>"000111000",
  28591=>"010000000",
  28592=>"011011011",
  28593=>"111011110",
  28594=>"010010110",
  28595=>"000000000",
  28596=>"111111111",
  28597=>"111011111",
  28598=>"110111100",
  28599=>"111000000",
  28600=>"000000111",
  28601=>"111101001",
  28602=>"110100100",
  28603=>"001000000",
  28604=>"000000001",
  28605=>"000000000",
  28606=>"000000001",
  28607=>"111000001",
  28608=>"000111111",
  28609=>"101111111",
  28610=>"001000000",
  28611=>"110111001",
  28612=>"000000000",
  28613=>"000000000",
  28614=>"000000110",
  28615=>"110010000",
  28616=>"000100100",
  28617=>"000010000",
  28618=>"000110100",
  28619=>"101111111",
  28620=>"000000000",
  28621=>"111111110",
  28622=>"111100000",
  28623=>"000000111",
  28624=>"000110001",
  28625=>"101111111",
  28626=>"000000110",
  28627=>"000000000",
  28628=>"000000000",
  28629=>"111001000",
  28630=>"110100111",
  28631=>"110111000",
  28632=>"001001000",
  28633=>"000000111",
  28634=>"011110000",
  28635=>"001000000",
  28636=>"010011000",
  28637=>"100011111",
  28638=>"010010000",
  28639=>"000111111",
  28640=>"111111111",
  28641=>"111100100",
  28642=>"000000000",
  28643=>"000000000",
  28644=>"000000111",
  28645=>"000001000",
  28646=>"100001111",
  28647=>"111111111",
  28648=>"111101111",
  28649=>"101101111",
  28650=>"010000000",
  28651=>"111111111",
  28652=>"011000000",
  28653=>"100100011",
  28654=>"011001001",
  28655=>"000000100",
  28656=>"111000000",
  28657=>"110111111",
  28658=>"111111111",
  28659=>"111001011",
  28660=>"101000111",
  28661=>"000110110",
  28662=>"100101101",
  28663=>"101000000",
  28664=>"111111000",
  28665=>"000100101",
  28666=>"111010000",
  28667=>"111011101",
  28668=>"101011011",
  28669=>"000000100",
  28670=>"000000100",
  28671=>"011100111",
  28672=>"000010011",
  28673=>"000000000",
  28674=>"001001111",
  28675=>"000000101",
  28676=>"100000001",
  28677=>"000000000",
  28678=>"000000000",
  28679=>"111111000",
  28680=>"100100001",
  28681=>"111100011",
  28682=>"001000000",
  28683=>"000011011",
  28684=>"001001001",
  28685=>"000000000",
  28686=>"000000100",
  28687=>"010010010",
  28688=>"000010110",
  28689=>"000000000",
  28690=>"000111111",
  28691=>"111101000",
  28692=>"000000000",
  28693=>"010001111",
  28694=>"001001101",
  28695=>"111111110",
  28696=>"011000110",
  28697=>"000001000",
  28698=>"000000000",
  28699=>"000111010",
  28700=>"110110000",
  28701=>"011000000",
  28702=>"000000111",
  28703=>"111110110",
  28704=>"010011000",
  28705=>"100100110",
  28706=>"000000110",
  28707=>"011001001",
  28708=>"000000000",
  28709=>"000001011",
  28710=>"001011000",
  28711=>"010110110",
  28712=>"111010000",
  28713=>"000000000",
  28714=>"110111000",
  28715=>"111110010",
  28716=>"001001001",
  28717=>"111001011",
  28718=>"000000001",
  28719=>"000000010",
  28720=>"001001111",
  28721=>"101101111",
  28722=>"011001000",
  28723=>"100111111",
  28724=>"100111111",
  28725=>"011111101",
  28726=>"000000000",
  28727=>"111000100",
  28728=>"001101111",
  28729=>"000000010",
  28730=>"000000000",
  28731=>"101111111",
  28732=>"101100000",
  28733=>"111111111",
  28734=>"000000100",
  28735=>"000000000",
  28736=>"010110000",
  28737=>"001001000",
  28738=>"000011111",
  28739=>"111110110",
  28740=>"011111111",
  28741=>"000010001",
  28742=>"000000000",
  28743=>"000000000",
  28744=>"011011001",
  28745=>"101111111",
  28746=>"111111111",
  28747=>"110011001",
  28748=>"111111111",
  28749=>"011110000",
  28750=>"000100110",
  28751=>"001000000",
  28752=>"000000000",
  28753=>"111111111",
  28754=>"000001000",
  28755=>"001001001",
  28756=>"110101000",
  28757=>"000000000",
  28758=>"111001000",
  28759=>"000000000",
  28760=>"110110111",
  28761=>"000000001",
  28762=>"001001000",
  28763=>"011011000",
  28764=>"000110111",
  28765=>"111110111",
  28766=>"000000010",
  28767=>"111010000",
  28768=>"000000010",
  28769=>"111111111",
  28770=>"000000000",
  28771=>"111111111",
  28772=>"111100000",
  28773=>"110110001",
  28774=>"110111111",
  28775=>"000111111",
  28776=>"000000000",
  28777=>"110100000",
  28778=>"111001101",
  28779=>"111111111",
  28780=>"001110001",
  28781=>"101001001",
  28782=>"110010010",
  28783=>"111011000",
  28784=>"110111011",
  28785=>"010000111",
  28786=>"100100000",
  28787=>"000111111",
  28788=>"000000000",
  28789=>"000001000",
  28790=>"111111111",
  28791=>"011001011",
  28792=>"000010010",
  28793=>"110110010",
  28794=>"001101111",
  28795=>"101001000",
  28796=>"100100000",
  28797=>"111111111",
  28798=>"100100111",
  28799=>"000001001",
  28800=>"000000000",
  28801=>"000000000",
  28802=>"110110010",
  28803=>"111111111",
  28804=>"000000000",
  28805=>"000000000",
  28806=>"000000000",
  28807=>"111011010",
  28808=>"001001001",
  28809=>"001000001",
  28810=>"111111110",
  28811=>"100000000",
  28812=>"110110110",
  28813=>"000001001",
  28814=>"000000110",
  28815=>"110110111",
  28816=>"111000101",
  28817=>"000001001",
  28818=>"110000000",
  28819=>"000110000",
  28820=>"000000000",
  28821=>"011011011",
  28822=>"000000000",
  28823=>"101001000",
  28824=>"001001110",
  28825=>"000001001",
  28826=>"001001001",
  28827=>"000010110",
  28828=>"111011000",
  28829=>"100110110",
  28830=>"111111000",
  28831=>"000000000",
  28832=>"000000000",
  28833=>"111100000",
  28834=>"111011000",
  28835=>"000000001",
  28836=>"001111111",
  28837=>"011110111",
  28838=>"101000000",
  28839=>"111110111",
  28840=>"111111010",
  28841=>"001001100",
  28842=>"111000000",
  28843=>"111111111",
  28844=>"000000000",
  28845=>"000000011",
  28846=>"111111111",
  28847=>"011011010",
  28848=>"111111011",
  28849=>"001110111",
  28850=>"110110000",
  28851=>"000001101",
  28852=>"111111111",
  28853=>"000000001",
  28854=>"000000101",
  28855=>"000001111",
  28856=>"001000000",
  28857=>"101100100",
  28858=>"000111101",
  28859=>"010110110",
  28860=>"111111111",
  28861=>"110110110",
  28862=>"000000000",
  28863=>"000111111",
  28864=>"111111111",
  28865=>"000000000",
  28866=>"000000101",
  28867=>"110110110",
  28868=>"110000000",
  28869=>"000011000",
  28870=>"111101011",
  28871=>"110111110",
  28872=>"001000000",
  28873=>"001101111",
  28874=>"111001000",
  28875=>"111111111",
  28876=>"111110000",
  28877=>"011001110",
  28878=>"110110000",
  28879=>"110111111",
  28880=>"000000011",
  28881=>"000000100",
  28882=>"111110000",
  28883=>"000001000",
  28884=>"000000000",
  28885=>"000001000",
  28886=>"101000001",
  28887=>"111010111",
  28888=>"010010000",
  28889=>"111111101",
  28890=>"111101001",
  28891=>"111010110",
  28892=>"111111111",
  28893=>"010110110",
  28894=>"100111111",
  28895=>"001000000",
  28896=>"000010000",
  28897=>"001010000",
  28898=>"001000111",
  28899=>"111111011",
  28900=>"000000010",
  28901=>"110110100",
  28902=>"000000000",
  28903=>"000001111",
  28904=>"000101101",
  28905=>"100111111",
  28906=>"111111001",
  28907=>"111111111",
  28908=>"011111111",
  28909=>"111011001",
  28910=>"000000011",
  28911=>"000111111",
  28912=>"111001001",
  28913=>"100110110",
  28914=>"000000001",
  28915=>"110111001",
  28916=>"000000010",
  28917=>"111110000",
  28918=>"011011110",
  28919=>"111111101",
  28920=>"010000000",
  28921=>"011000000",
  28922=>"000000001",
  28923=>"101011111",
  28924=>"111111111",
  28925=>"000000001",
  28926=>"111010011",
  28927=>"111111111",
  28928=>"110000000",
  28929=>"111111111",
  28930=>"000000100",
  28931=>"010010000",
  28932=>"111001111",
  28933=>"110110000",
  28934=>"001000000",
  28935=>"000000000",
  28936=>"000000000",
  28937=>"100100110",
  28938=>"110111110",
  28939=>"001101111",
  28940=>"100100110",
  28941=>"111110110",
  28942=>"000110110",
  28943=>"001001000",
  28944=>"000000000",
  28945=>"111100000",
  28946=>"001101111",
  28947=>"101101111",
  28948=>"001001100",
  28949=>"011000000",
  28950=>"111111000",
  28951=>"000000000",
  28952=>"111111000",
  28953=>"000000000",
  28954=>"000000000",
  28955=>"111111101",
  28956=>"100100100",
  28957=>"000010110",
  28958=>"111111111",
  28959=>"000000010",
  28960=>"001000000",
  28961=>"110111110",
  28962=>"001000111",
  28963=>"111000000",
  28964=>"001000110",
  28965=>"000000000",
  28966=>"111111111",
  28967=>"110100101",
  28968=>"011111111",
  28969=>"000000001",
  28970=>"011010000",
  28971=>"111111010",
  28972=>"001001000",
  28973=>"100100000",
  28974=>"000001000",
  28975=>"111111100",
  28976=>"001101101",
  28977=>"110100101",
  28978=>"000000000",
  28979=>"010000110",
  28980=>"111011000",
  28981=>"111010010",
  28982=>"011111000",
  28983=>"110111111",
  28984=>"011011000",
  28985=>"111000000",
  28986=>"000111111",
  28987=>"000101111",
  28988=>"110000000",
  28989=>"000000000",
  28990=>"000000010",
  28991=>"110001000",
  28992=>"100000000",
  28993=>"000000100",
  28994=>"100100101",
  28995=>"000000000",
  28996=>"000001000",
  28997=>"111011000",
  28998=>"000111111",
  28999=>"000000111",
  29000=>"000000001",
  29001=>"010010000",
  29002=>"000000000",
  29003=>"111110110",
  29004=>"110110111",
  29005=>"000111111",
  29006=>"101111110",
  29007=>"001001001",
  29008=>"001100000",
  29009=>"000000011",
  29010=>"000000000",
  29011=>"001000001",
  29012=>"000111111",
  29013=>"000000001",
  29014=>"001001001",
  29015=>"111110110",
  29016=>"111111111",
  29017=>"001111111",
  29018=>"010110110",
  29019=>"000000100",
  29020=>"110111111",
  29021=>"000000000",
  29022=>"000000001",
  29023=>"111101110",
  29024=>"001001001",
  29025=>"000000101",
  29026=>"000001101",
  29027=>"111100110",
  29028=>"000000000",
  29029=>"000001001",
  29030=>"011111011",
  29031=>"001011011",
  29032=>"110111110",
  29033=>"000000000",
  29034=>"000011011",
  29035=>"100001001",
  29036=>"001001101",
  29037=>"000100100",
  29038=>"111001000",
  29039=>"010000000",
  29040=>"100100000",
  29041=>"000001111",
  29042=>"000000000",
  29043=>"111111111",
  29044=>"010000000",
  29045=>"001000001",
  29046=>"111100000",
  29047=>"111011000",
  29048=>"101000000",
  29049=>"111001000",
  29050=>"001000000",
  29051=>"000000000",
  29052=>"000000100",
  29053=>"000000000",
  29054=>"000000000",
  29055=>"111111111",
  29056=>"110110110",
  29057=>"000000011",
  29058=>"001000000",
  29059=>"111111110",
  29060=>"111111111",
  29061=>"000000000",
  29062=>"100110111",
  29063=>"001000110",
  29064=>"100000111",
  29065=>"111111111",
  29066=>"101001001",
  29067=>"111101000",
  29068=>"000000111",
  29069=>"110111100",
  29070=>"011110111",
  29071=>"010110010",
  29072=>"111001000",
  29073=>"011010010",
  29074=>"111111110",
  29075=>"111100110",
  29076=>"000000000",
  29077=>"011011011",
  29078=>"101111111",
  29079=>"001111001",
  29080=>"000010000",
  29081=>"111110110",
  29082=>"110111111",
  29083=>"000011001",
  29084=>"000000000",
  29085=>"000111001",
  29086=>"000000000",
  29087=>"010110110",
  29088=>"000000101",
  29089=>"001001111",
  29090=>"101011001",
  29091=>"111111111",
  29092=>"001000000",
  29093=>"011001011",
  29094=>"111111000",
  29095=>"101110111",
  29096=>"000000000",
  29097=>"001010110",
  29098=>"000001111",
  29099=>"001000000",
  29100=>"001001001",
  29101=>"000010110",
  29102=>"111110100",
  29103=>"111111111",
  29104=>"111000100",
  29105=>"110110100",
  29106=>"100111111",
  29107=>"111101000",
  29108=>"110110110",
  29109=>"011000000",
  29110=>"101000100",
  29111=>"100110010",
  29112=>"110010011",
  29113=>"101110110",
  29114=>"001001111",
  29115=>"001001101",
  29116=>"000000001",
  29117=>"111110110",
  29118=>"001011111",
  29119=>"001000000",
  29120=>"000000001",
  29121=>"001001000",
  29122=>"001000111",
  29123=>"000000011",
  29124=>"101001101",
  29125=>"111111001",
  29126=>"000000001",
  29127=>"000001111",
  29128=>"000111101",
  29129=>"000000000",
  29130=>"101001001",
  29131=>"011001000",
  29132=>"000000000",
  29133=>"110111111",
  29134=>"011110110",
  29135=>"010010111",
  29136=>"000111111",
  29137=>"000000001",
  29138=>"111110110",
  29139=>"111011000",
  29140=>"011011110",
  29141=>"100100111",
  29142=>"001001011",
  29143=>"011010011",
  29144=>"100000000",
  29145=>"111011000",
  29146=>"001011000",
  29147=>"000000000",
  29148=>"000101100",
  29149=>"110110111",
  29150=>"111000000",
  29151=>"000000001",
  29152=>"011001000",
  29153=>"111111101",
  29154=>"111111011",
  29155=>"111011111",
  29156=>"110110111",
  29157=>"000000000",
  29158=>"000000110",
  29159=>"111001000",
  29160=>"001101111",
  29161=>"111111110",
  29162=>"100000010",
  29163=>"000101000",
  29164=>"000000000",
  29165=>"000010000",
  29166=>"101111111",
  29167=>"000000001",
  29168=>"000000100",
  29169=>"110111111",
  29170=>"000000000",
  29171=>"100111111",
  29172=>"111111110",
  29173=>"111111111",
  29174=>"110110111",
  29175=>"100110110",
  29176=>"111101001",
  29177=>"000000000",
  29178=>"001000000",
  29179=>"110110111",
  29180=>"011011001",
  29181=>"010010110",
  29182=>"000000000",
  29183=>"000000001",
  29184=>"001000000",
  29185=>"000000100",
  29186=>"001001001",
  29187=>"111111111",
  29188=>"001011111",
  29189=>"111111111",
  29190=>"100110110",
  29191=>"111111111",
  29192=>"110111111",
  29193=>"111011110",
  29194=>"001000000",
  29195=>"110000111",
  29196=>"000000100",
  29197=>"000000001",
  29198=>"001111110",
  29199=>"000010011",
  29200=>"010011010",
  29201=>"000000000",
  29202=>"000001111",
  29203=>"100100000",
  29204=>"111111111",
  29205=>"001000000",
  29206=>"101000000",
  29207=>"110111111",
  29208=>"111110110",
  29209=>"000001000",
  29210=>"111000000",
  29211=>"000011011",
  29212=>"111011000",
  29213=>"011000000",
  29214=>"010110110",
  29215=>"111111111",
  29216=>"000000001",
  29217=>"101100000",
  29218=>"000000000",
  29219=>"111111111",
  29220=>"100000000",
  29221=>"011111111",
  29222=>"000000000",
  29223=>"011011011",
  29224=>"000000001",
  29225=>"000100100",
  29226=>"000000000",
  29227=>"000000000",
  29228=>"100001111",
  29229=>"110101000",
  29230=>"111010100",
  29231=>"111001011",
  29232=>"100101111",
  29233=>"000000110",
  29234=>"100111000",
  29235=>"100110110",
  29236=>"111111111",
  29237=>"110100000",
  29238=>"000111111",
  29239=>"000100001",
  29240=>"111111001",
  29241=>"000000000",
  29242=>"000011111",
  29243=>"011111111",
  29244=>"000000000",
  29245=>"000000011",
  29246=>"111110111",
  29247=>"111111111",
  29248=>"000000111",
  29249=>"111100000",
  29250=>"000000100",
  29251=>"000001111",
  29252=>"000000000",
  29253=>"110100000",
  29254=>"111000000",
  29255=>"000000000",
  29256=>"000000001",
  29257=>"111101111",
  29258=>"111111000",
  29259=>"000000000",
  29260=>"011111111",
  29261=>"000000000",
  29262=>"000000000",
  29263=>"001001111",
  29264=>"000000000",
  29265=>"000000000",
  29266=>"000000000",
  29267=>"111111110",
  29268=>"111001111",
  29269=>"000010000",
  29270=>"111111111",
  29271=>"111111111",
  29272=>"000100111",
  29273=>"000000000",
  29274=>"111101111",
  29275=>"000010010",
  29276=>"100100100",
  29277=>"111011111",
  29278=>"000000000",
  29279=>"111111100",
  29280=>"000000111",
  29281=>"001000000",
  29282=>"000000000",
  29283=>"111000011",
  29284=>"000000000",
  29285=>"000000001",
  29286=>"000011111",
  29287=>"111111111",
  29288=>"111001000",
  29289=>"001000000",
  29290=>"000000000",
  29291=>"000000111",
  29292=>"111111101",
  29293=>"111110010",
  29294=>"011000001",
  29295=>"111011000",
  29296=>"011000000",
  29297=>"001101000",
  29298=>"011111010",
  29299=>"000100110",
  29300=>"111111111",
  29301=>"000110010",
  29302=>"000000000",
  29303=>"000000001",
  29304=>"001011111",
  29305=>"000000110",
  29306=>"110110111",
  29307=>"001111111",
  29308=>"000000000",
  29309=>"001001000",
  29310=>"111111111",
  29311=>"000000000",
  29312=>"111111101",
  29313=>"111111000",
  29314=>"111110100",
  29315=>"111111001",
  29316=>"000111111",
  29317=>"101001111",
  29318=>"111111011",
  29319=>"000000111",
  29320=>"001000000",
  29321=>"000000000",
  29322=>"000000111",
  29323=>"000000100",
  29324=>"111111111",
  29325=>"011001111",
  29326=>"011111011",
  29327=>"111111111",
  29328=>"111101101",
  29329=>"111111111",
  29330=>"011111111",
  29331=>"011011111",
  29332=>"111111101",
  29333=>"001001011",
  29334=>"011111111",
  29335=>"111010000",
  29336=>"001100000",
  29337=>"001000000",
  29338=>"000000000",
  29339=>"000000000",
  29340=>"000000000",
  29341=>"000010100",
  29342=>"111111111",
  29343=>"111111111",
  29344=>"100100000",
  29345=>"011111111",
  29346=>"011110100",
  29347=>"110111111",
  29348=>"110110111",
  29349=>"000111010",
  29350=>"000000000",
  29351=>"011001001",
  29352=>"000000000",
  29353=>"000000000",
  29354=>"111111110",
  29355=>"000000110",
  29356=>"110100100",
  29357=>"000110000",
  29358=>"111111111",
  29359=>"011001111",
  29360=>"000000001",
  29361=>"010110000",
  29362=>"110111010",
  29363=>"100000000",
  29364=>"000011001",
  29365=>"000000000",
  29366=>"001101111",
  29367=>"111111111",
  29368=>"000000000",
  29369=>"101000001",
  29370=>"111000010",
  29371=>"100000000",
  29372=>"111111111",
  29373=>"000000000",
  29374=>"100110111",
  29375=>"110100101",
  29376=>"011000000",
  29377=>"000100000",
  29378=>"110100110",
  29379=>"111111111",
  29380=>"000000000",
  29381=>"000000001",
  29382=>"010000100",
  29383=>"011011111",
  29384=>"000100100",
  29385=>"001000000",
  29386=>"111111011",
  29387=>"101001000",
  29388=>"001111111",
  29389=>"111111111",
  29390=>"000010111",
  29391=>"111111111",
  29392=>"111111111",
  29393=>"111100111",
  29394=>"011000001",
  29395=>"000100000",
  29396=>"001000001",
  29397=>"000110111",
  29398=>"000000101",
  29399=>"111111111",
  29400=>"111111000",
  29401=>"100110111",
  29402=>"011111010",
  29403=>"000001000",
  29404=>"000010010",
  29405=>"111011111",
  29406=>"000000100",
  29407=>"000010000",
  29408=>"110100000",
  29409=>"111111110",
  29410=>"101000001",
  29411=>"000110110",
  29412=>"110110010",
  29413=>"110000001",
  29414=>"111011011",
  29415=>"000001001",
  29416=>"111111111",
  29417=>"000000000",
  29418=>"000000000",
  29419=>"000000100",
  29420=>"111000001",
  29421=>"100000001",
  29422=>"001111111",
  29423=>"001001001",
  29424=>"011001000",
  29425=>"110110100",
  29426=>"000000000",
  29427=>"000000000",
  29428=>"111101000",
  29429=>"011111110",
  29430=>"000000000",
  29431=>"111110100",
  29432=>"111111111",
  29433=>"000000000",
  29434=>"000001000",
  29435=>"100100100",
  29436=>"011011001",
  29437=>"001001000",
  29438=>"111111111",
  29439=>"010111111",
  29440=>"000000000",
  29441=>"011011010",
  29442=>"000000000",
  29443=>"011010000",
  29444=>"000000000",
  29445=>"000100100",
  29446=>"111111111",
  29447=>"001000000",
  29448=>"000010011",
  29449=>"110000111",
  29450=>"000000001",
  29451=>"111110000",
  29452=>"001000001",
  29453=>"111011100",
  29454=>"101100000",
  29455=>"010000000",
  29456=>"001010110",
  29457=>"000111111",
  29458=>"000000000",
  29459=>"011011111",
  29460=>"000000000",
  29461=>"111111101",
  29462=>"000000000",
  29463=>"000001111",
  29464=>"001000100",
  29465=>"111100100",
  29466=>"001000011",
  29467=>"100000010",
  29468=>"000000000",
  29469=>"000000000",
  29470=>"000000000",
  29471=>"001100111",
  29472=>"100000110",
  29473=>"111111111",
  29474=>"111011000",
  29475=>"111100000",
  29476=>"100100100",
  29477=>"000000111",
  29478=>"001111011",
  29479=>"001111110",
  29480=>"111111111",
  29481=>"000000000",
  29482=>"000100100",
  29483=>"111110110",
  29484=>"110111011",
  29485=>"010010111",
  29486=>"000011000",
  29487=>"000000000",
  29488=>"000100110",
  29489=>"111111011",
  29490=>"001000000",
  29491=>"111011000",
  29492=>"000000111",
  29493=>"000000100",
  29494=>"000000001",
  29495=>"111000000",
  29496=>"000000000",
  29497=>"111111100",
  29498=>"110000000",
  29499=>"000001001",
  29500=>"100100000",
  29501=>"000100000",
  29502=>"111111111",
  29503=>"100111001",
  29504=>"000111111",
  29505=>"000010111",
  29506=>"111111111",
  29507=>"101011011",
  29508=>"011011000",
  29509=>"010110111",
  29510=>"000010010",
  29511=>"000000000",
  29512=>"111101000",
  29513=>"111111111",
  29514=>"011111111",
  29515=>"111111111",
  29516=>"111111110",
  29517=>"101100000",
  29518=>"000001011",
  29519=>"111111111",
  29520=>"100000000",
  29521=>"000111111",
  29522=>"000000000",
  29523=>"000000000",
  29524=>"111111111",
  29525=>"011001011",
  29526=>"111111111",
  29527=>"011000000",
  29528=>"111111111",
  29529=>"001001010",
  29530=>"000000000",
  29531=>"111111110",
  29532=>"000000000",
  29533=>"111111111",
  29534=>"011111000",
  29535=>"110111101",
  29536=>"000000000",
  29537=>"001000000",
  29538=>"000000011",
  29539=>"111111111",
  29540=>"000000000",
  29541=>"011010110",
  29542=>"111101111",
  29543=>"111111111",
  29544=>"011011000",
  29545=>"111111110",
  29546=>"111111011",
  29547=>"111011000",
  29548=>"000000000",
  29549=>"001011111",
  29550=>"000000000",
  29551=>"111111111",
  29552=>"000000000",
  29553=>"000000000",
  29554=>"111000000",
  29555=>"001000001",
  29556=>"111110110",
  29557=>"110110110",
  29558=>"011111111",
  29559=>"000010010",
  29560=>"000000100",
  29561=>"111111111",
  29562=>"000000000",
  29563=>"110011111",
  29564=>"110010000",
  29565=>"111110111",
  29566=>"011001000",
  29567=>"000000000",
  29568=>"000000000",
  29569=>"001111111",
  29570=>"111111011",
  29571=>"100110111",
  29572=>"110111111",
  29573=>"000000000",
  29574=>"110111100",
  29575=>"000000100",
  29576=>"000000000",
  29577=>"011010001",
  29578=>"000001001",
  29579=>"111000000",
  29580=>"111111111",
  29581=>"001111010",
  29582=>"000000000",
  29583=>"111000000",
  29584=>"100000000",
  29585=>"111111111",
  29586=>"000010110",
  29587=>"001001111",
  29588=>"000000001",
  29589=>"000000000",
  29590=>"111111111",
  29591=>"111111111",
  29592=>"000000000",
  29593=>"011010010",
  29594=>"100010000",
  29595=>"000000110",
  29596=>"000000001",
  29597=>"111111111",
  29598=>"000000000",
  29599=>"000000011",
  29600=>"110000000",
  29601=>"000000010",
  29602=>"111011001",
  29603=>"010100100",
  29604=>"000000000",
  29605=>"111111011",
  29606=>"000001000",
  29607=>"111100110",
  29608=>"010001001",
  29609=>"111111111",
  29610=>"000000001",
  29611=>"000000101",
  29612=>"000000000",
  29613=>"001111111",
  29614=>"000111111",
  29615=>"000101111",
  29616=>"000100111",
  29617=>"111000000",
  29618=>"000110110",
  29619=>"100100100",
  29620=>"111110111",
  29621=>"111111111",
  29622=>"000100111",
  29623=>"111111111",
  29624=>"111111111",
  29625=>"111111111",
  29626=>"100000000",
  29627=>"001000000",
  29628=>"111111110",
  29629=>"111111111",
  29630=>"100000000",
  29631=>"011011010",
  29632=>"000000000",
  29633=>"111111111",
  29634=>"000000000",
  29635=>"000100111",
  29636=>"000010000",
  29637=>"110100000",
  29638=>"000000000",
  29639=>"111101001",
  29640=>"001100000",
  29641=>"111111000",
  29642=>"000000000",
  29643=>"111111111",
  29644=>"111111000",
  29645=>"001001001",
  29646=>"000000000",
  29647=>"110110111",
  29648=>"111111111",
  29649=>"000000101",
  29650=>"001000000",
  29651=>"000000000",
  29652=>"000000110",
  29653=>"000110111",
  29654=>"000000011",
  29655=>"001111011",
  29656=>"000111010",
  29657=>"011111100",
  29658=>"100110110",
  29659=>"000000000",
  29660=>"000111111",
  29661=>"011011000",
  29662=>"111111001",
  29663=>"001011011",
  29664=>"111101001",
  29665=>"111100100",
  29666=>"000000000",
  29667=>"111111111",
  29668=>"000000100",
  29669=>"110010000",
  29670=>"100100100",
  29671=>"010111111",
  29672=>"111111111",
  29673=>"111011001",
  29674=>"011101100",
  29675=>"111111011",
  29676=>"000010110",
  29677=>"001111111",
  29678=>"000000000",
  29679=>"000010111",
  29680=>"111100101",
  29681=>"000000000",
  29682=>"111111000",
  29683=>"000000000",
  29684=>"011010100",
  29685=>"000111111",
  29686=>"111111111",
  29687=>"000000000",
  29688=>"001101111",
  29689=>"111111011",
  29690=>"011011110",
  29691=>"111100000",
  29692=>"000110111",
  29693=>"011101111",
  29694=>"011011010",
  29695=>"000000000",
  29696=>"111111000",
  29697=>"000000000",
  29698=>"111111111",
  29699=>"111111111",
  29700=>"110111110",
  29701=>"000000000",
  29702=>"111111111",
  29703=>"111111111",
  29704=>"000000000",
  29705=>"111111111",
  29706=>"000100111",
  29707=>"100100000",
  29708=>"100110000",
  29709=>"001111111",
  29710=>"000000111",
  29711=>"000000000",
  29712=>"000000110",
  29713=>"111011011",
  29714=>"000000001",
  29715=>"100011111",
  29716=>"111111111",
  29717=>"001011001",
  29718=>"111101000",
  29719=>"000000110",
  29720=>"001011111",
  29721=>"000000000",
  29722=>"000000001",
  29723=>"100000000",
  29724=>"000000000",
  29725=>"000000000",
  29726=>"000000000",
  29727=>"111000000",
  29728=>"111000000",
  29729=>"000000000",
  29730=>"000000000",
  29731=>"111110010",
  29732=>"010111100",
  29733=>"000000000",
  29734=>"000000000",
  29735=>"100110000",
  29736=>"111111111",
  29737=>"000000000",
  29738=>"000000000",
  29739=>"011111011",
  29740=>"111111111",
  29741=>"111010000",
  29742=>"001001001",
  29743=>"001000000",
  29744=>"111111111",
  29745=>"000000000",
  29746=>"000000000",
  29747=>"000000000",
  29748=>"111111111",
  29749=>"100110000",
  29750=>"101101001",
  29751=>"001001101",
  29752=>"111000001",
  29753=>"000011111",
  29754=>"000011101",
  29755=>"000000000",
  29756=>"000101111",
  29757=>"111111101",
  29758=>"111011110",
  29759=>"001001101",
  29760=>"000000000",
  29761=>"000000000",
  29762=>"000000000",
  29763=>"111111111",
  29764=>"111001101",
  29765=>"011011011",
  29766=>"000000000",
  29767=>"000111111",
  29768=>"011011111",
  29769=>"000001111",
  29770=>"111111111",
  29771=>"111111010",
  29772=>"111111101",
  29773=>"111111000",
  29774=>"111111000",
  29775=>"000000000",
  29776=>"000010110",
  29777=>"001101111",
  29778=>"110111111",
  29779=>"111111111",
  29780=>"000000000",
  29781=>"111111010",
  29782=>"000011000",
  29783=>"111111111",
  29784=>"001111000",
  29785=>"111000000",
  29786=>"111100100",
  29787=>"100100100",
  29788=>"000010000",
  29789=>"001010011",
  29790=>"100100111",
  29791=>"000000100",
  29792=>"111111111",
  29793=>"000000000",
  29794=>"000000000",
  29795=>"110111000",
  29796=>"111111011",
  29797=>"111111000",
  29798=>"111101111",
  29799=>"000000000",
  29800=>"000000000",
  29801=>"000000000",
  29802=>"000000111",
  29803=>"000000000",
  29804=>"011111111",
  29805=>"111111111",
  29806=>"101111111",
  29807=>"111111111",
  29808=>"000000000",
  29809=>"010000000",
  29810=>"111111111",
  29811=>"000000000",
  29812=>"000000100",
  29813=>"000000101",
  29814=>"111000001",
  29815=>"001111111",
  29816=>"000000000",
  29817=>"111001000",
  29818=>"000000000",
  29819=>"111110100",
  29820=>"000000000",
  29821=>"111111100",
  29822=>"111101000",
  29823=>"000000000",
  29824=>"111111111",
  29825=>"000000000",
  29826=>"001000000",
  29827=>"000000000",
  29828=>"111111111",
  29829=>"000000001",
  29830=>"110110000",
  29831=>"000000000",
  29832=>"111011111",
  29833=>"000000001",
  29834=>"111000000",
  29835=>"111000000",
  29836=>"000000000",
  29837=>"000000000",
  29838=>"100000000",
  29839=>"110110110",
  29840=>"111111111",
  29841=>"011111110",
  29842=>"000000000",
  29843=>"000111011",
  29844=>"000001111",
  29845=>"001000000",
  29846=>"000000111",
  29847=>"111111111",
  29848=>"110111111",
  29849=>"111111111",
  29850=>"111111001",
  29851=>"000000000",
  29852=>"000110011",
  29853=>"000000000",
  29854=>"011010110",
  29855=>"000000111",
  29856=>"000000101",
  29857=>"001000000",
  29858=>"001111111",
  29859=>"010111111",
  29860=>"110100000",
  29861=>"110000000",
  29862=>"000000111",
  29863=>"111111111",
  29864=>"111111111",
  29865=>"001000000",
  29866=>"000011010",
  29867=>"111111111",
  29868=>"101111111",
  29869=>"011001000",
  29870=>"000000000",
  29871=>"000000111",
  29872=>"000000000",
  29873=>"000000000",
  29874=>"111011000",
  29875=>"000000100",
  29876=>"100100000",
  29877=>"000000000",
  29878=>"000000000",
  29879=>"000000001",
  29880=>"111110011",
  29881=>"111111101",
  29882=>"111000000",
  29883=>"111111001",
  29884=>"111111110",
  29885=>"001011001",
  29886=>"000000001",
  29887=>"000000000",
  29888=>"101101111",
  29889=>"000000000",
  29890=>"111110011",
  29891=>"000000000",
  29892=>"000000001",
  29893=>"111111111",
  29894=>"000101111",
  29895=>"111111111",
  29896=>"111001001",
  29897=>"000000000",
  29898=>"001011111",
  29899=>"111001001",
  29900=>"001111111",
  29901=>"010001011",
  29902=>"000000000",
  29903=>"000000000",
  29904=>"000000000",
  29905=>"010000000",
  29906=>"000111100",
  29907=>"000110110",
  29908=>"011111111",
  29909=>"000000100",
  29910=>"111111111",
  29911=>"000000000",
  29912=>"000000110",
  29913=>"110100100",
  29914=>"000001111",
  29915=>"011000000",
  29916=>"000000101",
  29917=>"000000000",
  29918=>"000000000",
  29919=>"101000111",
  29920=>"010010110",
  29921=>"000000000",
  29922=>"000000000",
  29923=>"111110000",
  29924=>"100000000",
  29925=>"010011001",
  29926=>"111100100",
  29927=>"100110111",
  29928=>"111111111",
  29929=>"000000000",
  29930=>"111111111",
  29931=>"111000000",
  29932=>"111111111",
  29933=>"110000100",
  29934=>"110101000",
  29935=>"111111101",
  29936=>"000000000",
  29937=>"111111111",
  29938=>"000000000",
  29939=>"111000100",
  29940=>"000100100",
  29941=>"000000000",
  29942=>"000000000",
  29943=>"111111010",
  29944=>"111111111",
  29945=>"000000000",
  29946=>"000000000",
  29947=>"111010000",
  29948=>"000110110",
  29949=>"100000111",
  29950=>"010111110",
  29951=>"101101111",
  29952=>"110111111",
  29953=>"000000000",
  29954=>"111111111",
  29955=>"111000000",
  29956=>"111111111",
  29957=>"000011001",
  29958=>"101000000",
  29959=>"111110011",
  29960=>"110111011",
  29961=>"000011000",
  29962=>"001001000",
  29963=>"011010000",
  29964=>"000000000",
  29965=>"111111111",
  29966=>"111111111",
  29967=>"111111111",
  29968=>"001110111",
  29969=>"100101111",
  29970=>"111000111",
  29971=>"001000000",
  29972=>"000001000",
  29973=>"000000110",
  29974=>"100000000",
  29975=>"111111110",
  29976=>"011011000",
  29977=>"111110010",
  29978=>"001001001",
  29979=>"000000001",
  29980=>"000000000",
  29981=>"011000000",
  29982=>"010100000",
  29983=>"011001001",
  29984=>"000000100",
  29985=>"111111101",
  29986=>"111111111",
  29987=>"111111111",
  29988=>"000010010",
  29989=>"000000111",
  29990=>"001001111",
  29991=>"011010010",
  29992=>"000000000",
  29993=>"000001000",
  29994=>"001000000",
  29995=>"100000000",
  29996=>"000000000",
  29997=>"010111110",
  29998=>"111111111",
  29999=>"000000110",
  30000=>"000000000",
  30001=>"000000000",
  30002=>"110000000",
  30003=>"111110111",
  30004=>"111011000",
  30005=>"001001000",
  30006=>"011111111",
  30007=>"111001000",
  30008=>"000001111",
  30009=>"000000000",
  30010=>"111110001",
  30011=>"111111111",
  30012=>"000000000",
  30013=>"001000100",
  30014=>"000100111",
  30015=>"111111111",
  30016=>"111111111",
  30017=>"000100000",
  30018=>"000000000",
  30019=>"011000000",
  30020=>"000000000",
  30021=>"001001000",
  30022=>"000000000",
  30023=>"111111111",
  30024=>"000000000",
  30025=>"000000000",
  30026=>"111110000",
  30027=>"000000000",
  30028=>"001000000",
  30029=>"000000111",
  30030=>"011001111",
  30031=>"111111111",
  30032=>"010110110",
  30033=>"110000100",
  30034=>"111111111",
  30035=>"111111110",
  30036=>"110111111",
  30037=>"011111111",
  30038=>"111101000",
  30039=>"000000111",
  30040=>"001001001",
  30041=>"000000000",
  30042=>"001000000",
  30043=>"000000000",
  30044=>"110110110",
  30045=>"001001001",
  30046=>"111111111",
  30047=>"111111111",
  30048=>"010000110",
  30049=>"111111111",
  30050=>"000000000",
  30051=>"000000000",
  30052=>"100101101",
  30053=>"111111110",
  30054=>"111110111",
  30055=>"111111111",
  30056=>"000100100",
  30057=>"000000100",
  30058=>"001000000",
  30059=>"100000001",
  30060=>"110000110",
  30061=>"111001101",
  30062=>"000000001",
  30063=>"011010000",
  30064=>"000000000",
  30065=>"111111011",
  30066=>"111000100",
  30067=>"001000000",
  30068=>"000000000",
  30069=>"111111001",
  30070=>"110110111",
  30071=>"111001000",
  30072=>"000000000",
  30073=>"000101000",
  30074=>"111100111",
  30075=>"010000111",
  30076=>"000000010",
  30077=>"110000000",
  30078=>"111111000",
  30079=>"011111111",
  30080=>"001001001",
  30081=>"111011111",
  30082=>"110110110",
  30083=>"000000000",
  30084=>"000111111",
  30085=>"000000000",
  30086=>"000000000",
  30087=>"000000000",
  30088=>"111111111",
  30089=>"000000000",
  30090=>"000000000",
  30091=>"111111111",
  30092=>"001000000",
  30093=>"001000000",
  30094=>"000000000",
  30095=>"111111011",
  30096=>"000000000",
  30097=>"111100000",
  30098=>"011111111",
  30099=>"000100100",
  30100=>"001000000",
  30101=>"000000000",
  30102=>"000010011",
  30103=>"111111111",
  30104=>"101111111",
  30105=>"000000001",
  30106=>"000000101",
  30107=>"001111111",
  30108=>"000101111",
  30109=>"001001001",
  30110=>"101001111",
  30111=>"010010000",
  30112=>"111111000",
  30113=>"001111111",
  30114=>"111111111",
  30115=>"111111111",
  30116=>"000000000",
  30117=>"010010010",
  30118=>"111101000",
  30119=>"001001000",
  30120=>"000000000",
  30121=>"111111111",
  30122=>"110100000",
  30123=>"000000000",
  30124=>"000000000",
  30125=>"000100111",
  30126=>"000000010",
  30127=>"010010000",
  30128=>"111001111",
  30129=>"000000000",
  30130=>"010000000",
  30131=>"111111111",
  30132=>"111110110",
  30133=>"111111111",
  30134=>"000000001",
  30135=>"000000000",
  30136=>"000000000",
  30137=>"000000000",
  30138=>"000000000",
  30139=>"111111111",
  30140=>"111000000",
  30141=>"111111101",
  30142=>"111011000",
  30143=>"100000000",
  30144=>"000000000",
  30145=>"000000111",
  30146=>"111111111",
  30147=>"110100001",
  30148=>"000011001",
  30149=>"001000100",
  30150=>"000000000",
  30151=>"111111111",
  30152=>"100000000",
  30153=>"000110100",
  30154=>"000000111",
  30155=>"000000000",
  30156=>"100100111",
  30157=>"000000000",
  30158=>"111111101",
  30159=>"111111111",
  30160=>"111111001",
  30161=>"000000111",
  30162=>"000000000",
  30163=>"000111010",
  30164=>"111000000",
  30165=>"100111111",
  30166=>"110000000",
  30167=>"001000000",
  30168=>"010000101",
  30169=>"110010111",
  30170=>"111110000",
  30171=>"111111111",
  30172=>"011111000",
  30173=>"111111010",
  30174=>"111011000",
  30175=>"000000011",
  30176=>"111111100",
  30177=>"111111111",
  30178=>"000000000",
  30179=>"111111111",
  30180=>"111001100",
  30181=>"000000001",
  30182=>"011000011",
  30183=>"111111111",
  30184=>"011011111",
  30185=>"111111111",
  30186=>"000000000",
  30187=>"111111111",
  30188=>"111111111",
  30189=>"111100100",
  30190=>"100000000",
  30191=>"111111111",
  30192=>"100101100",
  30193=>"000000001",
  30194=>"100100111",
  30195=>"111100100",
  30196=>"000000000",
  30197=>"110000000",
  30198=>"001101000",
  30199=>"101111101",
  30200=>"000000000",
  30201=>"000011111",
  30202=>"100110000",
  30203=>"111111111",
  30204=>"111101111",
  30205=>"010000000",
  30206=>"111111111",
  30207=>"100000111",
  30208=>"000000000",
  30209=>"000000000",
  30210=>"101110010",
  30211=>"111111101",
  30212=>"000000111",
  30213=>"001001100",
  30214=>"000000000",
  30215=>"111111111",
  30216=>"111111111",
  30217=>"111111111",
  30218=>"000000000",
  30219=>"011111111",
  30220=>"000000000",
  30221=>"100000000",
  30222=>"000000000",
  30223=>"000000000",
  30224=>"011000111",
  30225=>"000000000",
  30226=>"000000000",
  30227=>"011011111",
  30228=>"111111111",
  30229=>"000001001",
  30230=>"111111111",
  30231=>"111111010",
  30232=>"000000000",
  30233=>"011000000",
  30234=>"000000000",
  30235=>"111011001",
  30236=>"111100100",
  30237=>"011000000",
  30238=>"000100000",
  30239=>"111100000",
  30240=>"000000000",
  30241=>"111111111",
  30242=>"111111101",
  30243=>"001110111",
  30244=>"111100000",
  30245=>"011111111",
  30246=>"111110111",
  30247=>"111111111",
  30248=>"101111111",
  30249=>"000000000",
  30250=>"000000001",
  30251=>"111001100",
  30252=>"111111111",
  30253=>"000101001",
  30254=>"101101101",
  30255=>"000000011",
  30256=>"000000000",
  30257=>"000000000",
  30258=>"100110110",
  30259=>"000000000",
  30260=>"000001000",
  30261=>"000000000",
  30262=>"011001100",
  30263=>"001101111",
  30264=>"000000111",
  30265=>"101111111",
  30266=>"000111000",
  30267=>"000000000",
  30268=>"110000100",
  30269=>"111101111",
  30270=>"000000111",
  30271=>"011111111",
  30272=>"100100000",
  30273=>"111110110",
  30274=>"000000000",
  30275=>"111111110",
  30276=>"110110110",
  30277=>"000000000",
  30278=>"111101001",
  30279=>"000000000",
  30280=>"011011011",
  30281=>"111111100",
  30282=>"001100111",
  30283=>"111111000",
  30284=>"000000100",
  30285=>"111111000",
  30286=>"100101101",
  30287=>"000000000",
  30288=>"111000000",
  30289=>"100111111",
  30290=>"110111111",
  30291=>"011011111",
  30292=>"110000000",
  30293=>"000000000",
  30294=>"110000100",
  30295=>"111110110",
  30296=>"111111111",
  30297=>"111101111",
  30298=>"000000000",
  30299=>"110100001",
  30300=>"000000000",
  30301=>"000000000",
  30302=>"001001000",
  30303=>"000111111",
  30304=>"111111111",
  30305=>"001000000",
  30306=>"111111111",
  30307=>"000010000",
  30308=>"010110011",
  30309=>"001111111",
  30310=>"000000000",
  30311=>"000000000",
  30312=>"111111011",
  30313=>"110100000",
  30314=>"000110000",
  30315=>"111111111",
  30316=>"111111100",
  30317=>"111111111",
  30318=>"000101111",
  30319=>"011000000",
  30320=>"001111011",
  30321=>"000000000",
  30322=>"111111111",
  30323=>"001001000",
  30324=>"111111111",
  30325=>"111111111",
  30326=>"000000001",
  30327=>"000000100",
  30328=>"001111111",
  30329=>"111111000",
  30330=>"101000000",
  30331=>"111001000",
  30332=>"111111000",
  30333=>"000000000",
  30334=>"111111111",
  30335=>"111101111",
  30336=>"111111111",
  30337=>"111111111",
  30338=>"111111111",
  30339=>"011011011",
  30340=>"111111111",
  30341=>"011101111",
  30342=>"110100101",
  30343=>"111111000",
  30344=>"100111111",
  30345=>"000000000",
  30346=>"000000000",
  30347=>"111111111",
  30348=>"001000000",
  30349=>"000000001",
  30350=>"000000000",
  30351=>"000000000",
  30352=>"110111111",
  30353=>"000000000",
  30354=>"000011011",
  30355=>"000011111",
  30356=>"000010111",
  30357=>"110000001",
  30358=>"000000000",
  30359=>"111000111",
  30360=>"100000000",
  30361=>"100100001",
  30362=>"111111111",
  30363=>"001000110",
  30364=>"011111111",
  30365=>"111111111",
  30366=>"111110111",
  30367=>"000000000",
  30368=>"010010100",
  30369=>"000110111",
  30370=>"111111111",
  30371=>"000000000",
  30372=>"111100000",
  30373=>"000000000",
  30374=>"110111111",
  30375=>"011111111",
  30376=>"111111111",
  30377=>"111111111",
  30378=>"001000001",
  30379=>"111111111",
  30380=>"000000000",
  30381=>"000011110",
  30382=>"000000000",
  30383=>"000111000",
  30384=>"100111000",
  30385=>"000000110",
  30386=>"110110110",
  30387=>"111111111",
  30388=>"111111111",
  30389=>"101001000",
  30390=>"000000111",
  30391=>"000000001",
  30392=>"101001000",
  30393=>"111111111",
  30394=>"100000000",
  30395=>"111011000",
  30396=>"111101111",
  30397=>"000001000",
  30398=>"111111111",
  30399=>"000000000",
  30400=>"110110010",
  30401=>"111111111",
  30402=>"111111111",
  30403=>"111101000",
  30404=>"111111111",
  30405=>"111111000",
  30406=>"111001000",
  30407=>"000000000",
  30408=>"000000000",
  30409=>"111101111",
  30410=>"011001101",
  30411=>"000000000",
  30412=>"111111111",
  30413=>"000111000",
  30414=>"010111000",
  30415=>"000000000",
  30416=>"011111000",
  30417=>"000111111",
  30418=>"111111001",
  30419=>"000000000",
  30420=>"000111111",
  30421=>"001000000",
  30422=>"111111111",
  30423=>"000100000",
  30424=>"111111111",
  30425=>"111111111",
  30426=>"001001111",
  30427=>"001000100",
  30428=>"000000000",
  30429=>"111111110",
  30430=>"111101000",
  30431=>"000101111",
  30432=>"000000000",
  30433=>"100000000",
  30434=>"011011111",
  30435=>"000000000",
  30436=>"000000000",
  30437=>"111111110",
  30438=>"111000000",
  30439=>"000101111",
  30440=>"111111000",
  30441=>"110011111",
  30442=>"000000000",
  30443=>"000000111",
  30444=>"000000000",
  30445=>"000001111",
  30446=>"110110100",
  30447=>"110000000",
  30448=>"000010010",
  30449=>"000000000",
  30450=>"111111101",
  30451=>"111111000",
  30452=>"011011011",
  30453=>"011111111",
  30454=>"111111110",
  30455=>"111111000",
  30456=>"000111111",
  30457=>"000000000",
  30458=>"111111111",
  30459=>"111111111",
  30460=>"111111111",
  30461=>"000000000",
  30462=>"110111110",
  30463=>"111100001",
  30464=>"111111110",
  30465=>"101111111",
  30466=>"111111111",
  30467=>"111111011",
  30468=>"000000000",
  30469=>"111111111",
  30470=>"000000000",
  30471=>"100000000",
  30472=>"111001101",
  30473=>"011110010",
  30474=>"000000000",
  30475=>"111111111",
  30476=>"110110000",
  30477=>"111111111",
  30478=>"111111111",
  30479=>"000111111",
  30480=>"001001011",
  30481=>"000001111",
  30482=>"111111111",
  30483=>"111111111",
  30484=>"110111111",
  30485=>"001101111",
  30486=>"000000000",
  30487=>"000010000",
  30488=>"000000000",
  30489=>"100000000",
  30490=>"000000000",
  30491=>"111111111",
  30492=>"000000110",
  30493=>"011000000",
  30494=>"111111111",
  30495=>"000000000",
  30496=>"011000011",
  30497=>"000000000",
  30498=>"000000000",
  30499=>"110111111",
  30500=>"111111111",
  30501=>"000000000",
  30502=>"000000001",
  30503=>"111110100",
  30504=>"111111001",
  30505=>"000100111",
  30506=>"111111101",
  30507=>"111111111",
  30508=>"111000000",
  30509=>"110100100",
  30510=>"110010111",
  30511=>"111111111",
  30512=>"111111111",
  30513=>"000000000",
  30514=>"111111111",
  30515=>"000000000",
  30516=>"000000000",
  30517=>"111001000",
  30518=>"111001001",
  30519=>"111011000",
  30520=>"000000000",
  30521=>"001000000",
  30522=>"111111111",
  30523=>"010000000",
  30524=>"000000000",
  30525=>"011111111",
  30526=>"000000000",
  30527=>"000000000",
  30528=>"111111000",
  30529=>"001111010",
  30530=>"101001001",
  30531=>"111000000",
  30532=>"101001000",
  30533=>"111000000",
  30534=>"000000000",
  30535=>"000000111",
  30536=>"100000000",
  30537=>"000111111",
  30538=>"111111001",
  30539=>"100101101",
  30540=>"111011000",
  30541=>"111111111",
  30542=>"100110111",
  30543=>"000100110",
  30544=>"001011011",
  30545=>"000000000",
  30546=>"100000000",
  30547=>"100000111",
  30548=>"100100111",
  30549=>"001001001",
  30550=>"111011111",
  30551=>"101111101",
  30552=>"111100101",
  30553=>"110010000",
  30554=>"000000000",
  30555=>"111010000",
  30556=>"010111110",
  30557=>"111111000",
  30558=>"101111111",
  30559=>"000000000",
  30560=>"111111111",
  30561=>"000000000",
  30562=>"000000000",
  30563=>"110011111",
  30564=>"100100110",
  30565=>"100000000",
  30566=>"100111000",
  30567=>"011011111",
  30568=>"100000110",
  30569=>"000000000",
  30570=>"011111111",
  30571=>"110110000",
  30572=>"110111111",
  30573=>"000000000",
  30574=>"000000000",
  30575=>"101000000",
  30576=>"000000000",
  30577=>"111111001",
  30578=>"000111000",
  30579=>"000000001",
  30580=>"111011001",
  30581=>"111111111",
  30582=>"111111111",
  30583=>"111111111",
  30584=>"111101000",
  30585=>"111111111",
  30586=>"111111111",
  30587=>"100101111",
  30588=>"001001001",
  30589=>"000000111",
  30590=>"000000000",
  30591=>"100100100",
  30592=>"100000000",
  30593=>"111111010",
  30594=>"000000000",
  30595=>"111111111",
  30596=>"111111010",
  30597=>"110110000",
  30598=>"000000000",
  30599=>"000000000",
  30600=>"000000100",
  30601=>"111111111",
  30602=>"000011111",
  30603=>"111111111",
  30604=>"111111111",
  30605=>"000110000",
  30606=>"000000000",
  30607=>"000000000",
  30608=>"111111111",
  30609=>"000000000",
  30610=>"000000000",
  30611=>"110011001",
  30612=>"111111111",
  30613=>"010111111",
  30614=>"111101101",
  30615=>"000000000",
  30616=>"011001111",
  30617=>"001111011",
  30618=>"000000000",
  30619=>"000000100",
  30620=>"001111111",
  30621=>"111111111",
  30622=>"000000000",
  30623=>"111011001",
  30624=>"000000000",
  30625=>"110100000",
  30626=>"001000000",
  30627=>"000000000",
  30628=>"011000000",
  30629=>"111111111",
  30630=>"111111111",
  30631=>"000000000",
  30632=>"000000000",
  30633=>"111011111",
  30634=>"111111111",
  30635=>"111111001",
  30636=>"100000001",
  30637=>"010010010",
  30638=>"111111111",
  30639=>"000000000",
  30640=>"000111111",
  30641=>"111010000",
  30642=>"000000000",
  30643=>"000000000",
  30644=>"000011111",
  30645=>"111111101",
  30646=>"000000110",
  30647=>"111011001",
  30648=>"000000000",
  30649=>"000000000",
  30650=>"111111111",
  30651=>"011111110",
  30652=>"000000001",
  30653=>"111111111",
  30654=>"110110000",
  30655=>"100000000",
  30656=>"000000100",
  30657=>"111011011",
  30658=>"111111111",
  30659=>"111111111",
  30660=>"000000000",
  30661=>"000000000",
  30662=>"111000000",
  30663=>"011111001",
  30664=>"110000000",
  30665=>"111111111",
  30666=>"111111111",
  30667=>"000000110",
  30668=>"111110111",
  30669=>"000000001",
  30670=>"110000000",
  30671=>"001011000",
  30672=>"110111111",
  30673=>"111111110",
  30674=>"111111111",
  30675=>"000000111",
  30676=>"111100000",
  30677=>"000000000",
  30678=>"100111111",
  30679=>"001011000",
  30680=>"000000000",
  30681=>"000000000",
  30682=>"110110100",
  30683=>"101001111",
  30684=>"111110000",
  30685=>"111111000",
  30686=>"000000000",
  30687=>"110111111",
  30688=>"000010010",
  30689=>"110000010",
  30690=>"000000100",
  30691=>"100001001",
  30692=>"000001000",
  30693=>"111111000",
  30694=>"100000000",
  30695=>"000000001",
  30696=>"111111110",
  30697=>"000000000",
  30698=>"110000000",
  30699=>"111111111",
  30700=>"111111111",
  30701=>"000000000",
  30702=>"000000000",
  30703=>"111101111",
  30704=>"000010110",
  30705=>"000101000",
  30706=>"011000000",
  30707=>"000010111",
  30708=>"000000000",
  30709=>"111111111",
  30710=>"100100010",
  30711=>"111110110",
  30712=>"111111111",
  30713=>"000000000",
  30714=>"000000000",
  30715=>"000000000",
  30716=>"000000000",
  30717=>"001000000",
  30718=>"000000000",
  30719=>"111111111",
  30720=>"110010010",
  30721=>"001000000",
  30722=>"101111111",
  30723=>"000000001",
  30724=>"001001111",
  30725=>"111111111",
  30726=>"000000000",
  30727=>"111111111",
  30728=>"111100100",
  30729=>"111001000",
  30730=>"111001001",
  30731=>"001101000",
  30732=>"000000001",
  30733=>"000000100",
  30734=>"111001100",
  30735=>"000000101",
  30736=>"110110111",
  30737=>"010011111",
  30738=>"010110110",
  30739=>"100000000",
  30740=>"010000010",
  30741=>"111000000",
  30742=>"000000000",
  30743=>"011011001",
  30744=>"111111111",
  30745=>"000111100",
  30746=>"000110000",
  30747=>"110100110",
  30748=>"001001001",
  30749=>"011110100",
  30750=>"110100100",
  30751=>"000000111",
  30752=>"000000000",
  30753=>"000000001",
  30754=>"111100000",
  30755=>"111011101",
  30756=>"010011010",
  30757=>"000100000",
  30758=>"101100000",
  30759=>"111111010",
  30760=>"111111111",
  30761=>"010010010",
  30762=>"111101111",
  30763=>"000100100",
  30764=>"101101101",
  30765=>"111111001",
  30766=>"111000000",
  30767=>"111111110",
  30768=>"101100000",
  30769=>"000000000",
  30770=>"100100100",
  30771=>"011111111",
  30772=>"000000000",
  30773=>"001011011",
  30774=>"111000000",
  30775=>"000000111",
  30776=>"001001000",
  30777=>"110110111",
  30778=>"111001000",
  30779=>"001000001",
  30780=>"111111111",
  30781=>"101101100",
  30782=>"100100000",
  30783=>"111111111",
  30784=>"000000000",
  30785=>"000000000",
  30786=>"000111111",
  30787=>"010011010",
  30788=>"111011000",
  30789=>"000000000",
  30790=>"000001000",
  30791=>"001000100",
  30792=>"110110110",
  30793=>"101000111",
  30794=>"011011010",
  30795=>"000000001",
  30796=>"100000000",
  30797=>"000000111",
  30798=>"001000101",
  30799=>"101001111",
  30800=>"101001001",
  30801=>"111111101",
  30802=>"111001000",
  30803=>"101001000",
  30804=>"000000000",
  30805=>"110110110",
  30806=>"111100000",
  30807=>"111111111",
  30808=>"000000000",
  30809=>"001001001",
  30810=>"000000110",
  30811=>"011000100",
  30812=>"000000000",
  30813=>"001000000",
  30814=>"010010110",
  30815=>"111011010",
  30816=>"110010000",
  30817=>"100100100",
  30818=>"001100101",
  30819=>"001000001",
  30820=>"000000000",
  30821=>"010000000",
  30822=>"110110000",
  30823=>"010110111",
  30824=>"000000111",
  30825=>"111101000",
  30826=>"000110111",
  30827=>"110111111",
  30828=>"011011011",
  30829=>"001000000",
  30830=>"100111111",
  30831=>"000000010",
  30832=>"001111110",
  30833=>"001001001",
  30834=>"101100100",
  30835=>"110000011",
  30836=>"011000000",
  30837=>"110110110",
  30838=>"110100011",
  30839=>"111101101",
  30840=>"000000001",
  30841=>"110110111",
  30842=>"010000000",
  30843=>"000000000",
  30844=>"100100100",
  30845=>"110010000",
  30846=>"010000000",
  30847=>"111111111",
  30848=>"111011000",
  30849=>"100110110",
  30850=>"011011111",
  30851=>"011101101",
  30852=>"011111111",
  30853=>"100001111",
  30854=>"111111000",
  30855=>"111111010",
  30856=>"010011011",
  30857=>"000000001",
  30858=>"100000000",
  30859=>"000011010",
  30860=>"000000010",
  30861=>"110100000",
  30862=>"001001001",
  30863=>"001001001",
  30864=>"111111111",
  30865=>"001000000",
  30866=>"011001001",
  30867=>"000000001",
  30868=>"010010010",
  30869=>"011111011",
  30870=>"000000100",
  30871=>"111111111",
  30872=>"001001001",
  30873=>"011011011",
  30874=>"000000000",
  30875=>"000000111",
  30876=>"010000010",
  30877=>"001000101",
  30878=>"110110110",
  30879=>"000000000",
  30880=>"011110010",
  30881=>"111111001",
  30882=>"000000000",
  30883=>"111111111",
  30884=>"000000001",
  30885=>"110111111",
  30886=>"111111110",
  30887=>"000000000",
  30888=>"001100100",
  30889=>"000101101",
  30890=>"000010111",
  30891=>"111011111",
  30892=>"100000000",
  30893=>"110110110",
  30894=>"000101101",
  30895=>"111111001",
  30896=>"000111111",
  30897=>"000001000",
  30898=>"111111111",
  30899=>"000000010",
  30900=>"000000111",
  30901=>"100110000",
  30902=>"000000110",
  30903=>"000000111",
  30904=>"001011111",
  30905=>"000000000",
  30906=>"100000001",
  30907=>"111110111",
  30908=>"001001001",
  30909=>"001000000",
  30910=>"000000000",
  30911=>"110111110",
  30912=>"000000000",
  30913=>"001000000",
  30914=>"111111111",
  30915=>"000101111",
  30916=>"011111100",
  30917=>"111111111",
  30918=>"000000000",
  30919=>"000100000",
  30920=>"001101101",
  30921=>"001000000",
  30922=>"111101101",
  30923=>"001000001",
  30924=>"110111100",
  30925=>"111111101",
  30926=>"110001001",
  30927=>"000000000",
  30928=>"111010111",
  30929=>"101101101",
  30930=>"011010011",
  30931=>"100100100",
  30932=>"111111111",
  30933=>"000001001",
  30934=>"000000000",
  30935=>"010000111",
  30936=>"110110110",
  30937=>"000100011",
  30938=>"000000101",
  30939=>"110111111",
  30940=>"000000011",
  30941=>"110111110",
  30942=>"111111110",
  30943=>"100100101",
  30944=>"000001001",
  30945=>"101001000",
  30946=>"101001001",
  30947=>"110110010",
  30948=>"110000000",
  30949=>"100100100",
  30950=>"000000000",
  30951=>"111001000",
  30952=>"111101000",
  30953=>"111101101",
  30954=>"111000000",
  30955=>"000000000",
  30956=>"111101101",
  30957=>"001111111",
  30958=>"111100001",
  30959=>"000000000",
  30960=>"011000001",
  30961=>"100100000",
  30962=>"000000100",
  30963=>"111111010",
  30964=>"011011001",
  30965=>"111111100",
  30966=>"011011011",
  30967=>"100000011",
  30968=>"111111111",
  30969=>"100100001",
  30970=>"000000001",
  30971=>"001001111",
  30972=>"111111100",
  30973=>"001001001",
  30974=>"110100000",
  30975=>"111111111",
  30976=>"000000000",
  30977=>"001001001",
  30978=>"111111000",
  30979=>"011000000",
  30980=>"101000000",
  30981=>"000001111",
  30982=>"111111101",
  30983=>"110111111",
  30984=>"110110110",
  30985=>"111101001",
  30986=>"101001101",
  30987=>"000000100",
  30988=>"001001001",
  30989=>"111000000",
  30990=>"111111111",
  30991=>"111001000",
  30992=>"111001011",
  30993=>"110110111",
  30994=>"001001000",
  30995=>"110100100",
  30996=>"000000000",
  30997=>"001011111",
  30998=>"110100100",
  30999=>"000000101",
  31000=>"001001001",
  31001=>"111111011",
  31002=>"111111111",
  31003=>"001001111",
  31004=>"001011011",
  31005=>"010011111",
  31006=>"111101001",
  31007=>"001001111",
  31008=>"001001000",
  31009=>"000100100",
  31010=>"111010111",
  31011=>"011011011",
  31012=>"111111111",
  31013=>"001000000",
  31014=>"101100000",
  31015=>"000000111",
  31016=>"101001000",
  31017=>"000000100",
  31018=>"101100111",
  31019=>"101101000",
  31020=>"001000000",
  31021=>"000001000",
  31022=>"111001111",
  31023=>"000100111",
  31024=>"100111110",
  31025=>"111001110",
  31026=>"001000000",
  31027=>"000000010",
  31028=>"011001011",
  31029=>"100111101",
  31030=>"010010010",
  31031=>"000000000",
  31032=>"100101111",
  31033=>"100110111",
  31034=>"000000000",
  31035=>"111010000",
  31036=>"000010111",
  31037=>"100110101",
  31038=>"111110110",
  31039=>"111100000",
  31040=>"000101101",
  31041=>"101101101",
  31042=>"111111111",
  31043=>"000001001",
  31044=>"000100111",
  31045=>"000001001",
  31046=>"111110111",
  31047=>"000000101",
  31048=>"101101101",
  31049=>"011011011",
  31050=>"111100101",
  31051=>"001001011",
  31052=>"011001011",
  31053=>"010000001",
  31054=>"111110001",
  31055=>"011001001",
  31056=>"011011111",
  31057=>"000111111",
  31058=>"001010110",
  31059=>"110110110",
  31060=>"000101101",
  31061=>"001001001",
  31062=>"111111011",
  31063=>"111111000",
  31064=>"111111011",
  31065=>"111111000",
  31066=>"110001111",
  31067=>"000000111",
  31068=>"100000000",
  31069=>"011001001",
  31070=>"101001101",
  31071=>"110110111",
  31072=>"010010000",
  31073=>"000010000",
  31074=>"011011011",
  31075=>"111111000",
  31076=>"011011011",
  31077=>"001001101",
  31078=>"010010110",
  31079=>"110110110",
  31080=>"101101101",
  31081=>"000000000",
  31082=>"001001001",
  31083=>"101001000",
  31084=>"111111100",
  31085=>"101000011",
  31086=>"101001000",
  31087=>"000101101",
  31088=>"111111110",
  31089=>"000011111",
  31090=>"111010111",
  31091=>"100100100",
  31092=>"000000010",
  31093=>"000000000",
  31094=>"011111111",
  31095=>"111111111",
  31096=>"111000000",
  31097=>"011010110",
  31098=>"111110110",
  31099=>"010110110",
  31100=>"000000000",
  31101=>"100100000",
  31102=>"111111011",
  31103=>"000000101",
  31104=>"100000100",
  31105=>"100000000",
  31106=>"000000000",
  31107=>"101101001",
  31108=>"111011010",
  31109=>"000000000",
  31110=>"100100111",
  31111=>"001000000",
  31112=>"000000111",
  31113=>"001001000",
  31114=>"111111110",
  31115=>"000111111",
  31116=>"110111111",
  31117=>"110100110",
  31118=>"000000000",
  31119=>"111111111",
  31120=>"011111011",
  31121=>"111111000",
  31122=>"000011000",
  31123=>"111111111",
  31124=>"000111111",
  31125=>"010010000",
  31126=>"011001001",
  31127=>"100100101",
  31128=>"111111111",
  31129=>"111111101",
  31130=>"110110110",
  31131=>"111111111",
  31132=>"000000000",
  31133=>"000000011",
  31134=>"000000000",
  31135=>"101101001",
  31136=>"010010000",
  31137=>"100100111",
  31138=>"111111111",
  31139=>"000000000",
  31140=>"100000001",
  31141=>"010010111",
  31142=>"010010011",
  31143=>"111110110",
  31144=>"000100101",
  31145=>"010111001",
  31146=>"000000000",
  31147=>"000001000",
  31148=>"000000000",
  31149=>"110110110",
  31150=>"111111100",
  31151=>"111111000",
  31152=>"001001000",
  31153=>"000000111",
  31154=>"111001001",
  31155=>"000010110",
  31156=>"000000001",
  31157=>"111111111",
  31158=>"111001101",
  31159=>"011000010",
  31160=>"011111101",
  31161=>"010110111",
  31162=>"000001000",
  31163=>"001011011",
  31164=>"001101101",
  31165=>"110110100",
  31166=>"101101100",
  31167=>"100100101",
  31168=>"111110110",
  31169=>"001001111",
  31170=>"001001000",
  31171=>"010001011",
  31172=>"111000000",
  31173=>"010110111",
  31174=>"100110110",
  31175=>"101000000",
  31176=>"000111111",
  31177=>"011010000",
  31178=>"000000000",
  31179=>"111101001",
  31180=>"000000011",
  31181=>"001001000",
  31182=>"110110110",
  31183=>"001000000",
  31184=>"101001101",
  31185=>"000111101",
  31186=>"110110110",
  31187=>"001111001",
  31188=>"001110011",
  31189=>"001001000",
  31190=>"010111111",
  31191=>"101000100",
  31192=>"111111111",
  31193=>"011111100",
  31194=>"001011111",
  31195=>"000000010",
  31196=>"000001111",
  31197=>"001001000",
  31198=>"111001011",
  31199=>"101000000",
  31200=>"110111110",
  31201=>"101111001",
  31202=>"101100000",
  31203=>"111111111",
  31204=>"001010111",
  31205=>"010010010",
  31206=>"101001101",
  31207=>"010010010",
  31208=>"000100001",
  31209=>"111111111",
  31210=>"011111110",
  31211=>"001101111",
  31212=>"000000000",
  31213=>"011011011",
  31214=>"001101101",
  31215=>"011000100",
  31216=>"000000001",
  31217=>"000000100",
  31218=>"001101101",
  31219=>"000100101",
  31220=>"111110110",
  31221=>"011010010",
  31222=>"111111001",
  31223=>"110100000",
  31224=>"001001000",
  31225=>"001001001",
  31226=>"111111111",
  31227=>"000000001",
  31228=>"000000101",
  31229=>"010110010",
  31230=>"000000000",
  31231=>"000001001",
  31232=>"111111111",
  31233=>"111111000",
  31234=>"111111000",
  31235=>"111011111",
  31236=>"011111111",
  31237=>"000101101",
  31238=>"000000000",
  31239=>"111111111",
  31240=>"001111100",
  31241=>"111000001",
  31242=>"100100000",
  31243=>"110000000",
  31244=>"000010000",
  31245=>"100000000",
  31246=>"000100100",
  31247=>"000000000",
  31248=>"001001000",
  31249=>"000000111",
  31250=>"100110111",
  31251=>"111111111",
  31252=>"000100000",
  31253=>"100000000",
  31254=>"000000000",
  31255=>"111111111",
  31256=>"110111111",
  31257=>"011110001",
  31258=>"111111011",
  31259=>"111011010",
  31260=>"000000000",
  31261=>"000000000",
  31262=>"000000001",
  31263=>"000101111",
  31264=>"000000000",
  31265=>"001001111",
  31266=>"110000000",
  31267=>"111001000",
  31268=>"000000000",
  31269=>"000010011",
  31270=>"111111111",
  31271=>"111111111",
  31272=>"000000111",
  31273=>"000000000",
  31274=>"000000000",
  31275=>"000000000",
  31276=>"111111001",
  31277=>"111111111",
  31278=>"000000000",
  31279=>"000000000",
  31280=>"111111111",
  31281=>"000000000",
  31282=>"111111000",
  31283=>"000011111",
  31284=>"110110111",
  31285=>"001010000",
  31286=>"000000001",
  31287=>"001001111",
  31288=>"111000000",
  31289=>"010010110",
  31290=>"000000000",
  31291=>"111111111",
  31292=>"000110111",
  31293=>"111111111",
  31294=>"110100100",
  31295=>"111000000",
  31296=>"110111000",
  31297=>"000000001",
  31298=>"110111111",
  31299=>"111110111",
  31300=>"110100001",
  31301=>"000000000",
  31302=>"111111111",
  31303=>"000000000",
  31304=>"111111011",
  31305=>"000000000",
  31306=>"111111111",
  31307=>"000011011",
  31308=>"111111101",
  31309=>"110100110",
  31310=>"010000000",
  31311=>"000000111",
  31312=>"100000100",
  31313=>"000101111",
  31314=>"000001001",
  31315=>"001001111",
  31316=>"000000000",
  31317=>"000000000",
  31318=>"000100000",
  31319=>"111111111",
  31320=>"000000000",
  31321=>"000000000",
  31322=>"100000000",
  31323=>"111000110",
  31324=>"000010010",
  31325=>"111111111",
  31326=>"110110100",
  31327=>"111001000",
  31328=>"110110110",
  31329=>"010111011",
  31330=>"111000101",
  31331=>"010000000",
  31332=>"001000000",
  31333=>"110111111",
  31334=>"000000100",
  31335=>"111000100",
  31336=>"110000000",
  31337=>"110110111",
  31338=>"011011111",
  31339=>"100110000",
  31340=>"111111101",
  31341=>"000000000",
  31342=>"001001001",
  31343=>"101111111",
  31344=>"000100000",
  31345=>"111000111",
  31346=>"011010010",
  31347=>"001001000",
  31348=>"000000000",
  31349=>"111001101",
  31350=>"000000000",
  31351=>"000000000",
  31352=>"111111001",
  31353=>"110111111",
  31354=>"110111110",
  31355=>"000000000",
  31356=>"011011111",
  31357=>"111001111",
  31358=>"000000001",
  31359=>"000000000",
  31360=>"101000111",
  31361=>"000000000",
  31362=>"000000111",
  31363=>"111011011",
  31364=>"111111110",
  31365=>"111000000",
  31366=>"001010011",
  31367=>"111111110",
  31368=>"100000000",
  31369=>"111001000",
  31370=>"011000000",
  31371=>"010110110",
  31372=>"111111111",
  31373=>"110010000",
  31374=>"111111111",
  31375=>"000000000",
  31376=>"000000000",
  31377=>"000000000",
  31378=>"000000000",
  31379=>"001010010",
  31380=>"000000111",
  31381=>"111000111",
  31382=>"111111111",
  31383=>"000000000",
  31384=>"111101111",
  31385=>"000000100",
  31386=>"001000000",
  31387=>"000011001",
  31388=>"110011000",
  31389=>"000001001",
  31390=>"000001001",
  31391=>"000011111",
  31392=>"000000000",
  31393=>"000000000",
  31394=>"111111000",
  31395=>"000000000",
  31396=>"101111000",
  31397=>"110100000",
  31398=>"111111000",
  31399=>"100100111",
  31400=>"011001111",
  31401=>"000000001",
  31402=>"100001111",
  31403=>"111111111",
  31404=>"000000010",
  31405=>"000010000",
  31406=>"000000000",
  31407=>"000000100",
  31408=>"111111101",
  31409=>"011111000",
  31410=>"111111111",
  31411=>"111000000",
  31412=>"111101101",
  31413=>"111001001",
  31414=>"111011000",
  31415=>"000100010",
  31416=>"000000100",
  31417=>"111111000",
  31418=>"100111111",
  31419=>"110111111",
  31420=>"001001111",
  31421=>"111111111",
  31422=>"111111101",
  31423=>"000000000",
  31424=>"000000000",
  31425=>"111011001",
  31426=>"111111111",
  31427=>"011001011",
  31428=>"000000000",
  31429=>"000000000",
  31430=>"101001000",
  31431=>"000000000",
  31432=>"111111111",
  31433=>"001011111",
  31434=>"111111110",
  31435=>"111110000",
  31436=>"011010000",
  31437=>"111000111",
  31438=>"011111111",
  31439=>"111111000",
  31440=>"010111101",
  31441=>"101000000",
  31442=>"000000000",
  31443=>"000111011",
  31444=>"000000110",
  31445=>"111011111",
  31446=>"101101111",
  31447=>"111111111",
  31448=>"111011011",
  31449=>"011001001",
  31450=>"001000000",
  31451=>"011111111",
  31452=>"110000111",
  31453=>"000010111",
  31454=>"111111111",
  31455=>"000000000",
  31456=>"010110110",
  31457=>"000000010",
  31458=>"000000000",
  31459=>"011111001",
  31460=>"100111000",
  31461=>"111101111",
  31462=>"001000000",
  31463=>"100000000",
  31464=>"011001000",
  31465=>"001000000",
  31466=>"111111111",
  31467=>"111110111",
  31468=>"001000000",
  31469=>"111100111",
  31470=>"011000000",
  31471=>"101101000",
  31472=>"000000011",
  31473=>"100111111",
  31474=>"000000100",
  31475=>"110010111",
  31476=>"101000111",
  31477=>"111111111",
  31478=>"100100100",
  31479=>"000000000",
  31480=>"111100100",
  31481=>"000000000",
  31482=>"110000000",
  31483=>"100100110",
  31484=>"111101111",
  31485=>"111111001",
  31486=>"111111111",
  31487=>"000000000",
  31488=>"011001000",
  31489=>"111111011",
  31490=>"010000000",
  31491=>"000000100",
  31492=>"111111001",
  31493=>"001111001",
  31494=>"000000000",
  31495=>"000000000",
  31496=>"111111000",
  31497=>"010010111",
  31498=>"111111101",
  31499=>"111111111",
  31500=>"110111111",
  31501=>"000000001",
  31502=>"010011111",
  31503=>"000000000",
  31504=>"100100000",
  31505=>"011000000",
  31506=>"000000000",
  31507=>"111111101",
  31508=>"000000001",
  31509=>"000000111",
  31510=>"000010000",
  31511=>"111111111",
  31512=>"000000110",
  31513=>"001000110",
  31514=>"000000000",
  31515=>"111111111",
  31516=>"000001000",
  31517=>"000000000",
  31518=>"111111011",
  31519=>"111000000",
  31520=>"100100110",
  31521=>"000110110",
  31522=>"000000000",
  31523=>"111111111",
  31524=>"100000000",
  31525=>"111011111",
  31526=>"100000010",
  31527=>"000001001",
  31528=>"000000110",
  31529=>"011000000",
  31530=>"111111000",
  31531=>"110110011",
  31532=>"110111111",
  31533=>"111001011",
  31534=>"100000000",
  31535=>"001000001",
  31536=>"011111111",
  31537=>"110100111",
  31538=>"001000000",
  31539=>"111111111",
  31540=>"100000000",
  31541=>"000000001",
  31542=>"111111100",
  31543=>"100101000",
  31544=>"111111111",
  31545=>"111111111",
  31546=>"110111111",
  31547=>"111111001",
  31548=>"000000000",
  31549=>"010000110",
  31550=>"000010111",
  31551=>"000000000",
  31552=>"111111110",
  31553=>"100111101",
  31554=>"011111100",
  31555=>"000000000",
  31556=>"111000011",
  31557=>"001000000",
  31558=>"111111111",
  31559=>"000001111",
  31560=>"000000000",
  31561=>"000000000",
  31562=>"000000100",
  31563=>"110111011",
  31564=>"101101111",
  31565=>"011101111",
  31566=>"111111111",
  31567=>"100100100",
  31568=>"001001000",
  31569=>"000000100",
  31570=>"001111111",
  31571=>"000000111",
  31572=>"000000011",
  31573=>"110100100",
  31574=>"011011110",
  31575=>"011001011",
  31576=>"000000010",
  31577=>"000000000",
  31578=>"110110110",
  31579=>"011111111",
  31580=>"000111001",
  31581=>"110001111",
  31582=>"111101001",
  31583=>"001001111",
  31584=>"000111111",
  31585=>"111111111",
  31586=>"100100100",
  31587=>"000000000",
  31588=>"110111111",
  31589=>"001111111",
  31590=>"111111000",
  31591=>"110011111",
  31592=>"111111111",
  31593=>"011111000",
  31594=>"011010110",
  31595=>"100110000",
  31596=>"111011011",
  31597=>"111111111",
  31598=>"000000000",
  31599=>"011111011",
  31600=>"101000000",
  31601=>"000000000",
  31602=>"000011000",
  31603=>"111011000",
  31604=>"111111111",
  31605=>"111111101",
  31606=>"000000100",
  31607=>"010000000",
  31608=>"000110010",
  31609=>"111111000",
  31610=>"111111111",
  31611=>"000000110",
  31612=>"000000000",
  31613=>"110111111",
  31614=>"001001111",
  31615=>"000000000",
  31616=>"111111111",
  31617=>"010011000",
  31618=>"000000000",
  31619=>"000100000",
  31620=>"001000000",
  31621=>"000000000",
  31622=>"110000011",
  31623=>"111110111",
  31624=>"000000000",
  31625=>"000000000",
  31626=>"000000000",
  31627=>"000000000",
  31628=>"110111111",
  31629=>"011001000",
  31630=>"000000000",
  31631=>"010000110",
  31632=>"111111111",
  31633=>"111111011",
  31634=>"111010000",
  31635=>"000000000",
  31636=>"000100100",
  31637=>"000000000",
  31638=>"111111111",
  31639=>"100100111",
  31640=>"000000000",
  31641=>"011000000",
  31642=>"111111111",
  31643=>"111000000",
  31644=>"000000111",
  31645=>"111111000",
  31646=>"000000111",
  31647=>"000000000",
  31648=>"111100101",
  31649=>"111111111",
  31650=>"000011111",
  31651=>"111111111",
  31652=>"100000111",
  31653=>"000000000",
  31654=>"000000000",
  31655=>"000000000",
  31656=>"000000000",
  31657=>"110000000",
  31658=>"111001111",
  31659=>"000110111",
  31660=>"000000000",
  31661=>"011000000",
  31662=>"000001111",
  31663=>"111111111",
  31664=>"000001000",
  31665=>"110110000",
  31666=>"000000000",
  31667=>"111111001",
  31668=>"100001011",
  31669=>"010010101",
  31670=>"111111000",
  31671=>"001110111",
  31672=>"010110000",
  31673=>"100111111",
  31674=>"111100010",
  31675=>"111100100",
  31676=>"111111111",
  31677=>"100110111",
  31678=>"111110111",
  31679=>"111111111",
  31680=>"011011011",
  31681=>"000000101",
  31682=>"000000000",
  31683=>"111111011",
  31684=>"111110000",
  31685=>"111110011",
  31686=>"000011000",
  31687=>"110111111",
  31688=>"111001111",
  31689=>"111011000",
  31690=>"000001000",
  31691=>"111111010",
  31692=>"011000010",
  31693=>"101000000",
  31694=>"000000000",
  31695=>"111111001",
  31696=>"111111111",
  31697=>"100110110",
  31698=>"111111111",
  31699=>"000000000",
  31700=>"111111111",
  31701=>"111001000",
  31702=>"000000110",
  31703=>"011000000",
  31704=>"111111010",
  31705=>"000000000",
  31706=>"000111000",
  31707=>"111101100",
  31708=>"101100100",
  31709=>"111111111",
  31710=>"001011011",
  31711=>"001001001",
  31712=>"111111111",
  31713=>"111111110",
  31714=>"111111101",
  31715=>"111111111",
  31716=>"111111111",
  31717=>"100100011",
  31718=>"100000000",
  31719=>"101101111",
  31720=>"000000000",
  31721=>"111111111",
  31722=>"000000000",
  31723=>"111111111",
  31724=>"000100000",
  31725=>"110111111",
  31726=>"000000010",
  31727=>"111111000",
  31728=>"001011111",
  31729=>"000100100",
  31730=>"111100110",
  31731=>"110110100",
  31732=>"101001001",
  31733=>"111101111",
  31734=>"111111111",
  31735=>"000000001",
  31736=>"000000111",
  31737=>"101111000",
  31738=>"110110111",
  31739=>"111111111",
  31740=>"111100111",
  31741=>"110000010",
  31742=>"111010110",
  31743=>"000000000",
  31744=>"000000000",
  31745=>"000000101",
  31746=>"000000000",
  31747=>"000000000",
  31748=>"000000000",
  31749=>"110110111",
  31750=>"000110111",
  31751=>"111111000",
  31752=>"111111111",
  31753=>"110100000",
  31754=>"111111101",
  31755=>"011010010",
  31756=>"000100100",
  31757=>"111111000",
  31758=>"111010010",
  31759=>"111111000",
  31760=>"111000100",
  31761=>"111111111",
  31762=>"000000000",
  31763=>"110100111",
  31764=>"000000111",
  31765=>"000000000",
  31766=>"000110000",
  31767=>"000000100",
  31768=>"000001111",
  31769=>"000000000",
  31770=>"100111001",
  31771=>"000000000",
  31772=>"111111111",
  31773=>"111011111",
  31774=>"001011111",
  31775=>"111111101",
  31776=>"101101101",
  31777=>"111111111",
  31778=>"111111111",
  31779=>"000000001",
  31780=>"000010010",
  31781=>"011000000",
  31782=>"011111111",
  31783=>"000000100",
  31784=>"000000011",
  31785=>"000000111",
  31786=>"000000000",
  31787=>"000011000",
  31788=>"000010111",
  31789=>"101100110",
  31790=>"000000011",
  31791=>"000000111",
  31792=>"011111000",
  31793=>"111011110",
  31794=>"001011111",
  31795=>"011011010",
  31796=>"010000001",
  31797=>"111111001",
  31798=>"111111000",
  31799=>"111001001",
  31800=>"000111100",
  31801=>"000000111",
  31802=>"000000011",
  31803=>"000010010",
  31804=>"000000111",
  31805=>"110111110",
  31806=>"010110100",
  31807=>"111111111",
  31808=>"111111000",
  31809=>"110100101",
  31810=>"111000000",
  31811=>"000000000",
  31812=>"011011000",
  31813=>"111000100",
  31814=>"000000000",
  31815=>"111111111",
  31816=>"000000000",
  31817=>"000000011",
  31818=>"111010000",
  31819=>"111101111",
  31820=>"000000000",
  31821=>"001000000",
  31822=>"011000000",
  31823=>"000111111",
  31824=>"100110100",
  31825=>"111110000",
  31826=>"001111111",
  31827=>"111111110",
  31828=>"000000000",
  31829=>"000110011",
  31830=>"000111111",
  31831=>"000000111",
  31832=>"111111001",
  31833=>"000111011",
  31834=>"011011000",
  31835=>"111111111",
  31836=>"000000000",
  31837=>"101111111",
  31838=>"000000000",
  31839=>"110000110",
  31840=>"111000000",
  31841=>"101101001",
  31842=>"000000000",
  31843=>"111000000",
  31844=>"111001011",
  31845=>"111111001",
  31846=>"111111011",
  31847=>"111111111",
  31848=>"100000000",
  31849=>"000000000",
  31850=>"110110111",
  31851=>"000011111",
  31852=>"111111111",
  31853=>"111111111",
  31854=>"111010010",
  31855=>"100000000",
  31856=>"000010010",
  31857=>"000000000",
  31858=>"000000000",
  31859=>"111111111",
  31860=>"100000001",
  31861=>"100110000",
  31862=>"000001111",
  31863=>"000000001",
  31864=>"111000001",
  31865=>"110111011",
  31866=>"000111111",
  31867=>"000000000",
  31868=>"011011001",
  31869=>"100100100",
  31870=>"001111111",
  31871=>"000000101",
  31872=>"110000000",
  31873=>"000000000",
  31874=>"000111110",
  31875=>"111111000",
  31876=>"100101000",
  31877=>"111100100",
  31878=>"111001110",
  31879=>"001001000",
  31880=>"000000000",
  31881=>"111000000",
  31882=>"000000000",
  31883=>"000110010",
  31884=>"110000001",
  31885=>"000111111",
  31886=>"110000000",
  31887=>"000000000",
  31888=>"001001001",
  31889=>"111111101",
  31890=>"111000000",
  31891=>"111110000",
  31892=>"000100011",
  31893=>"000000000",
  31894=>"000000000",
  31895=>"000000111",
  31896=>"100111000",
  31897=>"011101100",
  31898=>"111111111",
  31899=>"111111000",
  31900=>"000000001",
  31901=>"100000101",
  31902=>"000110111",
  31903=>"001001000",
  31904=>"000000100",
  31905=>"010110000",
  31906=>"111111111",
  31907=>"111111110",
  31908=>"000000110",
  31909=>"111111111",
  31910=>"111110110",
  31911=>"111110100",
  31912=>"000011101",
  31913=>"111111011",
  31914=>"111100000",
  31915=>"000000000",
  31916=>"111000110",
  31917=>"001011011",
  31918=>"111111101",
  31919=>"000000011",
  31920=>"000111111",
  31921=>"001011111",
  31922=>"111011111",
  31923=>"000000101",
  31924=>"010000111",
  31925=>"100110111",
  31926=>"000000111",
  31927=>"110110000",
  31928=>"011000000",
  31929=>"000000111",
  31930=>"000000111",
  31931=>"110100000",
  31932=>"000000010",
  31933=>"000000100",
  31934=>"110100000",
  31935=>"111001001",
  31936=>"011111111",
  31937=>"110111111",
  31938=>"100110111",
  31939=>"111111111",
  31940=>"111111111",
  31941=>"000111111",
  31942=>"111111111",
  31943=>"000000101",
  31944=>"110111000",
  31945=>"000000001",
  31946=>"000000001",
  31947=>"000100000",
  31948=>"010010000",
  31949=>"111111100",
  31950=>"111110000",
  31951=>"000000110",
  31952=>"000000000",
  31953=>"100000010",
  31954=>"111111001",
  31955=>"000000000",
  31956=>"010010011",
  31957=>"111110000",
  31958=>"000000111",
  31959=>"111111011",
  31960=>"110111111",
  31961=>"110110111",
  31962=>"000111011",
  31963=>"000000111",
  31964=>"111101100",
  31965=>"000111111",
  31966=>"111001000",
  31967=>"000001001",
  31968=>"000000001",
  31969=>"111000110",
  31970=>"000000100",
  31971=>"111111110",
  31972=>"111000110",
  31973=>"111111111",
  31974=>"000000111",
  31975=>"001000000",
  31976=>"100000000",
  31977=>"001001111",
  31978=>"110000100",
  31979=>"111100101",
  31980=>"000011000",
  31981=>"010110000",
  31982=>"011111000",
  31983=>"110000000",
  31984=>"100101111",
  31985=>"000000011",
  31986=>"000110110",
  31987=>"000100000",
  31988=>"000000000",
  31989=>"011001000",
  31990=>"111111110",
  31991=>"001000000",
  31992=>"000000000",
  31993=>"100000111",
  31994=>"010111111",
  31995=>"111001111",
  31996=>"000000001",
  31997=>"000000001",
  31998=>"111111001",
  31999=>"000001111",
  32000=>"111111111",
  32001=>"001011110",
  32002=>"001111000",
  32003=>"110110110",
  32004=>"000000000",
  32005=>"110100000",
  32006=>"000101111",
  32007=>"000111000",
  32008=>"010000000",
  32009=>"101111111",
  32010=>"111111010",
  32011=>"110111110",
  32012=>"100100000",
  32013=>"001100100",
  32014=>"000000000",
  32015=>"110000000",
  32016=>"110101111",
  32017=>"000111111",
  32018=>"000000110",
  32019=>"000000100",
  32020=>"000000000",
  32021=>"111000111",
  32022=>"011011011",
  32023=>"101100111",
  32024=>"111000111",
  32025=>"011111111",
  32026=>"000111111",
  32027=>"110100100",
  32028=>"000111111",
  32029=>"000000000",
  32030=>"111111000",
  32031=>"000011001",
  32032=>"000111001",
  32033=>"011000000",
  32034=>"000000001",
  32035=>"011000000",
  32036=>"000010111",
  32037=>"000111111",
  32038=>"110111011",
  32039=>"110000111",
  32040=>"111000000",
  32041=>"000100100",
  32042=>"000000011",
  32043=>"011000101",
  32044=>"010111001",
  32045=>"100000111",
  32046=>"000000000",
  32047=>"011000000",
  32048=>"111111111",
  32049=>"111111111",
  32050=>"111111111",
  32051=>"011000111",
  32052=>"101111111",
  32053=>"111111000",
  32054=>"000001001",
  32055=>"100110110",
  32056=>"000000000",
  32057=>"111111000",
  32058=>"000000100",
  32059=>"111110110",
  32060=>"000110110",
  32061=>"000000000",
  32062=>"000000000",
  32063=>"111111111",
  32064=>"010000000",
  32065=>"111111011",
  32066=>"110100000",
  32067=>"001000000",
  32068=>"111101111",
  32069=>"000000000",
  32070=>"000000000",
  32071=>"001000000",
  32072=>"000001111",
  32073=>"110100000",
  32074=>"010110111",
  32075=>"110000000",
  32076=>"000000000",
  32077=>"101000000",
  32078=>"010101111",
  32079=>"000000000",
  32080=>"111111111",
  32081=>"110111111",
  32082=>"111111111",
  32083=>"110100111",
  32084=>"000010000",
  32085=>"111111101",
  32086=>"111111111",
  32087=>"000001000",
  32088=>"000000000",
  32089=>"110010000",
  32090=>"011010111",
  32091=>"111111011",
  32092=>"110110110",
  32093=>"101000000",
  32094=>"011100100",
  32095=>"111101001",
  32096=>"111111111",
  32097=>"001000000",
  32098=>"100101101",
  32099=>"011000000",
  32100=>"111111100",
  32101=>"000000100",
  32102=>"000011111",
  32103=>"000000010",
  32104=>"011001000",
  32105=>"000111011",
  32106=>"111111111",
  32107=>"110111111",
  32108=>"011110000",
  32109=>"110010001",
  32110=>"000000000",
  32111=>"000000000",
  32112=>"001001001",
  32113=>"111111111",
  32114=>"010000000",
  32115=>"111111011",
  32116=>"111000000",
  32117=>"111110111",
  32118=>"000000001",
  32119=>"111111111",
  32120=>"111111100",
  32121=>"000000000",
  32122=>"000111111",
  32123=>"111111111",
  32124=>"111000000",
  32125=>"100111111",
  32126=>"111111101",
  32127=>"000000111",
  32128=>"011011011",
  32129=>"000001001",
  32130=>"001000011",
  32131=>"000000000",
  32132=>"110111111",
  32133=>"000000000",
  32134=>"111000011",
  32135=>"001110110",
  32136=>"000000000",
  32137=>"100100101",
  32138=>"001000100",
  32139=>"010100000",
  32140=>"111111111",
  32141=>"110111000",
  32142=>"111011000",
  32143=>"000000000",
  32144=>"111111111",
  32145=>"000011001",
  32146=>"111110100",
  32147=>"001011011",
  32148=>"000000000",
  32149=>"000000000",
  32150=>"000000111",
  32151=>"001001000",
  32152=>"000000000",
  32153=>"111101111",
  32154=>"000111000",
  32155=>"101100110",
  32156=>"111111111",
  32157=>"111111111",
  32158=>"100000101",
  32159=>"000111111",
  32160=>"100101111",
  32161=>"011000100",
  32162=>"110110000",
  32163=>"000111111",
  32164=>"111111100",
  32165=>"001111111",
  32166=>"000000011",
  32167=>"111111011",
  32168=>"110000010",
  32169=>"111100111",
  32170=>"001000000",
  32171=>"000000000",
  32172=>"000000000",
  32173=>"000100000",
  32174=>"111011010",
  32175=>"101101100",
  32176=>"111111001",
  32177=>"100111111",
  32178=>"000100000",
  32179=>"000000000",
  32180=>"111111111",
  32181=>"000110001",
  32182=>"110000000",
  32183=>"111101111",
  32184=>"000000111",
  32185=>"100111000",
  32186=>"001001000",
  32187=>"000000110",
  32188=>"000000000",
  32189=>"100110100",
  32190=>"000010111",
  32191=>"000010011",
  32192=>"001000110",
  32193=>"100000000",
  32194=>"110000000",
  32195=>"000000111",
  32196=>"010110000",
  32197=>"111111011",
  32198=>"000100111",
  32199=>"111111010",
  32200=>"000000000",
  32201=>"001101111",
  32202=>"111101111",
  32203=>"000000000",
  32204=>"010000000",
  32205=>"110111110",
  32206=>"111111111",
  32207=>"111111111",
  32208=>"000000000",
  32209=>"010110000",
  32210=>"111000000",
  32211=>"111001001",
  32212=>"000111111",
  32213=>"000100111",
  32214=>"000000100",
  32215=>"000000011",
  32216=>"000010111",
  32217=>"111100100",
  32218=>"111001000",
  32219=>"100000000",
  32220=>"000000010",
  32221=>"010100101",
  32222=>"111001000",
  32223=>"001111011",
  32224=>"110110110",
  32225=>"011000110",
  32226=>"100000000",
  32227=>"000000000",
  32228=>"000111111",
  32229=>"111111111",
  32230=>"011000000",
  32231=>"000000011",
  32232=>"000000000",
  32233=>"111111111",
  32234=>"001001111",
  32235=>"111100001",
  32236=>"000000111",
  32237=>"110100110",
  32238=>"011000000",
  32239=>"111111011",
  32240=>"001000011",
  32241=>"111000000",
  32242=>"011001011",
  32243=>"111100100",
  32244=>"000010010",
  32245=>"000001001",
  32246=>"000111111",
  32247=>"111110000",
  32248=>"111110110",
  32249=>"100100100",
  32250=>"111111111",
  32251=>"000000100",
  32252=>"111111111",
  32253=>"111111000",
  32254=>"010111111",
  32255=>"111111111",
  32256=>"000001001",
  32257=>"000000001",
  32258=>"010000111",
  32259=>"111111111",
  32260=>"111110100",
  32261=>"111111011",
  32262=>"100000000",
  32263=>"011011111",
  32264=>"000100110",
  32265=>"100011111",
  32266=>"111110100",
  32267=>"000000011",
  32268=>"110110110",
  32269=>"111111111",
  32270=>"111111011",
  32271=>"111001000",
  32272=>"000000111",
  32273=>"111110111",
  32274=>"000001000",
  32275=>"011011011",
  32276=>"000111111",
  32277=>"000100111",
  32278=>"111010000",
  32279=>"111111111",
  32280=>"111011111",
  32281=>"101101101",
  32282=>"000001111",
  32283=>"000001011",
  32284=>"111111001",
  32285=>"110000000",
  32286=>"111010110",
  32287=>"111000000",
  32288=>"101100111",
  32289=>"111100110",
  32290=>"111001000",
  32291=>"111011000",
  32292=>"110000000",
  32293=>"111001110",
  32294=>"111000000",
  32295=>"000111111",
  32296=>"111111111",
  32297=>"010111111",
  32298=>"001000111",
  32299=>"011010000",
  32300=>"100111111",
  32301=>"111111111",
  32302=>"111000000",
  32303=>"001001011",
  32304=>"001000000",
  32305=>"111001000",
  32306=>"011000011",
  32307=>"000110110",
  32308=>"101000000",
  32309=>"011001000",
  32310=>"000000000",
  32311=>"001000001",
  32312=>"111110100",
  32313=>"111110111",
  32314=>"000000000",
  32315=>"111110111",
  32316=>"011000000",
  32317=>"110000100",
  32318=>"111111111",
  32319=>"000000000",
  32320=>"000000000",
  32321=>"000011010",
  32322=>"110001111",
  32323=>"000000000",
  32324=>"001000000",
  32325=>"100110000",
  32326=>"100100111",
  32327=>"111111101",
  32328=>"000000000",
  32329=>"000000001",
  32330=>"000000111",
  32331=>"001101111",
  32332=>"111111001",
  32333=>"001011111",
  32334=>"010010111",
  32335=>"111111111",
  32336=>"000011001",
  32337=>"110000100",
  32338=>"001001111",
  32339=>"101101110",
  32340=>"111111011",
  32341=>"110000000",
  32342=>"111100000",
  32343=>"111000000",
  32344=>"110110000",
  32345=>"000100100",
  32346=>"000000000",
  32347=>"111010000",
  32348=>"111111101",
  32349=>"010111010",
  32350=>"111111000",
  32351=>"111000101",
  32352=>"000000000",
  32353=>"000111111",
  32354=>"000000000",
  32355=>"101101001",
  32356=>"000000100",
  32357=>"000100101",
  32358=>"010000111",
  32359=>"100101111",
  32360=>"111111100",
  32361=>"111111110",
  32362=>"000000000",
  32363=>"111010000",
  32364=>"000000000",
  32365=>"000000000",
  32366=>"111111111",
  32367=>"111000000",
  32368=>"000000011",
  32369=>"000011111",
  32370=>"000000000",
  32371=>"100111111",
  32372=>"001001000",
  32373=>"000000000",
  32374=>"000111111",
  32375=>"000010111",
  32376=>"000111111",
  32377=>"000000011",
  32378=>"111000100",
  32379=>"000111111",
  32380=>"011011111",
  32381=>"110000010",
  32382=>"111110000",
  32383=>"111111111",
  32384=>"111111100",
  32385=>"010111111",
  32386=>"110111111",
  32387=>"011001000",
  32388=>"010000000",
  32389=>"000000110",
  32390=>"111111101",
  32391=>"111111111",
  32392=>"110100000",
  32393=>"000000001",
  32394=>"111111000",
  32395=>"000000011",
  32396=>"100100100",
  32397=>"111011000",
  32398=>"010001001",
  32399=>"000001101",
  32400=>"000000111",
  32401=>"101101101",
  32402=>"111101001",
  32403=>"001001111",
  32404=>"111100100",
  32405=>"101000111",
  32406=>"111111000",
  32407=>"110110111",
  32408=>"111111110",
  32409=>"001000000",
  32410=>"111000000",
  32411=>"011000000",
  32412=>"000000001",
  32413=>"000001111",
  32414=>"111011000",
  32415=>"000000000",
  32416=>"110111011",
  32417=>"000111111",
  32418=>"000000001",
  32419=>"101000001",
  32420=>"111111111",
  32421=>"110100000",
  32422=>"000011111",
  32423=>"111111000",
  32424=>"110000111",
  32425=>"000000111",
  32426=>"000000000",
  32427=>"000000100",
  32428=>"011011001",
  32429=>"000000001",
  32430=>"000100110",
  32431=>"101111011",
  32432=>"000000000",
  32433=>"011011001",
  32434=>"000001001",
  32435=>"111111111",
  32436=>"111100100",
  32437=>"000000000",
  32438=>"111000001",
  32439=>"000000000",
  32440=>"111100110",
  32441=>"011111000",
  32442=>"101100011",
  32443=>"110100001",
  32444=>"000010000",
  32445=>"000000000",
  32446=>"110100000",
  32447=>"000000001",
  32448=>"000000001",
  32449=>"111110100",
  32450=>"100100111",
  32451=>"010111000",
  32452=>"111100100",
  32453=>"000000111",
  32454=>"000000000",
  32455=>"101111111",
  32456=>"000001001",
  32457=>"111111100",
  32458=>"000001011",
  32459=>"111111111",
  32460=>"010111111",
  32461=>"100110100",
  32462=>"111011001",
  32463=>"011100011",
  32464=>"111110001",
  32465=>"001001011",
  32466=>"000000000",
  32467=>"011001000",
  32468=>"111111000",
  32469=>"101111111",
  32470=>"000111111",
  32471=>"000001011",
  32472=>"000000111",
  32473=>"111111111",
  32474=>"000111110",
  32475=>"111000000",
  32476=>"111101001",
  32477=>"010000111",
  32478=>"000000000",
  32479=>"000000000",
  32480=>"000110110",
  32481=>"000111111",
  32482=>"000000000",
  32483=>"111101000",
  32484=>"110000000",
  32485=>"111100101",
  32486=>"110000001",
  32487=>"110111111",
  32488=>"000000110",
  32489=>"000001111",
  32490=>"111111001",
  32491=>"110010011",
  32492=>"100110100",
  32493=>"000111111",
  32494=>"111100110",
  32495=>"111100111",
  32496=>"101101111",
  32497=>"101101111",
  32498=>"000000000",
  32499=>"110110011",
  32500=>"111011001",
  32501=>"111111000",
  32502=>"000001000",
  32503=>"111110100",
  32504=>"000111111",
  32505=>"111000000",
  32506=>"011111001",
  32507=>"110110110",
  32508=>"111111000",
  32509=>"001000000",
  32510=>"011111000",
  32511=>"000000001",
  32512=>"000000110",
  32513=>"001111010",
  32514=>"111111111",
  32515=>"000000000",
  32516=>"001100101",
  32517=>"000000000",
  32518=>"000000011",
  32519=>"000011101",
  32520=>"110110111",
  32521=>"111111000",
  32522=>"111110000",
  32523=>"111111011",
  32524=>"000000110",
  32525=>"100101000",
  32526=>"111100100",
  32527=>"111110000",
  32528=>"000000000",
  32529=>"110100000",
  32530=>"111000000",
  32531=>"111000000",
  32532=>"000000000",
  32533=>"000100100",
  32534=>"011001001",
  32535=>"001101011",
  32536=>"111111001",
  32537=>"000111111",
  32538=>"000000001",
  32539=>"000000000",
  32540=>"001001000",
  32541=>"111110001",
  32542=>"000000000",
  32543=>"111111001",
  32544=>"110100110",
  32545=>"111111111",
  32546=>"000011000",
  32547=>"110100011",
  32548=>"000011111",
  32549=>"000000000",
  32550=>"110111010",
  32551=>"010111111",
  32552=>"111100000",
  32553=>"000001000",
  32554=>"110111111",
  32555=>"000000100",
  32556=>"111111000",
  32557=>"000101111",
  32558=>"000000111",
  32559=>"000000000",
  32560=>"111111111",
  32561=>"111111111",
  32562=>"010000000",
  32563=>"000000111",
  32564=>"110110110",
  32565=>"000110111",
  32566=>"000000001",
  32567=>"100110110",
  32568=>"000111100",
  32569=>"110110111",
  32570=>"101001001",
  32571=>"000000000",
  32572=>"100110111",
  32573=>"000000111",
  32574=>"111111101",
  32575=>"111000001",
  32576=>"000000000",
  32577=>"001001001",
  32578=>"000001000",
  32579=>"000000110",
  32580=>"101001111",
  32581=>"100111111",
  32582=>"111000000",
  32583=>"000000001",
  32584=>"000111001",
  32585=>"111100101",
  32586=>"111110000",
  32587=>"011111111",
  32588=>"000000000",
  32589=>"000100110",
  32590=>"111111001",
  32591=>"000001111",
  32592=>"111001001",
  32593=>"111111110",
  32594=>"000001000",
  32595=>"111110111",
  32596=>"001000000",
  32597=>"111111111",
  32598=>"110000000",
  32599=>"010011111",
  32600=>"001001111",
  32601=>"001011111",
  32602=>"111111011",
  32603=>"000111111",
  32604=>"000111110",
  32605=>"101111111",
  32606=>"000000111",
  32607=>"001111000",
  32608=>"001101111",
  32609=>"000000110",
  32610=>"001001011",
  32611=>"000011111",
  32612=>"111100000",
  32613=>"111100110",
  32614=>"100111111",
  32615=>"011000111",
  32616=>"000110110",
  32617=>"011000011",
  32618=>"111111111",
  32619=>"000001001",
  32620=>"101000100",
  32621=>"010000000",
  32622=>"000000001",
  32623=>"111001000",
  32624=>"001001011",
  32625=>"001001011",
  32626=>"000000001",
  32627=>"100101100",
  32628=>"001000111",
  32629=>"000000011",
  32630=>"001100111",
  32631=>"111001100",
  32632=>"011000111",
  32633=>"000100111",
  32634=>"010011011",
  32635=>"111000000",
  32636=>"101001101",
  32637=>"101110000",
  32638=>"111110000",
  32639=>"111111100",
  32640=>"110010000",
  32641=>"111011001",
  32642=>"011011001",
  32643=>"000001001",
  32644=>"000000000",
  32645=>"110110110",
  32646=>"111001001",
  32647=>"100111111",
  32648=>"110111111",
  32649=>"001111011",
  32650=>"110000011",
  32651=>"000000110",
  32652=>"101111111",
  32653=>"000000110",
  32654=>"000000000",
  32655=>"011001000",
  32656=>"111110000",
  32657=>"111111000",
  32658=>"000000100",
  32659=>"011101101",
  32660=>"000100110",
  32661=>"000000010",
  32662=>"100000000",
  32663=>"001001111",
  32664=>"000010110",
  32665=>"111001001",
  32666=>"000000011",
  32667=>"001000000",
  32668=>"000000111",
  32669=>"000111111",
  32670=>"001000000",
  32671=>"000001100",
  32672=>"101001000",
  32673=>"000000110",
  32674=>"110110011",
  32675=>"011111111",
  32676=>"000000000",
  32677=>"111101100",
  32678=>"100111111",
  32679=>"000000000",
  32680=>"110100000",
  32681=>"000001011",
  32682=>"000110111",
  32683=>"111100000",
  32684=>"110110111",
  32685=>"100000000",
  32686=>"000111001",
  32687=>"111111111",
  32688=>"000111000",
  32689=>"111110100",
  32690=>"100000000",
  32691=>"010000000",
  32692=>"110101001",
  32693=>"111110111",
  32694=>"000100111",
  32695=>"110000000",
  32696=>"000000111",
  32697=>"111111111",
  32698=>"111111101",
  32699=>"000110110",
  32700=>"011111000",
  32701=>"111111111",
  32702=>"011000000",
  32703=>"000010000",
  32704=>"110111001",
  32705=>"000000111",
  32706=>"000000111",
  32707=>"111111001",
  32708=>"111110111",
  32709=>"001011011",
  32710=>"000000111",
  32711=>"100100000",
  32712=>"010110110",
  32713=>"110010000",
  32714=>"111011111",
  32715=>"010010000",
  32716=>"010111100",
  32717=>"111111011",
  32718=>"111010000",
  32719=>"111000111",
  32720=>"000111111",
  32721=>"110110111",
  32722=>"000000000",
  32723=>"111111101",
  32724=>"110001001",
  32725=>"000000001",
  32726=>"111000000",
  32727=>"000000000",
  32728=>"000000001",
  32729=>"111011000",
  32730=>"101101111",
  32731=>"000000000",
  32732=>"001000000",
  32733=>"101111111",
  32734=>"111110111",
  32735=>"110000000",
  32736=>"100000111",
  32737=>"000000111",
  32738=>"000111010",
  32739=>"011000100",
  32740=>"001001001",
  32741=>"100100110",
  32742=>"000000101",
  32743=>"000101111",
  32744=>"111011001",
  32745=>"000110111",
  32746=>"000111111",
  32747=>"111000000",
  32748=>"000001101",
  32749=>"111000100",
  32750=>"000000110",
  32751=>"111011011",
  32752=>"111100001",
  32753=>"000001001",
  32754=>"111111111",
  32755=>"001000000",
  32756=>"111110000",
  32757=>"001111111",
  32758=>"000010011",
  32759=>"100000001",
  32760=>"000010000",
  32761=>"100000001",
  32762=>"110011001",
  32763=>"000000000",
  32764=>"001001000",
  32765=>"101111111",
  32766=>"000000000",
  32767=>"000000001",
  32768=>"111011001",
  32769=>"000110111",
  32770=>"111111111",
  32771=>"111111111",
  32772=>"010001000",
  32773=>"000011010",
  32774=>"000000000",
  32775=>"111111111",
  32776=>"111111000",
  32777=>"111101101",
  32778=>"111111111",
  32779=>"111111111",
  32780=>"011011000",
  32781=>"001001000",
  32782=>"111101111",
  32783=>"000000000",
  32784=>"100100000",
  32785=>"000000111",
  32786=>"000011011",
  32787=>"111111000",
  32788=>"000000000",
  32789=>"001001000",
  32790=>"000011000",
  32791=>"100000000",
  32792=>"011000000",
  32793=>"111111110",
  32794=>"000000000",
  32795=>"001111011",
  32796=>"111111110",
  32797=>"000000000",
  32798=>"110111010",
  32799=>"011000000",
  32800=>"110000010",
  32801=>"000110111",
  32802=>"000100110",
  32803=>"111111111",
  32804=>"000000001",
  32805=>"000111110",
  32806=>"111110010",
  32807=>"000011000",
  32808=>"110000111",
  32809=>"000000111",
  32810=>"000101000",
  32811=>"011011000",
  32812=>"111111111",
  32813=>"000111000",
  32814=>"000111111",
  32815=>"001000100",
  32816=>"111110000",
  32817=>"000000000",
  32818=>"100100100",
  32819=>"000111011",
  32820=>"100111101",
  32821=>"111011110",
  32822=>"011011000",
  32823=>"000011111",
  32824=>"000011011",
  32825=>"111001001",
  32826=>"000000001",
  32827=>"111000000",
  32828=>"111111111",
  32829=>"111011001",
  32830=>"110000000",
  32831=>"000101111",
  32832=>"111100000",
  32833=>"000000000",
  32834=>"000001111",
  32835=>"111110111",
  32836=>"011000110",
  32837=>"011011000",
  32838=>"000000000",
  32839=>"000000000",
  32840=>"110110000",
  32841=>"111101001",
  32842=>"101111101",
  32843=>"001000000",
  32844=>"111111111",
  32845=>"111000000",
  32846=>"111000000",
  32847=>"111101001",
  32848=>"110000000",
  32849=>"000010110",
  32850=>"111111111",
  32851=>"000000100",
  32852=>"000000001",
  32853=>"100000000",
  32854=>"001111111",
  32855=>"111111000",
  32856=>"000000000",
  32857=>"111011001",
  32858=>"000111001",
  32859=>"000000000",
  32860=>"000111111",
  32861=>"111110111",
  32862=>"111111111",
  32863=>"111000001",
  32864=>"011110111",
  32865=>"110111000",
  32866=>"000111111",
  32867=>"000110000",
  32868=>"111010000",
  32869=>"000010111",
  32870=>"000101111",
  32871=>"000011111",
  32872=>"000000000",
  32873=>"111111000",
  32874=>"001111010",
  32875=>"111101111",
  32876=>"011111111",
  32877=>"111000110",
  32878=>"111101101",
  32879=>"000000100",
  32880=>"001001011",
  32881=>"000110110",
  32882=>"111011001",
  32883=>"111111111",
  32884=>"000000001",
  32885=>"111111000",
  32886=>"011111111",
  32887=>"111010000",
  32888=>"100000000",
  32889=>"000000110",
  32890=>"000000000",
  32891=>"000000000",
  32892=>"111111111",
  32893=>"110111000",
  32894=>"111000000",
  32895=>"111000000",
  32896=>"111010000",
  32897=>"000111111",
  32898=>"111011011",
  32899=>"100111111",
  32900=>"100100111",
  32901=>"111111000",
  32902=>"111000100",
  32903=>"010111111",
  32904=>"000000111",
  32905=>"111101000",
  32906=>"011000000",
  32907=>"111000011",
  32908=>"111000101",
  32909=>"000000000",
  32910=>"000111111",
  32911=>"111111111",
  32912=>"001111101",
  32913=>"111111000",
  32914=>"100111111",
  32915=>"111000111",
  32916=>"001000000",
  32917=>"000000111",
  32918=>"111111100",
  32919=>"111000000",
  32920=>"100100000",
  32921=>"110000000",
  32922=>"000000111",
  32923=>"111000000",
  32924=>"111100111",
  32925=>"000111111",
  32926=>"001111111",
  32927=>"000000000",
  32928=>"111111111",
  32929=>"111001000",
  32930=>"000011111",
  32931=>"111111000",
  32932=>"100000000",
  32933=>"111111100",
  32934=>"001111110",
  32935=>"011111011",
  32936=>"110111000",
  32937=>"000000000",
  32938=>"000000111",
  32939=>"000111111",
  32940=>"100101000",
  32941=>"000110111",
  32942=>"111111110",
  32943=>"111000101",
  32944=>"000000111",
  32945=>"011011011",
  32946=>"111111111",
  32947=>"111000000",
  32948=>"111001000",
  32949=>"000001000",
  32950=>"000000001",
  32951=>"000000111",
  32952=>"111110100",
  32953=>"111000000",
  32954=>"001000000",
  32955=>"100000111",
  32956=>"111110111",
  32957=>"011000000",
  32958=>"111111111",
  32959=>"111111010",
  32960=>"111000111",
  32961=>"000110000",
  32962=>"000010011",
  32963=>"111111110",
  32964=>"110111111",
  32965=>"011111111",
  32966=>"010111011",
  32967=>"110111111",
  32968=>"111111111",
  32969=>"111011111",
  32970=>"110000000",
  32971=>"110000001",
  32972=>"001001001",
  32973=>"111111010",
  32974=>"000000000",
  32975=>"000110110",
  32976=>"110000000",
  32977=>"000110111",
  32978=>"000000111",
  32979=>"000000111",
  32980=>"110111000",
  32981=>"001001111",
  32982=>"111111111",
  32983=>"011010111",
  32984=>"111101000",
  32985=>"111111111",
  32986=>"111111011",
  32987=>"111000110",
  32988=>"111101101",
  32989=>"111011001",
  32990=>"010111111",
  32991=>"100000111",
  32992=>"000000000",
  32993=>"000000000",
  32994=>"101111001",
  32995=>"000000011",
  32996=>"010111111",
  32997=>"000000000",
  32998=>"100100000",
  32999=>"111110000",
  33000=>"111111111",
  33001=>"100000000",
  33002=>"000000100",
  33003=>"000101001",
  33004=>"001000000",
  33005=>"001111111",
  33006=>"000000111",
  33007=>"110000000",
  33008=>"111111000",
  33009=>"111111011",
  33010=>"001111101",
  33011=>"000011111",
  33012=>"100111110",
  33013=>"111000101",
  33014=>"101110111",
  33015=>"000000000",
  33016=>"000000111",
  33017=>"000101000",
  33018=>"111111110",
  33019=>"001111010",
  33020=>"111011000",
  33021=>"001001111",
  33022=>"000000001",
  33023=>"011011001",
  33024=>"010000010",
  33025=>"011011001",
  33026=>"000111111",
  33027=>"111000000",
  33028=>"000000000",
  33029=>"111111111",
  33030=>"000111111",
  33031=>"000000111",
  33032=>"000111111",
  33033=>"000000000",
  33034=>"110000001",
  33035=>"000000111",
  33036=>"000000101",
  33037=>"010010010",
  33038=>"111011000",
  33039=>"111111111",
  33040=>"000111011",
  33041=>"000000000",
  33042=>"110100000",
  33043=>"000010111",
  33044=>"001000000",
  33045=>"111111000",
  33046=>"000000101",
  33047=>"100000000",
  33048=>"111111000",
  33049=>"111111000",
  33050=>"100101001",
  33051=>"011000000",
  33052=>"111111100",
  33053=>"111111111",
  33054=>"000000001",
  33055=>"000111111",
  33056=>"100111111",
  33057=>"011000000",
  33058=>"000111111",
  33059=>"000100111",
  33060=>"000011111",
  33061=>"111000000",
  33062=>"110011001",
  33063=>"100000000",
  33064=>"100011001",
  33065=>"000000000",
  33066=>"111101000",
  33067=>"111111111",
  33068=>"110000000",
  33069=>"000111011",
  33070=>"000010000",
  33071=>"100111111",
  33072=>"000011111",
  33073=>"111010000",
  33074=>"000111111",
  33075=>"000000000",
  33076=>"111101111",
  33077=>"110000001",
  33078=>"100001111",
  33079=>"000000000",
  33080=>"000110011",
  33081=>"111110010",
  33082=>"000000000",
  33083=>"111111111",
  33084=>"000111111",
  33085=>"000000000",
  33086=>"000111110",
  33087=>"000000000",
  33088=>"000000000",
  33089=>"000000111",
  33090=>"000000000",
  33091=>"110010000",
  33092=>"111011111",
  33093=>"000111111",
  33094=>"000000000",
  33095=>"000000000",
  33096=>"000000111",
  33097=>"000000000",
  33098=>"100000000",
  33099=>"101101011",
  33100=>"100000000",
  33101=>"111000000",
  33102=>"000000000",
  33103=>"111111100",
  33104=>"000111111",
  33105=>"111000000",
  33106=>"111000000",
  33107=>"111100000",
  33108=>"100000000",
  33109=>"011011011",
  33110=>"011000010",
  33111=>"111111111",
  33112=>"000000000",
  33113=>"111011000",
  33114=>"000000110",
  33115=>"000000111",
  33116=>"000000000",
  33117=>"000000000",
  33118=>"000000000",
  33119=>"100101111",
  33120=>"001001000",
  33121=>"010111111",
  33122=>"111011000",
  33123=>"100000000",
  33124=>"111111111",
  33125=>"000111111",
  33126=>"000100101",
  33127=>"000000000",
  33128=>"001101101",
  33129=>"100000000",
  33130=>"111111111",
  33131=>"111101000",
  33132=>"000111111",
  33133=>"001000000",
  33134=>"111111001",
  33135=>"000000000",
  33136=>"100111111",
  33137=>"000011111",
  33138=>"111000100",
  33139=>"000011000",
  33140=>"111111111",
  33141=>"111100000",
  33142=>"100111111",
  33143=>"000000000",
  33144=>"111011000",
  33145=>"000100110",
  33146=>"000111111",
  33147=>"000101111",
  33148=>"001000111",
  33149=>"011000000",
  33150=>"100000111",
  33151=>"000111100",
  33152=>"111000000",
  33153=>"111111000",
  33154=>"100110000",
  33155=>"001000000",
  33156=>"000000000",
  33157=>"000000000",
  33158=>"100000000",
  33159=>"111001101",
  33160=>"111000011",
  33161=>"000000011",
  33162=>"111010001",
  33163=>"000000101",
  33164=>"000001111",
  33165=>"111000000",
  33166=>"000000001",
  33167=>"111111111",
  33168=>"000000000",
  33169=>"001000000",
  33170=>"111111101",
  33171=>"000111111",
  33172=>"111101001",
  33173=>"010010000",
  33174=>"010010011",
  33175=>"110110110",
  33176=>"011111111",
  33177=>"000011011",
  33178=>"111011001",
  33179=>"110110100",
  33180=>"000000000",
  33181=>"000000010",
  33182=>"000000000",
  33183=>"000100110",
  33184=>"000001110",
  33185=>"001100000",
  33186=>"000101101",
  33187=>"110111110",
  33188=>"111111000",
  33189=>"000000000",
  33190=>"110000000",
  33191=>"000000111",
  33192=>"110000000",
  33193=>"111101111",
  33194=>"111111111",
  33195=>"111001001",
  33196=>"000000000",
  33197=>"011111100",
  33198=>"100110000",
  33199=>"000000000",
  33200=>"000100000",
  33201=>"000000000",
  33202=>"111100110",
  33203=>"111111111",
  33204=>"000111011",
  33205=>"111111001",
  33206=>"110111111",
  33207=>"111110000",
  33208=>"111111101",
  33209=>"100111111",
  33210=>"111011000",
  33211=>"100111111",
  33212=>"111111011",
  33213=>"000000000",
  33214=>"010000000",
  33215=>"100111111",
  33216=>"011111111",
  33217=>"010000000",
  33218=>"000000011",
  33219=>"101001000",
  33220=>"000011111",
  33221=>"001000000",
  33222=>"111010000",
  33223=>"000000000",
  33224=>"000000000",
  33225=>"111111000",
  33226=>"100100000",
  33227=>"000101000",
  33228=>"001000101",
  33229=>"111000000",
  33230=>"000000111",
  33231=>"111111000",
  33232=>"000000110",
  33233=>"110000001",
  33234=>"111111111",
  33235=>"000100100",
  33236=>"111000100",
  33237=>"011111111",
  33238=>"000010110",
  33239=>"000000000",
  33240=>"111111000",
  33241=>"000010011",
  33242=>"111000111",
  33243=>"011111111",
  33244=>"000001001",
  33245=>"010000100",
  33246=>"000100111",
  33247=>"000011111",
  33248=>"000111111",
  33249=>"011111001",
  33250=>"000000110",
  33251=>"011000000",
  33252=>"111111111",
  33253=>"000000100",
  33254=>"000100111",
  33255=>"101000000",
  33256=>"111111010",
  33257=>"111111111",
  33258=>"000000011",
  33259=>"111111111",
  33260=>"111101111",
  33261=>"001001111",
  33262=>"111111111",
  33263=>"001000000",
  33264=>"000000000",
  33265=>"111111000",
  33266=>"110100000",
  33267=>"000001011",
  33268=>"000000000",
  33269=>"111110000",
  33270=>"000110000",
  33271=>"000000011",
  33272=>"000000000",
  33273=>"000001001",
  33274=>"000111111",
  33275=>"111001111",
  33276=>"000000111",
  33277=>"000000001",
  33278=>"111111111",
  33279=>"000000000",
  33280=>"111111111",
  33281=>"111111011",
  33282=>"000111111",
  33283=>"111111111",
  33284=>"001011011",
  33285=>"001011011",
  33286=>"100100110",
  33287=>"011110111",
  33288=>"111000000",
  33289=>"000000000",
  33290=>"111111111",
  33291=>"111111111",
  33292=>"011111111",
  33293=>"111111111",
  33294=>"000110011",
  33295=>"000100110",
  33296=>"000000000",
  33297=>"011011000",
  33298=>"000000001",
  33299=>"111111111",
  33300=>"000000000",
  33301=>"111011111",
  33302=>"000000011",
  33303=>"111111111",
  33304=>"100000000",
  33305=>"000001000",
  33306=>"111111111",
  33307=>"111110110",
  33308=>"000000000",
  33309=>"000111111",
  33310=>"111111011",
  33311=>"011000111",
  33312=>"000001001",
  33313=>"000011010",
  33314=>"100110000",
  33315=>"000000000",
  33316=>"000000000",
  33317=>"111000001",
  33318=>"000001000",
  33319=>"111110111",
  33320=>"000100101",
  33321=>"111100111",
  33322=>"111111100",
  33323=>"000011011",
  33324=>"011011111",
  33325=>"000100101",
  33326=>"011011111",
  33327=>"100100100",
  33328=>"111111111",
  33329=>"000001101",
  33330=>"011001000",
  33331=>"000100100",
  33332=>"111111101",
  33333=>"101111110",
  33334=>"101111000",
  33335=>"111111111",
  33336=>"111000111",
  33337=>"111111011",
  33338=>"101111111",
  33339=>"011010000",
  33340=>"000000000",
  33341=>"111000000",
  33342=>"110110110",
  33343=>"000000000",
  33344=>"000000000",
  33345=>"111111111",
  33346=>"111100000",
  33347=>"000000100",
  33348=>"110110111",
  33349=>"000000000",
  33350=>"111100000",
  33351=>"111111111",
  33352=>"000100100",
  33353=>"101001111",
  33354=>"111111111",
  33355=>"111111111",
  33356=>"100100000",
  33357=>"000000111",
  33358=>"000000000",
  33359=>"111111101",
  33360=>"000000001",
  33361=>"111110111",
  33362=>"000000000",
  33363=>"111111000",
  33364=>"000000000",
  33365=>"111111111",
  33366=>"001000001",
  33367=>"000000000",
  33368=>"111111111",
  33369=>"000000000",
  33370=>"000000000",
  33371=>"001000000",
  33372=>"111111111",
  33373=>"010000000",
  33374=>"001000000",
  33375=>"000000000",
  33376=>"110100000",
  33377=>"000000001",
  33378=>"000100100",
  33379=>"111111111",
  33380=>"111110000",
  33381=>"000000000",
  33382=>"000111000",
  33383=>"110011000",
  33384=>"001111111",
  33385=>"111111000",
  33386=>"000000010",
  33387=>"001001000",
  33388=>"011011011",
  33389=>"000010110",
  33390=>"000010000",
  33391=>"001001001",
  33392=>"011111111",
  33393=>"000000000",
  33394=>"111111111",
  33395=>"001001101",
  33396=>"000000000",
  33397=>"111111011",
  33398=>"000000000",
  33399=>"111111111",
  33400=>"000111111",
  33401=>"000111101",
  33402=>"111111000",
  33403=>"111111111",
  33404=>"000001000",
  33405=>"111111110",
  33406=>"000000000",
  33407=>"000000011",
  33408=>"000000000",
  33409=>"111111010",
  33410=>"000110000",
  33411=>"011111111",
  33412=>"100000000",
  33413=>"101000000",
  33414=>"111111111",
  33415=>"000000000",
  33416=>"000111111",
  33417=>"000000111",
  33418=>"100100111",
  33419=>"111100000",
  33420=>"111110000",
  33421=>"011001001",
  33422=>"000100000",
  33423=>"000000010",
  33424=>"111111111",
  33425=>"001001011",
  33426=>"000000000",
  33427=>"000000000",
  33428=>"111111000",
  33429=>"111111110",
  33430=>"000000000",
  33431=>"000111000",
  33432=>"111101111",
  33433=>"111000000",
  33434=>"000000000",
  33435=>"000000000",
  33436=>"011111111",
  33437=>"000000000",
  33438=>"011110111",
  33439=>"100110110",
  33440=>"000000111",
  33441=>"000000000",
  33442=>"000100000",
  33443=>"000000000",
  33444=>"111000001",
  33445=>"111110100",
  33446=>"110111010",
  33447=>"011011011",
  33448=>"111011000",
  33449=>"000000000",
  33450=>"111111111",
  33451=>"111111111",
  33452=>"111100111",
  33453=>"000000111",
  33454=>"111111011",
  33455=>"000000111",
  33456=>"000000011",
  33457=>"100000111",
  33458=>"111111010",
  33459=>"111111111",
  33460=>"001111000",
  33461=>"111111001",
  33462=>"000000000",
  33463=>"000000000",
  33464=>"000111111",
  33465=>"000001001",
  33466=>"001000000",
  33467=>"000000000",
  33468=>"000100100",
  33469=>"010000000",
  33470=>"000100000",
  33471=>"110011000",
  33472=>"001000000",
  33473=>"000000000",
  33474=>"001011110",
  33475=>"000000000",
  33476=>"000000000",
  33477=>"000000110",
  33478=>"010000000",
  33479=>"000010011",
  33480=>"000000000",
  33481=>"100100101",
  33482=>"000110000",
  33483=>"001101111",
  33484=>"000000000",
  33485=>"011000000",
  33486=>"000000100",
  33487=>"000000000",
  33488=>"111000000",
  33489=>"001001111",
  33490=>"011111000",
  33491=>"000000000",
  33492=>"000100000",
  33493=>"001001000",
  33494=>"000000000",
  33495=>"000000000",
  33496=>"111111111",
  33497=>"110100001",
  33498=>"100000001",
  33499=>"000000110",
  33500=>"000000001",
  33501=>"111011111",
  33502=>"000000000",
  33503=>"011111000",
  33504=>"000000000",
  33505=>"011011011",
  33506=>"111111100",
  33507=>"011111111",
  33508=>"000010010",
  33509=>"111001111",
  33510=>"100110111",
  33511=>"000000001",
  33512=>"000000111",
  33513=>"001111011",
  33514=>"110111111",
  33515=>"110111111",
  33516=>"000000000",
  33517=>"000000110",
  33518=>"111100000",
  33519=>"100000111",
  33520=>"000111111",
  33521=>"111000101",
  33522=>"000000000",
  33523=>"000100111",
  33524=>"100001111",
  33525=>"001000001",
  33526=>"011111111",
  33527=>"111111111",
  33528=>"000000000",
  33529=>"000000000",
  33530=>"000000000",
  33531=>"000000000",
  33532=>"001000000",
  33533=>"001000000",
  33534=>"111111011",
  33535=>"000011000",
  33536=>"000000000",
  33537=>"111100101",
  33538=>"001000000",
  33539=>"111111111",
  33540=>"000110110",
  33541=>"000010000",
  33542=>"111001111",
  33543=>"000000000",
  33544=>"111111011",
  33545=>"000001001",
  33546=>"000000000",
  33547=>"001001001",
  33548=>"000000000",
  33549=>"010000000",
  33550=>"100110110",
  33551=>"100101000",
  33552=>"000111111",
  33553=>"000000111",
  33554=>"000000000",
  33555=>"000000000",
  33556=>"111111111",
  33557=>"111111100",
  33558=>"100110100",
  33559=>"000000000",
  33560=>"010110010",
  33561=>"000111111",
  33562=>"011111111",
  33563=>"111111010",
  33564=>"111111001",
  33565=>"111111001",
  33566=>"111111111",
  33567=>"000111011",
  33568=>"000100101",
  33569=>"111111111",
  33570=>"110010111",
  33571=>"001111111",
  33572=>"000000001",
  33573=>"001011010",
  33574=>"000000000",
  33575=>"000000001",
  33576=>"000000000",
  33577=>"000000000",
  33578=>"101111111",
  33579=>"000111001",
  33580=>"000000000",
  33581=>"000011111",
  33582=>"101000000",
  33583=>"000000111",
  33584=>"010110110",
  33585=>"000000000",
  33586=>"000111111",
  33587=>"111001000",
  33588=>"000100111",
  33589=>"000000000",
  33590=>"011111111",
  33591=>"111110111",
  33592=>"000000000",
  33593=>"000000101",
  33594=>"111000000",
  33595=>"000000111",
  33596=>"000000111",
  33597=>"100110110",
  33598=>"111111111",
  33599=>"010110110",
  33600=>"011001111",
  33601=>"111111111",
  33602=>"111111111",
  33603=>"111111101",
  33604=>"000000000",
  33605=>"000000000",
  33606=>"011111101",
  33607=>"111111111",
  33608=>"111111111",
  33609=>"111111111",
  33610=>"000000000",
  33611=>"100110110",
  33612=>"000111010",
  33613=>"011000000",
  33614=>"111100100",
  33615=>"110100110",
  33616=>"100110110",
  33617=>"000001111",
  33618=>"000000000",
  33619=>"111111111",
  33620=>"111100101",
  33621=>"011011111",
  33622=>"111111111",
  33623=>"000000000",
  33624=>"000001001",
  33625=>"100111111",
  33626=>"000000010",
  33627=>"111111010",
  33628=>"000000010",
  33629=>"011010000",
  33630=>"000000000",
  33631=>"110110111",
  33632=>"111111111",
  33633=>"110111111",
  33634=>"111111100",
  33635=>"011000111",
  33636=>"110110000",
  33637=>"000111111",
  33638=>"111111111",
  33639=>"110111100",
  33640=>"001111011",
  33641=>"111111100",
  33642=>"111111100",
  33643=>"000111001",
  33644=>"111111111",
  33645=>"111001111",
  33646=>"111111111",
  33647=>"000000000",
  33648=>"111111111",
  33649=>"111111111",
  33650=>"111111111",
  33651=>"111111010",
  33652=>"000000000",
  33653=>"000000111",
  33654=>"011011111",
  33655=>"000011011",
  33656=>"000000000",
  33657=>"000000100",
  33658=>"000001001",
  33659=>"111100110",
  33660=>"000100110",
  33661=>"111111111",
  33662=>"000110000",
  33663=>"000000100",
  33664=>"000100111",
  33665=>"001000000",
  33666=>"000000000",
  33667=>"111111111",
  33668=>"000000001",
  33669=>"100000000",
  33670=>"000000000",
  33671=>"000000000",
  33672=>"000000000",
  33673=>"100100111",
  33674=>"000000000",
  33675=>"000000000",
  33676=>"001001111",
  33677=>"100100110",
  33678=>"000011011",
  33679=>"110110100",
  33680=>"000010000",
  33681=>"111001001",
  33682=>"000111111",
  33683=>"111110000",
  33684=>"111101101",
  33685=>"000000010",
  33686=>"111111000",
  33687=>"000000000",
  33688=>"000000001",
  33689=>"000000000",
  33690=>"000000000",
  33691=>"111111111",
  33692=>"111111000",
  33693=>"000000000",
  33694=>"000000001",
  33695=>"111111000",
  33696=>"110000000",
  33697=>"000100110",
  33698=>"111111111",
  33699=>"111011111",
  33700=>"111111111",
  33701=>"000000000",
  33702=>"111111011",
  33703=>"000000000",
  33704=>"111111111",
  33705=>"001011000",
  33706=>"110111111",
  33707=>"000101000",
  33708=>"000000000",
  33709=>"000000110",
  33710=>"000000000",
  33711=>"111011010",
  33712=>"110111111",
  33713=>"111111111",
  33714=>"111111111",
  33715=>"000111111",
  33716=>"000110000",
  33717=>"001001111",
  33718=>"110110111",
  33719=>"000000000",
  33720=>"110110111",
  33721=>"110110111",
  33722=>"000000100",
  33723=>"111111101",
  33724=>"000000000",
  33725=>"100110111",
  33726=>"000000000",
  33727=>"111101011",
  33728=>"111111111",
  33729=>"001111111",
  33730=>"111111111",
  33731=>"000000000",
  33732=>"111001001",
  33733=>"111111111",
  33734=>"000000111",
  33735=>"000000000",
  33736=>"101001001",
  33737=>"100000011",
  33738=>"000000011",
  33739=>"000000000",
  33740=>"000110000",
  33741=>"011111011",
  33742=>"000000000",
  33743=>"111000000",
  33744=>"010011001",
  33745=>"000111111",
  33746=>"111111111",
  33747=>"111111111",
  33748=>"000100100",
  33749=>"111110000",
  33750=>"000000000",
  33751=>"111111111",
  33752=>"110110000",
  33753=>"010010110",
  33754=>"111111111",
  33755=>"111000010",
  33756=>"111001000",
  33757=>"100110100",
  33758=>"000000000",
  33759=>"111111011",
  33760=>"100111111",
  33761=>"111111111",
  33762=>"100111111",
  33763=>"110111111",
  33764=>"000000000",
  33765=>"010000000",
  33766=>"000000000",
  33767=>"000000000",
  33768=>"010110110",
  33769=>"111110110",
  33770=>"111000000",
  33771=>"000000010",
  33772=>"001111111",
  33773=>"000000000",
  33774=>"111111111",
  33775=>"111000000",
  33776=>"000000000",
  33777=>"100110000",
  33778=>"000000000",
  33779=>"000000000",
  33780=>"000000001",
  33781=>"000000000",
  33782=>"111001000",
  33783=>"110110111",
  33784=>"000000000",
  33785=>"111111111",
  33786=>"111111111",
  33787=>"110110110",
  33788=>"111000000",
  33789=>"111111111",
  33790=>"000000000",
  33791=>"000001001",
  33792=>"101111111",
  33793=>"000000111",
  33794=>"000000111",
  33795=>"111111111",
  33796=>"001000100",
  33797=>"100100000",
  33798=>"000001001",
  33799=>"100111111",
  33800=>"110111011",
  33801=>"000011111",
  33802=>"111110011",
  33803=>"001001001",
  33804=>"000110111",
  33805=>"111111111",
  33806=>"011000000",
  33807=>"000000000",
  33808=>"111111010",
  33809=>"000000000",
  33810=>"001000000",
  33811=>"111111011",
  33812=>"111111111",
  33813=>"111111110",
  33814=>"100001101",
  33815=>"110111100",
  33816=>"111111111",
  33817=>"000100110",
  33818=>"000000000",
  33819=>"011011000",
  33820=>"000000000",
  33821=>"101000000",
  33822=>"000000100",
  33823=>"111111111",
  33824=>"011000000",
  33825=>"000100100",
  33826=>"110110000",
  33827=>"001001001",
  33828=>"110000000",
  33829=>"000110111",
  33830=>"000000000",
  33831=>"000000000",
  33832=>"000010000",
  33833=>"000000000",
  33834=>"011001001",
  33835=>"100111111",
  33836=>"000111111",
  33837=>"100000000",
  33838=>"001000000",
  33839=>"001111111",
  33840=>"000000111",
  33841=>"000000000",
  33842=>"000000000",
  33843=>"011011011",
  33844=>"001001100",
  33845=>"000000000",
  33846=>"100000000",
  33847=>"100010000",
  33848=>"000101000",
  33849=>"000000000",
  33850=>"000111111",
  33851=>"111101000",
  33852=>"101101111",
  33853=>"000011011",
  33854=>"001001011",
  33855=>"000000001",
  33856=>"000000101",
  33857=>"000100110",
  33858=>"100110111",
  33859=>"111111010",
  33860=>"110110100",
  33861=>"011011011",
  33862=>"000000000",
  33863=>"110111110",
  33864=>"001111111",
  33865=>"101111101",
  33866=>"000000000",
  33867=>"111111111",
  33868=>"000010000",
  33869=>"011111010",
  33870=>"000100101",
  33871=>"010011110",
  33872=>"001011111",
  33873=>"100000000",
  33874=>"000000000",
  33875=>"111111001",
  33876=>"011010000",
  33877=>"000011111",
  33878=>"001111111",
  33879=>"000000101",
  33880=>"000110111",
  33881=>"101000101",
  33882=>"111101101",
  33883=>"110000001",
  33884=>"011011000",
  33885=>"111111111",
  33886=>"000000000",
  33887=>"011001000",
  33888=>"000000000",
  33889=>"011111100",
  33890=>"110110111",
  33891=>"000000111",
  33892=>"110111111",
  33893=>"000010000",
  33894=>"000000000",
  33895=>"111001000",
  33896=>"000000110",
  33897=>"000101101",
  33898=>"010000111",
  33899=>"001000011",
  33900=>"000000000",
  33901=>"111011000",
  33902=>"111111111",
  33903=>"000000000",
  33904=>"000000000",
  33905=>"000000000",
  33906=>"101000000",
  33907=>"000000000",
  33908=>"000001000",
  33909=>"000000000",
  33910=>"100001000",
  33911=>"111111011",
  33912=>"000111111",
  33913=>"000000100",
  33914=>"111010000",
  33915=>"100100100",
  33916=>"100110111",
  33917=>"001000001",
  33918=>"000000000",
  33919=>"011111011",
  33920=>"000001111",
  33921=>"000000000",
  33922=>"111010000",
  33923=>"000000000",
  33924=>"000111111",
  33925=>"111001000",
  33926=>"110110100",
  33927=>"010110000",
  33928=>"000000000",
  33929=>"101101010",
  33930=>"000100001",
  33931=>"000111111",
  33932=>"000000110",
  33933=>"000000111",
  33934=>"110110110",
  33935=>"000011000",
  33936=>"000000000",
  33937=>"100000000",
  33938=>"000000000",
  33939=>"110110000",
  33940=>"101000100",
  33941=>"111111111",
  33942=>"000000111",
  33943=>"110100100",
  33944=>"000000101",
  33945=>"000000001",
  33946=>"110000000",
  33947=>"000111011",
  33948=>"111011011",
  33949=>"011111000",
  33950=>"000000011",
  33951=>"000001000",
  33952=>"011111111",
  33953=>"000111111",
  33954=>"000000000",
  33955=>"111000000",
  33956=>"000000000",
  33957=>"111111111",
  33958=>"111111110",
  33959=>"000000000",
  33960=>"001001111",
  33961=>"011111111",
  33962=>"111101111",
  33963=>"011000000",
  33964=>"000001001",
  33965=>"111111111",
  33966=>"000000100",
  33967=>"111111110",
  33968=>"000000110",
  33969=>"011110000",
  33970=>"000110110",
  33971=>"111111111",
  33972=>"111000000",
  33973=>"111111111",
  33974=>"011010000",
  33975=>"000011111",
  33976=>"010000000",
  33977=>"111100000",
  33978=>"111111111",
  33979=>"110111111",
  33980=>"111000000",
  33981=>"110111111",
  33982=>"000100000",
  33983=>"111111111",
  33984=>"000000000",
  33985=>"000000100",
  33986=>"111011001",
  33987=>"111111111",
  33988=>"111111111",
  33989=>"000111111",
  33990=>"111111111",
  33991=>"000010000",
  33992=>"100111111",
  33993=>"000000000",
  33994=>"111111100",
  33995=>"000000000",
  33996=>"000100000",
  33997=>"010110000",
  33998=>"000000000",
  33999=>"001011111",
  34000=>"100000000",
  34001=>"111111100",
  34002=>"000111111",
  34003=>"100000000",
  34004=>"000000000",
  34005=>"001111110",
  34006=>"000000101",
  34007=>"111111001",
  34008=>"000001011",
  34009=>"010100100",
  34010=>"111111111",
  34011=>"110010000",
  34012=>"000110110",
  34013=>"000101111",
  34014=>"000000000",
  34015=>"000010111",
  34016=>"111111111",
  34017=>"000000000",
  34018=>"111001111",
  34019=>"011111111",
  34020=>"111111101",
  34021=>"111100000",
  34022=>"000000001",
  34023=>"111111111",
  34024=>"111111110",
  34025=>"111001000",
  34026=>"110110000",
  34027=>"000000111",
  34028=>"011111111",
  34029=>"111111111",
  34030=>"000111100",
  34031=>"000100111",
  34032=>"111111001",
  34033=>"111111111",
  34034=>"011110000",
  34035=>"110110000",
  34036=>"000111111",
  34037=>"100000000",
  34038=>"010110110",
  34039=>"111111111",
  34040=>"000000001",
  34041=>"000000000",
  34042=>"000111111",
  34043=>"111000000",
  34044=>"001001001",
  34045=>"001111111",
  34046=>"000000000",
  34047=>"111111111",
  34048=>"000010000",
  34049=>"111100000",
  34050=>"010000000",
  34051=>"001111111",
  34052=>"000000000",
  34053=>"000100111",
  34054=>"001010111",
  34055=>"000111101",
  34056=>"010100000",
  34057=>"001001111",
  34058=>"110000000",
  34059=>"011000000",
  34060=>"111110100",
  34061=>"000011111",
  34062=>"110110000",
  34063=>"111111110",
  34064=>"001001000",
  34065=>"011111111",
  34066=>"111001111",
  34067=>"010111111",
  34068=>"000111111",
  34069=>"000000000",
  34070=>"110110001",
  34071=>"000000000",
  34072=>"000000110",
  34073=>"111111111",
  34074=>"001011010",
  34075=>"111111111",
  34076=>"000111000",
  34077=>"011011010",
  34078=>"111111111",
  34079=>"001111111",
  34080=>"010010000",
  34081=>"010100100",
  34082=>"111111111",
  34083=>"000000000",
  34084=>"000110110",
  34085=>"000010110",
  34086=>"000011000",
  34087=>"011011111",
  34088=>"000000000",
  34089=>"001011111",
  34090=>"011111110",
  34091=>"000000111",
  34092=>"110111111",
  34093=>"000000000",
  34094=>"111001000",
  34095=>"100000001",
  34096=>"111100000",
  34097=>"000010111",
  34098=>"111111111",
  34099=>"000000000",
  34100=>"011000000",
  34101=>"000011001",
  34102=>"000000000",
  34103=>"011110111",
  34104=>"000000100",
  34105=>"100100101",
  34106=>"000000101",
  34107=>"000111111",
  34108=>"000001011",
  34109=>"111111111",
  34110=>"000001001",
  34111=>"111111011",
  34112=>"000100101",
  34113=>"010000000",
  34114=>"111111110",
  34115=>"000000000",
  34116=>"110100000",
  34117=>"011011111",
  34118=>"111000001",
  34119=>"000000000",
  34120=>"000111111",
  34121=>"000000110",
  34122=>"010111111",
  34123=>"000000000",
  34124=>"000000000",
  34125=>"110111010",
  34126=>"111111111",
  34127=>"111011000",
  34128=>"111111011",
  34129=>"000000101",
  34130=>"010110111",
  34131=>"001011000",
  34132=>"111000000",
  34133=>"011011011",
  34134=>"110111111",
  34135=>"000000111",
  34136=>"111111111",
  34137=>"000000000",
  34138=>"000000000",
  34139=>"111111001",
  34140=>"011111111",
  34141=>"111011000",
  34142=>"000000111",
  34143=>"000000000",
  34144=>"100000000",
  34145=>"111111111",
  34146=>"000000000",
  34147=>"111111000",
  34148=>"000000000",
  34149=>"001000000",
  34150=>"000000111",
  34151=>"000100000",
  34152=>"000000000",
  34153=>"111000000",
  34154=>"000010000",
  34155=>"011010000",
  34156=>"100100000",
  34157=>"000100111",
  34158=>"111001001",
  34159=>"000000000",
  34160=>"011000000",
  34161=>"010010111",
  34162=>"000000010",
  34163=>"011011000",
  34164=>"000000000",
  34165=>"110100110",
  34166=>"000000000",
  34167=>"111011000",
  34168=>"111111111",
  34169=>"011100101",
  34170=>"100100000",
  34171=>"000000011",
  34172=>"000000010",
  34173=>"111110111",
  34174=>"011011011",
  34175=>"111111111",
  34176=>"100100000",
  34177=>"110110111",
  34178=>"100110110",
  34179=>"110100000",
  34180=>"000100111",
  34181=>"000000101",
  34182=>"000000000",
  34183=>"110111111",
  34184=>"001000000",
  34185=>"000001011",
  34186=>"111101000",
  34187=>"000000000",
  34188=>"111111111",
  34189=>"000111111",
  34190=>"000000000",
  34191=>"011011010",
  34192=>"000110000",
  34193=>"000000101",
  34194=>"111110110",
  34195=>"000000100",
  34196=>"110110000",
  34197=>"000000000",
  34198=>"000110110",
  34199=>"000000101",
  34200=>"011111000",
  34201=>"000000000",
  34202=>"111111100",
  34203=>"100100100",
  34204=>"011001000",
  34205=>"011111111",
  34206=>"000000101",
  34207=>"000000101",
  34208=>"000011000",
  34209=>"011000100",
  34210=>"010110100",
  34211=>"111111111",
  34212=>"000111101",
  34213=>"101000000",
  34214=>"000000001",
  34215=>"111111111",
  34216=>"000001100",
  34217=>"000000001",
  34218=>"000000000",
  34219=>"000000000",
  34220=>"111111010",
  34221=>"000001001",
  34222=>"000000000",
  34223=>"011111011",
  34224=>"111111100",
  34225=>"111111101",
  34226=>"000001000",
  34227=>"000010011",
  34228=>"111010110",
  34229=>"001100111",
  34230=>"111111111",
  34231=>"010010111",
  34232=>"111110111",
  34233=>"110111000",
  34234=>"000000010",
  34235=>"000000101",
  34236=>"011111111",
  34237=>"111111101",
  34238=>"100100100",
  34239=>"110011000",
  34240=>"000000000",
  34241=>"011011000",
  34242=>"000110111",
  34243=>"001101111",
  34244=>"000111111",
  34245=>"000000110",
  34246=>"000000000",
  34247=>"000000111",
  34248=>"100000000",
  34249=>"111111011",
  34250=>"000000000",
  34251=>"111111000",
  34252=>"111111111",
  34253=>"000100101",
  34254=>"000110100",
  34255=>"111111101",
  34256=>"000000000",
  34257=>"111001011",
  34258=>"000000111",
  34259=>"111111111",
  34260=>"000000000",
  34261=>"110110100",
  34262=>"111111111",
  34263=>"000001011",
  34264=>"111110111",
  34265=>"000000000",
  34266=>"010011111",
  34267=>"000110111",
  34268=>"000001011",
  34269=>"011011111",
  34270=>"111111111",
  34271=>"110000000",
  34272=>"100000111",
  34273=>"111111001",
  34274=>"110011111",
  34275=>"001010000",
  34276=>"110110011",
  34277=>"011011111",
  34278=>"100100101",
  34279=>"001010011",
  34280=>"010110111",
  34281=>"001001001",
  34282=>"101000000",
  34283=>"011111011",
  34284=>"110111111",
  34285=>"000011111",
  34286=>"111000000",
  34287=>"111111111",
  34288=>"000000000",
  34289=>"001111011",
  34290=>"001011000",
  34291=>"111111111",
  34292=>"000111111",
  34293=>"101001111",
  34294=>"011111110",
  34295=>"111111010",
  34296=>"100000000",
  34297=>"000001001",
  34298=>"110000000",
  34299=>"011111001",
  34300=>"110110100",
  34301=>"000000000",
  34302=>"111111000",
  34303=>"000111111",
  34304=>"111110110",
  34305=>"010010000",
  34306=>"101000001",
  34307=>"000000110",
  34308=>"111110001",
  34309=>"000000000",
  34310=>"000000000",
  34311=>"111111111",
  34312=>"111111110",
  34313=>"000000000",
  34314=>"001000000",
  34315=>"111011110",
  34316=>"000100000",
  34317=>"100111111",
  34318=>"000000000",
  34319=>"111111111",
  34320=>"111111111",
  34321=>"000100111",
  34322=>"000000000",
  34323=>"000000000",
  34324=>"000111001",
  34325=>"000010011",
  34326=>"110111000",
  34327=>"000100100",
  34328=>"111110000",
  34329=>"110001111",
  34330=>"000000111",
  34331=>"110111000",
  34332=>"111111101",
  34333=>"100000001",
  34334=>"111001000",
  34335=>"111111000",
  34336=>"111100100",
  34337=>"111111111",
  34338=>"001001000",
  34339=>"001111111",
  34340=>"111111111",
  34341=>"101011011",
  34342=>"001000000",
  34343=>"000101111",
  34344=>"111111011",
  34345=>"000000000",
  34346=>"001001101",
  34347=>"111100000",
  34348=>"001111111",
  34349=>"000001011",
  34350=>"101010010",
  34351=>"000000000",
  34352=>"111000100",
  34353=>"111000000",
  34354=>"000101111",
  34355=>"110100100",
  34356=>"001000001",
  34357=>"010011011",
  34358=>"011111011",
  34359=>"000000001",
  34360=>"000110100",
  34361=>"000000110",
  34362=>"000000000",
  34363=>"000000000",
  34364=>"000000000",
  34365=>"000101000",
  34366=>"110111111",
  34367=>"111111000",
  34368=>"000111111",
  34369=>"000110110",
  34370=>"000111111",
  34371=>"000000100",
  34372=>"110110110",
  34373=>"111111010",
  34374=>"100000000",
  34375=>"111111111",
  34376=>"011111111",
  34377=>"111001111",
  34378=>"000000000",
  34379=>"100111111",
  34380=>"111111010",
  34381=>"000000100",
  34382=>"011000000",
  34383=>"000000000",
  34384=>"000000000",
  34385=>"000000111",
  34386=>"000000000",
  34387=>"111111001",
  34388=>"000101111",
  34389=>"111111111",
  34390=>"000001001",
  34391=>"100110110",
  34392=>"100000000",
  34393=>"000000101",
  34394=>"000000100",
  34395=>"000010010",
  34396=>"000000000",
  34397=>"111111110",
  34398=>"110111000",
  34399=>"000100000",
  34400=>"000000011",
  34401=>"000000111",
  34402=>"011001001",
  34403=>"000000000",
  34404=>"111001000",
  34405=>"000000111",
  34406=>"000000000",
  34407=>"111101100",
  34408=>"000000000",
  34409=>"000000010",
  34410=>"000000010",
  34411=>"110000110",
  34412=>"111111111",
  34413=>"111100000",
  34414=>"000000000",
  34415=>"100000000",
  34416=>"000000000",
  34417=>"110111111",
  34418=>"011000000",
  34419=>"001000000",
  34420=>"111111111",
  34421=>"101111111",
  34422=>"000000000",
  34423=>"001000110",
  34424=>"111000100",
  34425=>"000000000",
  34426=>"111000111",
  34427=>"000000100",
  34428=>"001010000",
  34429=>"111111111",
  34430=>"111000000",
  34431=>"001100000",
  34432=>"110111110",
  34433=>"000110110",
  34434=>"000110000",
  34435=>"000001101",
  34436=>"111110111",
  34437=>"000000000",
  34438=>"111111001",
  34439=>"111010011",
  34440=>"111100000",
  34441=>"110000000",
  34442=>"100100000",
  34443=>"011001111",
  34444=>"000001001",
  34445=>"000000000",
  34446=>"111000000",
  34447=>"111111001",
  34448=>"000000001",
  34449=>"111111111",
  34450=>"111111000",
  34451=>"111111001",
  34452=>"010111111",
  34453=>"111111000",
  34454=>"000010000",
  34455=>"000000000",
  34456=>"000000000",
  34457=>"111111110",
  34458=>"111111111",
  34459=>"100011000",
  34460=>"111111111",
  34461=>"001011000",
  34462=>"111111111",
  34463=>"000100000",
  34464=>"000111111",
  34465=>"111111110",
  34466=>"000110000",
  34467=>"111011111",
  34468=>"111011111",
  34469=>"111111001",
  34470=>"001000111",
  34471=>"101101101",
  34472=>"011011000",
  34473=>"111111111",
  34474=>"011000000",
  34475=>"000100101",
  34476=>"000000000",
  34477=>"111111001",
  34478=>"000110000",
  34479=>"111111001",
  34480=>"000111000",
  34481=>"111111011",
  34482=>"011111111",
  34483=>"111001111",
  34484=>"111110110",
  34485=>"000000100",
  34486=>"011111011",
  34487=>"011111111",
  34488=>"111111111",
  34489=>"001000000",
  34490=>"111000011",
  34491=>"001001011",
  34492=>"110111110",
  34493=>"000000000",
  34494=>"111111110",
  34495=>"111111110",
  34496=>"111111111",
  34497=>"111111111",
  34498=>"010010110",
  34499=>"000000111",
  34500=>"011001001",
  34501=>"000000100",
  34502=>"000000100",
  34503=>"100100111",
  34504=>"011010111",
  34505=>"101111111",
  34506=>"001000000",
  34507=>"111010000",
  34508=>"000001111",
  34509=>"100100101",
  34510=>"000111111",
  34511=>"111100100",
  34512=>"100010011",
  34513=>"111111000",
  34514=>"111000000",
  34515=>"110111111",
  34516=>"100100111",
  34517=>"111111111",
  34518=>"000000000",
  34519=>"110011001",
  34520=>"111110000",
  34521=>"101000000",
  34522=>"000000000",
  34523=>"111111111",
  34524=>"000000000",
  34525=>"111111111",
  34526=>"000000000",
  34527=>"000000000",
  34528=>"011111000",
  34529=>"000000000",
  34530=>"000000010",
  34531=>"111111000",
  34532=>"111000010",
  34533=>"001000101",
  34534=>"111111100",
  34535=>"011100001",
  34536=>"000000111",
  34537=>"111101101",
  34538=>"000100110",
  34539=>"100101111",
  34540=>"000000000",
  34541=>"000000000",
  34542=>"110111000",
  34543=>"000000000",
  34544=>"111001000",
  34545=>"011000000",
  34546=>"111000000",
  34547=>"000111111",
  34548=>"111111111",
  34549=>"000111011",
  34550=>"101101000",
  34551=>"000000111",
  34552=>"001101111",
  34553=>"000000000",
  34554=>"000111110",
  34555=>"001111111",
  34556=>"000000000",
  34557=>"011010100",
  34558=>"000000100",
  34559=>"111111000",
  34560=>"000111111",
  34561=>"111011000",
  34562=>"111111111",
  34563=>"111101100",
  34564=>"110100100",
  34565=>"110111111",
  34566=>"000000001",
  34567=>"000000000",
  34568=>"000000111",
  34569=>"110000000",
  34570=>"000000001",
  34571=>"111111111",
  34572=>"101000000",
  34573=>"000000000",
  34574=>"100100011",
  34575=>"000111111",
  34576=>"111111110",
  34577=>"010111000",
  34578=>"000000101",
  34579=>"001001111",
  34580=>"111000000",
  34581=>"110110111",
  34582=>"100100000",
  34583=>"100110111",
  34584=>"111111111",
  34585=>"111111010",
  34586=>"111111111",
  34587=>"111001000",
  34588=>"111111000",
  34589=>"010010110",
  34590=>"000000000",
  34591=>"000000000",
  34592=>"111111000",
  34593=>"000010110",
  34594=>"000000111",
  34595=>"000001001",
  34596=>"011000000",
  34597=>"100110110",
  34598=>"100000000",
  34599=>"110110000",
  34600=>"000000100",
  34601=>"111111111",
  34602=>"111111010",
  34603=>"000000000",
  34604=>"000100111",
  34605=>"101111111",
  34606=>"000000111",
  34607=>"000000000",
  34608=>"000000001",
  34609=>"001001011",
  34610=>"111111111",
  34611=>"111000000",
  34612=>"000000000",
  34613=>"000011011",
  34614=>"010111000",
  34615=>"111000001",
  34616=>"000000000",
  34617=>"000000000",
  34618=>"111101101",
  34619=>"111101000",
  34620=>"000100100",
  34621=>"011111000",
  34622=>"111100000",
  34623=>"111111000",
  34624=>"000110000",
  34625=>"110111100",
  34626=>"000000000",
  34627=>"000000110",
  34628=>"111111111",
  34629=>"000001000",
  34630=>"111101100",
  34631=>"000000000",
  34632=>"100000000",
  34633=>"111000010",
  34634=>"110000000",
  34635=>"110100100",
  34636=>"000100111",
  34637=>"010000001",
  34638=>"111111111",
  34639=>"111111011",
  34640=>"011011111",
  34641=>"101111110",
  34642=>"111111111",
  34643=>"100110111",
  34644=>"111001011",
  34645=>"011011011",
  34646=>"000100111",
  34647=>"111001000",
  34648=>"000001000",
  34649=>"000000000",
  34650=>"111111111",
  34651=>"000000000",
  34652=>"111110100",
  34653=>"010011000",
  34654=>"111011011",
  34655=>"100000000",
  34656=>"000000000",
  34657=>"111111111",
  34658=>"000001001",
  34659=>"100000000",
  34660=>"000011011",
  34661=>"000000000",
  34662=>"000000101",
  34663=>"111100101",
  34664=>"000111110",
  34665=>"111111111",
  34666=>"000100100",
  34667=>"101111111",
  34668=>"100111110",
  34669=>"000011111",
  34670=>"010111111",
  34671=>"001000000",
  34672=>"000000000",
  34673=>"111100100",
  34674=>"000000000",
  34675=>"111111111",
  34676=>"111110001",
  34677=>"011000000",
  34678=>"000001000",
  34679=>"000000110",
  34680=>"011111111",
  34681=>"000110000",
  34682=>"000000011",
  34683=>"000000000",
  34684=>"000000100",
  34685=>"001000100",
  34686=>"000000000",
  34687=>"100000001",
  34688=>"000101000",
  34689=>"110111110",
  34690=>"110110110",
  34691=>"100000000",
  34692=>"000001111",
  34693=>"001011110",
  34694=>"011001101",
  34695=>"110000000",
  34696=>"000000001",
  34697=>"010111011",
  34698=>"111000000",
  34699=>"000000000",
  34700=>"111111111",
  34701=>"000100000",
  34702=>"000000000",
  34703=>"000000100",
  34704=>"000000000",
  34705=>"000000000",
  34706=>"000000000",
  34707=>"001001001",
  34708=>"011111111",
  34709=>"000000000",
  34710=>"001001111",
  34711=>"000000010",
  34712=>"000000000",
  34713=>"000100100",
  34714=>"000000000",
  34715=>"111111110",
  34716=>"100110000",
  34717=>"111111110",
  34718=>"111101111",
  34719=>"111111111",
  34720=>"000000000",
  34721=>"111101100",
  34722=>"000100101",
  34723=>"000000000",
  34724=>"000000000",
  34725=>"110110111",
  34726=>"111111111",
  34727=>"111100000",
  34728=>"000100000",
  34729=>"001000000",
  34730=>"000000111",
  34731=>"111000001",
  34732=>"000000000",
  34733=>"000000000",
  34734=>"000010100",
  34735=>"111111101",
  34736=>"000100111",
  34737=>"000000000",
  34738=>"111111010",
  34739=>"011001010",
  34740=>"111111010",
  34741=>"000000111",
  34742=>"111100111",
  34743=>"010000000",
  34744=>"000111110",
  34745=>"000011001",
  34746=>"000000110",
  34747=>"000110110",
  34748=>"000111111",
  34749=>"000000000",
  34750=>"000000000",
  34751=>"100111000",
  34752=>"111111011",
  34753=>"100000001",
  34754=>"110111000",
  34755=>"000000000",
  34756=>"000110110",
  34757=>"001000011",
  34758=>"000110110",
  34759=>"001000000",
  34760=>"000000000",
  34761=>"100000000",
  34762=>"000000000",
  34763=>"000111011",
  34764=>"111111001",
  34765=>"001001111",
  34766=>"111001000",
  34767=>"001000110",
  34768=>"111011000",
  34769=>"111111011",
  34770=>"100100111",
  34771=>"100000000",
  34772=>"110111011",
  34773=>"000000000",
  34774=>"000000111",
  34775=>"001001000",
  34776=>"000111111",
  34777=>"001111111",
  34778=>"111110110",
  34779=>"001011111",
  34780=>"111111111",
  34781=>"000001011",
  34782=>"111111101",
  34783=>"110101001",
  34784=>"001111111",
  34785=>"100000000",
  34786=>"011111111",
  34787=>"000001111",
  34788=>"010111100",
  34789=>"111100100",
  34790=>"000000000",
  34791=>"000000000",
  34792=>"001111110",
  34793=>"001001000",
  34794=>"000111111",
  34795=>"001000000",
  34796=>"111011001",
  34797=>"101111111",
  34798=>"001001111",
  34799=>"011011111",
  34800=>"111111111",
  34801=>"111111111",
  34802=>"100111111",
  34803=>"000000000",
  34804=>"001011000",
  34805=>"000000011",
  34806=>"000000001",
  34807=>"011000000",
  34808=>"000100000",
  34809=>"000000001",
  34810=>"001000000",
  34811=>"000000011",
  34812=>"001000000",
  34813=>"010000000",
  34814=>"000000000",
  34815=>"111111111",
  34816=>"100111111",
  34817=>"111001001",
  34818=>"001111111",
  34819=>"000000000",
  34820=>"000000000",
  34821=>"001001011",
  34822=>"110110111",
  34823=>"111000000",
  34824=>"100000000",
  34825=>"010111000",
  34826=>"000100111",
  34827=>"111111111",
  34828=>"001111111",
  34829=>"100111001",
  34830=>"000010000",
  34831=>"111011111",
  34832=>"110000100",
  34833=>"000000000",
  34834=>"000000111",
  34835=>"011000000",
  34836=>"000000000",
  34837=>"111111000",
  34838=>"110110110",
  34839=>"000000011",
  34840=>"110110000",
  34841=>"000010011",
  34842=>"111111000",
  34843=>"011011111",
  34844=>"000000110",
  34845=>"011001111",
  34846=>"110000000",
  34847=>"000000000",
  34848=>"100111111",
  34849=>"110110111",
  34850=>"111011000",
  34851=>"111101101",
  34852=>"100100111",
  34853=>"111111111",
  34854=>"111111000",
  34855=>"110100000",
  34856=>"100101111",
  34857=>"000000000",
  34858=>"111111111",
  34859=>"100110111",
  34860=>"111100000",
  34861=>"111111001",
  34862=>"110010001",
  34863=>"111001011",
  34864=>"100100000",
  34865=>"000001111",
  34866=>"110110111",
  34867=>"100101001",
  34868=>"011011111",
  34869=>"111011001",
  34870=>"000100110",
  34871=>"011001000",
  34872=>"000000111",
  34873=>"110100000",
  34874=>"000000000",
  34875=>"011011000",
  34876=>"000000001",
  34877=>"000000111",
  34878=>"000000000",
  34879=>"000000100",
  34880=>"000000100",
  34881=>"111111111",
  34882=>"100100111",
  34883=>"111001001",
  34884=>"000000111",
  34885=>"100000001",
  34886=>"111111000",
  34887=>"111111111",
  34888=>"011011111",
  34889=>"000000000",
  34890=>"111111110",
  34891=>"000000000",
  34892=>"110111000",
  34893=>"111111111",
  34894=>"111100111",
  34895=>"110000000",
  34896=>"111110010",
  34897=>"000001000",
  34898=>"000000000",
  34899=>"001101000",
  34900=>"000000001",
  34901=>"100000000",
  34902=>"111000100",
  34903=>"000000000",
  34904=>"001000000",
  34905=>"000000000",
  34906=>"000000000",
  34907=>"011001001",
  34908=>"000111110",
  34909=>"111001000",
  34910=>"111110111",
  34911=>"101101100",
  34912=>"100100110",
  34913=>"000000000",
  34914=>"111111000",
  34915=>"000001000",
  34916=>"110111000",
  34917=>"000000111",
  34918=>"000000011",
  34919=>"000000000",
  34920=>"111000000",
  34921=>"100110000",
  34922=>"111111110",
  34923=>"001000000",
  34924=>"000001000",
  34925=>"111000111",
  34926=>"000111000",
  34927=>"111010000",
  34928=>"000000011",
  34929=>"001001111",
  34930=>"111111001",
  34931=>"111010010",
  34932=>"000000111",
  34933=>"001111100",
  34934=>"010111011",
  34935=>"000000000",
  34936=>"000000000",
  34937=>"000110111",
  34938=>"111000111",
  34939=>"111110000",
  34940=>"000000011",
  34941=>"100101110",
  34942=>"101111101",
  34943=>"111110000",
  34944=>"000000000",
  34945=>"111000000",
  34946=>"111110000",
  34947=>"110011111",
  34948=>"111000000",
  34949=>"010001111",
  34950=>"000000100",
  34951=>"000001000",
  34952=>"000111111",
  34953=>"011011000",
  34954=>"100100111",
  34955=>"111100000",
  34956=>"001101011",
  34957=>"001001001",
  34958=>"001111111",
  34959=>"000001111",
  34960=>"010111111",
  34961=>"000110010",
  34962=>"001000111",
  34963=>"000111111",
  34964=>"000000100",
  34965=>"111111000",
  34966=>"000000110",
  34967=>"111111000",
  34968=>"001000011",
  34969=>"011110111",
  34970=>"000001000",
  34971=>"000110000",
  34972=>"001111111",
  34973=>"100000000",
  34974=>"000100000",
  34975=>"111110000",
  34976=>"001000000",
  34977=>"001000000",
  34978=>"000000000",
  34979=>"001111011",
  34980=>"111101101",
  34981=>"100111101",
  34982=>"111111111",
  34983=>"111001000",
  34984=>"100100001",
  34985=>"000000000",
  34986=>"000000000",
  34987=>"000000001",
  34988=>"000010110",
  34989=>"000001111",
  34990=>"000100100",
  34991=>"110000000",
  34992=>"111011000",
  34993=>"100000111",
  34994=>"111111111",
  34995=>"000001111",
  34996=>"110111110",
  34997=>"011000000",
  34998=>"000000010",
  34999=>"110111100",
  35000=>"111001001",
  35001=>"111011111",
  35002=>"111110110",
  35003=>"100111111",
  35004=>"000000100",
  35005=>"000000100",
  35006=>"111000111",
  35007=>"110111000",
  35008=>"010010000",
  35009=>"111000110",
  35010=>"000100100",
  35011=>"111001111",
  35012=>"000111111",
  35013=>"000000000",
  35014=>"000000000",
  35015=>"110110000",
  35016=>"000000010",
  35017=>"111111111",
  35018=>"111111000",
  35019=>"000000000",
  35020=>"011000000",
  35021=>"110110000",
  35022=>"111111000",
  35023=>"111000001",
  35024=>"101101000",
  35025=>"100000100",
  35026=>"110111001",
  35027=>"111111111",
  35028=>"000000000",
  35029=>"001001000",
  35030=>"000000011",
  35031=>"000000010",
  35032=>"000011000",
  35033=>"101000101",
  35034=>"001011000",
  35035=>"101111000",
  35036=>"001000000",
  35037=>"010000001",
  35038=>"110111111",
  35039=>"000111000",
  35040=>"110100100",
  35041=>"000100100",
  35042=>"111001101",
  35043=>"000000000",
  35044=>"101111111",
  35045=>"101111111",
  35046=>"111100110",
  35047=>"001000000",
  35048=>"000011001",
  35049=>"111111000",
  35050=>"110100000",
  35051=>"111001111",
  35052=>"010110010",
  35053=>"011001000",
  35054=>"000000001",
  35055=>"000000000",
  35056=>"110110000",
  35057=>"100111001",
  35058=>"001001100",
  35059=>"101101001",
  35060=>"000000110",
  35061=>"001001101",
  35062=>"011000000",
  35063=>"011000000",
  35064=>"111111111",
  35065=>"111010011",
  35066=>"100100111",
  35067=>"000000001",
  35068=>"100101001",
  35069=>"101001000",
  35070=>"111111111",
  35071=>"111111101",
  35072=>"110000000",
  35073=>"111111111",
  35074=>"111101101",
  35075=>"110000000",
  35076=>"101000000",
  35077=>"111111110",
  35078=>"100000000",
  35079=>"111000100",
  35080=>"111100111",
  35081=>"000000111",
  35082=>"111000000",
  35083=>"100001000",
  35084=>"000010111",
  35085=>"000011011",
  35086=>"100111000",
  35087=>"111111000",
  35088=>"000000100",
  35089=>"010000000",
  35090=>"000000000",
  35091=>"111000000",
  35092=>"000000000",
  35093=>"000000111",
  35094=>"011000001",
  35095=>"000000011",
  35096=>"111111111",
  35097=>"100100111",
  35098=>"010000010",
  35099=>"001011000",
  35100=>"110001001",
  35101=>"000000000",
  35102=>"100000000",
  35103=>"000000110",
  35104=>"110100000",
  35105=>"100111111",
  35106=>"000001011",
  35107=>"100111111",
  35108=>"000001001",
  35109=>"011000000",
  35110=>"000111111",
  35111=>"000000000",
  35112=>"000111000",
  35113=>"000000000",
  35114=>"001011111",
  35115=>"000110111",
  35116=>"001001001",
  35117=>"000011011",
  35118=>"000000000",
  35119=>"111110111",
  35120=>"001001011",
  35121=>"111100100",
  35122=>"001000111",
  35123=>"110000000",
  35124=>"100000100",
  35125=>"000010011",
  35126=>"101000000",
  35127=>"100000110",
  35128=>"011000000",
  35129=>"001000101",
  35130=>"000000110",
  35131=>"000111111",
  35132=>"111111111",
  35133=>"001001011",
  35134=>"111111000",
  35135=>"110111110",
  35136=>"000000000",
  35137=>"111111110",
  35138=>"111000111",
  35139=>"000111000",
  35140=>"111101000",
  35141=>"110100101",
  35142=>"001001101",
  35143=>"101111111",
  35144=>"000000000",
  35145=>"000000000",
  35146=>"001111111",
  35147=>"100100110",
  35148=>"011101000",
  35149=>"000000000",
  35150=>"000100001",
  35151=>"100111111",
  35152=>"111111100",
  35153=>"111001111",
  35154=>"010000000",
  35155=>"111000000",
  35156=>"000110111",
  35157=>"000000101",
  35158=>"000001100",
  35159=>"110000111",
  35160=>"000000000",
  35161=>"000000000",
  35162=>"000111110",
  35163=>"000100111",
  35164=>"111010000",
  35165=>"000000000",
  35166=>"001101100",
  35167=>"000100101",
  35168=>"001111011",
  35169=>"111000000",
  35170=>"000000000",
  35171=>"000000000",
  35172=>"110101000",
  35173=>"000000000",
  35174=>"000000000",
  35175=>"111111111",
  35176=>"011001001",
  35177=>"000001001",
  35178=>"000011011",
  35179=>"000100111",
  35180=>"001001111",
  35181=>"111110110",
  35182=>"100000110",
  35183=>"000000000",
  35184=>"001001010",
  35185=>"110000111",
  35186=>"111010000",
  35187=>"011111011",
  35188=>"000111111",
  35189=>"000100000",
  35190=>"111110000",
  35191=>"111001000",
  35192=>"111001001",
  35193=>"111001001",
  35194=>"111000010",
  35195=>"101101111",
  35196=>"111101111",
  35197=>"000000100",
  35198=>"100111100",
  35199=>"100110111",
  35200=>"000000000",
  35201=>"000000000",
  35202=>"001000000",
  35203=>"000000000",
  35204=>"000000011",
  35205=>"001101111",
  35206=>"110111110",
  35207=>"111101000",
  35208=>"000111010",
  35209=>"111011111",
  35210=>"111111111",
  35211=>"000001110",
  35212=>"111101111",
  35213=>"000011000",
  35214=>"100100111",
  35215=>"111111000",
  35216=>"110000111",
  35217=>"101101100",
  35218=>"111010011",
  35219=>"111110111",
  35220=>"101000000",
  35221=>"000010001",
  35222=>"101111111",
  35223=>"101100100",
  35224=>"000011111",
  35225=>"000011111",
  35226=>"111000011",
  35227=>"111111011",
  35228=>"111111000",
  35229=>"111011000",
  35230=>"000111111",
  35231=>"000001001",
  35232=>"100000000",
  35233=>"011110000",
  35234=>"111111111",
  35235=>"000101001",
  35236=>"111110100",
  35237=>"101100000",
  35238=>"100100000",
  35239=>"011111111",
  35240=>"000000001",
  35241=>"000100101",
  35242=>"111111011",
  35243=>"000111111",
  35244=>"111100010",
  35245=>"011000000",
  35246=>"000000111",
  35247=>"111110111",
  35248=>"000000111",
  35249=>"000010011",
  35250=>"100100000",
  35251=>"000000000",
  35252=>"000010111",
  35253=>"111111000",
  35254=>"111111111",
  35255=>"111111000",
  35256=>"011001011",
  35257=>"011111111",
  35258=>"001001000",
  35259=>"111111111",
  35260=>"011000111",
  35261=>"111111111",
  35262=>"111111111",
  35263=>"111101111",
  35264=>"111111011",
  35265=>"110111111",
  35266=>"000100111",
  35267=>"111000000",
  35268=>"000000001",
  35269=>"101001000",
  35270=>"110011011",
  35271=>"000101111",
  35272=>"111111111",
  35273=>"000000111",
  35274=>"001000001",
  35275=>"111000000",
  35276=>"000000000",
  35277=>"111111000",
  35278=>"111000000",
  35279=>"011011111",
  35280=>"110000111",
  35281=>"000111110",
  35282=>"000111100",
  35283=>"111111000",
  35284=>"010000000",
  35285=>"111101001",
  35286=>"000011111",
  35287=>"110111111",
  35288=>"000000111",
  35289=>"111000111",
  35290=>"111111110",
  35291=>"000000000",
  35292=>"000000000",
  35293=>"100111111",
  35294=>"111111000",
  35295=>"111100111",
  35296=>"011000000",
  35297=>"001000000",
  35298=>"110110000",
  35299=>"001010111",
  35300=>"000111111",
  35301=>"111111111",
  35302=>"111111111",
  35303=>"111111111",
  35304=>"111111011",
  35305=>"000000111",
  35306=>"111001000",
  35307=>"000000000",
  35308=>"100111110",
  35309=>"001000001",
  35310=>"010111110",
  35311=>"111011111",
  35312=>"001111111",
  35313=>"000100100",
  35314=>"100100000",
  35315=>"000010000",
  35316=>"101111111",
  35317=>"101001001",
  35318=>"000000100",
  35319=>"101001111",
  35320=>"000001111",
  35321=>"101001001",
  35322=>"101001001",
  35323=>"011111111",
  35324=>"111000000",
  35325=>"011111110",
  35326=>"111000111",
  35327=>"110110000",
  35328=>"111111111",
  35329=>"111111111",
  35330=>"000000000",
  35331=>"111111011",
  35332=>"000000000",
  35333=>"111111010",
  35334=>"001000001",
  35335=>"100111101",
  35336=>"000110111",
  35337=>"000001111",
  35338=>"000000000",
  35339=>"110111000",
  35340=>"111111110",
  35341=>"000100111",
  35342=>"000100000",
  35343=>"100111110",
  35344=>"000100111",
  35345=>"000011000",
  35346=>"011111111",
  35347=>"000000000",
  35348=>"000000000",
  35349=>"110000011",
  35350=>"110110100",
  35351=>"000001000",
  35352=>"111001001",
  35353=>"000000000",
  35354=>"100100000",
  35355=>"000100111",
  35356=>"100000000",
  35357=>"111111111",
  35358=>"110011000",
  35359=>"000000101",
  35360=>"111000000",
  35361=>"111111111",
  35362=>"011111111",
  35363=>"000000000",
  35364=>"111111000",
  35365=>"000001001",
  35366=>"110110100",
  35367=>"001101111",
  35368=>"111111000",
  35369=>"000000000",
  35370=>"111111110",
  35371=>"111111111",
  35372=>"111001011",
  35373=>"010011111",
  35374=>"001001111",
  35375=>"000000000",
  35376=>"000000111",
  35377=>"110110100",
  35378=>"001001001",
  35379=>"101000001",
  35380=>"110110111",
  35381=>"000001001",
  35382=>"000000000",
  35383=>"000000000",
  35384=>"000000001",
  35385=>"111111111",
  35386=>"111010001",
  35387=>"000000000",
  35388=>"101000111",
  35389=>"101000000",
  35390=>"111100111",
  35391=>"001001000",
  35392=>"000000000",
  35393=>"000000000",
  35394=>"111111111",
  35395=>"000011111",
  35396=>"110111000",
  35397=>"111111001",
  35398=>"111111111",
  35399=>"111111111",
  35400=>"111111011",
  35401=>"110000011",
  35402=>"000001000",
  35403=>"000000000",
  35404=>"111000000",
  35405=>"111000000",
  35406=>"111010110",
  35407=>"001000111",
  35408=>"000000000",
  35409=>"111000000",
  35410=>"001111000",
  35411=>"101101000",
  35412=>"011000001",
  35413=>"100001011",
  35414=>"110000000",
  35415=>"100100111",
  35416=>"111100100",
  35417=>"001000000",
  35418=>"000000000",
  35419=>"000000000",
  35420=>"000000110",
  35421=>"101101000",
  35422=>"111000111",
  35423=>"000000100",
  35424=>"000000000",
  35425=>"000000000",
  35426=>"000000011",
  35427=>"000000000",
  35428=>"111111111",
  35429=>"111001111",
  35430=>"000000011",
  35431=>"000000000",
  35432=>"110100000",
  35433=>"000000001",
  35434=>"111111000",
  35435=>"000010111",
  35436=>"000111111",
  35437=>"100000000",
  35438=>"111101000",
  35439=>"000110000",
  35440=>"000000001",
  35441=>"010010010",
  35442=>"000000000",
  35443=>"101000010",
  35444=>"001000100",
  35445=>"000010010",
  35446=>"000000000",
  35447=>"000000011",
  35448=>"110000010",
  35449=>"111111100",
  35450=>"000000101",
  35451=>"000000001",
  35452=>"110110111",
  35453=>"001000100",
  35454=>"000000000",
  35455=>"000000000",
  35456=>"000000000",
  35457=>"011011011",
  35458=>"111101001",
  35459=>"011011000",
  35460=>"111111111",
  35461=>"100000111",
  35462=>"000000111",
  35463=>"110000000",
  35464=>"000000100",
  35465=>"011111111",
  35466=>"000000000",
  35467=>"000000000",
  35468=>"111000111",
  35469=>"100111111",
  35470=>"010010110",
  35471=>"111000000",
  35472=>"000001011",
  35473=>"010110111",
  35474=>"011000000",
  35475=>"111001000",
  35476=>"011010111",
  35477=>"000000000",
  35478=>"000100111",
  35479=>"100100000",
  35480=>"000000000",
  35481=>"111111111",
  35482=>"000000000",
  35483=>"111000000",
  35484=>"000000010",
  35485=>"100000001",
  35486=>"000000101",
  35487=>"000000000",
  35488=>"111111111",
  35489=>"010111000",
  35490=>"000011000",
  35491=>"011010010",
  35492=>"100110111",
  35493=>"111111111",
  35494=>"111111111",
  35495=>"001111001",
  35496=>"111110100",
  35497=>"000010001",
  35498=>"111000000",
  35499=>"000000001",
  35500=>"011000000",
  35501=>"000011111",
  35502=>"111111000",
  35503=>"000000001",
  35504=>"010000000",
  35505=>"111111000",
  35506=>"111111111",
  35507=>"110111111",
  35508=>"000000111",
  35509=>"100101100",
  35510=>"111111111",
  35511=>"000000111",
  35512=>"111111111",
  35513=>"000000110",
  35514=>"000010011",
  35515=>"011100110",
  35516=>"101111001",
  35517=>"001000000",
  35518=>"110111000",
  35519=>"111000000",
  35520=>"000000000",
  35521=>"100111111",
  35522=>"110110110",
  35523=>"000000000",
  35524=>"110000000",
  35525=>"111111111",
  35526=>"111000010",
  35527=>"000111111",
  35528=>"000000000",
  35529=>"000000101",
  35530=>"001000111",
  35531=>"000000000",
  35532=>"111111001",
  35533=>"000000000",
  35534=>"111000001",
  35535=>"000000000",
  35536=>"000111111",
  35537=>"000000000",
  35538=>"000001000",
  35539=>"111111011",
  35540=>"111111011",
  35541=>"111111111",
  35542=>"000000000",
  35543=>"000010000",
  35544=>"000000001",
  35545=>"000000001",
  35546=>"000000111",
  35547=>"001000111",
  35548=>"111111111",
  35549=>"000100111",
  35550=>"110000000",
  35551=>"000000110",
  35552=>"000000011",
  35553=>"000100000",
  35554=>"000000010",
  35555=>"101000000",
  35556=>"000000011",
  35557=>"000000000",
  35558=>"011000001",
  35559=>"000000100",
  35560=>"111111000",
  35561=>"111111111",
  35562=>"000111011",
  35563=>"000000000",
  35564=>"000000010",
  35565=>"000000011",
  35566=>"000110111",
  35567=>"000001111",
  35568=>"110111101",
  35569=>"100000011",
  35570=>"000000011",
  35571=>"111111010",
  35572=>"111111100",
  35573=>"000100001",
  35574=>"000101111",
  35575=>"000111000",
  35576=>"111111110",
  35577=>"010110111",
  35578=>"000110111",
  35579=>"000001011",
  35580=>"000000000",
  35581=>"101001001",
  35582=>"000000000",
  35583=>"111111111",
  35584=>"011000000",
  35585=>"111100111",
  35586=>"000000011",
  35587=>"000000001",
  35588=>"111000100",
  35589=>"000000000",
  35590=>"000000111",
  35591=>"000100111",
  35592=>"000000000",
  35593=>"000000000",
  35594=>"111111100",
  35595=>"000000000",
  35596=>"111010011",
  35597=>"000000001",
  35598=>"000000111",
  35599=>"000000110",
  35600=>"100111101",
  35601=>"111111111",
  35602=>"000011111",
  35603=>"111111100",
  35604=>"111111000",
  35605=>"001000000",
  35606=>"001000111",
  35607=>"000000100",
  35608=>"111111000",
  35609=>"000000000",
  35610=>"000000100",
  35611=>"000000000",
  35612=>"111111110",
  35613=>"111110100",
  35614=>"000000111",
  35615=>"011000000",
  35616=>"001001001",
  35617=>"000000000",
  35618=>"011011000",
  35619=>"000110111",
  35620=>"101101111",
  35621=>"100111111",
  35622=>"000111111",
  35623=>"011100000",
  35624=>"000000100",
  35625=>"111111100",
  35626=>"111000000",
  35627=>"001000000",
  35628=>"000000000",
  35629=>"000000000",
  35630=>"101100111",
  35631=>"111111100",
  35632=>"000111011",
  35633=>"111011101",
  35634=>"000000000",
  35635=>"111010000",
  35636=>"001001111",
  35637=>"000000111",
  35638=>"000111001",
  35639=>"111111111",
  35640=>"000000000",
  35641=>"111111111",
  35642=>"111111111",
  35643=>"110110110",
  35644=>"111111011",
  35645=>"110010111",
  35646=>"111100101",
  35647=>"000000101",
  35648=>"110000000",
  35649=>"011110000",
  35650=>"111111010",
  35651=>"000000010",
  35652=>"111111111",
  35653=>"000011111",
  35654=>"000001111",
  35655=>"000000111",
  35656=>"000000100",
  35657=>"000000000",
  35658=>"100111111",
  35659=>"000011001",
  35660=>"001001001",
  35661=>"111000000",
  35662=>"000000011",
  35663=>"001111111",
  35664=>"111111111",
  35665=>"000000001",
  35666=>"111011111",
  35667=>"000010000",
  35668=>"101111000",
  35669=>"011011001",
  35670=>"100000111",
  35671=>"000000111",
  35672=>"000001101",
  35673=>"011000101",
  35674=>"111111111",
  35675=>"000000111",
  35676=>"111000000",
  35677=>"111111100",
  35678=>"000110111",
  35679=>"111111000",
  35680=>"110111001",
  35681=>"001000000",
  35682=>"111110100",
  35683=>"001001101",
  35684=>"101111001",
  35685=>"000000010",
  35686=>"111111111",
  35687=>"111000001",
  35688=>"000000000",
  35689=>"000011011",
  35690=>"110110000",
  35691=>"111110000",
  35692=>"000000000",
  35693=>"111111010",
  35694=>"000100111",
  35695=>"000000001",
  35696=>"000100001",
  35697=>"000000000",
  35698=>"000000111",
  35699=>"111111101",
  35700=>"000000000",
  35701=>"000000111",
  35702=>"000100111",
  35703=>"000000000",
  35704=>"000001001",
  35705=>"011111111",
  35706=>"111111110",
  35707=>"111111111",
  35708=>"000100100",
  35709=>"100000100",
  35710=>"111000000",
  35711=>"101101100",
  35712=>"111011000",
  35713=>"111111111",
  35714=>"111111111",
  35715=>"000000000",
  35716=>"111111111",
  35717=>"000000010",
  35718=>"000000000",
  35719=>"000111111",
  35720=>"000011111",
  35721=>"100100101",
  35722=>"000000000",
  35723=>"111111000",
  35724=>"111111111",
  35725=>"000100110",
  35726=>"000000001",
  35727=>"111111100",
  35728=>"010010000",
  35729=>"000001111",
  35730=>"110111111",
  35731=>"111111110",
  35732=>"011111111",
  35733=>"000010000",
  35734=>"111010000",
  35735=>"000000111",
  35736=>"110110111",
  35737=>"000000100",
  35738=>"111111111",
  35739=>"111001000",
  35740=>"111111110",
  35741=>"110110000",
  35742=>"111000101",
  35743=>"111000000",
  35744=>"111111000",
  35745=>"011011011",
  35746=>"000000000",
  35747=>"000000011",
  35748=>"111111000",
  35749=>"010111111",
  35750=>"001001111",
  35751=>"110111000",
  35752=>"100000100",
  35753=>"000000010",
  35754=>"111111110",
  35755=>"011010000",
  35756=>"000000000",
  35757=>"000000000",
  35758=>"000111111",
  35759=>"101000000",
  35760=>"110111111",
  35761=>"000001111",
  35762=>"000000111",
  35763=>"000000000",
  35764=>"110000000",
  35765=>"000000111",
  35766=>"000000000",
  35767=>"000000111",
  35768=>"000000001",
  35769=>"111100110",
  35770=>"111111000",
  35771=>"011111100",
  35772=>"000000000",
  35773=>"111111111",
  35774=>"111101000",
  35775=>"000100110",
  35776=>"111111111",
  35777=>"111101000",
  35778=>"111111111",
  35779=>"001001111",
  35780=>"000000001",
  35781=>"101111111",
  35782=>"000000100",
  35783=>"010011111",
  35784=>"000100100",
  35785=>"000100111",
  35786=>"000000001",
  35787=>"001111111",
  35788=>"111111100",
  35789=>"000000000",
  35790=>"000000001",
  35791=>"000111011",
  35792=>"000110000",
  35793=>"100100000",
  35794=>"000110110",
  35795=>"111111111",
  35796=>"101101101",
  35797=>"111001110",
  35798=>"011011000",
  35799=>"111111111",
  35800=>"001000011",
  35801=>"110010010",
  35802=>"111111000",
  35803=>"001000111",
  35804=>"111000001",
  35805=>"111111110",
  35806=>"111111101",
  35807=>"000000101",
  35808=>"111000000",
  35809=>"000000111",
  35810=>"000000000",
  35811=>"000000111",
  35812=>"111000000",
  35813=>"000000100",
  35814=>"000000100",
  35815=>"000110000",
  35816=>"000000111",
  35817=>"101111111",
  35818=>"111010000",
  35819=>"111111000",
  35820=>"000000000",
  35821=>"000000001",
  35822=>"100000110",
  35823=>"000110110",
  35824=>"111111111",
  35825=>"011111010",
  35826=>"000110111",
  35827=>"000000001",
  35828=>"010000010",
  35829=>"000000000",
  35830=>"111001100",
  35831=>"111111100",
  35832=>"111111111",
  35833=>"000000001",
  35834=>"000000010",
  35835=>"001101111",
  35836=>"111111000",
  35837=>"111000011",
  35838=>"111111110",
  35839=>"111111111",
  35840=>"001011111",
  35841=>"000000000",
  35842=>"111111111",
  35843=>"000000000",
  35844=>"100100100",
  35845=>"011111111",
  35846=>"000000000",
  35847=>"111000000",
  35848=>"111010100",
  35849=>"011011011",
  35850=>"111111111",
  35851=>"111100000",
  35852=>"000101111",
  35853=>"000010111",
  35854=>"101111111",
  35855=>"111111111",
  35856=>"111111111",
  35857=>"000000000",
  35858=>"010011000",
  35859=>"111000000",
  35860=>"111111000",
  35861=>"010000111",
  35862=>"000000010",
  35863=>"110111111",
  35864=>"111110111",
  35865=>"000010000",
  35866=>"111111111",
  35867=>"001000111",
  35868=>"000111111",
  35869=>"000000000",
  35870=>"111110100",
  35871=>"000000100",
  35872=>"010010000",
  35873=>"111111111",
  35874=>"000100000",
  35875=>"000000000",
  35876=>"011011011",
  35877=>"000000100",
  35878=>"111111010",
  35879=>"000111111",
  35880=>"111010000",
  35881=>"000000000",
  35882=>"000000111",
  35883=>"111111111",
  35884=>"000000000",
  35885=>"101101001",
  35886=>"001000000",
  35887=>"111111111",
  35888=>"010000000",
  35889=>"000000000",
  35890=>"000100111",
  35891=>"000100111",
  35892=>"000000000",
  35893=>"000000000",
  35894=>"011111110",
  35895=>"110111111",
  35896=>"111111111",
  35897=>"111101111",
  35898=>"000001001",
  35899=>"000000000",
  35900=>"100000000",
  35901=>"010000100",
  35902=>"011110111",
  35903=>"001101111",
  35904=>"111101111",
  35905=>"100100000",
  35906=>"000000000",
  35907=>"111111101",
  35908=>"110110110",
  35909=>"011111111",
  35910=>"111111111",
  35911=>"111111111",
  35912=>"110100100",
  35913=>"000000001",
  35914=>"111111111",
  35915=>"111110100",
  35916=>"000000000",
  35917=>"010000000",
  35918=>"000000000",
  35919=>"111111111",
  35920=>"111000000",
  35921=>"111111111",
  35922=>"011010000",
  35923=>"000000000",
  35924=>"000000111",
  35925=>"010110110",
  35926=>"111111111",
  35927=>"100000000",
  35928=>"001011111",
  35929=>"000000000",
  35930=>"111011001",
  35931=>"000000000",
  35932=>"000100111",
  35933=>"111111111",
  35934=>"111111111",
  35935=>"000000000",
  35936=>"000000000",
  35937=>"000000000",
  35938=>"010000000",
  35939=>"100110111",
  35940=>"000000000",
  35941=>"000010111",
  35942=>"111111110",
  35943=>"000000000",
  35944=>"111111111",
  35945=>"000000000",
  35946=>"110000000",
  35947=>"000000000",
  35948=>"111111111",
  35949=>"011000000",
  35950=>"111111111",
  35951=>"000000000",
  35952=>"000000000",
  35953=>"101110000",
  35954=>"111001001",
  35955=>"100111101",
  35956=>"110111111",
  35957=>"000000110",
  35958=>"001000000",
  35959=>"011000000",
  35960=>"000000000",
  35961=>"111000000",
  35962=>"100100000",
  35963=>"111000111",
  35964=>"111001111",
  35965=>"000000000",
  35966=>"100000000",
  35967=>"000000000",
  35968=>"111011001",
  35969=>"111111111",
  35970=>"111111111",
  35971=>"000000011",
  35972=>"111111111",
  35973=>"000000000",
  35974=>"111111110",
  35975=>"011111000",
  35976=>"111001000",
  35977=>"110011000",
  35978=>"000000000",
  35979=>"111111111",
  35980=>"001000011",
  35981=>"010010000",
  35982=>"100100110",
  35983=>"000000000",
  35984=>"000111111",
  35985=>"000000100",
  35986=>"011000000",
  35987=>"111011111",
  35988=>"000000111",
  35989=>"111010000",
  35990=>"111000111",
  35991=>"101100000",
  35992=>"000000000",
  35993=>"111111111",
  35994=>"000000111",
  35995=>"111111111",
  35996=>"010111111",
  35997=>"001001101",
  35998=>"000000111",
  35999=>"111111111",
  36000=>"011000000",
  36001=>"100100000",
  36002=>"000000000",
  36003=>"111000111",
  36004=>"000000000",
  36005=>"000000000",
  36006=>"101101101",
  36007=>"010110111",
  36008=>"111111110",
  36009=>"101100100",
  36010=>"111111111",
  36011=>"111010110",
  36012=>"011011000",
  36013=>"101101111",
  36014=>"011001000",
  36015=>"000100110",
  36016=>"100111111",
  36017=>"000000000",
  36018=>"101111000",
  36019=>"100000001",
  36020=>"000000000",
  36021=>"000000000",
  36022=>"000100100",
  36023=>"000000001",
  36024=>"111111110",
  36025=>"110111111",
  36026=>"000110110",
  36027=>"110000100",
  36028=>"111001001",
  36029=>"100111111",
  36030=>"111111011",
  36031=>"111110010",
  36032=>"111111111",
  36033=>"000000000",
  36034=>"111001000",
  36035=>"111000000",
  36036=>"000000001",
  36037=>"000001011",
  36038=>"000000000",
  36039=>"011111110",
  36040=>"000010000",
  36041=>"110100111",
  36042=>"010000000",
  36043=>"000011000",
  36044=>"101111101",
  36045=>"000111101",
  36046=>"000000101",
  36047=>"000000000",
  36048=>"011011111",
  36049=>"000110111",
  36050=>"111111111",
  36051=>"011111111",
  36052=>"000000011",
  36053=>"111101100",
  36054=>"111111111",
  36055=>"000000000",
  36056=>"001000000",
  36057=>"111100000",
  36058=>"010011011",
  36059=>"101001111",
  36060=>"000000000",
  36061=>"111110111",
  36062=>"001001000",
  36063=>"111111011",
  36064=>"101000000",
  36065=>"000000000",
  36066=>"000000001",
  36067=>"110111111",
  36068=>"000000000",
  36069=>"110110111",
  36070=>"010110110",
  36071=>"011111000",
  36072=>"011111111",
  36073=>"001000111",
  36074=>"000000000",
  36075=>"111000100",
  36076=>"000111111",
  36077=>"111011011",
  36078=>"111111111",
  36079=>"101101000",
  36080=>"110111111",
  36081=>"111101000",
  36082=>"110111111",
  36083=>"101000000",
  36084=>"000000000",
  36085=>"100000011",
  36086=>"110111000",
  36087=>"000000000",
  36088=>"111111000",
  36089=>"000100100",
  36090=>"111111111",
  36091=>"111111111",
  36092=>"000001001",
  36093=>"111011111",
  36094=>"111111111",
  36095=>"011000000",
  36096=>"100000000",
  36097=>"111000000",
  36098=>"000000000",
  36099=>"111111111",
  36100=>"111111011",
  36101=>"111111111",
  36102=>"111110000",
  36103=>"001101111",
  36104=>"110111111",
  36105=>"000100100",
  36106=>"111111111",
  36107=>"111111111",
  36108=>"000011101",
  36109=>"001000101",
  36110=>"000000000",
  36111=>"100000000",
  36112=>"111111111",
  36113=>"010111111",
  36114=>"000000000",
  36115=>"111111100",
  36116=>"111000011",
  36117=>"000111111",
  36118=>"101100111",
  36119=>"000000110",
  36120=>"000101110",
  36121=>"111100110",
  36122=>"001101101",
  36123=>"000000000",
  36124=>"101101111",
  36125=>"000010000",
  36126=>"000000000",
  36127=>"000010010",
  36128=>"000100001",
  36129=>"111111111",
  36130=>"000100111",
  36131=>"011011110",
  36132=>"111111011",
  36133=>"000000000",
  36134=>"001100100",
  36135=>"101001001",
  36136=>"000000110",
  36137=>"000000010",
  36138=>"000000000",
  36139=>"100110001",
  36140=>"100000000",
  36141=>"001001111",
  36142=>"000000000",
  36143=>"000000000",
  36144=>"101101111",
  36145=>"000000000",
  36146=>"111111111",
  36147=>"000011111",
  36148=>"001000000",
  36149=>"111100101",
  36150=>"111111000",
  36151=>"110011011",
  36152=>"000000000",
  36153=>"010000000",
  36154=>"000111111",
  36155=>"100011111",
  36156=>"011111110",
  36157=>"000100111",
  36158=>"000000000",
  36159=>"111111111",
  36160=>"000000000",
  36161=>"000000000",
  36162=>"011001000",
  36163=>"110000110",
  36164=>"111110100",
  36165=>"100000110",
  36166=>"011111111",
  36167=>"111010000",
  36168=>"000000000",
  36169=>"111000000",
  36170=>"000000000",
  36171=>"111100000",
  36172=>"110010011",
  36173=>"011110000",
  36174=>"110000000",
  36175=>"011011000",
  36176=>"000000000",
  36177=>"011000000",
  36178=>"001001101",
  36179=>"110111111",
  36180=>"001000000",
  36181=>"011011011",
  36182=>"000000000",
  36183=>"100100111",
  36184=>"111111111",
  36185=>"100000000",
  36186=>"000000010",
  36187=>"000000000",
  36188=>"100111111",
  36189=>"000111111",
  36190=>"101001000",
  36191=>"000000000",
  36192=>"101000000",
  36193=>"000000100",
  36194=>"101101100",
  36195=>"000000001",
  36196=>"000000000",
  36197=>"111111001",
  36198=>"111111000",
  36199=>"010100100",
  36200=>"011000001",
  36201=>"110110110",
  36202=>"000000010",
  36203=>"111111100",
  36204=>"000000000",
  36205=>"111111101",
  36206=>"111000000",
  36207=>"000000000",
  36208=>"000000100",
  36209=>"100001000",
  36210=>"000000100",
  36211=>"000000000",
  36212=>"110001001",
  36213=>"011000000",
  36214=>"000110110",
  36215=>"111111111",
  36216=>"000000000",
  36217=>"111111111",
  36218=>"111111111",
  36219=>"000001010",
  36220=>"011111111",
  36221=>"111111111",
  36222=>"000000001",
  36223=>"000000000",
  36224=>"110000000",
  36225=>"011111100",
  36226=>"100011011",
  36227=>"100110000",
  36228=>"000000000",
  36229=>"000000000",
  36230=>"011000000",
  36231=>"111111011",
  36232=>"000000001",
  36233=>"011111111",
  36234=>"111000110",
  36235=>"100000100",
  36236=>"111111111",
  36237=>"001010100",
  36238=>"000000010",
  36239=>"000000000",
  36240=>"000100100",
  36241=>"100000000",
  36242=>"100000000",
  36243=>"111111111",
  36244=>"111111111",
  36245=>"000000000",
  36246=>"001111111",
  36247=>"111001111",
  36248=>"000111001",
  36249=>"000000000",
  36250=>"111111111",
  36251=>"001111111",
  36252=>"011111111",
  36253=>"001000000",
  36254=>"000000000",
  36255=>"000000000",
  36256=>"111111001",
  36257=>"100001111",
  36258=>"101110110",
  36259=>"000010111",
  36260=>"111111110",
  36261=>"000000000",
  36262=>"111111111",
  36263=>"000000000",
  36264=>"100000111",
  36265=>"111111100",
  36266=>"011111110",
  36267=>"100100001",
  36268=>"011000000",
  36269=>"000100110",
  36270=>"010111111",
  36271=>"111111111",
  36272=>"000000000",
  36273=>"110100110",
  36274=>"000001001",
  36275=>"000000000",
  36276=>"011111111",
  36277=>"011010001",
  36278=>"110000000",
  36279=>"000000000",
  36280=>"000110110",
  36281=>"111111111",
  36282=>"110000110",
  36283=>"110010011",
  36284=>"111101111",
  36285=>"000110100",
  36286=>"111101000",
  36287=>"000000000",
  36288=>"110000111",
  36289=>"000000000",
  36290=>"001000000",
  36291=>"111110111",
  36292=>"101100000",
  36293=>"001000000",
  36294=>"000000000",
  36295=>"000001111",
  36296=>"000000000",
  36297=>"000000111",
  36298=>"101000111",
  36299=>"000000000",
  36300=>"000000000",
  36301=>"111011111",
  36302=>"000000000",
  36303=>"111101101",
  36304=>"100111111",
  36305=>"000000010",
  36306=>"111111111",
  36307=>"000000000",
  36308=>"000000001",
  36309=>"111011000",
  36310=>"100000011",
  36311=>"001011011",
  36312=>"001000000",
  36313=>"010000000",
  36314=>"110111111",
  36315=>"111111111",
  36316=>"110110010",
  36317=>"111100100",
  36318=>"000000000",
  36319=>"001101111",
  36320=>"111111111",
  36321=>"000111111",
  36322=>"111111111",
  36323=>"111111110",
  36324=>"111111111",
  36325=>"000000110",
  36326=>"000000111",
  36327=>"111111111",
  36328=>"000000000",
  36329=>"111111000",
  36330=>"111101100",
  36331=>"100100000",
  36332=>"111001111",
  36333=>"100100111",
  36334=>"000000001",
  36335=>"011011001",
  36336=>"000110110",
  36337=>"000010000",
  36338=>"111111111",
  36339=>"000000000",
  36340=>"000000000",
  36341=>"000000000",
  36342=>"001111111",
  36343=>"111011111",
  36344=>"000000000",
  36345=>"001001001",
  36346=>"111110100",
  36347=>"011001001",
  36348=>"110111111",
  36349=>"011001000",
  36350=>"111111111",
  36351=>"000000000",
  36352=>"001011011",
  36353=>"111111101",
  36354=>"111111111",
  36355=>"110111111",
  36356=>"111111111",
  36357=>"001100110",
  36358=>"001001000",
  36359=>"000000001",
  36360=>"000011001",
  36361=>"010011011",
  36362=>"111111111",
  36363=>"001011111",
  36364=>"000000000",
  36365=>"100111110",
  36366=>"000001011",
  36367=>"010110011",
  36368=>"111100111",
  36369=>"000011101",
  36370=>"000000100",
  36371=>"100111111",
  36372=>"000000011",
  36373=>"011011011",
  36374=>"000000011",
  36375=>"000000000",
  36376=>"111111111",
  36377=>"000110110",
  36378=>"111010111",
  36379=>"010000011",
  36380=>"111111100",
  36381=>"111111011",
  36382=>"100011000",
  36383=>"100100110",
  36384=>"000000001",
  36385=>"000010110",
  36386=>"000000001",
  36387=>"111111111",
  36388=>"111111111",
  36389=>"101111111",
  36390=>"111011011",
  36391=>"000000000",
  36392=>"000000011",
  36393=>"000000000",
  36394=>"111111111",
  36395=>"000100110",
  36396=>"111100101",
  36397=>"111111011",
  36398=>"100100100",
  36399=>"000000000",
  36400=>"010000000",
  36401=>"000000000",
  36402=>"111000000",
  36403=>"101101101",
  36404=>"100000000",
  36405=>"000010010",
  36406=>"111111111",
  36407=>"001001000",
  36408=>"101000110",
  36409=>"000110111",
  36410=>"000000000",
  36411=>"111111111",
  36412=>"100000001",
  36413=>"000000011",
  36414=>"000100100",
  36415=>"000000001",
  36416=>"000000111",
  36417=>"010100001",
  36418=>"111111111",
  36419=>"011011000",
  36420=>"111001011",
  36421=>"000000000",
  36422=>"001000000",
  36423=>"011001000",
  36424=>"110000011",
  36425=>"010000000",
  36426=>"111111101",
  36427=>"111111111",
  36428=>"000000000",
  36429=>"111111111",
  36430=>"000001111",
  36431=>"000000000",
  36432=>"100000100",
  36433=>"010011011",
  36434=>"001001100",
  36435=>"000000010",
  36436=>"100000000",
  36437=>"111111000",
  36438=>"111111101",
  36439=>"111101111",
  36440=>"000000110",
  36441=>"111111000",
  36442=>"011110000",
  36443=>"111011000",
  36444=>"000000000",
  36445=>"110000001",
  36446=>"111000110",
  36447=>"101101001",
  36448=>"000000001",
  36449=>"000000000",
  36450=>"000000000",
  36451=>"111111111",
  36452=>"011111110",
  36453=>"000000111",
  36454=>"000111100",
  36455=>"010010111",
  36456=>"110000000",
  36457=>"111111011",
  36458=>"000000010",
  36459=>"010111111",
  36460=>"000011110",
  36461=>"000000000",
  36462=>"100000000",
  36463=>"010000011",
  36464=>"100101111",
  36465=>"111111111",
  36466=>"111100000",
  36467=>"000000000",
  36468=>"000000000",
  36469=>"000000000",
  36470=>"011000000",
  36471=>"001000110",
  36472=>"000110100",
  36473=>"000001111",
  36474=>"111111001",
  36475=>"111111111",
  36476=>"110110110",
  36477=>"111100001",
  36478=>"111111001",
  36479=>"000110000",
  36480=>"000000000",
  36481=>"000001001",
  36482=>"000110000",
  36483=>"010111011",
  36484=>"111000001",
  36485=>"111111111",
  36486=>"011111100",
  36487=>"000010111",
  36488=>"111101001",
  36489=>"111000000",
  36490=>"000010000",
  36491=>"111111111",
  36492=>"001011110",
  36493=>"000000000",
  36494=>"111100111",
  36495=>"100000011",
  36496=>"001001001",
  36497=>"000100100",
  36498=>"011000000",
  36499=>"010000000",
  36500=>"111111111",
  36501=>"000000111",
  36502=>"111111111",
  36503=>"000000000",
  36504=>"000000000",
  36505=>"000010011",
  36506=>"000000000",
  36507=>"011011011",
  36508=>"110101100",
  36509=>"000000000",
  36510=>"000000011",
  36511=>"111111011",
  36512=>"001000000",
  36513=>"001101101",
  36514=>"000000000",
  36515=>"101100011",
  36516=>"011111111",
  36517=>"011000000",
  36518=>"111111101",
  36519=>"100110111",
  36520=>"001001000",
  36521=>"000010000",
  36522=>"000000000",
  36523=>"111110111",
  36524=>"000000111",
  36525=>"111000000",
  36526=>"000000000",
  36527=>"011001111",
  36528=>"000011000",
  36529=>"000000000",
  36530=>"011011000",
  36531=>"101000111",
  36532=>"011000000",
  36533=>"101001000",
  36534=>"011000001",
  36535=>"100000000",
  36536=>"111111111",
  36537=>"110000011",
  36538=>"000000010",
  36539=>"000001111",
  36540=>"111111111",
  36541=>"000000000",
  36542=>"100000000",
  36543=>"000000011",
  36544=>"000000100",
  36545=>"011011111",
  36546=>"111111111",
  36547=>"011100111",
  36548=>"000000000",
  36549=>"000000000",
  36550=>"000011111",
  36551=>"111111111",
  36552=>"000000110",
  36553=>"000000110",
  36554=>"100011011",
  36555=>"000000000",
  36556=>"000001001",
  36557=>"110111000",
  36558=>"000000100",
  36559=>"000100011",
  36560=>"000000000",
  36561=>"011111111",
  36562=>"111111110",
  36563=>"000000100",
  36564=>"110100110",
  36565=>"010110010",
  36566=>"001011111",
  36567=>"000000011",
  36568=>"111111110",
  36569=>"001000000",
  36570=>"111011110",
  36571=>"111111110",
  36572=>"101000000",
  36573=>"111111111",
  36574=>"111111111",
  36575=>"100111111",
  36576=>"000000000",
  36577=>"110100100",
  36578=>"111111111",
  36579=>"111111111",
  36580=>"111111111",
  36581=>"001000000",
  36582=>"111000000",
  36583=>"000000011",
  36584=>"111001110",
  36585=>"010000000",
  36586=>"100100111",
  36587=>"000000000",
  36588=>"111111111",
  36589=>"111100000",
  36590=>"000000000",
  36591=>"111001000",
  36592=>"111111111",
  36593=>"000001011",
  36594=>"000001101",
  36595=>"100001011",
  36596=>"111000000",
  36597=>"000000000",
  36598=>"001001100",
  36599=>"000100111",
  36600=>"111111111",
  36601=>"111111111",
  36602=>"000111111",
  36603=>"100000000",
  36604=>"000001111",
  36605=>"001000000",
  36606=>"111011000",
  36607=>"011000000",
  36608=>"000000010",
  36609=>"000000000",
  36610=>"000000000",
  36611=>"110111111",
  36612=>"100100100",
  36613=>"110111111",
  36614=>"111000110",
  36615=>"011111100",
  36616=>"111111111",
  36617=>"000000000",
  36618=>"111111111",
  36619=>"111111110",
  36620=>"111011000",
  36621=>"111111110",
  36622=>"111111111",
  36623=>"000000000",
  36624=>"111101001",
  36625=>"000000000",
  36626=>"000000110",
  36627=>"001001110",
  36628=>"001011000",
  36629=>"011111100",
  36630=>"001001110",
  36631=>"001001111",
  36632=>"110111100",
  36633=>"111100000",
  36634=>"000000000",
  36635=>"111111111",
  36636=>"111001000",
  36637=>"110111111",
  36638=>"111111111",
  36639=>"000000111",
  36640=>"110111011",
  36641=>"110111111",
  36642=>"011001100",
  36643=>"000000000",
  36644=>"011001101",
  36645=>"111111001",
  36646=>"000111111",
  36647=>"101001111",
  36648=>"101111000",
  36649=>"100000111",
  36650=>"100100100",
  36651=>"111111111",
  36652=>"111010000",
  36653=>"000111101",
  36654=>"000000000",
  36655=>"110011011",
  36656=>"110000000",
  36657=>"000010011",
  36658=>"001100111",
  36659=>"010000000",
  36660=>"111111111",
  36661=>"100100111",
  36662=>"011001000",
  36663=>"000000000",
  36664=>"000000000",
  36665=>"111001111",
  36666=>"000111011",
  36667=>"111111000",
  36668=>"111111111",
  36669=>"111100100",
  36670=>"010100101",
  36671=>"000111011",
  36672=>"000000000",
  36673=>"100100000",
  36674=>"000000000",
  36675=>"010000000",
  36676=>"111111111",
  36677=>"000000000",
  36678=>"100100101",
  36679=>"100000000",
  36680=>"111011011",
  36681=>"000010000",
  36682=>"001101000",
  36683=>"011001001",
  36684=>"111001011",
  36685=>"011000000",
  36686=>"011011111",
  36687=>"101001001",
  36688=>"100100100",
  36689=>"000000000",
  36690=>"111010111",
  36691=>"100110111",
  36692=>"000000000",
  36693=>"001001001",
  36694=>"000110110",
  36695=>"110000000",
  36696=>"000000000",
  36697=>"000001111",
  36698=>"110111000",
  36699=>"100111111",
  36700=>"111111111",
  36701=>"000110111",
  36702=>"011111000",
  36703=>"000010111",
  36704=>"011000000",
  36705=>"110101111",
  36706=>"011110110",
  36707=>"110101101",
  36708=>"100001111",
  36709=>"000000111",
  36710=>"000110110",
  36711=>"000000000",
  36712=>"100100100",
  36713=>"110110000",
  36714=>"000000000",
  36715=>"111111100",
  36716=>"110000110",
  36717=>"100111111",
  36718=>"000100000",
  36719=>"111101111",
  36720=>"100100100",
  36721=>"111111111",
  36722=>"100000000",
  36723=>"000000011",
  36724=>"011011000",
  36725=>"001001000",
  36726=>"011000111",
  36727=>"111111000",
  36728=>"111111111",
  36729=>"111111111",
  36730=>"000111111",
  36731=>"110011011",
  36732=>"010111100",
  36733=>"111000001",
  36734=>"011000001",
  36735=>"000000000",
  36736=>"000000000",
  36737=>"011000000",
  36738=>"001001111",
  36739=>"000000111",
  36740=>"000010000",
  36741=>"101101100",
  36742=>"111111101",
  36743=>"000001011",
  36744=>"010111111",
  36745=>"111111011",
  36746=>"111111111",
  36747=>"000000000",
  36748=>"000000111",
  36749=>"000000000",
  36750=>"111001011",
  36751=>"111000000",
  36752=>"111111101",
  36753=>"111101111",
  36754=>"111111110",
  36755=>"111110110",
  36756=>"000001011",
  36757=>"010010000",
  36758=>"011011111",
  36759=>"000110111",
  36760=>"000000101",
  36761=>"101001111",
  36762=>"000111111",
  36763=>"000000000",
  36764=>"111011111",
  36765=>"001000000",
  36766=>"101100100",
  36767=>"111111111",
  36768=>"000001011",
  36769=>"000100000",
  36770=>"100111111",
  36771=>"011011001",
  36772=>"110110111",
  36773=>"000000000",
  36774=>"000000000",
  36775=>"010000000",
  36776=>"111000000",
  36777=>"110001001",
  36778=>"111111111",
  36779=>"000100111",
  36780=>"011000000",
  36781=>"000000000",
  36782=>"000000000",
  36783=>"111111111",
  36784=>"000010110",
  36785=>"111111111",
  36786=>"101111011",
  36787=>"111111101",
  36788=>"101111111",
  36789=>"000000010",
  36790=>"111111111",
  36791=>"111111000",
  36792=>"111111100",
  36793=>"001001001",
  36794=>"000001000",
  36795=>"000000100",
  36796=>"000001111",
  36797=>"000000000",
  36798=>"000100100",
  36799=>"111100100",
  36800=>"100111111",
  36801=>"000000000",
  36802=>"111101111",
  36803=>"000100111",
  36804=>"110000000",
  36805=>"100111001",
  36806=>"011111000",
  36807=>"111100101",
  36808=>"000100000",
  36809=>"000101000",
  36810=>"100110110",
  36811=>"111111111",
  36812=>"100100000",
  36813=>"101100110",
  36814=>"110000000",
  36815=>"101111111",
  36816=>"111111001",
  36817=>"000000000",
  36818=>"111010001",
  36819=>"011011111",
  36820=>"111111111",
  36821=>"111111111",
  36822=>"001101111",
  36823=>"000000000",
  36824=>"111111111",
  36825=>"111111111",
  36826=>"100000000",
  36827=>"000000000",
  36828=>"111111101",
  36829=>"001000000",
  36830=>"010000000",
  36831=>"011011111",
  36832=>"000000001",
  36833=>"011111111",
  36834=>"111111111",
  36835=>"101001111",
  36836=>"000000111",
  36837=>"111111001",
  36838=>"000000000",
  36839=>"010111011",
  36840=>"100101011",
  36841=>"000000000",
  36842=>"111100101",
  36843=>"000000001",
  36844=>"001111001",
  36845=>"100000111",
  36846=>"000110111",
  36847=>"111111111",
  36848=>"000000011",
  36849=>"100000000",
  36850=>"111100111",
  36851=>"110000111",
  36852=>"001011111",
  36853=>"100001000",
  36854=>"010000011",
  36855=>"000000000",
  36856=>"111101011",
  36857=>"000001000",
  36858=>"000110110",
  36859=>"111111111",
  36860=>"100111111",
  36861=>"111100111",
  36862=>"100100000",
  36863=>"110111011",
  36864=>"111111111",
  36865=>"011001111",
  36866=>"111111111",
  36867=>"000000000",
  36868=>"000111111",
  36869=>"101111111",
  36870=>"000000000",
  36871=>"000000111",
  36872=>"111101000",
  36873=>"000000000",
  36874=>"110100000",
  36875=>"100100110",
  36876=>"000111001",
  36877=>"110100000",
  36878=>"000100010",
  36879=>"111011111",
  36880=>"000010110",
  36881=>"011100000",
  36882=>"111111111",
  36883=>"000000110",
  36884=>"110111111",
  36885=>"111101000",
  36886=>"110000111",
  36887=>"110000111",
  36888=>"010000100",
  36889=>"011011111",
  36890=>"000000000",
  36891=>"111011000",
  36892=>"111010000",
  36893=>"111000000",
  36894=>"000000000",
  36895=>"110100100",
  36896=>"000000000",
  36897=>"000000100",
  36898=>"111111111",
  36899=>"010111111",
  36900=>"000000000",
  36901=>"100101011",
  36902=>"000000001",
  36903=>"111000000",
  36904=>"000000000",
  36905=>"111111000",
  36906=>"111011111",
  36907=>"110000000",
  36908=>"000000000",
  36909=>"111111111",
  36910=>"000000001",
  36911=>"011001000",
  36912=>"000000001",
  36913=>"011111111",
  36914=>"000000000",
  36915=>"111011000",
  36916=>"011111111",
  36917=>"000000001",
  36918=>"000000000",
  36919=>"101111000",
  36920=>"010000000",
  36921=>"000011111",
  36922=>"110110110",
  36923=>"000000010",
  36924=>"000001011",
  36925=>"000000000",
  36926=>"110100100",
  36927=>"110000000",
  36928=>"000001001",
  36929=>"100100000",
  36930=>"001001000",
  36931=>"000000000",
  36932=>"000000000",
  36933=>"000000000",
  36934=>"000000111",
  36935=>"111111110",
  36936=>"010010011",
  36937=>"000000001",
  36938=>"111111111",
  36939=>"110011011",
  36940=>"000001001",
  36941=>"111111101",
  36942=>"111000011",
  36943=>"000000000",
  36944=>"111111111",
  36945=>"000000000",
  36946=>"000010000",
  36947=>"000001011",
  36948=>"111111111",
  36949=>"110110000",
  36950=>"011010000",
  36951=>"000000100",
  36952=>"011011000",
  36953=>"111000000",
  36954=>"000000000",
  36955=>"000010001",
  36956=>"000000000",
  36957=>"000000101",
  36958=>"111100001",
  36959=>"000000000",
  36960=>"010110000",
  36961=>"000000000",
  36962=>"000011010",
  36963=>"000000000",
  36964=>"110100110",
  36965=>"111111001",
  36966=>"111001000",
  36967=>"110111001",
  36968=>"111111111",
  36969=>"111111111",
  36970=>"000110111",
  36971=>"100111111",
  36972=>"011011001",
  36973=>"000000000",
  36974=>"000000101",
  36975=>"000000001",
  36976=>"111111000",
  36977=>"001001000",
  36978=>"011111111",
  36979=>"000000000",
  36980=>"111111111",
  36981=>"000110000",
  36982=>"110000000",
  36983=>"000000000",
  36984=>"111111111",
  36985=>"100001111",
  36986=>"000000000",
  36987=>"110111111",
  36988=>"001011001",
  36989=>"111111000",
  36990=>"000000000",
  36991=>"000000000",
  36992=>"111111111",
  36993=>"111111111",
  36994=>"000000111",
  36995=>"100110100",
  36996=>"011000000",
  36997=>"111111100",
  36998=>"111111001",
  36999=>"000000000",
  37000=>"010010110",
  37001=>"001110000",
  37002=>"000000000",
  37003=>"111011000",
  37004=>"111111100",
  37005=>"011111111",
  37006=>"001000100",
  37007=>"000000000",
  37008=>"111011000",
  37009=>"111111111",
  37010=>"000010000",
  37011=>"111110111",
  37012=>"100111011",
  37013=>"000000111",
  37014=>"000000000",
  37015=>"000000000",
  37016=>"111111001",
  37017=>"101100100",
  37018=>"000000000",
  37019=>"100000000",
  37020=>"111111111",
  37021=>"000000000",
  37022=>"001001111",
  37023=>"111011011",
  37024=>"000011010",
  37025=>"111101110",
  37026=>"111000001",
  37027=>"100000000",
  37028=>"000000000",
  37029=>"001000000",
  37030=>"111111011",
  37031=>"100100100",
  37032=>"000000000",
  37033=>"001000001",
  37034=>"001000000",
  37035=>"111111111",
  37036=>"000000000",
  37037=>"000100000",
  37038=>"111110000",
  37039=>"111101000",
  37040=>"111111111",
  37041=>"000100101",
  37042=>"111111111",
  37043=>"111000000",
  37044=>"011000000",
  37045=>"111111111",
  37046=>"111100100",
  37047=>"111111111",
  37048=>"111111111",
  37049=>"111111111",
  37050=>"000000000",
  37051=>"011111111",
  37052=>"010010111",
  37053=>"111110000",
  37054=>"111111000",
  37055=>"111111111",
  37056=>"111011011",
  37057=>"110110111",
  37058=>"111000110",
  37059=>"111111111",
  37060=>"001000110",
  37061=>"000000000",
  37062=>"001001101",
  37063=>"111111111",
  37064=>"111111111",
  37065=>"000000001",
  37066=>"111111011",
  37067=>"110111111",
  37068=>"000000100",
  37069=>"111111100",
  37070=>"000000000",
  37071=>"100111111",
  37072=>"110111111",
  37073=>"000000001",
  37074=>"011000011",
  37075=>"000010111",
  37076=>"011000000",
  37077=>"000000000",
  37078=>"000100100",
  37079=>"111111000",
  37080=>"100100000",
  37081=>"010110110",
  37082=>"111100000",
  37083=>"111111111",
  37084=>"001001011",
  37085=>"000000000",
  37086=>"000111111",
  37087=>"001110100",
  37088=>"111110100",
  37089=>"111111111",
  37090=>"001000001",
  37091=>"001000000",
  37092=>"111100100",
  37093=>"000000000",
  37094=>"101101101",
  37095=>"000110111",
  37096=>"000000000",
  37097=>"000010110",
  37098=>"001000000",
  37099=>"111111111",
  37100=>"001000100",
  37101=>"111111111",
  37102=>"111111111",
  37103=>"111010000",
  37104=>"111111111",
  37105=>"000100111",
  37106=>"000000001",
  37107=>"001001100",
  37108=>"111111000",
  37109=>"000000000",
  37110=>"111101100",
  37111=>"111011001",
  37112=>"111111111",
  37113=>"111111111",
  37114=>"111111111",
  37115=>"000111111",
  37116=>"000001000",
  37117=>"111010000",
  37118=>"000101111",
  37119=>"000100110",
  37120=>"010110100",
  37121=>"000010011",
  37122=>"000000000",
  37123=>"111111111",
  37124=>"111111111",
  37125=>"011111111",
  37126=>"111011000",
  37127=>"000000100",
  37128=>"000000000",
  37129=>"000000000",
  37130=>"111111011",
  37131=>"000111000",
  37132=>"001001111",
  37133=>"111111000",
  37134=>"111111111",
  37135=>"000111011",
  37136=>"111111111",
  37137=>"111011000",
  37138=>"110100100",
  37139=>"000000000",
  37140=>"000000110",
  37141=>"011111001",
  37142=>"001001100",
  37143=>"000111111",
  37144=>"111111111",
  37145=>"111111100",
  37146=>"000111111",
  37147=>"101111111",
  37148=>"110100100",
  37149=>"111110000",
  37150=>"111111111",
  37151=>"011001001",
  37152=>"100110111",
  37153=>"111111111",
  37154=>"011000001",
  37155=>"000111011",
  37156=>"100111000",
  37157=>"111111111",
  37158=>"111110110",
  37159=>"000000011",
  37160=>"000000001",
  37161=>"111101000",
  37162=>"101000111",
  37163=>"111111111",
  37164=>"000100110",
  37165=>"110010110",
  37166=>"000000100",
  37167=>"011000000",
  37168=>"111001111",
  37169=>"111011111",
  37170=>"111111110",
  37171=>"000000001",
  37172=>"111000000",
  37173=>"000000000",
  37174=>"111111111",
  37175=>"000000000",
  37176=>"001000111",
  37177=>"100001111",
  37178=>"000000000",
  37179=>"000000000",
  37180=>"000000100",
  37181=>"111111111",
  37182=>"111000000",
  37183=>"000000110",
  37184=>"000000000",
  37185=>"100111111",
  37186=>"111111001",
  37187=>"111111111",
  37188=>"110111001",
  37189=>"011000000",
  37190=>"110111111",
  37191=>"111111111",
  37192=>"000000000",
  37193=>"111111000",
  37194=>"111111111",
  37195=>"111111110",
  37196=>"100101100",
  37197=>"000000011",
  37198=>"110110010",
  37199=>"000110110",
  37200=>"000010110",
  37201=>"111111000",
  37202=>"000000000",
  37203=>"001001011",
  37204=>"011111111",
  37205=>"110100100",
  37206=>"000100100",
  37207=>"000000001",
  37208=>"101101000",
  37209=>"111111000",
  37210=>"001111111",
  37211=>"111000101",
  37212=>"000000000",
  37213=>"111111111",
  37214=>"001001111",
  37215=>"111111100",
  37216=>"100000000",
  37217=>"000000001",
  37218=>"000000010",
  37219=>"111111111",
  37220=>"000000000",
  37221=>"011000100",
  37222=>"000000111",
  37223=>"000000000",
  37224=>"111000001",
  37225=>"011111111",
  37226=>"001001111",
  37227=>"000011000",
  37228=>"001001001",
  37229=>"000000110",
  37230=>"111001111",
  37231=>"111111111",
  37232=>"000000000",
  37233=>"000001000",
  37234=>"011000000",
  37235=>"000000110",
  37236=>"100110100",
  37237=>"000111111",
  37238=>"010111000",
  37239=>"100101111",
  37240=>"110100000",
  37241=>"000000100",
  37242=>"000000111",
  37243=>"011011001",
  37244=>"100100110",
  37245=>"011000000",
  37246=>"111111000",
  37247=>"111011011",
  37248=>"011111100",
  37249=>"101000000",
  37250=>"000000000",
  37251=>"100000001",
  37252=>"000000000",
  37253=>"111111111",
  37254=>"110000000",
  37255=>"101101000",
  37256=>"101100000",
  37257=>"110000000",
  37258=>"001101111",
  37259=>"000001111",
  37260=>"001000001",
  37261=>"001001001",
  37262=>"111111111",
  37263=>"001000000",
  37264=>"100111111",
  37265=>"000000000",
  37266=>"011000000",
  37267=>"111111001",
  37268=>"000000000",
  37269=>"100111111",
  37270=>"111110110",
  37271=>"011001011",
  37272=>"011000111",
  37273=>"000100000",
  37274=>"111110000",
  37275=>"000000111",
  37276=>"110111111",
  37277=>"111111001",
  37278=>"111111111",
  37279=>"000000010",
  37280=>"000000000",
  37281=>"001001001",
  37282=>"011000000",
  37283=>"000000111",
  37284=>"000000000",
  37285=>"111111111",
  37286=>"111000000",
  37287=>"111001001",
  37288=>"011100000",
  37289=>"000110111",
  37290=>"111111111",
  37291=>"111011111",
  37292=>"000000010",
  37293=>"110100101",
  37294=>"000011111",
  37295=>"000000100",
  37296=>"000000000",
  37297=>"000000111",
  37298=>"011000000",
  37299=>"000001000",
  37300=>"111111110",
  37301=>"111111111",
  37302=>"000000100",
  37303=>"111110010",
  37304=>"111111000",
  37305=>"111101011",
  37306=>"000000000",
  37307=>"111000000",
  37308=>"011000000",
  37309=>"111111111",
  37310=>"000100111",
  37311=>"111111111",
  37312=>"001000111",
  37313=>"111001101",
  37314=>"000000000",
  37315=>"111000000",
  37316=>"111111111",
  37317=>"000000100",
  37318=>"101111111",
  37319=>"111101101",
  37320=>"011111111",
  37321=>"111111100",
  37322=>"000000011",
  37323=>"000000100",
  37324=>"111111111",
  37325=>"111111111",
  37326=>"001001111",
  37327=>"111000000",
  37328=>"001000011",
  37329=>"101111111",
  37330=>"111111111",
  37331=>"000000000",
  37332=>"100110111",
  37333=>"000111110",
  37334=>"111111111",
  37335=>"100111111",
  37336=>"111001001",
  37337=>"000000000",
  37338=>"111111011",
  37339=>"011000000",
  37340=>"111111111",
  37341=>"001101110",
  37342=>"110001011",
  37343=>"011011111",
  37344=>"010000000",
  37345=>"000000100",
  37346=>"011000000",
  37347=>"011111111",
  37348=>"000000000",
  37349=>"000010010",
  37350=>"111111111",
  37351=>"000000111",
  37352=>"000000000",
  37353=>"111111000",
  37354=>"110111000",
  37355=>"101111111",
  37356=>"110111111",
  37357=>"111111111",
  37358=>"000100111",
  37359=>"000000110",
  37360=>"111111111",
  37361=>"010000000",
  37362=>"111000000",
  37363=>"000000000",
  37364=>"111111111",
  37365=>"111111111",
  37366=>"100000000",
  37367=>"100100110",
  37368=>"000000110",
  37369=>"011011011",
  37370=>"011111111",
  37371=>"111111111",
  37372=>"000000000",
  37373=>"000000001",
  37374=>"000000000",
  37375=>"111111111",
  37376=>"011011111",
  37377=>"011000111",
  37378=>"111111111",
  37379=>"000000000",
  37380=>"111110010",
  37381=>"111000100",
  37382=>"110111111",
  37383=>"000000000",
  37384=>"100000000",
  37385=>"111111000",
  37386=>"010000000",
  37387=>"101100100",
  37388=>"000001000",
  37389=>"111111111",
  37390=>"000000101",
  37391=>"000000000",
  37392=>"100111111",
  37393=>"000101000",
  37394=>"100101111",
  37395=>"010000000",
  37396=>"000000000",
  37397=>"000100100",
  37398=>"111111111",
  37399=>"000000000",
  37400=>"111111001",
  37401=>"010111111",
  37402=>"000000000",
  37403=>"111110110",
  37404=>"111111000",
  37405=>"000111110",
  37406=>"011110110",
  37407=>"111111111",
  37408=>"000001011",
  37409=>"111111111",
  37410=>"000000000",
  37411=>"110010111",
  37412=>"111011111",
  37413=>"001101000",
  37414=>"111110110",
  37415=>"000000111",
  37416=>"110110100",
  37417=>"011111111",
  37418=>"110110110",
  37419=>"111111000",
  37420=>"111100100",
  37421=>"111111000",
  37422=>"111111111",
  37423=>"001001101",
  37424=>"101001001",
  37425=>"000000000",
  37426=>"011011011",
  37427=>"001001111",
  37428=>"100011111",
  37429=>"001000000",
  37430=>"000110000",
  37431=>"000110110",
  37432=>"000000000",
  37433=>"001111000",
  37434=>"111111111",
  37435=>"000000000",
  37436=>"001000000",
  37437=>"111111011",
  37438=>"110100000",
  37439=>"001101111",
  37440=>"111111111",
  37441=>"111101000",
  37442=>"111111000",
  37443=>"111111111",
  37444=>"110000000",
  37445=>"111111110",
  37446=>"000000000",
  37447=>"111111111",
  37448=>"100100100",
  37449=>"111111111",
  37450=>"001111111",
  37451=>"001110100",
  37452=>"111001111",
  37453=>"111111000",
  37454=>"000000111",
  37455=>"000000111",
  37456=>"101111101",
  37457=>"111111101",
  37458=>"111111011",
  37459=>"010000100",
  37460=>"000000100",
  37461=>"100000000",
  37462=>"100000000",
  37463=>"110110110",
  37464=>"000000000",
  37465=>"111100100",
  37466=>"111111100",
  37467=>"111111111",
  37468=>"000001000",
  37469=>"111111111",
  37470=>"111111111",
  37471=>"100001001",
  37472=>"111111111",
  37473=>"100100111",
  37474=>"111000000",
  37475=>"011001100",
  37476=>"110100100",
  37477=>"000000111",
  37478=>"101101111",
  37479=>"000001011",
  37480=>"111111111",
  37481=>"111000000",
  37482=>"000100111",
  37483=>"101000000",
  37484=>"110111111",
  37485=>"000011011",
  37486=>"111111111",
  37487=>"110111111",
  37488=>"011001000",
  37489=>"001111111",
  37490=>"000001001",
  37491=>"001000111",
  37492=>"000000000",
  37493=>"111110100",
  37494=>"111111111",
  37495=>"000000000",
  37496=>"111111111",
  37497=>"000001111",
  37498=>"000000000",
  37499=>"000000000",
  37500=>"111001000",
  37501=>"111111000",
  37502=>"100111111",
  37503=>"110100000",
  37504=>"111111111",
  37505=>"101100000",
  37506=>"000000000",
  37507=>"111111111",
  37508=>"111111111",
  37509=>"001000000",
  37510=>"101001001",
  37511=>"000000000",
  37512=>"000000010",
  37513=>"111111111",
  37514=>"111111001",
  37515=>"111111111",
  37516=>"000100100",
  37517=>"000000000",
  37518=>"111100111",
  37519=>"111111101",
  37520=>"101000000",
  37521=>"111000011",
  37522=>"111111111",
  37523=>"111100110",
  37524=>"111111110",
  37525=>"110111110",
  37526=>"111101111",
  37527=>"111001000",
  37528=>"111100000",
  37529=>"111111111",
  37530=>"111010000",
  37531=>"100100110",
  37532=>"000110111",
  37533=>"000001001",
  37534=>"000000001",
  37535=>"100100100",
  37536=>"111010000",
  37537=>"100001111",
  37538=>"111110000",
  37539=>"001111111",
  37540=>"000100100",
  37541=>"011011100",
  37542=>"101001000",
  37543=>"111100000",
  37544=>"100111111",
  37545=>"000010000",
  37546=>"000000000",
  37547=>"111111111",
  37548=>"111111100",
  37549=>"111111111",
  37550=>"110100000",
  37551=>"100101111",
  37552=>"000000111",
  37553=>"111111011",
  37554=>"110111111",
  37555=>"000000000",
  37556=>"110001111",
  37557=>"000000000",
  37558=>"100110101",
  37559=>"000000100",
  37560=>"111100100",
  37561=>"000000000",
  37562=>"000000000",
  37563=>"101111111",
  37564=>"111000000",
  37565=>"000000011",
  37566=>"111111111",
  37567=>"000000001",
  37568=>"101100000",
  37569=>"111100100",
  37570=>"100000000",
  37571=>"011000111",
  37572=>"111111000",
  37573=>"000000000",
  37574=>"000001111",
  37575=>"111100111",
  37576=>"110000000",
  37577=>"111000000",
  37578=>"111001010",
  37579=>"111111100",
  37580=>"000101111",
  37581=>"000111000",
  37582=>"000001000",
  37583=>"000100100",
  37584=>"000000110",
  37585=>"110100110",
  37586=>"000000001",
  37587=>"100111111",
  37588=>"011001101",
  37589=>"011110110",
  37590=>"111101100",
  37591=>"111011111",
  37592=>"000000000",
  37593=>"111111110",
  37594=>"000000000",
  37595=>"111111101",
  37596=>"111100101",
  37597=>"101100110",
  37598=>"111111111",
  37599=>"000111111",
  37600=>"111111111",
  37601=>"111111111",
  37602=>"111001000",
  37603=>"000000000",
  37604=>"000000000",
  37605=>"111110110",
  37606=>"111111111",
  37607=>"111111111",
  37608=>"111111001",
  37609=>"111111100",
  37610=>"000000000",
  37611=>"001001101",
  37612=>"001000000",
  37613=>"011111100",
  37614=>"000000101",
  37615=>"000000000",
  37616=>"111111111",
  37617=>"000000000",
  37618=>"101000000",
  37619=>"000010111",
  37620=>"001001111",
  37621=>"001111110",
  37622=>"111010011",
  37623=>"111111111",
  37624=>"111110000",
  37625=>"000111111",
  37626=>"111111111",
  37627=>"110000010",
  37628=>"001001000",
  37629=>"111011001",
  37630=>"000000111",
  37631=>"100000100",
  37632=>"111110110",
  37633=>"111101111",
  37634=>"000000110",
  37635=>"000100000",
  37636=>"000000110",
  37637=>"001011111",
  37638=>"100000111",
  37639=>"111001001",
  37640=>"111000000",
  37641=>"111111101",
  37642=>"000111111",
  37643=>"111001000",
  37644=>"111111111",
  37645=>"001000100",
  37646=>"111101101",
  37647=>"001001100",
  37648=>"000000001",
  37649=>"000000000",
  37650=>"000000100",
  37651=>"011011000",
  37652=>"001111111",
  37653=>"111001000",
  37654=>"100001101",
  37655=>"000000001",
  37656=>"111011110",
  37657=>"111111111",
  37658=>"000000000",
  37659=>"110111100",
  37660=>"000000001",
  37661=>"111111111",
  37662=>"000111111",
  37663=>"111111111",
  37664=>"111110111",
  37665=>"101000001",
  37666=>"111011000",
  37667=>"000000100",
  37668=>"011111110",
  37669=>"100000000",
  37670=>"111001000",
  37671=>"101001000",
  37672=>"000110100",
  37673=>"100111000",
  37674=>"111111111",
  37675=>"010010111",
  37676=>"111110000",
  37677=>"110000110",
  37678=>"001000000",
  37679=>"100100001",
  37680=>"111000111",
  37681=>"111110110",
  37682=>"011110111",
  37683=>"100000011",
  37684=>"000000000",
  37685=>"111111111",
  37686=>"111111001",
  37687=>"000000000",
  37688=>"010110111",
  37689=>"000000101",
  37690=>"111101100",
  37691=>"111111101",
  37692=>"100000001",
  37693=>"001000000",
  37694=>"000000001",
  37695=>"001000000",
  37696=>"011011001",
  37697=>"101100101",
  37698=>"000000000",
  37699=>"000000000",
  37700=>"111111101",
  37701=>"111110000",
  37702=>"001001001",
  37703=>"000000000",
  37704=>"111110100",
  37705=>"000000110",
  37706=>"000000110",
  37707=>"111011011",
  37708=>"000110111",
  37709=>"111111001",
  37710=>"000100110",
  37711=>"010110000",
  37712=>"110111111",
  37713=>"010011001",
  37714=>"000111111",
  37715=>"000000000",
  37716=>"111100000",
  37717=>"111000000",
  37718=>"000000101",
  37719=>"100000000",
  37720=>"011111111",
  37721=>"000000000",
  37722=>"000000000",
  37723=>"000000000",
  37724=>"000000000",
  37725=>"000100100",
  37726=>"000011010",
  37727=>"111111111",
  37728=>"000000000",
  37729=>"000000001",
  37730=>"100011011",
  37731=>"111111111",
  37732=>"110110010",
  37733=>"000000000",
  37734=>"100100110",
  37735=>"111110000",
  37736=>"000100110",
  37737=>"101001001",
  37738=>"011111111",
  37739=>"111010000",
  37740=>"110010110",
  37741=>"000000000",
  37742=>"100100000",
  37743=>"100101001",
  37744=>"111111111",
  37745=>"000000000",
  37746=>"111111111",
  37747=>"010000000",
  37748=>"000010111",
  37749=>"110000000",
  37750=>"111111011",
  37751=>"000000111",
  37752=>"111001000",
  37753=>"011011000",
  37754=>"111000000",
  37755=>"101111111",
  37756=>"011001001",
  37757=>"111001001",
  37758=>"111011001",
  37759=>"000000000",
  37760=>"110111111",
  37761=>"001000000",
  37762=>"111111111",
  37763=>"000000000",
  37764=>"011110110",
  37765=>"111111000",
  37766=>"000010110",
  37767=>"101001111",
  37768=>"000000000",
  37769=>"110111111",
  37770=>"111111110",
  37771=>"000111111",
  37772=>"000000000",
  37773=>"000100110",
  37774=>"111110111",
  37775=>"111011101",
  37776=>"001000100",
  37777=>"000000111",
  37778=>"111100100",
  37779=>"111111111",
  37780=>"000000000",
  37781=>"000100000",
  37782=>"111011001",
  37783=>"011010010",
  37784=>"111111111",
  37785=>"001101000",
  37786=>"011000000",
  37787=>"100111111",
  37788=>"000000110",
  37789=>"000011011",
  37790=>"111111000",
  37791=>"011111111",
  37792=>"000111111",
  37793=>"011001001",
  37794=>"111011000",
  37795=>"111111111",
  37796=>"001000000",
  37797=>"000000000",
  37798=>"000000000",
  37799=>"001001101",
  37800=>"000000100",
  37801=>"100110111",
  37802=>"000010111",
  37803=>"111111111",
  37804=>"000111111",
  37805=>"111111111",
  37806=>"100100100",
  37807=>"100100001",
  37808=>"101111100",
  37809=>"000000110",
  37810=>"111111111",
  37811=>"111110110",
  37812=>"001000101",
  37813=>"000000110",
  37814=>"111000000",
  37815=>"000001000",
  37816=>"000000011",
  37817=>"001111111",
  37818=>"000000000",
  37819=>"100110000",
  37820=>"000000111",
  37821=>"111011001",
  37822=>"111000011",
  37823=>"100101101",
  37824=>"111111111",
  37825=>"111111111",
  37826=>"000000000",
  37827=>"111111000",
  37828=>"111011111",
  37829=>"110110100",
  37830=>"111111100",
  37831=>"111110000",
  37832=>"000011111",
  37833=>"000000000",
  37834=>"111101100",
  37835=>"000000111",
  37836=>"011101111",
  37837=>"111111111",
  37838=>"101100101",
  37839=>"001000000",
  37840=>"111111111",
  37841=>"001110000",
  37842=>"001001111",
  37843=>"000000000",
  37844=>"011111111",
  37845=>"111111111",
  37846=>"111001000",
  37847=>"000000000",
  37848=>"000000000",
  37849=>"000000010",
  37850=>"111111011",
  37851=>"011011111",
  37852=>"000110100",
  37853=>"100100111",
  37854=>"100000000",
  37855=>"100100111",
  37856=>"111000000",
  37857=>"111111000",
  37858=>"111111111",
  37859=>"001001011",
  37860=>"000000111",
  37861=>"111001000",
  37862=>"001001111",
  37863=>"011111111",
  37864=>"111001000",
  37865=>"111111111",
  37866=>"011111111",
  37867=>"100000000",
  37868=>"101101111",
  37869=>"100101111",
  37870=>"000000010",
  37871=>"011000000",
  37872=>"100100000",
  37873=>"000000000",
  37874=>"011011011",
  37875=>"000001111",
  37876=>"000011111",
  37877=>"000000110",
  37878=>"111100100",
  37879=>"111100100",
  37880=>"111111110",
  37881=>"001000001",
  37882=>"111111000",
  37883=>"111000000",
  37884=>"111111111",
  37885=>"111000110",
  37886=>"111111111",
  37887=>"000000100",
  37888=>"000000000",
  37889=>"111111001",
  37890=>"100110010",
  37891=>"111101101",
  37892=>"100000000",
  37893=>"000000000",
  37894=>"000011000",
  37895=>"000000000",
  37896=>"101111111",
  37897=>"000111111",
  37898=>"111111111",
  37899=>"000000000",
  37900=>"000100100",
  37901=>"000001101",
  37902=>"000000000",
  37903=>"000011011",
  37904=>"100111111",
  37905=>"000111000",
  37906=>"000000011",
  37907=>"010010010",
  37908=>"111111000",
  37909=>"010110111",
  37910=>"000110010",
  37911=>"111111111",
  37912=>"111111001",
  37913=>"010010000",
  37914=>"111100000",
  37915=>"010000000",
  37916=>"111101000",
  37917=>"000100000",
  37918=>"111011011",
  37919=>"110100100",
  37920=>"100110000",
  37921=>"011011111",
  37922=>"111111110",
  37923=>"111100100",
  37924=>"001011011",
  37925=>"010010000",
  37926=>"000111000",
  37927=>"000000000",
  37928=>"111111101",
  37929=>"000000000",
  37930=>"111111011",
  37931=>"110000000",
  37932=>"111111111",
  37933=>"001101101",
  37934=>"111111111",
  37935=>"001001001",
  37936=>"111101101",
  37937=>"000000001",
  37938=>"011111110",
  37939=>"000000000",
  37940=>"111111111",
  37941=>"000100110",
  37942=>"000000000",
  37943=>"000000000",
  37944=>"110111100",
  37945=>"000000110",
  37946=>"011000001",
  37947=>"000000110",
  37948=>"001000000",
  37949=>"000000011",
  37950=>"110111111",
  37951=>"101000001",
  37952=>"110110110",
  37953=>"001001111",
  37954=>"111111111",
  37955=>"000100000",
  37956=>"011011000",
  37957=>"110010011",
  37958=>"000000000",
  37959=>"111111111",
  37960=>"011000110",
  37961=>"001000101",
  37962=>"000000000",
  37963=>"011011011",
  37964=>"000001111",
  37965=>"111111010",
  37966=>"011111001",
  37967=>"110111111",
  37968=>"000000011",
  37969=>"111111110",
  37970=>"000000010",
  37971=>"110111011",
  37972=>"000000010",
  37973=>"111111111",
  37974=>"000000100",
  37975=>"100011001",
  37976=>"111111111",
  37977=>"100000000",
  37978=>"111110110",
  37979=>"101111001",
  37980=>"111111010",
  37981=>"111111111",
  37982=>"001000001",
  37983=>"111110110",
  37984=>"000000000",
  37985=>"000001111",
  37986=>"111100100",
  37987=>"000000010",
  37988=>"000000000",
  37989=>"110110010",
  37990=>"111011111",
  37991=>"111000000",
  37992=>"000111111",
  37993=>"110111111",
  37994=>"001001000",
  37995=>"000100101",
  37996=>"111111111",
  37997=>"000000000",
  37998=>"111111000",
  37999=>"100000000",
  38000=>"101111111",
  38001=>"111111111",
  38002=>"010111001",
  38003=>"001000100",
  38004=>"010000000",
  38005=>"000000001",
  38006=>"111111111",
  38007=>"000000011",
  38008=>"111111111",
  38009=>"111111110",
  38010=>"000000000",
  38011=>"111011010",
  38012=>"111111111",
  38013=>"110000001",
  38014=>"011000000",
  38015=>"010000010",
  38016=>"000000111",
  38017=>"111111111",
  38018=>"110000111",
  38019=>"000001001",
  38020=>"101000000",
  38021=>"000101111",
  38022=>"000000000",
  38023=>"000000000",
  38024=>"000000000",
  38025=>"001000000",
  38026=>"000000000",
  38027=>"111111111",
  38028=>"111111110",
  38029=>"111111111",
  38030=>"010000111",
  38031=>"010111011",
  38032=>"000000010",
  38033=>"100000000",
  38034=>"010110010",
  38035=>"011001000",
  38036=>"111111111",
  38037=>"100111011",
  38038=>"000000000",
  38039=>"000000100",
  38040=>"000001101",
  38041=>"000000000",
  38042=>"001001000",
  38043=>"001001000",
  38044=>"111001100",
  38045=>"110000000",
  38046=>"111001000",
  38047=>"111000000",
  38048=>"000000000",
  38049=>"000000000",
  38050=>"000000111",
  38051=>"000001000",
  38052=>"000000000",
  38053=>"111111111",
  38054=>"111111111",
  38055=>"111111111",
  38056=>"000000000",
  38057=>"000000000",
  38058=>"000001001",
  38059=>"000000100",
  38060=>"100000110",
  38061=>"100001001",
  38062=>"111111111",
  38063=>"000001111",
  38064=>"111110111",
  38065=>"000000110",
  38066=>"101101111",
  38067=>"000000000",
  38068=>"110000101",
  38069=>"000000000",
  38070=>"000000000",
  38071=>"010111111",
  38072=>"011011001",
  38073=>"011111111",
  38074=>"000010000",
  38075=>"000000000",
  38076=>"111111111",
  38077=>"010000000",
  38078=>"000000000",
  38079=>"000011111",
  38080=>"000001000",
  38081=>"000000010",
  38082=>"111111111",
  38083=>"111111111",
  38084=>"001001111",
  38085=>"111111111",
  38086=>"001001001",
  38087=>"000000000",
  38088=>"110100000",
  38089=>"110000111",
  38090=>"001000000",
  38091=>"000100100",
  38092=>"000000100",
  38093=>"001111111",
  38094=>"000010111",
  38095=>"000000000",
  38096=>"101001001",
  38097=>"001000000",
  38098=>"000000000",
  38099=>"101000101",
  38100=>"111111111",
  38101=>"000000101",
  38102=>"111101100",
  38103=>"001001101",
  38104=>"000000000",
  38105=>"100110111",
  38106=>"000000000",
  38107=>"000011111",
  38108=>"101101111",
  38109=>"111111110",
  38110=>"000101111",
  38111=>"111111111",
  38112=>"111111001",
  38113=>"000000000",
  38114=>"111100000",
  38115=>"111000000",
  38116=>"000001001",
  38117=>"001000000",
  38118=>"000000000",
  38119=>"100110100",
  38120=>"001111000",
  38121=>"000000000",
  38122=>"101111111",
  38123=>"111111011",
  38124=>"111111011",
  38125=>"010110000",
  38126=>"000000000",
  38127=>"111111111",
  38128=>"110110100",
  38129=>"010000111",
  38130=>"000111111",
  38131=>"110110000",
  38132=>"110110110",
  38133=>"011111011",
  38134=>"111111110",
  38135=>"101100100",
  38136=>"101001001",
  38137=>"100100111",
  38138=>"000010111",
  38139=>"000000001",
  38140=>"100000000",
  38141=>"100000110",
  38142=>"001000111",
  38143=>"000111111",
  38144=>"000001111",
  38145=>"000100111",
  38146=>"000001000",
  38147=>"000001111",
  38148=>"111001111",
  38149=>"001000000",
  38150=>"000100111",
  38151=>"000010000",
  38152=>"000001000",
  38153=>"000010110",
  38154=>"100001001",
  38155=>"000000000",
  38156=>"000000001",
  38157=>"000111110",
  38158=>"000001111",
  38159=>"000001000",
  38160=>"111000000",
  38161=>"000000111",
  38162=>"111000001",
  38163=>"001001000",
  38164=>"110110100",
  38165=>"101101101",
  38166=>"011011111",
  38167=>"000000001",
  38168=>"111111111",
  38169=>"111110110",
  38170=>"111110010",
  38171=>"101001011",
  38172=>"000011111",
  38173=>"111110111",
  38174=>"000000000",
  38175=>"111111110",
  38176=>"000000010",
  38177=>"000000001",
  38178=>"101101101",
  38179=>"111111001",
  38180=>"110010010",
  38181=>"111001001",
  38182=>"000000000",
  38183=>"010000000",
  38184=>"110000000",
  38185=>"111111111",
  38186=>"110000000",
  38187=>"111111111",
  38188=>"111111010",
  38189=>"110110110",
  38190=>"000000000",
  38191=>"001010110",
  38192=>"111111111",
  38193=>"010010010",
  38194=>"111111000",
  38195=>"111001000",
  38196=>"001000001",
  38197=>"001001000",
  38198=>"010001111",
  38199=>"111111100",
  38200=>"101101101",
  38201=>"111100000",
  38202=>"000001001",
  38203=>"101111000",
  38204=>"000000100",
  38205=>"001101111",
  38206=>"010011011",
  38207=>"000000000",
  38208=>"011111111",
  38209=>"101111100",
  38210=>"000000000",
  38211=>"111111000",
  38212=>"000000010",
  38213=>"001001101",
  38214=>"000000000",
  38215=>"001111111",
  38216=>"000000000",
  38217=>"111001000",
  38218=>"110010000",
  38219=>"110110110",
  38220=>"000000000",
  38221=>"000100111",
  38222=>"001001000",
  38223=>"001001001",
  38224=>"100100110",
  38225=>"000010011",
  38226=>"010001000",
  38227=>"101001000",
  38228=>"100111110",
  38229=>"111110111",
  38230=>"010010111",
  38231=>"000000000",
  38232=>"100000111",
  38233=>"111111111",
  38234=>"000000000",
  38235=>"010111111",
  38236=>"000111111",
  38237=>"000000011",
  38238=>"111111111",
  38239=>"111001001",
  38240=>"000000000",
  38241=>"000000010",
  38242=>"000110110",
  38243=>"000000000",
  38244=>"110111111",
  38245=>"101111111",
  38246=>"000000111",
  38247=>"111111101",
  38248=>"111111111",
  38249=>"010000000",
  38250=>"000111111",
  38251=>"111000110",
  38252=>"011000000",
  38253=>"111111111",
  38254=>"111111111",
  38255=>"000000000",
  38256=>"110111110",
  38257=>"001101111",
  38258=>"101111011",
  38259=>"000000000",
  38260=>"111011011",
  38261=>"111100101",
  38262=>"010011011",
  38263=>"000000000",
  38264=>"000000000",
  38265=>"111111000",
  38266=>"011000000",
  38267=>"100000000",
  38268=>"010000000",
  38269=>"000000000",
  38270=>"111111111",
  38271=>"000010000",
  38272=>"011001011",
  38273=>"000010000",
  38274=>"111110110",
  38275=>"011011011",
  38276=>"001000000",
  38277=>"111111111",
  38278=>"000100111",
  38279=>"111100000",
  38280=>"000001111",
  38281=>"000000100",
  38282=>"111111101",
  38283=>"110100100",
  38284=>"101111111",
  38285=>"000000001",
  38286=>"111111111",
  38287=>"000010111",
  38288=>"001000000",
  38289=>"111111110",
  38290=>"111101111",
  38291=>"001001001",
  38292=>"000000000",
  38293=>"000001001",
  38294=>"001001000",
  38295=>"111111111",
  38296=>"110111111",
  38297=>"000000000",
  38298=>"000110000",
  38299=>"011011111",
  38300=>"011111100",
  38301=>"001101111",
  38302=>"100100100",
  38303=>"011111011",
  38304=>"011111111",
  38305=>"000000100",
  38306=>"000001101",
  38307=>"000100110",
  38308=>"001111101",
  38309=>"001000101",
  38310=>"010001000",
  38311=>"001000000",
  38312=>"001000000",
  38313=>"000000000",
  38314=>"000000110",
  38315=>"000100000",
  38316=>"111111111",
  38317=>"000001111",
  38318=>"111111111",
  38319=>"011011000",
  38320=>"011011111",
  38321=>"000000000",
  38322=>"000000000",
  38323=>"011011101",
  38324=>"011000000",
  38325=>"110111100",
  38326=>"111111001",
  38327=>"110111111",
  38328=>"000101111",
  38329=>"100111111",
  38330=>"000000000",
  38331=>"100100000",
  38332=>"111001000",
  38333=>"000101000",
  38334=>"000000000",
  38335=>"111111111",
  38336=>"101000000",
  38337=>"111111101",
  38338=>"000000000",
  38339=>"001000001",
  38340=>"110100000",
  38341=>"001000111",
  38342=>"011111101",
  38343=>"111111111",
  38344=>"000000000",
  38345=>"000011111",
  38346=>"000000100",
  38347=>"101101001",
  38348=>"111111011",
  38349=>"000000100",
  38350=>"001000000",
  38351=>"011111111",
  38352=>"000000000",
  38353=>"010111000",
  38354=>"000000000",
  38355=>"111100000",
  38356=>"111011111",
  38357=>"111011001",
  38358=>"111111111",
  38359=>"011011011",
  38360=>"111001000",
  38361=>"111111111",
  38362=>"110011000",
  38363=>"111111101",
  38364=>"000000001",
  38365=>"000011000",
  38366=>"000000000",
  38367=>"001011111",
  38368=>"000000000",
  38369=>"111111000",
  38370=>"111111110",
  38371=>"010010000",
  38372=>"100100111",
  38373=>"110110000",
  38374=>"000000000",
  38375=>"000000010",
  38376=>"000000010",
  38377=>"000111111",
  38378=>"000111111",
  38379=>"000000000",
  38380=>"110110000",
  38381=>"110110110",
  38382=>"100110000",
  38383=>"000001000",
  38384=>"000000000",
  38385=>"000000000",
  38386=>"100001101",
  38387=>"111000000",
  38388=>"111111100",
  38389=>"011111111",
  38390=>"000000110",
  38391=>"000000000",
  38392=>"011111011",
  38393=>"100111110",
  38394=>"111111111",
  38395=>"110110000",
  38396=>"101111111",
  38397=>"111001001",
  38398=>"000000000",
  38399=>"000000111",
  38400=>"011011101",
  38401=>"000000111",
  38402=>"000000000",
  38403=>"000111111",
  38404=>"000000000",
  38405=>"111101001",
  38406=>"100000000",
  38407=>"000000111",
  38408=>"000010000",
  38409=>"101111111",
  38410=>"011000001",
  38411=>"111111111",
  38412=>"000000000",
  38413=>"100101111",
  38414=>"000001111",
  38415=>"001001001",
  38416=>"001011111",
  38417=>"000100000",
  38418=>"001001011",
  38419=>"000000000",
  38420=>"000000000",
  38421=>"111111001",
  38422=>"011011011",
  38423=>"100000001",
  38424=>"111111111",
  38425=>"000001001",
  38426=>"100001000",
  38427=>"000000000",
  38428=>"110110100",
  38429=>"001011011",
  38430=>"001001000",
  38431=>"111110010",
  38432=>"000000000",
  38433=>"111111111",
  38434=>"011001011",
  38435=>"111011001",
  38436=>"000000001",
  38437=>"000000100",
  38438=>"111111111",
  38439=>"000000110",
  38440=>"011001111",
  38441=>"000000000",
  38442=>"000000000",
  38443=>"111111101",
  38444=>"111111000",
  38445=>"001001111",
  38446=>"010110111",
  38447=>"100110110",
  38448=>"011111100",
  38449=>"000000000",
  38450=>"110110100",
  38451=>"111111111",
  38452=>"011011011",
  38453=>"010011000",
  38454=>"000000000",
  38455=>"100000001",
  38456=>"111111100",
  38457=>"111111111",
  38458=>"001001111",
  38459=>"010000000",
  38460=>"111111111",
  38461=>"000000000",
  38462=>"000000011",
  38463=>"001000111",
  38464=>"011000000",
  38465=>"000000000",
  38466=>"110110111",
  38467=>"111001111",
  38468=>"111001001",
  38469=>"011010000",
  38470=>"100100011",
  38471=>"000000000",
  38472=>"011111000",
  38473=>"001001011",
  38474=>"000100100",
  38475=>"111010010",
  38476=>"111111111",
  38477=>"000111000",
  38478=>"111100101",
  38479=>"001001111",
  38480=>"001000000",
  38481=>"011011000",
  38482=>"000000000",
  38483=>"001000101",
  38484=>"110111111",
  38485=>"100100111",
  38486=>"111100000",
  38487=>"111111001",
  38488=>"111111111",
  38489=>"001000000",
  38490=>"011111110",
  38491=>"100111010",
  38492=>"000000000",
  38493=>"111111111",
  38494=>"111111111",
  38495=>"011111111",
  38496=>"000001011",
  38497=>"101001001",
  38498=>"011010001",
  38499=>"100100100",
  38500=>"111111111",
  38501=>"100100100",
  38502=>"100000000",
  38503=>"100100000",
  38504=>"111110110",
  38505=>"111101001",
  38506=>"000000000",
  38507=>"111111111",
  38508=>"000000000",
  38509=>"000000000",
  38510=>"111111011",
  38511=>"001001001",
  38512=>"001000111",
  38513=>"111110000",
  38514=>"001000000",
  38515=>"111011111",
  38516=>"110110110",
  38517=>"000000000",
  38518=>"000000000",
  38519=>"111111111",
  38520=>"001000111",
  38521=>"111101101",
  38522=>"110110110",
  38523=>"000000000",
  38524=>"000000000",
  38525=>"111111111",
  38526=>"111111000",
  38527=>"110110000",
  38528=>"000011111",
  38529=>"000000011",
  38530=>"011111010",
  38531=>"111011000",
  38532=>"001000000",
  38533=>"000000010",
  38534=>"000000000",
  38535=>"011000011",
  38536=>"111101111",
  38537=>"111101111",
  38538=>"000000000",
  38539=>"000100111",
  38540=>"001000100",
  38541=>"111111001",
  38542=>"011011011",
  38543=>"000011010",
  38544=>"111111111",
  38545=>"111111100",
  38546=>"001000000",
  38547=>"110000100",
  38548=>"111111000",
  38549=>"100101110",
  38550=>"001001001",
  38551=>"001001111",
  38552=>"000000001",
  38553=>"000000000",
  38554=>"100110111",
  38555=>"000000000",
  38556=>"111111111",
  38557=>"100100111",
  38558=>"001110110",
  38559=>"111111111",
  38560=>"111100000",
  38561=>"100001001",
  38562=>"100100001",
  38563=>"111111111",
  38564=>"111111110",
  38565=>"000000000",
  38566=>"101100111",
  38567=>"101101101",
  38568=>"111111000",
  38569=>"111111111",
  38570=>"111111111",
  38571=>"111111111",
  38572=>"111111111",
  38573=>"000000000",
  38574=>"000000101",
  38575=>"001001011",
  38576=>"111111111",
  38577=>"000000000",
  38578=>"111111111",
  38579=>"000000000",
  38580=>"110110111",
  38581=>"111111110",
  38582=>"000001000",
  38583=>"100100111",
  38584=>"000000100",
  38585=>"000000000",
  38586=>"010110000",
  38587=>"001011111",
  38588=>"111111111",
  38589=>"001000000",
  38590=>"111110111",
  38591=>"000000011",
  38592=>"111100100",
  38593=>"111111111",
  38594=>"011111111",
  38595=>"000000000",
  38596=>"111111011",
  38597=>"001001011",
  38598=>"011100110",
  38599=>"001001000",
  38600=>"000000011",
  38601=>"111101000",
  38602=>"110111011",
  38603=>"000000000",
  38604=>"111001111",
  38605=>"110111111",
  38606=>"111111111",
  38607=>"000000000",
  38608=>"000000100",
  38609=>"100000001",
  38610=>"110110111",
  38611=>"010110110",
  38612=>"101111111",
  38613=>"001011111",
  38614=>"000000000",
  38615=>"100000110",
  38616=>"001000000",
  38617=>"110101111",
  38618=>"111011111",
  38619=>"111111111",
  38620=>"111111111",
  38621=>"100000011",
  38622=>"000000000",
  38623=>"001001000",
  38624=>"000000000",
  38625=>"000000010",
  38626=>"001001111",
  38627=>"001011111",
  38628=>"110110111",
  38629=>"011011011",
  38630=>"011001001",
  38631=>"000000000",
  38632=>"000000000",
  38633=>"000000000",
  38634=>"000000000",
  38635=>"001000000",
  38636=>"111101001",
  38637=>"000111010",
  38638=>"100110111",
  38639=>"110000000",
  38640=>"111111111",
  38641=>"111001001",
  38642=>"000000000",
  38643=>"011111111",
  38644=>"011111111",
  38645=>"111111111",
  38646=>"111011011",
  38647=>"111001000",
  38648=>"111011001",
  38649=>"000000000",
  38650=>"101101111",
  38651=>"000000000",
  38652=>"110111001",
  38653=>"000000110",
  38654=>"111101011",
  38655=>"110000000",
  38656=>"010000000",
  38657=>"000001000",
  38658=>"000000000",
  38659=>"011011111",
  38660=>"001001001",
  38661=>"000000000",
  38662=>"111111111",
  38663=>"111010010",
  38664=>"111101101",
  38665=>"000000000",
  38666=>"101000111",
  38667=>"000000110",
  38668=>"111101111",
  38669=>"001100100",
  38670=>"111111111",
  38671=>"000000000",
  38672=>"100111000",
  38673=>"110000000",
  38674=>"100100100",
  38675=>"001000000",
  38676=>"000000100",
  38677=>"000000000",
  38678=>"100111111",
  38679=>"100100100",
  38680=>"100100111",
  38681=>"100100000",
  38682=>"000000000",
  38683=>"001001001",
  38684=>"111111111",
  38685=>"111000000",
  38686=>"000000011",
  38687=>"000000011",
  38688=>"111111111",
  38689=>"000000000",
  38690=>"100000000",
  38691=>"111000100",
  38692=>"000000010",
  38693=>"001111111",
  38694=>"000100111",
  38695=>"100110110",
  38696=>"100000000",
  38697=>"111001001",
  38698=>"101101100",
  38699=>"000000000",
  38700=>"111111111",
  38701=>"001111111",
  38702=>"000000111",
  38703=>"000000000",
  38704=>"111111111",
  38705=>"011011101",
  38706=>"001000000",
  38707=>"000000111",
  38708=>"000000000",
  38709=>"101000101",
  38710=>"000000000",
  38711=>"100100110",
  38712=>"000000000",
  38713=>"111111111",
  38714=>"111111111",
  38715=>"111111111",
  38716=>"110100110",
  38717=>"001101111",
  38718=>"110111111",
  38719=>"111111111",
  38720=>"000000000",
  38721=>"001000000",
  38722=>"000000111",
  38723=>"100100001",
  38724=>"001000000",
  38725=>"000001111",
  38726=>"000000100",
  38727=>"000000001",
  38728=>"000000000",
  38729=>"010000111",
  38730=>"110110110",
  38731=>"011001011",
  38732=>"000001111",
  38733=>"100111111",
  38734=>"010000110",
  38735=>"000000111",
  38736=>"011001000",
  38737=>"110110100",
  38738=>"000000000",
  38739=>"100110111",
  38740=>"001000001",
  38741=>"011011011",
  38742=>"000001101",
  38743=>"101000000",
  38744=>"000000000",
  38745=>"000000000",
  38746=>"000000100",
  38747=>"111111111",
  38748=>"000000000",
  38749=>"111111111",
  38750=>"111110111",
  38751=>"000000000",
  38752=>"111111100",
  38753=>"111111111",
  38754=>"111011001",
  38755=>"011000000",
  38756=>"110111111",
  38757=>"000000001",
  38758=>"111001000",
  38759=>"000000000",
  38760=>"000000000",
  38761=>"000000000",
  38762=>"100100000",
  38763=>"000000000",
  38764=>"000000000",
  38765=>"001101000",
  38766=>"111111111",
  38767=>"000010000",
  38768=>"000000000",
  38769=>"000101111",
  38770=>"011011111",
  38771=>"101000001",
  38772=>"000000000",
  38773=>"111000100",
  38774=>"110110000",
  38775=>"000000000",
  38776=>"000000000",
  38777=>"000000000",
  38778=>"111011011",
  38779=>"111111111",
  38780=>"100110110",
  38781=>"111001000",
  38782=>"110000000",
  38783=>"111111001",
  38784=>"000000000",
  38785=>"001001000",
  38786=>"111111101",
  38787=>"000000000",
  38788=>"101111111",
  38789=>"000000000",
  38790=>"111111110",
  38791=>"000000111",
  38792=>"111011011",
  38793=>"000011011",
  38794=>"111111111",
  38795=>"000000111",
  38796=>"111111011",
  38797=>"000001101",
  38798=>"011011000",
  38799=>"000000000",
  38800=>"000000000",
  38801=>"000000000",
  38802=>"111000000",
  38803=>"111111111",
  38804=>"001001001",
  38805=>"000010000",
  38806=>"000000000",
  38807=>"000011000",
  38808=>"110000001",
  38809=>"100000000",
  38810=>"111111111",
  38811=>"100000000",
  38812=>"111011011",
  38813=>"100000000",
  38814=>"010011001",
  38815=>"000000000",
  38816=>"111100110",
  38817=>"001000111",
  38818=>"111111110",
  38819=>"010110010",
  38820=>"011111111",
  38821=>"111111111",
  38822=>"000000101",
  38823=>"000000111",
  38824=>"000000000",
  38825=>"000000001",
  38826=>"110111111",
  38827=>"000000000",
  38828=>"100100101",
  38829=>"000000101",
  38830=>"101001111",
  38831=>"110110110",
  38832=>"111111001",
  38833=>"111111110",
  38834=>"000001111",
  38835=>"000000000",
  38836=>"000000111",
  38837=>"011011111",
  38838=>"111111111",
  38839=>"110011011",
  38840=>"111011000",
  38841=>"001100100",
  38842=>"000000010",
  38843=>"111000000",
  38844=>"111111111",
  38845=>"000000000",
  38846=>"000000000",
  38847=>"000000000",
  38848=>"000000101",
  38849=>"100000101",
  38850=>"100100111",
  38851=>"000100100",
  38852=>"101111111",
  38853=>"111011001",
  38854=>"111100100",
  38855=>"000100100",
  38856=>"011011000",
  38857=>"010000000",
  38858=>"111000101",
  38859=>"111111111",
  38860=>"111111001",
  38861=>"000000001",
  38862=>"111111111",
  38863=>"110110100",
  38864=>"100100110",
  38865=>"111111111",
  38866=>"111111111",
  38867=>"000110111",
  38868=>"001000000",
  38869=>"000000000",
  38870=>"000011111",
  38871=>"000000000",
  38872=>"111111111",
  38873=>"011111111",
  38874=>"111010110",
  38875=>"111100111",
  38876=>"110100001",
  38877=>"000000110",
  38878=>"111111111",
  38879=>"100100100",
  38880=>"001001101",
  38881=>"110111111",
  38882=>"111111000",
  38883=>"000000000",
  38884=>"100100110",
  38885=>"111111110",
  38886=>"000000111",
  38887=>"111000000",
  38888=>"101100100",
  38889=>"111111111",
  38890=>"000000000",
  38891=>"111111111",
  38892=>"110000100",
  38893=>"011000001",
  38894=>"000000000",
  38895=>"000000000",
  38896=>"111000100",
  38897=>"000111111",
  38898=>"111110111",
  38899=>"000000000",
  38900=>"111111111",
  38901=>"110000100",
  38902=>"000000000",
  38903=>"100000100",
  38904=>"000000000",
  38905=>"001000001",
  38906=>"000100000",
  38907=>"001001011",
  38908=>"011011000",
  38909=>"000000000",
  38910=>"100100000",
  38911=>"000000011",
  38912=>"111111111",
  38913=>"111111100",
  38914=>"111111111",
  38915=>"000000000",
  38916=>"111111111",
  38917=>"011000110",
  38918=>"000000000",
  38919=>"111111111",
  38920=>"000011011",
  38921=>"000000000",
  38922=>"111111111",
  38923=>"111111111",
  38924=>"111101000",
  38925=>"000000000",
  38926=>"000100000",
  38927=>"111111111",
  38928=>"111111011",
  38929=>"011011111",
  38930=>"111111000",
  38931=>"001001000",
  38932=>"111101001",
  38933=>"001001111",
  38934=>"000000000",
  38935=>"110110110",
  38936=>"000001001",
  38937=>"011011011",
  38938=>"111111111",
  38939=>"110110111",
  38940=>"111111111",
  38941=>"111111111",
  38942=>"011000000",
  38943=>"010111000",
  38944=>"101100111",
  38945=>"111111111",
  38946=>"111001111",
  38947=>"000000111",
  38948=>"111110000",
  38949=>"000000000",
  38950=>"011101000",
  38951=>"111111001",
  38952=>"111111111",
  38953=>"101000000",
  38954=>"111111111",
  38955=>"100100100",
  38956=>"100110111",
  38957=>"000000000",
  38958=>"000000000",
  38959=>"101111001",
  38960=>"000000000",
  38961=>"111111000",
  38962=>"011011001",
  38963=>"001111101",
  38964=>"111111111",
  38965=>"110110110",
  38966=>"111100100",
  38967=>"000100100",
  38968=>"111111001",
  38969=>"001000001",
  38970=>"000000000",
  38971=>"000000101",
  38972=>"001111111",
  38973=>"011111111",
  38974=>"011011011",
  38975=>"000000000",
  38976=>"111010000",
  38977=>"000000000",
  38978=>"000110111",
  38979=>"001001011",
  38980=>"011001001",
  38981=>"001001011",
  38982=>"000000000",
  38983=>"111111111",
  38984=>"011011011",
  38985=>"000000111",
  38986=>"000000100",
  38987=>"111000111",
  38988=>"111111111",
  38989=>"110000000",
  38990=>"000000100",
  38991=>"111111111",
  38992=>"111111111",
  38993=>"000000000",
  38994=>"100000000",
  38995=>"110110011",
  38996=>"000000111",
  38997=>"000000000",
  38998=>"000000111",
  38999=>"001000001",
  39000=>"000000000",
  39001=>"111111111",
  39002=>"001111111",
  39003=>"000011111",
  39004=>"000000000",
  39005=>"001001010",
  39006=>"001000111",
  39007=>"000010000",
  39008=>"001000111",
  39009=>"001001000",
  39010=>"111101101",
  39011=>"111111011",
  39012=>"111111001",
  39013=>"000000000",
  39014=>"000000000",
  39015=>"011111111",
  39016=>"000000000",
  39017=>"111011000",
  39018=>"000000000",
  39019=>"111111011",
  39020=>"110110111",
  39021=>"011000000",
  39022=>"000001011",
  39023=>"000000000",
  39024=>"000000100",
  39025=>"001000000",
  39026=>"111111111",
  39027=>"000000000",
  39028=>"000000000",
  39029=>"010000000",
  39030=>"100000101",
  39031=>"111111100",
  39032=>"000100000",
  39033=>"000000100",
  39034=>"010000011",
  39035=>"000000000",
  39036=>"000000000",
  39037=>"010000000",
  39038=>"000000010",
  39039=>"111111101",
  39040=>"000011011",
  39041=>"111111000",
  39042=>"000110111",
  39043=>"000000000",
  39044=>"111111110",
  39045=>"000000011",
  39046=>"000000000",
  39047=>"000000001",
  39048=>"111000000",
  39049=>"101000100",
  39050=>"000000000",
  39051=>"011000000",
  39052=>"111111111",
  39053=>"111000000",
  39054=>"000000000",
  39055=>"011011001",
  39056=>"000000000",
  39057=>"000000000",
  39058=>"000000000",
  39059=>"100000111",
  39060=>"000000000",
  39061=>"111011111",
  39062=>"110100111",
  39063=>"000000000",
  39064=>"000000000",
  39065=>"011000001",
  39066=>"000000000",
  39067=>"000000000",
  39068=>"111110111",
  39069=>"110100000",
  39070=>"011111111",
  39071=>"000000010",
  39072=>"000000100",
  39073=>"011000000",
  39074=>"000000000",
  39075=>"100100000",
  39076=>"110110100",
  39077=>"010011111",
  39078=>"111111111",
  39079=>"000000000",
  39080=>"011111111",
  39081=>"111111111",
  39082=>"111111011",
  39083=>"011011010",
  39084=>"111101111",
  39085=>"100110100",
  39086=>"111110000",
  39087=>"100000001",
  39088=>"111000000",
  39089=>"111111111",
  39090=>"111111111",
  39091=>"111010111",
  39092=>"110000000",
  39093=>"111111111",
  39094=>"000000000",
  39095=>"000000000",
  39096=>"111111111",
  39097=>"111110110",
  39098=>"000000000",
  39099=>"110110100",
  39100=>"011000000",
  39101=>"110111111",
  39102=>"001100000",
  39103=>"111111111",
  39104=>"111111111",
  39105=>"111111111",
  39106=>"011000000",
  39107=>"111100000",
  39108=>"001011111",
  39109=>"000000000",
  39110=>"000000001",
  39111=>"000000000",
  39112=>"111111011",
  39113=>"001101001",
  39114=>"111111001",
  39115=>"111111011",
  39116=>"111111111",
  39117=>"000000111",
  39118=>"111111111",
  39119=>"111111111",
  39120=>"110111111",
  39121=>"000000000",
  39122=>"000001000",
  39123=>"000000010",
  39124=>"000000000",
  39125=>"111111111",
  39126=>"000000000",
  39127=>"110110100",
  39128=>"111110000",
  39129=>"111110111",
  39130=>"111000000",
  39131=>"111111111",
  39132=>"000011111",
  39133=>"000011011",
  39134=>"011111111",
  39135=>"111110000",
  39136=>"000000000",
  39137=>"101001000",
  39138=>"100100110",
  39139=>"111111111",
  39140=>"111011000",
  39141=>"111111111",
  39142=>"110110000",
  39143=>"111011111",
  39144=>"000000111",
  39145=>"111111111",
  39146=>"111101101",
  39147=>"111100100",
  39148=>"011011000",
  39149=>"000000000",
  39150=>"111111111",
  39151=>"111111111",
  39152=>"000000000",
  39153=>"000110000",
  39154=>"000000000",
  39155=>"000110000",
  39156=>"110100000",
  39157=>"100110111",
  39158=>"000000100",
  39159=>"001000000",
  39160=>"110110010",
  39161=>"001000000",
  39162=>"001011001",
  39163=>"111011111",
  39164=>"111101000",
  39165=>"001100000",
  39166=>"000000000",
  39167=>"011111111",
  39168=>"000000000",
  39169=>"001011001",
  39170=>"000000000",
  39171=>"000000000",
  39172=>"000000111",
  39173=>"000000101",
  39174=>"111111111",
  39175=>"111111011",
  39176=>"010000000",
  39177=>"000001001",
  39178=>"001100000",
  39179=>"000000111",
  39180=>"001000000",
  39181=>"111110111",
  39182=>"111111000",
  39183=>"111111111",
  39184=>"011000100",
  39185=>"111111111",
  39186=>"000000000",
  39187=>"000000000",
  39188=>"110001000",
  39189=>"011010000",
  39190=>"111111111",
  39191=>"111111000",
  39192=>"000000011",
  39193=>"110110000",
  39194=>"000000001",
  39195=>"011101111",
  39196=>"111111111",
  39197=>"000000000",
  39198=>"011000000",
  39199=>"010011001",
  39200=>"110110100",
  39201=>"110001011",
  39202=>"110111110",
  39203=>"111100111",
  39204=>"111111111",
  39205=>"000100111",
  39206=>"111111111",
  39207=>"110111101",
  39208=>"111111100",
  39209=>"111111111",
  39210=>"111011110",
  39211=>"000000000",
  39212=>"011111111",
  39213=>"000001001",
  39214=>"000000000",
  39215=>"111001001",
  39216=>"011000001",
  39217=>"111111101",
  39218=>"100111000",
  39219=>"111100010",
  39220=>"000000000",
  39221=>"011011111",
  39222=>"100000000",
  39223=>"111111111",
  39224=>"100100110",
  39225=>"000000000",
  39226=>"000111010",
  39227=>"111111111",
  39228=>"011111000",
  39229=>"111100000",
  39230=>"111111111",
  39231=>"000000111",
  39232=>"101000000",
  39233=>"111000000",
  39234=>"111110100",
  39235=>"111111111",
  39236=>"001000000",
  39237=>"111111111",
  39238=>"111111111",
  39239=>"111100100",
  39240=>"011111000",
  39241=>"000000110",
  39242=>"111100101",
  39243=>"110000000",
  39244=>"000000000",
  39245=>"001001101",
  39246=>"111011111",
  39247=>"111011001",
  39248=>"011001011",
  39249=>"111111111",
  39250=>"111111111",
  39251=>"111101000",
  39252=>"000000000",
  39253=>"011011001",
  39254=>"110110111",
  39255=>"011011000",
  39256=>"110110010",
  39257=>"111110000",
  39258=>"111111111",
  39259=>"000000000",
  39260=>"000000000",
  39261=>"000000000",
  39262=>"111100000",
  39263=>"001000001",
  39264=>"010010111",
  39265=>"000000000",
  39266=>"111110110",
  39267=>"111111100",
  39268=>"000000000",
  39269=>"111111101",
  39270=>"111001111",
  39271=>"111110110",
  39272=>"111001101",
  39273=>"111111100",
  39274=>"111111111",
  39275=>"000000000",
  39276=>"000001001",
  39277=>"000111111",
  39278=>"000000000",
  39279=>"000000001",
  39280=>"000000000",
  39281=>"111111011",
  39282=>"000000000",
  39283=>"011011011",
  39284=>"000011111",
  39285=>"000000000",
  39286=>"111010000",
  39287=>"000000000",
  39288=>"000000110",
  39289=>"111111111",
  39290=>"100101111",
  39291=>"111111010",
  39292=>"011111000",
  39293=>"110000000",
  39294=>"111111111",
  39295=>"111111111",
  39296=>"111111111",
  39297=>"011111111",
  39298=>"100100111",
  39299=>"000100000",
  39300=>"111001010",
  39301=>"000000000",
  39302=>"010110111",
  39303=>"111111111",
  39304=>"000000101",
  39305=>"110111111",
  39306=>"000001111",
  39307=>"111110000",
  39308=>"111111111",
  39309=>"011011011",
  39310=>"111111001",
  39311=>"000000000",
  39312=>"000000000",
  39313=>"000000011",
  39314=>"011111111",
  39315=>"110000000",
  39316=>"000100000",
  39317=>"000000010",
  39318=>"011001001",
  39319=>"111110000",
  39320=>"111100000",
  39321=>"000100110",
  39322=>"100111111",
  39323=>"111111111",
  39324=>"000010000",
  39325=>"000000000",
  39326=>"110111001",
  39327=>"000000000",
  39328=>"000000000",
  39329=>"111110110",
  39330=>"001111111",
  39331=>"111111111",
  39332=>"001110000",
  39333=>"000001011",
  39334=>"111111001",
  39335=>"100111111",
  39336=>"110111111",
  39337=>"000000000",
  39338=>"001101111",
  39339=>"000000000",
  39340=>"000000000",
  39341=>"000000011",
  39342=>"000000000",
  39343=>"111111000",
  39344=>"111111111",
  39345=>"111111111",
  39346=>"010000000",
  39347=>"100100000",
  39348=>"111101000",
  39349=>"111011001",
  39350=>"000000000",
  39351=>"000000000",
  39352=>"010110111",
  39353=>"111110000",
  39354=>"111110000",
  39355=>"110000000",
  39356=>"111000000",
  39357=>"100111111",
  39358=>"001001100",
  39359=>"000100110",
  39360=>"000000000",
  39361=>"111101111",
  39362=>"000000000",
  39363=>"110111111",
  39364=>"111000000",
  39365=>"011001001",
  39366=>"100100000",
  39367=>"000000000",
  39368=>"011000000",
  39369=>"111111011",
  39370=>"001000000",
  39371=>"000000000",
  39372=>"111101001",
  39373=>"111111111",
  39374=>"101000000",
  39375=>"111111111",
  39376=>"100000000",
  39377=>"111001001",
  39378=>"000000000",
  39379=>"111111010",
  39380=>"000000111",
  39381=>"111111111",
  39382=>"000000000",
  39383=>"011011111",
  39384=>"001100100",
  39385=>"011000000",
  39386=>"011001000",
  39387=>"001000111",
  39388=>"100000000",
  39389=>"111111001",
  39390=>"110110000",
  39391=>"010011111",
  39392=>"111111111",
  39393=>"000000000",
  39394=>"000011011",
  39395=>"111111101",
  39396=>"001000111",
  39397=>"000000100",
  39398=>"101101000",
  39399=>"000000110",
  39400=>"111000000",
  39401=>"100110000",
  39402=>"001000000",
  39403=>"000000000",
  39404=>"111101100",
  39405=>"110110100",
  39406=>"111111111",
  39407=>"000000000",
  39408=>"000000000",
  39409=>"001111111",
  39410=>"001000100",
  39411=>"111010000",
  39412=>"000000110",
  39413=>"000000011",
  39414=>"111111111",
  39415=>"111011001",
  39416=>"111111011",
  39417=>"001001001",
  39418=>"000000000",
  39419=>"000100100",
  39420=>"110111111",
  39421=>"011111111",
  39422=>"000000000",
  39423=>"000110000",
  39424=>"011001100",
  39425=>"000111111",
  39426=>"000000010",
  39427=>"001001001",
  39428=>"110110110",
  39429=>"001001011",
  39430=>"110111110",
  39431=>"111100101",
  39432=>"111000000",
  39433=>"000000000",
  39434=>"000100111",
  39435=>"100110110",
  39436=>"100110110",
  39437=>"110100000",
  39438=>"010011000",
  39439=>"011111000",
  39440=>"110000000",
  39441=>"111111111",
  39442=>"000000000",
  39443=>"001000000",
  39444=>"000000000",
  39445=>"111010010",
  39446=>"010010010",
  39447=>"000110110",
  39448=>"001001010",
  39449=>"111001001",
  39450=>"111000000",
  39451=>"001111101",
  39452=>"110110110",
  39453=>"111011001",
  39454=>"001001001",
  39455=>"110110111",
  39456=>"000110110",
  39457=>"000000000",
  39458=>"111111000",
  39459=>"000000111",
  39460=>"000001111",
  39461=>"001111111",
  39462=>"001000011",
  39463=>"000000110",
  39464=>"000010111",
  39465=>"111111111",
  39466=>"000000111",
  39467=>"111111111",
  39468=>"111111111",
  39469=>"011111111",
  39470=>"000000000",
  39471=>"000000000",
  39472=>"000000000",
  39473=>"000000000",
  39474=>"100100100",
  39475=>"000000000",
  39476=>"011011010",
  39477=>"100101011",
  39478=>"111111111",
  39479=>"110110000",
  39480=>"110100100",
  39481=>"100110000",
  39482=>"000111110",
  39483=>"001111111",
  39484=>"101000000",
  39485=>"010000000",
  39486=>"100000000",
  39487=>"000011111",
  39488=>"000000000",
  39489=>"011001001",
  39490=>"111111001",
  39491=>"001001001",
  39492=>"011010000",
  39493=>"000000000",
  39494=>"101110110",
  39495=>"000000100",
  39496=>"000001001",
  39497=>"000000011",
  39498=>"000010000",
  39499=>"000000010",
  39500=>"111011000",
  39501=>"000110111",
  39502=>"000110110",
  39503=>"001011000",
  39504=>"000100111",
  39505=>"111011000",
  39506=>"000000001",
  39507=>"001001000",
  39508=>"111111111",
  39509=>"110110111",
  39510=>"111101111",
  39511=>"110110100",
  39512=>"010111110",
  39513=>"111000101",
  39514=>"011001111",
  39515=>"110110111",
  39516=>"111111111",
  39517=>"001000000",
  39518=>"111011111",
  39519=>"110000000",
  39520=>"000010011",
  39521=>"010110010",
  39522=>"000000000",
  39523=>"000001000",
  39524=>"111010110",
  39525=>"100100000",
  39526=>"111100111",
  39527=>"111111111",
  39528=>"011011000",
  39529=>"111101011",
  39530=>"011010111",
  39531=>"111000111",
  39532=>"001000000",
  39533=>"010111110",
  39534=>"111001111",
  39535=>"011001101",
  39536=>"000000111",
  39537=>"100101011",
  39538=>"101101001",
  39539=>"000000010",
  39540=>"110000100",
  39541=>"000000100",
  39542=>"001001000",
  39543=>"000000000",
  39544=>"000000000",
  39545=>"100111111",
  39546=>"000100100",
  39547=>"100000110",
  39548=>"011001001",
  39549=>"000010000",
  39550=>"100110111",
  39551=>"001001001",
  39552=>"111111000",
  39553=>"111000000",
  39554=>"000110111",
  39555=>"100100000",
  39556=>"110000000",
  39557=>"111111101",
  39558=>"001000110",
  39559=>"110110110",
  39560=>"001111111",
  39561=>"010000010",
  39562=>"010000000",
  39563=>"111111111",
  39564=>"000110000",
  39565=>"001101001",
  39566=>"111111110",
  39567=>"010110110",
  39568=>"001001111",
  39569=>"111111111",
  39570=>"101100000",
  39571=>"000000100",
  39572=>"000111011",
  39573=>"111111111",
  39574=>"111010010",
  39575=>"000000100",
  39576=>"001001111",
  39577=>"000000111",
  39578=>"010010011",
  39579=>"101101000",
  39580=>"110010000",
  39581=>"010000000",
  39582=>"111110100",
  39583=>"000001111",
  39584=>"000000011",
  39585=>"111111001",
  39586=>"111111111",
  39587=>"011111111",
  39588=>"100111111",
  39589=>"111110010",
  39590=>"001001100",
  39591=>"101111001",
  39592=>"110100100",
  39593=>"000000000",
  39594=>"000001000",
  39595=>"000000100",
  39596=>"011010001",
  39597=>"101101001",
  39598=>"111111010",
  39599=>"000111001",
  39600=>"011001111",
  39601=>"110110110",
  39602=>"001111110",
  39603=>"111111100",
  39604=>"100000000",
  39605=>"111110000",
  39606=>"110110111",
  39607=>"111111111",
  39608=>"111101010",
  39609=>"011111111",
  39610=>"110100000",
  39611=>"111110110",
  39612=>"111000000",
  39613=>"111011000",
  39614=>"011010111",
  39615=>"001000000",
  39616=>"001000111",
  39617=>"000100001",
  39618=>"001111111",
  39619=>"001111111",
  39620=>"011100000",
  39621=>"000010111",
  39622=>"000111111",
  39623=>"110111101",
  39624=>"001001001",
  39625=>"000110100",
  39626=>"010001000",
  39627=>"000011011",
  39628=>"111010000",
  39629=>"000000000",
  39630=>"100010000",
  39631=>"110110000",
  39632=>"101100111",
  39633=>"000001001",
  39634=>"000110000",
  39635=>"000000111",
  39636=>"110101111",
  39637=>"110111011",
  39638=>"001001111",
  39639=>"000001000",
  39640=>"110100100",
  39641=>"010000000",
  39642=>"111111111",
  39643=>"111101111",
  39644=>"111000000",
  39645=>"111110000",
  39646=>"000010000",
  39647=>"110110000",
  39648=>"001001000",
  39649=>"001001111",
  39650=>"111001111",
  39651=>"111111000",
  39652=>"111110000",
  39653=>"111011011",
  39654=>"001111111",
  39655=>"111111000",
  39656=>"001101111",
  39657=>"110110000",
  39658=>"000000000",
  39659=>"111110111",
  39660=>"000000000",
  39661=>"111111111",
  39662=>"000110111",
  39663=>"000111111",
  39664=>"110110000",
  39665=>"110100000",
  39666=>"100000010",
  39667=>"000100100",
  39668=>"111111111",
  39669=>"111100000",
  39670=>"111111000",
  39671=>"001111111",
  39672=>"011111111",
  39673=>"101111111",
  39674=>"111011001",
  39675=>"000000110",
  39676=>"100000111",
  39677=>"011010110",
  39678=>"110110110",
  39679=>"000000000",
  39680=>"100000000",
  39681=>"101101000",
  39682=>"001001001",
  39683=>"100011001",
  39684=>"000110111",
  39685=>"000111000",
  39686=>"000000001",
  39687=>"111111001",
  39688=>"110000001",
  39689=>"111101000",
  39690=>"010000111",
  39691=>"111111000",
  39692=>"001000000",
  39693=>"001000001",
  39694=>"000000111",
  39695=>"111011111",
  39696=>"111110000",
  39697=>"000110000",
  39698=>"111111000",
  39699=>"101110110",
  39700=>"111111111",
  39701=>"101111001",
  39702=>"101111111",
  39703=>"100110100",
  39704=>"010111010",
  39705=>"110010000",
  39706=>"110111000",
  39707=>"010110110",
  39708=>"000000000",
  39709=>"000101000",
  39710=>"000000100",
  39711=>"111111111",
  39712=>"111111000",
  39713=>"100110110",
  39714=>"111011111",
  39715=>"000111000",
  39716=>"111111010",
  39717=>"000000000",
  39718=>"011111000",
  39719=>"000111000",
  39720=>"011011101",
  39721=>"000010000",
  39722=>"111110000",
  39723=>"001111000",
  39724=>"110110111",
  39725=>"000000001",
  39726=>"111111000",
  39727=>"000000111",
  39728=>"101111001",
  39729=>"111111011",
  39730=>"110000000",
  39731=>"111000001",
  39732=>"000010000",
  39733=>"000000100",
  39734=>"111101001",
  39735=>"100110111",
  39736=>"001111000",
  39737=>"001000101",
  39738=>"111100100",
  39739=>"000000111",
  39740=>"000000000",
  39741=>"110111000",
  39742=>"110110000",
  39743=>"000000000",
  39744=>"111111111",
  39745=>"000000100",
  39746=>"111111111",
  39747=>"100110101",
  39748=>"100000001",
  39749=>"100111111",
  39750=>"110110100",
  39751=>"001001011",
  39752=>"111001001",
  39753=>"000111101",
  39754=>"000110000",
  39755=>"010000000",
  39756=>"100110010",
  39757=>"111001111",
  39758=>"110000000",
  39759=>"001011111",
  39760=>"111101100",
  39761=>"101111110",
  39762=>"110111111",
  39763=>"000000011",
  39764=>"001111100",
  39765=>"101000000",
  39766=>"000000000",
  39767=>"000011010",
  39768=>"111000000",
  39769=>"000111001",
  39770=>"111111001",
  39771=>"111011111",
  39772=>"001000111",
  39773=>"000000110",
  39774=>"001111011",
  39775=>"000001000",
  39776=>"001111001",
  39777=>"000110111",
  39778=>"000011110",
  39779=>"001001111",
  39780=>"000000010",
  39781=>"000000000",
  39782=>"000111111",
  39783=>"100110101",
  39784=>"001000001",
  39785=>"000000000",
  39786=>"011111100",
  39787=>"100000000",
  39788=>"100111111",
  39789=>"000100000",
  39790=>"110110000",
  39791=>"110111111",
  39792=>"000000000",
  39793=>"000000000",
  39794=>"100000000",
  39795=>"111111000",
  39796=>"110110010",
  39797=>"000000101",
  39798=>"100000110",
  39799=>"001001011",
  39800=>"000000000",
  39801=>"111111001",
  39802=>"110010000",
  39803=>"001001001",
  39804=>"111111100",
  39805=>"000000000",
  39806=>"111000000",
  39807=>"111111000",
  39808=>"101101110",
  39809=>"010110101",
  39810=>"000000001",
  39811=>"000001111",
  39812=>"111110000",
  39813=>"111011000",
  39814=>"000000001",
  39815=>"111111000",
  39816=>"000111111",
  39817=>"000000100",
  39818=>"000001111",
  39819=>"000000010",
  39820=>"111110111",
  39821=>"000000000",
  39822=>"000100111",
  39823=>"111100100",
  39824=>"001001111",
  39825=>"100110000",
  39826=>"111111000",
  39827=>"010001001",
  39828=>"001000100",
  39829=>"000000000",
  39830=>"001110000",
  39831=>"101111000",
  39832=>"111111111",
  39833=>"110110111",
  39834=>"000000000",
  39835=>"111110000",
  39836=>"111101111",
  39837=>"001111010",
  39838=>"100000000",
  39839=>"000111110",
  39840=>"000000110",
  39841=>"000000000",
  39842=>"111011001",
  39843=>"111101111",
  39844=>"000011000",
  39845=>"001001000",
  39846=>"000000000",
  39847=>"111111111",
  39848=>"001000000",
  39849=>"001000001",
  39850=>"000000000",
  39851=>"000000010",
  39852=>"111111111",
  39853=>"001000000",
  39854=>"111000001",
  39855=>"000000100",
  39856=>"101100001",
  39857=>"111111100",
  39858=>"001110111",
  39859=>"000000000",
  39860=>"111110100",
  39861=>"000001111",
  39862=>"000100110",
  39863=>"000000101",
  39864=>"000000101",
  39865=>"111111000",
  39866=>"000000111",
  39867=>"011111011",
  39868=>"011011011",
  39869=>"110110000",
  39870=>"001011000",
  39871=>"100101001",
  39872=>"111011010",
  39873=>"000000000",
  39874=>"001101001",
  39875=>"001011111",
  39876=>"001000001",
  39877=>"111111001",
  39878=>"001001111",
  39879=>"000111111",
  39880=>"111101111",
  39881=>"000100111",
  39882=>"000001001",
  39883=>"000011000",
  39884=>"111001010",
  39885=>"101111111",
  39886=>"111110001",
  39887=>"111111111",
  39888=>"000111110",
  39889=>"111111011",
  39890=>"111011001",
  39891=>"000000000",
  39892=>"111111100",
  39893=>"001000011",
  39894=>"000001011",
  39895=>"011011001",
  39896=>"111111111",
  39897=>"111111000",
  39898=>"100100111",
  39899=>"111111000",
  39900=>"000111110",
  39901=>"111111000",
  39902=>"100110000",
  39903=>"000100111",
  39904=>"001000000",
  39905=>"111001000",
  39906=>"001111111",
  39907=>"011111111",
  39908=>"110000101",
  39909=>"011011000",
  39910=>"001101000",
  39911=>"000000111",
  39912=>"011111110",
  39913=>"000100110",
  39914=>"001111111",
  39915=>"000100111",
  39916=>"000110111",
  39917=>"111011011",
  39918=>"001000000",
  39919=>"011111111",
  39920=>"000000000",
  39921=>"000110110",
  39922=>"101000000",
  39923=>"001101000",
  39924=>"000000000",
  39925=>"011000000",
  39926=>"000000000",
  39927=>"111100100",
  39928=>"000000111",
  39929=>"011010011",
  39930=>"111111110",
  39931=>"011111000",
  39932=>"011001111",
  39933=>"001000000",
  39934=>"101000111",
  39935=>"000000110",
  39936=>"111100010",
  39937=>"000000111",
  39938=>"010010111",
  39939=>"000010010",
  39940=>"111111101",
  39941=>"000000001",
  39942=>"000000111",
  39943=>"111000000",
  39944=>"000101111",
  39945=>"101101001",
  39946=>"111100111",
  39947=>"000100111",
  39948=>"010111100",
  39949=>"100111111",
  39950=>"111010000",
  39951=>"111111111",
  39952=>"000010111",
  39953=>"100111011",
  39954=>"011111111",
  39955=>"111101111",
  39956=>"111111111",
  39957=>"000000001",
  39958=>"001110000",
  39959=>"011011000",
  39960=>"010000000",
  39961=>"001001001",
  39962=>"000000000",
  39963=>"000011001",
  39964=>"101100100",
  39965=>"101001001",
  39966=>"000000000",
  39967=>"000000111",
  39968=>"000111101",
  39969=>"000001011",
  39970=>"001100000",
  39971=>"110000100",
  39972=>"011000110",
  39973=>"000000000",
  39974=>"011000000",
  39975=>"111111111",
  39976=>"101100000",
  39977=>"000000000",
  39978=>"000000000",
  39979=>"111111111",
  39980=>"001111111",
  39981=>"111101000",
  39982=>"101000000",
  39983=>"001000000",
  39984=>"111111111",
  39985=>"111111101",
  39986=>"111111111",
  39987=>"111111100",
  39988=>"000110000",
  39989=>"010011000",
  39990=>"101101000",
  39991=>"100100000",
  39992=>"111111000",
  39993=>"111111001",
  39994=>"111111111",
  39995=>"000000000",
  39996=>"000000000",
  39997=>"000111111",
  39998=>"001001001",
  39999=>"111111111",
  40000=>"101111111",
  40001=>"001001101",
  40002=>"110111111",
  40003=>"011110111",
  40004=>"000000001",
  40005=>"111111110",
  40006=>"110010111",
  40007=>"000110000",
  40008=>"011011001",
  40009=>"000000000",
  40010=>"111111111",
  40011=>"111111111",
  40012=>"100111111",
  40013=>"100111111",
  40014=>"000000000",
  40015=>"000111111",
  40016=>"111111101",
  40017=>"111000000",
  40018=>"000010011",
  40019=>"001101100",
  40020=>"000001101",
  40021=>"111111100",
  40022=>"001000000",
  40023=>"111111111",
  40024=>"111111111",
  40025=>"110110000",
  40026=>"000000000",
  40027=>"011011011",
  40028=>"111111101",
  40029=>"111111111",
  40030=>"001000000",
  40031=>"001001011",
  40032=>"000000001",
  40033=>"000000000",
  40034=>"000000001",
  40035=>"101101111",
  40036=>"111100100",
  40037=>"111111011",
  40038=>"000111111",
  40039=>"111111111",
  40040=>"110001111",
  40041=>"111101000",
  40042=>"100100100",
  40043=>"000000010",
  40044=>"000000000",
  40045=>"111000110",
  40046=>"001000000",
  40047=>"100000000",
  40048=>"111000100",
  40049=>"001000000",
  40050=>"000010010",
  40051=>"001111111",
  40052=>"111111001",
  40053=>"000111111",
  40054=>"000000001",
  40055=>"101001001",
  40056=>"111111111",
  40057=>"000000000",
  40058=>"000000000",
  40059=>"000000111",
  40060=>"000000100",
  40061=>"000000000",
  40062=>"100000000",
  40063=>"000000000",
  40064=>"000000111",
  40065=>"111111100",
  40066=>"000100111",
  40067=>"111111000",
  40068=>"100000100",
  40069=>"000000110",
  40070=>"001000000",
  40071=>"000100101",
  40072=>"111111011",
  40073=>"101011000",
  40074=>"111101101",
  40075=>"111111111",
  40076=>"111000001",
  40077=>"111111000",
  40078=>"000000000",
  40079=>"111111000",
  40080=>"111111111",
  40081=>"101111111",
  40082=>"000000000",
  40083=>"110110110",
  40084=>"111111111",
  40085=>"001000111",
  40086=>"000001011",
  40087=>"111000000",
  40088=>"001001101",
  40089=>"111111100",
  40090=>"000000000",
  40091=>"010111111",
  40092=>"111111011",
  40093=>"000000100",
  40094=>"011111100",
  40095=>"111111111",
  40096=>"001000000",
  40097=>"100100101",
  40098=>"111101101",
  40099=>"011000010",
  40100=>"000111001",
  40101=>"111111111",
  40102=>"111111011",
  40103=>"000000000",
  40104=>"111111010",
  40105=>"001000100",
  40106=>"111000000",
  40107=>"001000001",
  40108=>"001000000",
  40109=>"000010110",
  40110=>"100110101",
  40111=>"111110110",
  40112=>"111111111",
  40113=>"110110110",
  40114=>"101111001",
  40115=>"111101000",
  40116=>"000000011",
  40117=>"000110100",
  40118=>"000000000",
  40119=>"001111111",
  40120=>"111111011",
  40121=>"111111111",
  40122=>"001111011",
  40123=>"001111110",
  40124=>"111111110",
  40125=>"001000110",
  40126=>"111100111",
  40127=>"111100000",
  40128=>"111110110",
  40129=>"000001111",
  40130=>"000000000",
  40131=>"111001111",
  40132=>"001000000",
  40133=>"000111111",
  40134=>"111001000",
  40135=>"000000101",
  40136=>"111010000",
  40137=>"001001001",
  40138=>"111110111",
  40139=>"111111111",
  40140=>"000011011",
  40141=>"111001000",
  40142=>"000000000",
  40143=>"000000000",
  40144=>"011111111",
  40145=>"000111111",
  40146=>"111111110",
  40147=>"000000000",
  40148=>"000100000",
  40149=>"111111110",
  40150=>"110110110",
  40151=>"111011001",
  40152=>"000000000",
  40153=>"111101111",
  40154=>"000000000",
  40155=>"000000111",
  40156=>"110111000",
  40157=>"001101100",
  40158=>"000011000",
  40159=>"000000000",
  40160=>"000000000",
  40161=>"111111111",
  40162=>"110011111",
  40163=>"000000000",
  40164=>"000000000",
  40165=>"100000000",
  40166=>"110110000",
  40167=>"111111011",
  40168=>"111011000",
  40169=>"111111111",
  40170=>"111001111",
  40171=>"000000000",
  40172=>"000111101",
  40173=>"000000000",
  40174=>"000000001",
  40175=>"100000000",
  40176=>"111111111",
  40177=>"001111111",
  40178=>"000000111",
  40179=>"000111001",
  40180=>"001001011",
  40181=>"000001011",
  40182=>"011000000",
  40183=>"111001000",
  40184=>"111111111",
  40185=>"111111111",
  40186=>"111111111",
  40187=>"100111110",
  40188=>"001100110",
  40189=>"001000110",
  40190=>"110111110",
  40191=>"000110000",
  40192=>"001000000",
  40193=>"000010000",
  40194=>"000000110",
  40195=>"001011111",
  40196=>"110110000",
  40197=>"100111111",
  40198=>"000000001",
  40199=>"000011111",
  40200=>"011010001",
  40201=>"010000100",
  40202=>"000000000",
  40203=>"111111111",
  40204=>"000000000",
  40205=>"000100111",
  40206=>"111111111",
  40207=>"000000000",
  40208=>"111110000",
  40209=>"111111111",
  40210=>"101000000",
  40211=>"000000000",
  40212=>"000000100",
  40213=>"000000000",
  40214=>"001000010",
  40215=>"101101111",
  40216=>"101111001",
  40217=>"111000000",
  40218=>"000000000",
  40219=>"101100110",
  40220=>"001001011",
  40221=>"101011011",
  40222=>"111111111",
  40223=>"000111111",
  40224=>"001000000",
  40225=>"111111101",
  40226=>"000000000",
  40227=>"111110000",
  40228=>"010011011",
  40229=>"111111111",
  40230=>"000111111",
  40231=>"111111101",
  40232=>"111011000",
  40233=>"111111111",
  40234=>"001111111",
  40235=>"000111010",
  40236=>"000000000",
  40237=>"000000000",
  40238=>"000000111",
  40239=>"000000000",
  40240=>"011000000",
  40241=>"000000000",
  40242=>"011111100",
  40243=>"000000011",
  40244=>"100000111",
  40245=>"000011011",
  40246=>"000000000",
  40247=>"000000000",
  40248=>"111100100",
  40249=>"111000000",
  40250=>"111100110",
  40251=>"000000100",
  40252=>"111111111",
  40253=>"110110111",
  40254=>"001000000",
  40255=>"100000000",
  40256=>"000000111",
  40257=>"000110001",
  40258=>"001001001",
  40259=>"111111000",
  40260=>"101111001",
  40261=>"111111100",
  40262=>"000000000",
  40263=>"111111111",
  40264=>"111111111",
  40265=>"111000101",
  40266=>"001111111",
  40267=>"000000111",
  40268=>"000000000",
  40269=>"000010100",
  40270=>"011111101",
  40271=>"000000001",
  40272=>"101000101",
  40273=>"110110111",
  40274=>"000110100",
  40275=>"111111111",
  40276=>"000001000",
  40277=>"111011111",
  40278=>"000000010",
  40279=>"000000100",
  40280=>"000000000",
  40281=>"001111111",
  40282=>"000000001",
  40283=>"011111001",
  40284=>"000000000",
  40285=>"111101000",
  40286=>"000110110",
  40287=>"000000000",
  40288=>"110100100",
  40289=>"111100000",
  40290=>"001000000",
  40291=>"001000000",
  40292=>"000000011",
  40293=>"000101000",
  40294=>"000111111",
  40295=>"001001111",
  40296=>"000011011",
  40297=>"010010000",
  40298=>"001101101",
  40299=>"000100111",
  40300=>"001001001",
  40301=>"001111111",
  40302=>"111111111",
  40303=>"111111111",
  40304=>"000000000",
  40305=>"001000001",
  40306=>"000111111",
  40307=>"111111100",
  40308=>"111110000",
  40309=>"110000001",
  40310=>"100000111",
  40311=>"000111001",
  40312=>"000000111",
  40313=>"000000001",
  40314=>"000000001",
  40315=>"111111111",
  40316=>"111111111",
  40317=>"111111111",
  40318=>"111111110",
  40319=>"101000000",
  40320=>"000000000",
  40321=>"000011001",
  40322=>"111111011",
  40323=>"111111111",
  40324=>"000010000",
  40325=>"000100100",
  40326=>"111110000",
  40327=>"000000000",
  40328=>"000000100",
  40329=>"001001000",
  40330=>"111111000",
  40331=>"000000001",
  40332=>"000111111",
  40333=>"000000000",
  40334=>"101100101",
  40335=>"111111110",
  40336=>"111111000",
  40337=>"111111110",
  40338=>"000000000",
  40339=>"111111111",
  40340=>"000000000",
  40341=>"000000000",
  40342=>"110100000",
  40343=>"000000100",
  40344=>"000011111",
  40345=>"001000000",
  40346=>"111111011",
  40347=>"111111000",
  40348=>"000100111",
  40349=>"000100100",
  40350=>"111111111",
  40351=>"110111111",
  40352=>"000000010",
  40353=>"000000000",
  40354=>"000111111",
  40355=>"111111000",
  40356=>"111110100",
  40357=>"000000000",
  40358=>"110111111",
  40359=>"111111111",
  40360=>"011011111",
  40361=>"111111101",
  40362=>"000100110",
  40363=>"111111111",
  40364=>"110110000",
  40365=>"000000000",
  40366=>"001001011",
  40367=>"111111111",
  40368=>"100100111",
  40369=>"000000000",
  40370=>"000111111",
  40371=>"101000000",
  40372=>"111111111",
  40373=>"110100000",
  40374=>"111011100",
  40375=>"100000000",
  40376=>"111111000",
  40377=>"111111111",
  40378=>"000000000",
  40379=>"000000000",
  40380=>"111111111",
  40381=>"111111111",
  40382=>"000000000",
  40383=>"001011111",
  40384=>"111111111",
  40385=>"100101111",
  40386=>"000000000",
  40387=>"001001001",
  40388=>"111111111",
  40389=>"000000001",
  40390=>"000000000",
  40391=>"000101111",
  40392=>"011001000",
  40393=>"111000000",
  40394=>"000110111",
  40395=>"111111000",
  40396=>"111000000",
  40397=>"111111111",
  40398=>"000000000",
  40399=>"001111111",
  40400=>"000100110",
  40401=>"111111111",
  40402=>"000001000",
  40403=>"011011000",
  40404=>"001000000",
  40405=>"111100000",
  40406=>"011100100",
  40407=>"110110110",
  40408=>"111111000",
  40409=>"000000111",
  40410=>"000000100",
  40411=>"000000000",
  40412=>"101101110",
  40413=>"000000000",
  40414=>"000000000",
  40415=>"000000001",
  40416=>"101101111",
  40417=>"111111111",
  40418=>"111111111",
  40419=>"111111111",
  40420=>"111111000",
  40421=>"110111111",
  40422=>"000100110",
  40423=>"111111111",
  40424=>"001000000",
  40425=>"000000000",
  40426=>"000000000",
  40427=>"011111000",
  40428=>"100111111",
  40429=>"100110110",
  40430=>"010111111",
  40431=>"000100000",
  40432=>"111111111",
  40433=>"100111111",
  40434=>"001000000",
  40435=>"111111111",
  40436=>"000000000",
  40437=>"000000000",
  40438=>"111111100",
  40439=>"000000000",
  40440=>"000000000",
  40441=>"111100100",
  40442=>"000000011",
  40443=>"000000000",
  40444=>"111111000",
  40445=>"000001011",
  40446=>"000000000",
  40447=>"111111111",
  40448=>"000000000",
  40449=>"111111111",
  40450=>"000000100",
  40451=>"110011011",
  40452=>"000001111",
  40453=>"101110000",
  40454=>"111111111",
  40455=>"111111111",
  40456=>"111111111",
  40457=>"000000111",
  40458=>"100101101",
  40459=>"000000000",
  40460=>"001011001",
  40461=>"110111111",
  40462=>"100100111",
  40463=>"000100111",
  40464=>"111111111",
  40465=>"111111101",
  40466=>"001001000",
  40467=>"110000111",
  40468=>"000011001",
  40469=>"010010111",
  40470=>"110100000",
  40471=>"100100110",
  40472=>"001111111",
  40473=>"000000000",
  40474=>"000000111",
  40475=>"111011011",
  40476=>"000000000",
  40477=>"000000000",
  40478=>"001001010",
  40479=>"001111111",
  40480=>"110110010",
  40481=>"111111110",
  40482=>"111111100",
  40483=>"000000001",
  40484=>"000100110",
  40485=>"000000000",
  40486=>"000000111",
  40487=>"111111111",
  40488=>"000000101",
  40489=>"101110111",
  40490=>"110011001",
  40491=>"100100100",
  40492=>"111101000",
  40493=>"111111001",
  40494=>"111111001",
  40495=>"111110000",
  40496=>"000000000",
  40497=>"010000000",
  40498=>"100100100",
  40499=>"100000000",
  40500=>"000000000",
  40501=>"000000000",
  40502=>"000000000",
  40503=>"110110100",
  40504=>"001100001",
  40505=>"111111000",
  40506=>"000001111",
  40507=>"101001000",
  40508=>"111001000",
  40509=>"110010111",
  40510=>"111111110",
  40511=>"101101111",
  40512=>"100000000",
  40513=>"010010110",
  40514=>"000000100",
  40515=>"000000000",
  40516=>"000000000",
  40517=>"001000110",
  40518=>"000111111",
  40519=>"000000000",
  40520=>"000000000",
  40521=>"000000111",
  40522=>"111111100",
  40523=>"000000001",
  40524=>"111111111",
  40525=>"000010010",
  40526=>"000110111",
  40527=>"111100100",
  40528=>"111111001",
  40529=>"001011000",
  40530=>"100000000",
  40531=>"100000001",
  40532=>"000000000",
  40533=>"111111111",
  40534=>"000000000",
  40535=>"110110100",
  40536=>"000011111",
  40537=>"111000100",
  40538=>"000000110",
  40539=>"000100111",
  40540=>"000000000",
  40541=>"000000000",
  40542=>"011011011",
  40543=>"111111111",
  40544=>"111010000",
  40545=>"100110110",
  40546=>"011111111",
  40547=>"000000000",
  40548=>"011011111",
  40549=>"111000000",
  40550=>"000000000",
  40551=>"111001000",
  40552=>"111111111",
  40553=>"000000000",
  40554=>"000011111",
  40555=>"000000000",
  40556=>"001011000",
  40557=>"000000000",
  40558=>"110010011",
  40559=>"011111111",
  40560=>"111110000",
  40561=>"000000000",
  40562=>"111000000",
  40563=>"000000000",
  40564=>"100100111",
  40565=>"110100110",
  40566=>"000000000",
  40567=>"000100000",
  40568=>"111111101",
  40569=>"110111111",
  40570=>"010000110",
  40571=>"000000000",
  40572=>"110110000",
  40573=>"000000000",
  40574=>"000000011",
  40575=>"111111111",
  40576=>"000000000",
  40577=>"111111111",
  40578=>"110111111",
  40579=>"110000000",
  40580=>"110111111",
  40581=>"001000111",
  40582=>"010000110",
  40583=>"111111000",
  40584=>"000101111",
  40585=>"111110110",
  40586=>"000001111",
  40587=>"110101001",
  40588=>"101101101",
  40589=>"111111111",
  40590=>"110000000",
  40591=>"110110011",
  40592=>"011011011",
  40593=>"111110010",
  40594=>"111111111",
  40595=>"111111111",
  40596=>"000000000",
  40597=>"100000000",
  40598=>"111111111",
  40599=>"000000011",
  40600=>"000000000",
  40601=>"000000001",
  40602=>"000100100",
  40603=>"000000000",
  40604=>"110111111",
  40605=>"111110110",
  40606=>"110000000",
  40607=>"100100111",
  40608=>"111010000",
  40609=>"111111111",
  40610=>"000000000",
  40611=>"111100010",
  40612=>"010111100",
  40613=>"111100111",
  40614=>"111111111",
  40615=>"111111010",
  40616=>"000000001",
  40617=>"011111111",
  40618=>"111111111",
  40619=>"011000000",
  40620=>"010110110",
  40621=>"111110000",
  40622=>"111110110",
  40623=>"011001000",
  40624=>"000111000",
  40625=>"100100000",
  40626=>"111111110",
  40627=>"010111111",
  40628=>"000000000",
  40629=>"111110100",
  40630=>"010110111",
  40631=>"000000000",
  40632=>"101000100",
  40633=>"111111011",
  40634=>"000000000",
  40635=>"111011000",
  40636=>"111111111",
  40637=>"000101111",
  40638=>"111111111",
  40639=>"000100000",
  40640=>"111111111",
  40641=>"100110111",
  40642=>"111111111",
  40643=>"001000111",
  40644=>"000000000",
  40645=>"000000000",
  40646=>"001111111",
  40647=>"000000000",
  40648=>"111010000",
  40649=>"100111111",
  40650=>"000000100",
  40651=>"000000000",
  40652=>"000111111",
  40653=>"000110110",
  40654=>"000000101",
  40655=>"111111111",
  40656=>"111111111",
  40657=>"001000000",
  40658=>"010110100",
  40659=>"000000000",
  40660=>"100101111",
  40661=>"111111110",
  40662=>"000000000",
  40663=>"001111101",
  40664=>"100111111",
  40665=>"000001011",
  40666=>"000000000",
  40667=>"101100101",
  40668=>"111100000",
  40669=>"001011001",
  40670=>"101111111",
  40671=>"000000000",
  40672=>"000001111",
  40673=>"000001000",
  40674=>"000000000",
  40675=>"111111111",
  40676=>"000100101",
  40677=>"000100000",
  40678=>"001011111",
  40679=>"111111111",
  40680=>"111111100",
  40681=>"111111111",
  40682=>"011000000",
  40683=>"000000100",
  40684=>"000000000",
  40685=>"000001001",
  40686=>"001111110",
  40687=>"000000100",
  40688=>"110110111",
  40689=>"110111011",
  40690=>"010000000",
  40691=>"000001011",
  40692=>"100101111",
  40693=>"001101111",
  40694=>"100000000",
  40695=>"111111111",
  40696=>"000101110",
  40697=>"111111111",
  40698=>"111111011",
  40699=>"111111010",
  40700=>"100110011",
  40701=>"111111111",
  40702=>"111111111",
  40703=>"100000000",
  40704=>"110111111",
  40705=>"000001001",
  40706=>"111111000",
  40707=>"111111110",
  40708=>"100000111",
  40709=>"000100100",
  40710=>"000000000",
  40711=>"000011101",
  40712=>"110111111",
  40713=>"111111001",
  40714=>"111111111",
  40715=>"000000000",
  40716=>"111000000",
  40717=>"100111111",
  40718=>"011001011",
  40719=>"110111000",
  40720=>"100000101",
  40721=>"111111111",
  40722=>"111111111",
  40723=>"000111111",
  40724=>"111111111",
  40725=>"110111001",
  40726=>"111001000",
  40727=>"000000000",
  40728=>"000100111",
  40729=>"111001111",
  40730=>"000000000",
  40731=>"111110111",
  40732=>"000000000",
  40733=>"111111111",
  40734=>"111111111",
  40735=>"111111100",
  40736=>"100110000",
  40737=>"000000000",
  40738=>"001000000",
  40739=>"011011111",
  40740=>"000000000",
  40741=>"000000111",
  40742=>"100110100",
  40743=>"001111111",
  40744=>"111111111",
  40745=>"111100000",
  40746=>"101000000",
  40747=>"111111111",
  40748=>"111111111",
  40749=>"111111111",
  40750=>"110111111",
  40751=>"000000000",
  40752=>"001000001",
  40753=>"000111111",
  40754=>"110010010",
  40755=>"111111011",
  40756=>"000000111",
  40757=>"000000000",
  40758=>"000000000",
  40759=>"000000101",
  40760=>"011011000",
  40761=>"111111000",
  40762=>"000000000",
  40763=>"000000000",
  40764=>"001000001",
  40765=>"000000110",
  40766=>"000110111",
  40767=>"010000100",
  40768=>"111111111",
  40769=>"000000100",
  40770=>"000000000",
  40771=>"111111111",
  40772=>"000000110",
  40773=>"000000110",
  40774=>"100000000",
  40775=>"100000000",
  40776=>"000000000",
  40777=>"110100111",
  40778=>"001111111",
  40779=>"011000110",
  40780=>"000000000",
  40781=>"001000000",
  40782=>"000000000",
  40783=>"000000000",
  40784=>"000000000",
  40785=>"111111111",
  40786=>"010000000",
  40787=>"000000000",
  40788=>"000000000",
  40789=>"011001011",
  40790=>"000000000",
  40791=>"111111111",
  40792=>"000000000",
  40793=>"111101111",
  40794=>"111111000",
  40795=>"000000011",
  40796=>"111011011",
  40797=>"100000000",
  40798=>"110110110",
  40799=>"011001001",
  40800=>"100111110",
  40801=>"000000000",
  40802=>"110110011",
  40803=>"111101101",
  40804=>"110100110",
  40805=>"111101000",
  40806=>"000000000",
  40807=>"111111111",
  40808=>"110010010",
  40809=>"111111111",
  40810=>"000000000",
  40811=>"111111111",
  40812=>"000000000",
  40813=>"000000100",
  40814=>"110111111",
  40815=>"000000000",
  40816=>"111000000",
  40817=>"111111111",
  40818=>"000110111",
  40819=>"001011000",
  40820=>"010001001",
  40821=>"100100111",
  40822=>"111001001",
  40823=>"001001001",
  40824=>"111111111",
  40825=>"111111110",
  40826=>"110110111",
  40827=>"010000100",
  40828=>"110000101",
  40829=>"111111111",
  40830=>"000000000",
  40831=>"000011111",
  40832=>"000000110",
  40833=>"111000000",
  40834=>"000000010",
  40835=>"000000101",
  40836=>"000001111",
  40837=>"101101111",
  40838=>"111111101",
  40839=>"001001011",
  40840=>"000000101",
  40841=>"111111100",
  40842=>"000000010",
  40843=>"011101001",
  40844=>"001001111",
  40845=>"111111111",
  40846=>"000000000",
  40847=>"000000010",
  40848=>"111010000",
  40849=>"111000000",
  40850=>"000000000",
  40851=>"100000100",
  40852=>"111111111",
  40853=>"000010000",
  40854=>"001001101",
  40855=>"110111110",
  40856=>"001001000",
  40857=>"000001001",
  40858=>"000000011",
  40859=>"000000000",
  40860=>"110001000",
  40861=>"000000000",
  40862=>"110100000",
  40863=>"001000000",
  40864=>"000000010",
  40865=>"010010010",
  40866=>"110000000",
  40867=>"111111111",
  40868=>"110111111",
  40869=>"111111111",
  40870=>"100111111",
  40871=>"000000110",
  40872=>"000000111",
  40873=>"011111111",
  40874=>"111111111",
  40875=>"110110000",
  40876=>"100100110",
  40877=>"111001000",
  40878=>"000001000",
  40879=>"001000101",
  40880=>"000000000",
  40881=>"110111111",
  40882=>"111111111",
  40883=>"100101111",
  40884=>"111111111",
  40885=>"100100110",
  40886=>"111100000",
  40887=>"001011111",
  40888=>"001000000",
  40889=>"111111111",
  40890=>"111111111",
  40891=>"000000100",
  40892=>"111111111",
  40893=>"100100001",
  40894=>"000001000",
  40895=>"000000000",
  40896=>"111101000",
  40897=>"000000000",
  40898=>"000000001",
  40899=>"000000000",
  40900=>"011011111",
  40901=>"110110100",
  40902=>"100000010",
  40903=>"000000100",
  40904=>"000011010",
  40905=>"100110111",
  40906=>"110010000",
  40907=>"111111111",
  40908=>"111111000",
  40909=>"111111111",
  40910=>"000000100",
  40911=>"000000011",
  40912=>"111111111",
  40913=>"110111111",
  40914=>"001000000",
  40915=>"000000011",
  40916=>"000000000",
  40917=>"100111111",
  40918=>"000000000",
  40919=>"100100100",
  40920=>"111111111",
  40921=>"000000010",
  40922=>"111111111",
  40923=>"111111111",
  40924=>"111111110",
  40925=>"100000100",
  40926=>"000000000",
  40927=>"000000000",
  40928=>"111000111",
  40929=>"111111111",
  40930=>"000000000",
  40931=>"111111111",
  40932=>"111111111",
  40933=>"111111000",
  40934=>"000011000",
  40935=>"111111101",
  40936=>"111111000",
  40937=>"000100100",
  40938=>"011011011",
  40939=>"100111111",
  40940=>"111111100",
  40941=>"111111010",
  40942=>"111111111",
  40943=>"111110111",
  40944=>"111100000",
  40945=>"111111110",
  40946=>"111111111",
  40947=>"101111110",
  40948=>"001001111",
  40949=>"111111111",
  40950=>"000000000",
  40951=>"110100110",
  40952=>"000000111",
  40953=>"100000000",
  40954=>"111100000",
  40955=>"000000000",
  40956=>"111111110",
  40957=>"111111000",
  40958=>"100111111",
  40959=>"111110110",
  40960=>"001000000",
  40961=>"110000000",
  40962=>"111111111",
  40963=>"111110011",
  40964=>"111000001",
  40965=>"111111000",
  40966=>"001000001",
  40967=>"111111111",
  40968=>"011000000",
  40969=>"000000000",
  40970=>"111010000",
  40971=>"011010110",
  40972=>"111111010",
  40973=>"111111001",
  40974=>"111111111",
  40975=>"000000000",
  40976=>"100000011",
  40977=>"000000000",
  40978=>"000000000",
  40979=>"000000001",
  40980=>"001000000",
  40981=>"111101111",
  40982=>"000000000",
  40983=>"000000000",
  40984=>"111111111",
  40985=>"000000000",
  40986=>"111111001",
  40987=>"000000000",
  40988=>"111111111",
  40989=>"111100000",
  40990=>"110011001",
  40991=>"000000001",
  40992=>"000000001",
  40993=>"110110110",
  40994=>"000000000",
  40995=>"111111101",
  40996=>"111111000",
  40997=>"000000000",
  40998=>"000000000",
  40999=>"000000011",
  41000=>"000101101",
  41001=>"000000000",
  41002=>"111111111",
  41003=>"111100111",
  41004=>"111111111",
  41005=>"000000010",
  41006=>"000000111",
  41007=>"111101011",
  41008=>"111111101",
  41009=>"000000000",
  41010=>"111111001",
  41011=>"100111101",
  41012=>"000001101",
  41013=>"000111111",
  41014=>"011001111",
  41015=>"110110110",
  41016=>"111110001",
  41017=>"110000000",
  41018=>"111001001",
  41019=>"000110110",
  41020=>"000000000",
  41021=>"000001111",
  41022=>"000000100",
  41023=>"000000000",
  41024=>"110110111",
  41025=>"000000000",
  41026=>"111111000",
  41027=>"111111000",
  41028=>"000000000",
  41029=>"011001111",
  41030=>"001000010",
  41031=>"111111110",
  41032=>"110110110",
  41033=>"000000000",
  41034=>"111111000",
  41035=>"010000001",
  41036=>"001000000",
  41037=>"111111110",
  41038=>"100110111",
  41039=>"000000000",
  41040=>"011111111",
  41041=>"001001011",
  41042=>"001011111",
  41043=>"000110111",
  41044=>"000000100",
  41045=>"000000110",
  41046=>"100000100",
  41047=>"000000111",
  41048=>"000101101",
  41049=>"111100001",
  41050=>"111111000",
  41051=>"110100000",
  41052=>"000110110",
  41053=>"111111111",
  41054=>"001001000",
  41055=>"111110111",
  41056=>"000010110",
  41057=>"000101000",
  41058=>"111110100",
  41059=>"000000000",
  41060=>"110000000",
  41061=>"000000111",
  41062=>"000000111",
  41063=>"111111111",
  41064=>"111111000",
  41065=>"001001011",
  41066=>"111111000",
  41067=>"000000001",
  41068=>"000000110",
  41069=>"111111111",
  41070=>"110111111",
  41071=>"010111111",
  41072=>"000000111",
  41073=>"100000000",
  41074=>"100111111",
  41075=>"000000000",
  41076=>"011011111",
  41077=>"011011000",
  41078=>"110100111",
  41079=>"110000010",
  41080=>"000000000",
  41081=>"000000000",
  41082=>"000000101",
  41083=>"000000000",
  41084=>"110110100",
  41085=>"000001100",
  41086=>"001001101",
  41087=>"000000000",
  41088=>"011011111",
  41089=>"111111111",
  41090=>"111000000",
  41091=>"000011111",
  41092=>"111111000",
  41093=>"111000000",
  41094=>"111011000",
  41095=>"110110010",
  41096=>"000000000",
  41097=>"000000000",
  41098=>"000000111",
  41099=>"000111111",
  41100=>"000100001",
  41101=>"000000000",
  41102=>"000000000",
  41103=>"000000000",
  41104=>"111111010",
  41105=>"000000110",
  41106=>"100000011",
  41107=>"000000000",
  41108=>"111111111",
  41109=>"000111111",
  41110=>"111000000",
  41111=>"111000000",
  41112=>"000000100",
  41113=>"111111011",
  41114=>"111111111",
  41115=>"011111111",
  41116=>"111111111",
  41117=>"000000000",
  41118=>"000000000",
  41119=>"000000111",
  41120=>"110000111",
  41121=>"000000000",
  41122=>"000000000",
  41123=>"000000011",
  41124=>"000100111",
  41125=>"111001000",
  41126=>"001000000",
  41127=>"110111111",
  41128=>"000000000",
  41129=>"000011000",
  41130=>"000111111",
  41131=>"111011111",
  41132=>"111111111",
  41133=>"100100100",
  41134=>"001001101",
  41135=>"010010000",
  41136=>"111000000",
  41137=>"000000000",
  41138=>"111111011",
  41139=>"011011000",
  41140=>"001001101",
  41141=>"111111001",
  41142=>"000000000",
  41143=>"100111000",
  41144=>"000000110",
  41145=>"010000000",
  41146=>"000000100",
  41147=>"000001011",
  41148=>"100000100",
  41149=>"000000000",
  41150=>"111111111",
  41151=>"001000000",
  41152=>"011011000",
  41153=>"011111111",
  41154=>"000000000",
  41155=>"111001000",
  41156=>"111000000",
  41157=>"000001000",
  41158=>"000000010",
  41159=>"111010111",
  41160=>"110000000",
  41161=>"000000100",
  41162=>"110111111",
  41163=>"111101100",
  41164=>"110101111",
  41165=>"000000011",
  41166=>"110111111",
  41167=>"100110100",
  41168=>"100000000",
  41169=>"000000000",
  41170=>"000110010",
  41171=>"111111111",
  41172=>"101101101",
  41173=>"000000000",
  41174=>"111111111",
  41175=>"110011111",
  41176=>"110010000",
  41177=>"111111111",
  41178=>"000110000",
  41179=>"111111000",
  41180=>"111111111",
  41181=>"000000100",
  41182=>"111111111",
  41183=>"111111001",
  41184=>"111111111",
  41185=>"001000111",
  41186=>"111111010",
  41187=>"111111111",
  41188=>"000100001",
  41189=>"001001001",
  41190=>"000000110",
  41191=>"000001011",
  41192=>"000000000",
  41193=>"100111011",
  41194=>"111111111",
  41195=>"111000000",
  41196=>"000001000",
  41197=>"110000000",
  41198=>"110111111",
  41199=>"000000000",
  41200=>"000001000",
  41201=>"000000000",
  41202=>"010000010",
  41203=>"000000111",
  41204=>"000000000",
  41205=>"011011111",
  41206=>"111110010",
  41207=>"000000000",
  41208=>"000000010",
  41209=>"000001001",
  41210=>"000000110",
  41211=>"000000011",
  41212=>"001001111",
  41213=>"000011111",
  41214=>"111101111",
  41215=>"111111111",
  41216=>"100111111",
  41217=>"000100111",
  41218=>"110111001",
  41219=>"111111111",
  41220=>"001001111",
  41221=>"000000000",
  41222=>"000000111",
  41223=>"110000000",
  41224=>"001101011",
  41225=>"010000000",
  41226=>"111011011",
  41227=>"000011111",
  41228=>"000010110",
  41229=>"000000100",
  41230=>"111111101",
  41231=>"101000000",
  41232=>"111111000",
  41233=>"111111111",
  41234=>"100100101",
  41235=>"000010111",
  41236=>"000001000",
  41237=>"110010000",
  41238=>"110110000",
  41239=>"000000001",
  41240=>"000110110",
  41241=>"000000011",
  41242=>"001000000",
  41243=>"111011000",
  41244=>"000100111",
  41245=>"100000000",
  41246=>"111111001",
  41247=>"000111110",
  41248=>"000010010",
  41249=>"111001011",
  41250=>"111111111",
  41251=>"001001001",
  41252=>"000100111",
  41253=>"011111111",
  41254=>"000000000",
  41255=>"110000100",
  41256=>"111111011",
  41257=>"011001111",
  41258=>"011000000",
  41259=>"101000101",
  41260=>"000000100",
  41261=>"001011011",
  41262=>"000000000",
  41263=>"000000010",
  41264=>"111011001",
  41265=>"101111111",
  41266=>"111111100",
  41267=>"010111111",
  41268=>"000000000",
  41269=>"111111111",
  41270=>"000000011",
  41271=>"000000000",
  41272=>"110000000",
  41273=>"111000000",
  41274=>"111101000",
  41275=>"101000000",
  41276=>"111000011",
  41277=>"111110010",
  41278=>"000000000",
  41279=>"000100101",
  41280=>"111001011",
  41281=>"000000000",
  41282=>"111111111",
  41283=>"001000000",
  41284=>"111011111",
  41285=>"000000000",
  41286=>"011000011",
  41287=>"111111111",
  41288=>"111101000",
  41289=>"000000000",
  41290=>"000011011",
  41291=>"000010110",
  41292=>"001000000",
  41293=>"010000000",
  41294=>"111111110",
  41295=>"000111111",
  41296=>"011011000",
  41297=>"111111000",
  41298=>"011001111",
  41299=>"111110000",
  41300=>"000111111",
  41301=>"011011011",
  41302=>"111111000",
  41303=>"010010111",
  41304=>"111111111",
  41305=>"111011000",
  41306=>"110010000",
  41307=>"000111111",
  41308=>"111111011",
  41309=>"100000100",
  41310=>"000000000",
  41311=>"011001000",
  41312=>"000000011",
  41313=>"111111111",
  41314=>"011111000",
  41315=>"111111111",
  41316=>"111011111",
  41317=>"000000000",
  41318=>"000101101",
  41319=>"100100100",
  41320=>"000000111",
  41321=>"000000011",
  41322=>"000000111",
  41323=>"010110100",
  41324=>"001111110",
  41325=>"111111111",
  41326=>"000000000",
  41327=>"110000000",
  41328=>"011111000",
  41329=>"010111000",
  41330=>"001000000",
  41331=>"000000001",
  41332=>"111100100",
  41333=>"001011001",
  41334=>"000000001",
  41335=>"110110111",
  41336=>"000000011",
  41337=>"111000000",
  41338=>"000000000",
  41339=>"000000000",
  41340=>"000000000",
  41341=>"100000000",
  41342=>"000000101",
  41343=>"000000000",
  41344=>"000000000",
  41345=>"011011011",
  41346=>"110110111",
  41347=>"000000000",
  41348=>"000000111",
  41349=>"001001011",
  41350=>"000000000",
  41351=>"000111111",
  41352=>"111111000",
  41353=>"111111000",
  41354=>"000000000",
  41355=>"111011001",
  41356=>"111001001",
  41357=>"000000111",
  41358=>"001000000",
  41359=>"000110100",
  41360=>"010111010",
  41361=>"111110110",
  41362=>"111111000",
  41363=>"100000010",
  41364=>"000000000",
  41365=>"000000000",
  41366=>"100000000",
  41367=>"000000000",
  41368=>"111000001",
  41369=>"000000110",
  41370=>"000000000",
  41371=>"110000000",
  41372=>"111100111",
  41373=>"001000011",
  41374=>"000000000",
  41375=>"101000000",
  41376=>"111000000",
  41377=>"111111111",
  41378=>"000000000",
  41379=>"111111000",
  41380=>"000001000",
  41381=>"110111000",
  41382=>"000111111",
  41383=>"111111010",
  41384=>"110010000",
  41385=>"000000110",
  41386=>"000100100",
  41387=>"100000000",
  41388=>"000000000",
  41389=>"001111111",
  41390=>"100110111",
  41391=>"000111111",
  41392=>"110111011",
  41393=>"000000000",
  41394=>"111111111",
  41395=>"111111110",
  41396=>"111111000",
  41397=>"111000000",
  41398=>"111011000",
  41399=>"000000000",
  41400=>"110000000",
  41401=>"000000000",
  41402=>"100000000",
  41403=>"011000111",
  41404=>"010000000",
  41405=>"001000000",
  41406=>"000010000",
  41407=>"101000110",
  41408=>"110100110",
  41409=>"111010000",
  41410=>"000000111",
  41411=>"100000000",
  41412=>"111100100",
  41413=>"110011011",
  41414=>"111110111",
  41415=>"111101101",
  41416=>"100000101",
  41417=>"111111001",
  41418=>"000011001",
  41419=>"000000011",
  41420=>"110000000",
  41421=>"111000000",
  41422=>"100000011",
  41423=>"000000000",
  41424=>"011000000",
  41425=>"000000001",
  41426=>"111111111",
  41427=>"000000111",
  41428=>"111101111",
  41429=>"111100100",
  41430=>"000000111",
  41431=>"000010000",
  41432=>"111011011",
  41433=>"111010110",
  41434=>"000111111",
  41435=>"000110110",
  41436=>"000000000",
  41437=>"000000100",
  41438=>"111111001",
  41439=>"111101111",
  41440=>"111001001",
  41441=>"111011000",
  41442=>"000000100",
  41443=>"011010001",
  41444=>"111011000",
  41445=>"000000001",
  41446=>"000000111",
  41447=>"000000110",
  41448=>"000111111",
  41449=>"111111111",
  41450=>"000000111",
  41451=>"000000000",
  41452=>"101000000",
  41453=>"001011011",
  41454=>"111100100",
  41455=>"000000000",
  41456=>"110110110",
  41457=>"000000000",
  41458=>"100111011",
  41459=>"111000000",
  41460=>"000111111",
  41461=>"000100000",
  41462=>"000000000",
  41463=>"110111111",
  41464=>"000000001",
  41465=>"001111111",
  41466=>"111111111",
  41467=>"111111001",
  41468=>"111111111",
  41469=>"000111111",
  41470=>"110000000",
  41471=>"000000000",
  41472=>"110111111",
  41473=>"111011011",
  41474=>"111000001",
  41475=>"110111011",
  41476=>"000000000",
  41477=>"100000001",
  41478=>"111111110",
  41479=>"000000000",
  41480=>"111111111",
  41481=>"110000000",
  41482=>"111001111",
  41483=>"111111111",
  41484=>"001000000",
  41485=>"000000000",
  41486=>"011011111",
  41487=>"101000100",
  41488=>"111000000",
  41489=>"000000011",
  41490=>"111001000",
  41491=>"000000000",
  41492=>"111110110",
  41493=>"000000111",
  41494=>"111001001",
  41495=>"111111001",
  41496=>"000000001",
  41497=>"111100000",
  41498=>"111110000",
  41499=>"111111111",
  41500=>"111111111",
  41501=>"100101000",
  41502=>"100100111",
  41503=>"111111000",
  41504=>"111111111",
  41505=>"001001000",
  41506=>"001111100",
  41507=>"110001111",
  41508=>"111111111",
  41509=>"111111110",
  41510=>"111111111",
  41511=>"100000000",
  41512=>"001000000",
  41513=>"000000001",
  41514=>"111111111",
  41515=>"000000000",
  41516=>"000110100",
  41517=>"111101111",
  41518=>"001001001",
  41519=>"110000010",
  41520=>"110111111",
  41521=>"100100111",
  41522=>"111111111",
  41523=>"000000011",
  41524=>"111010011",
  41525=>"111000000",
  41526=>"001001001",
  41527=>"011011000",
  41528=>"111111111",
  41529=>"100111111",
  41530=>"000111111",
  41531=>"000001000",
  41532=>"000000000",
  41533=>"000000111",
  41534=>"110110111",
  41535=>"110111110",
  41536=>"000110111",
  41537=>"111111100",
  41538=>"000100000",
  41539=>"010111111",
  41540=>"000000000",
  41541=>"000000000",
  41542=>"000100110",
  41543=>"111111100",
  41544=>"001010010",
  41545=>"001000000",
  41546=>"000000000",
  41547=>"101111111",
  41548=>"000010011",
  41549=>"000111000",
  41550=>"000000000",
  41551=>"111001001",
  41552=>"011110110",
  41553=>"010011011",
  41554=>"110110111",
  41555=>"110110110",
  41556=>"000000000",
  41557=>"111101100",
  41558=>"000000000",
  41559=>"111111111",
  41560=>"000000000",
  41561=>"001011111",
  41562=>"000000000",
  41563=>"001011000",
  41564=>"111111111",
  41565=>"000000000",
  41566=>"011111000",
  41567=>"110000111",
  41568=>"111111111",
  41569=>"000000000",
  41570=>"101001001",
  41571=>"111111111",
  41572=>"000000000",
  41573=>"110000010",
  41574=>"111000000",
  41575=>"111100000",
  41576=>"000000000",
  41577=>"000000000",
  41578=>"100111100",
  41579=>"111111110",
  41580=>"111111011",
  41581=>"101111111",
  41582=>"000011111",
  41583=>"000000110",
  41584=>"000001111",
  41585=>"011000000",
  41586=>"101000100",
  41587=>"111111101",
  41588=>"000111111",
  41589=>"111111111",
  41590=>"111111111",
  41591=>"000001111",
  41592=>"111000000",
  41593=>"110010111",
  41594=>"111001001",
  41595=>"000000000",
  41596=>"110110010",
  41597=>"000100000",
  41598=>"111111111",
  41599=>"000000000",
  41600=>"111111111",
  41601=>"101111001",
  41602=>"111110111",
  41603=>"010111111",
  41604=>"001000000",
  41605=>"000000000",
  41606=>"111111111",
  41607=>"110111111",
  41608=>"111111111",
  41609=>"111111000",
  41610=>"100101111",
  41611=>"100100110",
  41612=>"100000000",
  41613=>"111111111",
  41614=>"100010000",
  41615=>"100100101",
  41616=>"000000000",
  41617=>"000011010",
  41618=>"111110000",
  41619=>"000100100",
  41620=>"001111111",
  41621=>"000000000",
  41622=>"111111111",
  41623=>"111111011",
  41624=>"000000111",
  41625=>"111111000",
  41626=>"011111111",
  41627=>"111111111",
  41628=>"001101100",
  41629=>"101001011",
  41630=>"101000000",
  41631=>"000000000",
  41632=>"111111110",
  41633=>"110011000",
  41634=>"110110100",
  41635=>"111101100",
  41636=>"111001001",
  41637=>"111110100",
  41638=>"111000111",
  41639=>"001000000",
  41640=>"111111111",
  41641=>"111000101",
  41642=>"001000000",
  41643=>"011011111",
  41644=>"101101001",
  41645=>"000000010",
  41646=>"000000101",
  41647=>"000000000",
  41648=>"111111111",
  41649=>"000111111",
  41650=>"101100100",
  41651=>"000000000",
  41652=>"100110010",
  41653=>"000000000",
  41654=>"111111111",
  41655=>"111111100",
  41656=>"110100000",
  41657=>"111000111",
  41658=>"001100100",
  41659=>"101000000",
  41660=>"000000000",
  41661=>"100100100",
  41662=>"000000000",
  41663=>"111111111",
  41664=>"100110110",
  41665=>"000000000",
  41666=>"000100110",
  41667=>"111111111",
  41668=>"110000000",
  41669=>"111011111",
  41670=>"111111001",
  41671=>"110110110",
  41672=>"000000000",
  41673=>"000100111",
  41674=>"110100010",
  41675=>"000100111",
  41676=>"000011011",
  41677=>"110111111",
  41678=>"100000000",
  41679=>"100110000",
  41680=>"111001000",
  41681=>"111001101",
  41682=>"000000000",
  41683=>"001000000",
  41684=>"000010000",
  41685=>"000000000",
  41686=>"011000000",
  41687=>"110000000",
  41688=>"111111111",
  41689=>"111111111",
  41690=>"111111111",
  41691=>"000000100",
  41692=>"110110110",
  41693=>"000000000",
  41694=>"000000000",
  41695=>"111110110",
  41696=>"000000000",
  41697=>"111101110",
  41698=>"000111111",
  41699=>"100100100",
  41700=>"000000000",
  41701=>"000000000",
  41702=>"111111111",
  41703=>"111111111",
  41704=>"000000000",
  41705=>"011011111",
  41706=>"001011111",
  41707=>"000000011",
  41708=>"110110000",
  41709=>"100000000",
  41710=>"111111001",
  41711=>"000000000",
  41712=>"111111011",
  41713=>"111110110",
  41714=>"100111111",
  41715=>"011000000",
  41716=>"000000000",
  41717=>"001111110",
  41718=>"001001111",
  41719=>"000000111",
  41720=>"111001001",
  41721=>"111110100",
  41722=>"111111111",
  41723=>"000011011",
  41724=>"010110100",
  41725=>"101101001",
  41726=>"000000010",
  41727=>"111010000",
  41728=>"000000000",
  41729=>"110100111",
  41730=>"100011011",
  41731=>"111111110",
  41732=>"011001111",
  41733=>"010011000",
  41734=>"111111000",
  41735=>"111111110",
  41736=>"100111110",
  41737=>"100110110",
  41738=>"111110010",
  41739=>"101011111",
  41740=>"110110111",
  41741=>"001111111",
  41742=>"111011011",
  41743=>"110000000",
  41744=>"111000000",
  41745=>"001001001",
  41746=>"000111010",
  41747=>"000111111",
  41748=>"011101100",
  41749=>"000000111",
  41750=>"001000000",
  41751=>"011011000",
  41752=>"111111000",
  41753=>"100100011",
  41754=>"111100100",
  41755=>"000000110",
  41756=>"111011111",
  41757=>"111111111",
  41758=>"111111111",
  41759=>"000011111",
  41760=>"111111001",
  41761=>"111000000",
  41762=>"111111111",
  41763=>"111111000",
  41764=>"000101101",
  41765=>"111111111",
  41766=>"110010010",
  41767=>"111111001",
  41768=>"011111111",
  41769=>"000000000",
  41770=>"110011100",
  41771=>"111111111",
  41772=>"111111110",
  41773=>"110110110",
  41774=>"111110111",
  41775=>"100000000",
  41776=>"110110100",
  41777=>"000000010",
  41778=>"111111011",
  41779=>"111000000",
  41780=>"111110000",
  41781=>"110110011",
  41782=>"000000010",
  41783=>"111110000",
  41784=>"011001011",
  41785=>"001000100",
  41786=>"111111011",
  41787=>"110000111",
  41788=>"100100111",
  41789=>"110010000",
  41790=>"111110101",
  41791=>"000000000",
  41792=>"111111111",
  41793=>"111111100",
  41794=>"000000000",
  41795=>"000001011",
  41796=>"011111100",
  41797=>"000000010",
  41798=>"100000000",
  41799=>"001001001",
  41800=>"100110110",
  41801=>"111111011",
  41802=>"111111111",
  41803=>"111111010",
  41804=>"111000000",
  41805=>"111101000",
  41806=>"000000000",
  41807=>"010010111",
  41808=>"000010000",
  41809=>"110111101",
  41810=>"111100000",
  41811=>"111111111",
  41812=>"111111111",
  41813=>"001000001",
  41814=>"100000000",
  41815=>"110111000",
  41816=>"000011000",
  41817=>"011000000",
  41818=>"000110000",
  41819=>"111001001",
  41820=>"100000000",
  41821=>"011000000",
  41822=>"111101001",
  41823=>"011111000",
  41824=>"000000101",
  41825=>"000000000",
  41826=>"011011111",
  41827=>"111111111",
  41828=>"000111111",
  41829=>"001001000",
  41830=>"111111111",
  41831=>"001111111",
  41832=>"001101000",
  41833=>"000000000",
  41834=>"011000000",
  41835=>"110111111",
  41836=>"000110000",
  41837=>"100000000",
  41838=>"101100100",
  41839=>"111111111",
  41840=>"101101111",
  41841=>"000000000",
  41842=>"110000000",
  41843=>"110111111",
  41844=>"001111111",
  41845=>"000000000",
  41846=>"100100110",
  41847=>"000000000",
  41848=>"000000000",
  41849=>"000110111",
  41850=>"000000000",
  41851=>"011111110",
  41852=>"111111000",
  41853=>"000011111",
  41854=>"000000000",
  41855=>"100000100",
  41856=>"001000001",
  41857=>"011111111",
  41858=>"011010000",
  41859=>"001000000",
  41860=>"100100111",
  41861=>"000000000",
  41862=>"101001101",
  41863=>"101111111",
  41864=>"000000000",
  41865=>"100000000",
  41866=>"111111111",
  41867=>"001011111",
  41868=>"111110110",
  41869=>"101111111",
  41870=>"100000110",
  41871=>"100100001",
  41872=>"111111111",
  41873=>"111111111",
  41874=>"011011000",
  41875=>"011111111",
  41876=>"000000000",
  41877=>"011001011",
  41878=>"101100101",
  41879=>"000000000",
  41880=>"001001111",
  41881=>"111101001",
  41882=>"001000111",
  41883=>"001000000",
  41884=>"111100111",
  41885=>"110111111",
  41886=>"101101000",
  41887=>"000000111",
  41888=>"001001000",
  41889=>"110110111",
  41890=>"100111111",
  41891=>"000000000",
  41892=>"110110111",
  41893=>"111111000",
  41894=>"000000100",
  41895=>"000000000",
  41896=>"111111111",
  41897=>"010000000",
  41898=>"100100000",
  41899=>"011011010",
  41900=>"000000000",
  41901=>"000000000",
  41902=>"101101111",
  41903=>"000000000",
  41904=>"000000000",
  41905=>"000000000",
  41906=>"100100110",
  41907=>"111011010",
  41908=>"110111011",
  41909=>"111111111",
  41910=>"001001001",
  41911=>"110100000",
  41912=>"110110111",
  41913=>"000100000",
  41914=>"110110000",
  41915=>"010110000",
  41916=>"011000000",
  41917=>"111001001",
  41918=>"100010111",
  41919=>"011001011",
  41920=>"000000010",
  41921=>"001000000",
  41922=>"000000000",
  41923=>"111111111",
  41924=>"111111111",
  41925=>"100000000",
  41926=>"110111111",
  41927=>"110110010",
  41928=>"000000001",
  41929=>"111111111",
  41930=>"111111110",
  41931=>"111111111",
  41932=>"111111101",
  41933=>"010111111",
  41934=>"000110011",
  41935=>"101101111",
  41936=>"111111111",
  41937=>"000010000",
  41938=>"111111111",
  41939=>"100101101",
  41940=>"110110110",
  41941=>"001011001",
  41942=>"000000000",
  41943=>"100010010",
  41944=>"000000100",
  41945=>"000000000",
  41946=>"111000001",
  41947=>"110110110",
  41948=>"111101111",
  41949=>"111100111",
  41950=>"110000000",
  41951=>"111100110",
  41952=>"111111111",
  41953=>"111111001",
  41954=>"100101111",
  41955=>"000000000",
  41956=>"111111111",
  41957=>"000000001",
  41958=>"010111111",
  41959=>"111110110",
  41960=>"000000000",
  41961=>"000000000",
  41962=>"111110000",
  41963=>"000000110",
  41964=>"000000000",
  41965=>"000000000",
  41966=>"000000000",
  41967=>"111111000",
  41968=>"000000000",
  41969=>"111010110",
  41970=>"011011111",
  41971=>"111111111",
  41972=>"001011111",
  41973=>"000000000",
  41974=>"111111111",
  41975=>"001001010",
  41976=>"000111111",
  41977=>"000010010",
  41978=>"001001011",
  41979=>"000000000",
  41980=>"110111111",
  41981=>"111010110",
  41982=>"110111111",
  41983=>"000000000",
  41984=>"111111111",
  41985=>"111001001",
  41986=>"010000000",
  41987=>"000000110",
  41988=>"000000000",
  41989=>"111111001",
  41990=>"111111101",
  41991=>"000000000",
  41992=>"111000000",
  41993=>"000000001",
  41994=>"000000000",
  41995=>"111000000",
  41996=>"110110111",
  41997=>"111111111",
  41998=>"110111110",
  41999=>"000011001",
  42000=>"100111011",
  42001=>"000000000",
  42002=>"111111111",
  42003=>"000000011",
  42004=>"000101111",
  42005=>"000000000",
  42006=>"000000100",
  42007=>"100100100",
  42008=>"100100110",
  42009=>"111111111",
  42010=>"111101101",
  42011=>"111000000",
  42012=>"000000110",
  42013=>"101101101",
  42014=>"011010000",
  42015=>"101101001",
  42016=>"000010110",
  42017=>"000100111",
  42018=>"000111000",
  42019=>"111111010",
  42020=>"100100100",
  42021=>"111000000",
  42022=>"010011111",
  42023=>"001001100",
  42024=>"000000101",
  42025=>"000111101",
  42026=>"000000111",
  42027=>"001111111",
  42028=>"100000111",
  42029=>"011001000",
  42030=>"110111111",
  42031=>"010000011",
  42032=>"111111101",
  42033=>"101000101",
  42034=>"111111011",
  42035=>"000100111",
  42036=>"110111111",
  42037=>"110111111",
  42038=>"111001001",
  42039=>"111111011",
  42040=>"000111000",
  42041=>"011111111",
  42042=>"000101001",
  42043=>"000000100",
  42044=>"101000111",
  42045=>"011000000",
  42046=>"111111110",
  42047=>"000000100",
  42048=>"001011000",
  42049=>"000000110",
  42050=>"100111111",
  42051=>"111111111",
  42052=>"111111111",
  42053=>"100100111",
  42054=>"100000000",
  42055=>"100000000",
  42056=>"001111001",
  42057=>"000000101",
  42058=>"001101111",
  42059=>"001000000",
  42060=>"111110000",
  42061=>"101000000",
  42062=>"111111110",
  42063=>"100001001",
  42064=>"000001001",
  42065=>"110010000",
  42066=>"000000001",
  42067=>"110111110",
  42068=>"100000000",
  42069=>"000000000",
  42070=>"001000100",
  42071=>"000000001",
  42072=>"110010000",
  42073=>"111100000",
  42074=>"011011001",
  42075=>"000011111",
  42076=>"000000000",
  42077=>"000000101",
  42078=>"011001000",
  42079=>"000110110",
  42080=>"110010000",
  42081=>"111111000",
  42082=>"100101111",
  42083=>"111011001",
  42084=>"001000000",
  42085=>"000000000",
  42086=>"000000000",
  42087=>"111111111",
  42088=>"110100100",
  42089=>"101111111",
  42090=>"011000000",
  42091=>"110100111",
  42092=>"111011000",
  42093=>"111111111",
  42094=>"000000010",
  42095=>"110110111",
  42096=>"111011001",
  42097=>"101101101",
  42098=>"011011011",
  42099=>"000000000",
  42100=>"000000000",
  42101=>"110111000",
  42102=>"000111111",
  42103=>"111111010",
  42104=>"000001000",
  42105=>"111111111",
  42106=>"000000000",
  42107=>"111111111",
  42108=>"110110111",
  42109=>"001000000",
  42110=>"111111111",
  42111=>"001111011",
  42112=>"001001111",
  42113=>"000000000",
  42114=>"000100000",
  42115=>"111111111",
  42116=>"000000101",
  42117=>"101000100",
  42118=>"001000000",
  42119=>"111110000",
  42120=>"111000110",
  42121=>"001001111",
  42122=>"000000111",
  42123=>"111111111",
  42124=>"001100100",
  42125=>"000000000",
  42126=>"011111111",
  42127=>"111111111",
  42128=>"111101111",
  42129=>"001001001",
  42130=>"111111111",
  42131=>"011000000",
  42132=>"000000000",
  42133=>"110100110",
  42134=>"000000101",
  42135=>"000000000",
  42136=>"011001000",
  42137=>"111111111",
  42138=>"111111111",
  42139=>"011011011",
  42140=>"111111111",
  42141=>"101001000",
  42142=>"111111011",
  42143=>"000000000",
  42144=>"011011111",
  42145=>"011001011",
  42146=>"000000101",
  42147=>"100111110",
  42148=>"110111000",
  42149=>"010010000",
  42150=>"111001001",
  42151=>"011011011",
  42152=>"111101100",
  42153=>"111000000",
  42154=>"000001111",
  42155=>"111111000",
  42156=>"010110111",
  42157=>"110110110",
  42158=>"000000100",
  42159=>"101001000",
  42160=>"111011000",
  42161=>"000000110",
  42162=>"111111011",
  42163=>"000000000",
  42164=>"110010011",
  42165=>"001111111",
  42166=>"111100100",
  42167=>"101001000",
  42168=>"000000000",
  42169=>"011001000",
  42170=>"000000000",
  42171=>"011011111",
  42172=>"100100100",
  42173=>"110111111",
  42174=>"111111111",
  42175=>"000000000",
  42176=>"010000000",
  42177=>"000000000",
  42178=>"001111111",
  42179=>"100111111",
  42180=>"000000000",
  42181=>"000100000",
  42182=>"000000000",
  42183=>"000011011",
  42184=>"001001000",
  42185=>"000000000",
  42186=>"111101100",
  42187=>"000000000",
  42188=>"101101111",
  42189=>"111011000",
  42190=>"100111111",
  42191=>"000110001",
  42192=>"000000000",
  42193=>"101101000",
  42194=>"110100001",
  42195=>"110111001",
  42196=>"100110110",
  42197=>"000000000",
  42198=>"000000000",
  42199=>"101101111",
  42200=>"000000000",
  42201=>"010110010",
  42202=>"111111111",
  42203=>"000000111",
  42204=>"000100000",
  42205=>"000000000",
  42206=>"111111111",
  42207=>"000001111",
  42208=>"000000000",
  42209=>"011001001",
  42210=>"000000111",
  42211=>"011001001",
  42212=>"000100110",
  42213=>"111111111",
  42214=>"111111111",
  42215=>"101101111",
  42216=>"000000000",
  42217=>"111001000",
  42218=>"111111101",
  42219=>"100100101",
  42220=>"000000000",
  42221=>"000111111",
  42222=>"011000001",
  42223=>"111000000",
  42224=>"111111110",
  42225=>"010000000",
  42226=>"100000101",
  42227=>"000000100",
  42228=>"111100101",
  42229=>"001100111",
  42230=>"000000001",
  42231=>"100000100",
  42232=>"000000000",
  42233=>"000000000",
  42234=>"111111111",
  42235=>"111101000",
  42236=>"011111111",
  42237=>"100111111",
  42238=>"111111111",
  42239=>"010000000",
  42240=>"001000000",
  42241=>"000000001",
  42242=>"110110000",
  42243=>"000011011",
  42244=>"110111010",
  42245=>"011011011",
  42246=>"110110100",
  42247=>"000110000",
  42248=>"000000000",
  42249=>"011111011",
  42250=>"001101101",
  42251=>"110111010",
  42252=>"111001001",
  42253=>"000000000",
  42254=>"001000100",
  42255=>"011010110",
  42256=>"000100000",
  42257=>"001011111",
  42258=>"111001000",
  42259=>"000001101",
  42260=>"111111111",
  42261=>"100111111",
  42262=>"000001101",
  42263=>"000001000",
  42264=>"011001000",
  42265=>"000000111",
  42266=>"000010010",
  42267=>"011011000",
  42268=>"110110100",
  42269=>"000000001",
  42270=>"000000000",
  42271=>"110100101",
  42272=>"011010110",
  42273=>"000100101",
  42274=>"111100000",
  42275=>"111111101",
  42276=>"000000100",
  42277=>"111111111",
  42278=>"111111111",
  42279=>"111111101",
  42280=>"111111100",
  42281=>"111111111",
  42282=>"001000001",
  42283=>"110000111",
  42284=>"000000000",
  42285=>"011101000",
  42286=>"000000000",
  42287=>"111111011",
  42288=>"001000000",
  42289=>"000000100",
  42290=>"011000000",
  42291=>"111100000",
  42292=>"000000000",
  42293=>"100111111",
  42294=>"011111111",
  42295=>"000000000",
  42296=>"011001011",
  42297=>"000000101",
  42298=>"000000000",
  42299=>"000000100",
  42300=>"000000111",
  42301=>"001001000",
  42302=>"000000011",
  42303=>"000000000",
  42304=>"011011001",
  42305=>"000001000",
  42306=>"110110010",
  42307=>"000001001",
  42308=>"111110010",
  42309=>"111111111",
  42310=>"000111111",
  42311=>"111111111",
  42312=>"000000000",
  42313=>"000000000",
  42314=>"011111111",
  42315=>"111111111",
  42316=>"001000000",
  42317=>"111001001",
  42318=>"111111111",
  42319=>"110110100",
  42320=>"110111110",
  42321=>"100000101",
  42322=>"000111000",
  42323=>"000001111",
  42324=>"100000000",
  42325=>"011001011",
  42326=>"111011111",
  42327=>"000000000",
  42328=>"000000000",
  42329=>"111101101",
  42330=>"011011000",
  42331=>"110110110",
  42332=>"000000000",
  42333=>"000000010",
  42334=>"111010010",
  42335=>"111111111",
  42336=>"000011001",
  42337=>"111011001",
  42338=>"000000000",
  42339=>"100100000",
  42340=>"100100000",
  42341=>"111011111",
  42342=>"111111111",
  42343=>"001001111",
  42344=>"001011111",
  42345=>"110111001",
  42346=>"000001001",
  42347=>"010011111",
  42348=>"010000101",
  42349=>"000100111",
  42350=>"111111000",
  42351=>"011111011",
  42352=>"000000000",
  42353=>"011111110",
  42354=>"000000000",
  42355=>"100100000",
  42356=>"000000000",
  42357=>"000000000",
  42358=>"000000011",
  42359=>"000000000",
  42360=>"000000000",
  42361=>"111111111",
  42362=>"001000100",
  42363=>"000000000",
  42364=>"000000000",
  42365=>"111111111",
  42366=>"000010110",
  42367=>"111100111",
  42368=>"011001111",
  42369=>"111110111",
  42370=>"000001001",
  42371=>"011001000",
  42372=>"111111101",
  42373=>"100100111",
  42374=>"000110100",
  42375=>"111100111",
  42376=>"111011011",
  42377=>"011001000",
  42378=>"111111111",
  42379=>"000000100",
  42380=>"000100111",
  42381=>"111111010",
  42382=>"011111011",
  42383=>"000000000",
  42384=>"000011011",
  42385=>"111111111",
  42386=>"101001001",
  42387=>"010000001",
  42388=>"111101000",
  42389=>"000010010",
  42390=>"101000101",
  42391=>"000111111",
  42392=>"111111111",
  42393=>"110100010",
  42394=>"000000000",
  42395=>"000000110",
  42396=>"111111101",
  42397=>"001000000",
  42398=>"011011011",
  42399=>"111111111",
  42400=>"100100100",
  42401=>"000000100",
  42402=>"111011000",
  42403=>"111000011",
  42404=>"011111111",
  42405=>"000000000",
  42406=>"101000000",
  42407=>"111111110",
  42408=>"000000000",
  42409=>"100111111",
  42410=>"111111111",
  42411=>"100000011",
  42412=>"101101111",
  42413=>"111001000",
  42414=>"100111111",
  42415=>"111110111",
  42416=>"111111110",
  42417=>"111111111",
  42418=>"111111011",
  42419=>"001000000",
  42420=>"101001011",
  42421=>"001010111",
  42422=>"000000000",
  42423=>"111111111",
  42424=>"111111110",
  42425=>"100001000",
  42426=>"000000000",
  42427=>"111111111",
  42428=>"000000010",
  42429=>"111110110",
  42430=>"011100000",
  42431=>"001011010",
  42432=>"011011000",
  42433=>"111111111",
  42434=>"000000000",
  42435=>"111000001",
  42436=>"111111001",
  42437=>"000001001",
  42438=>"000001000",
  42439=>"111111111",
  42440=>"011000000",
  42441=>"110111111",
  42442=>"000000000",
  42443=>"111000001",
  42444=>"000000000",
  42445=>"000000101",
  42446=>"000001111",
  42447=>"111111010",
  42448=>"011011001",
  42449=>"111100000",
  42450=>"110111110",
  42451=>"000000111",
  42452=>"111111111",
  42453=>"101001001",
  42454=>"111111100",
  42455=>"011011010",
  42456=>"111111111",
  42457=>"100111110",
  42458=>"000000001",
  42459=>"111111111",
  42460=>"100110100",
  42461=>"110000000",
  42462=>"001000000",
  42463=>"000111111",
  42464=>"110011011",
  42465=>"010111000",
  42466=>"111111101",
  42467=>"101000000",
  42468=>"111111111",
  42469=>"000001001",
  42470=>"001011100",
  42471=>"000101100",
  42472=>"001000000",
  42473=>"111000000",
  42474=>"011000100",
  42475=>"111111111",
  42476=>"000000000",
  42477=>"010111011",
  42478=>"000110110",
  42479=>"111100101",
  42480=>"110111011",
  42481=>"010000110",
  42482=>"000100100",
  42483=>"000011001",
  42484=>"111111110",
  42485=>"110001011",
  42486=>"111111011",
  42487=>"111111001",
  42488=>"011010111",
  42489=>"111011001",
  42490=>"000000001",
  42491=>"111111111",
  42492=>"011011000",
  42493=>"001011001",
  42494=>"111100100",
  42495=>"001111111",
  42496=>"111111111",
  42497=>"000001111",
  42498=>"001001001",
  42499=>"000000000",
  42500=>"000011011",
  42501=>"110110111",
  42502=>"011000111",
  42503=>"111111111",
  42504=>"111111110",
  42505=>"000110001",
  42506=>"111010000",
  42507=>"111011011",
  42508=>"100110110",
  42509=>"000000110",
  42510=>"101111010",
  42511=>"000010010",
  42512=>"111010010",
  42513=>"000000000",
  42514=>"000000000",
  42515=>"000111111",
  42516=>"010000000",
  42517=>"111000000",
  42518=>"010000000",
  42519=>"010000000",
  42520=>"010011111",
  42521=>"011101100",
  42522=>"110000101",
  42523=>"000000010",
  42524=>"111101111",
  42525=>"000000100",
  42526=>"101111110",
  42527=>"000101001",
  42528=>"000010011",
  42529=>"111111100",
  42530=>"111111110",
  42531=>"001001110",
  42532=>"110000000",
  42533=>"010010011",
  42534=>"001111110",
  42535=>"000000000",
  42536=>"000000011",
  42537=>"000000000",
  42538=>"000000111",
  42539=>"111111111",
  42540=>"111000000",
  42541=>"111000000",
  42542=>"110100111",
  42543=>"001101111",
  42544=>"000000000",
  42545=>"011011101",
  42546=>"010010011",
  42547=>"111111111",
  42548=>"000000110",
  42549=>"010001001",
  42550=>"111000000",
  42551=>"000001011",
  42552=>"100000000",
  42553=>"000000000",
  42554=>"100000000",
  42555=>"000000000",
  42556=>"000000000",
  42557=>"001001011",
  42558=>"111111111",
  42559=>"111100110",
  42560=>"110000001",
  42561=>"100000101",
  42562=>"111111111",
  42563=>"001000010",
  42564=>"001001111",
  42565=>"011011111",
  42566=>"110111111",
  42567=>"110000000",
  42568=>"111111111",
  42569=>"111111111",
  42570=>"111111111",
  42571=>"111001001",
  42572=>"000000011",
  42573=>"001000000",
  42574=>"000000001",
  42575=>"000000000",
  42576=>"111111000",
  42577=>"111111000",
  42578=>"111111100",
  42579=>"101101111",
  42580=>"111111111",
  42581=>"000000000",
  42582=>"111000000",
  42583=>"100101111",
  42584=>"000000000",
  42585=>"111000000",
  42586=>"111110111",
  42587=>"111111111",
  42588=>"010000110",
  42589=>"111101011",
  42590=>"111111110",
  42591=>"010000000",
  42592=>"111000000",
  42593=>"000111010",
  42594=>"111011011",
  42595=>"000000011",
  42596=>"000000000",
  42597=>"110110111",
  42598=>"000000100",
  42599=>"111111111",
  42600=>"111111111",
  42601=>"111111111",
  42602=>"111111000",
  42603=>"111111111",
  42604=>"100110111",
  42605=>"001000001",
  42606=>"111111110",
  42607=>"111111111",
  42608=>"000000001",
  42609=>"000000000",
  42610=>"100100100",
  42611=>"111111000",
  42612=>"011111111",
  42613=>"000110100",
  42614=>"000000000",
  42615=>"000000000",
  42616=>"000001111",
  42617=>"000000011",
  42618=>"000000000",
  42619=>"011010000",
  42620=>"111111011",
  42621=>"111111100",
  42622=>"111111111",
  42623=>"111000000",
  42624=>"000000001",
  42625=>"001001001",
  42626=>"000000000",
  42627=>"110111111",
  42628=>"110110000",
  42629=>"111101111",
  42630=>"001111111",
  42631=>"011000000",
  42632=>"001000000",
  42633=>"111111111",
  42634=>"000000000",
  42635=>"111000000",
  42636=>"111111000",
  42637=>"110100110",
  42638=>"000000000",
  42639=>"000101111",
  42640=>"001001111",
  42641=>"111111111",
  42642=>"010000000",
  42643=>"000011010",
  42644=>"001001111",
  42645=>"110111111",
  42646=>"111111111",
  42647=>"111111000",
  42648=>"000000110",
  42649=>"111111111",
  42650=>"111111110",
  42651=>"000000010",
  42652=>"111000000",
  42653=>"110000001",
  42654=>"111100000",
  42655=>"000000010",
  42656=>"101111111",
  42657=>"000000000",
  42658=>"111111100",
  42659=>"000000000",
  42660=>"000000000",
  42661=>"001001011",
  42662=>"111111111",
  42663=>"010011000",
  42664=>"111111110",
  42665=>"000110111",
  42666=>"000000111",
  42667=>"000000101",
  42668=>"000000000",
  42669=>"111111111",
  42670=>"011111111",
  42671=>"111111110",
  42672=>"111111000",
  42673=>"000000000",
  42674=>"111110110",
  42675=>"111000100",
  42676=>"111111111",
  42677=>"111000000",
  42678=>"000001111",
  42679=>"101000001",
  42680=>"111111111",
  42681=>"111111111",
  42682=>"111001000",
  42683=>"111111111",
  42684=>"001001111",
  42685=>"000000000",
  42686=>"111001111",
  42687=>"100000000",
  42688=>"000000000",
  42689=>"000100100",
  42690=>"111100000",
  42691=>"000000000",
  42692=>"000000000",
  42693=>"000000111",
  42694=>"000000000",
  42695=>"000000101",
  42696=>"111111110",
  42697=>"001111111",
  42698=>"001001000",
  42699=>"111101001",
  42700=>"000000110",
  42701=>"000000110",
  42702=>"000000000",
  42703=>"110000001",
  42704=>"010111111",
  42705=>"011000000",
  42706=>"000000000",
  42707=>"111111111",
  42708=>"000000111",
  42709=>"010010000",
  42710=>"111111111",
  42711=>"000000001",
  42712=>"110000001",
  42713=>"000100000",
  42714=>"111011111",
  42715=>"000000011",
  42716=>"100000001",
  42717=>"000010000",
  42718=>"000111001",
  42719=>"111110110",
  42720=>"111000010",
  42721=>"110111111",
  42722=>"000000100",
  42723=>"111000000",
  42724=>"111111001",
  42725=>"110110111",
  42726=>"111111110",
  42727=>"011111000",
  42728=>"000000000",
  42729=>"000000000",
  42730=>"100100000",
  42731=>"000100111",
  42732=>"000000000",
  42733=>"111111111",
  42734=>"001000000",
  42735=>"111101101",
  42736=>"001000000",
  42737=>"000010010",
  42738=>"000001111",
  42739=>"111001111",
  42740=>"111011000",
  42741=>"000000000",
  42742=>"001011000",
  42743=>"110110111",
  42744=>"111111111",
  42745=>"000101111",
  42746=>"111000000",
  42747=>"010111111",
  42748=>"000011011",
  42749=>"001001001",
  42750=>"001001111",
  42751=>"111111110",
  42752=>"000000000",
  42753=>"000110111",
  42754=>"100000000",
  42755=>"000000110",
  42756=>"111111111",
  42757=>"001000000",
  42758=>"111111111",
  42759=>"001000110",
  42760=>"001000101",
  42761=>"000001001",
  42762=>"111111010",
  42763=>"110110110",
  42764=>"001000101",
  42765=>"111110111",
  42766=>"111000000",
  42767=>"000000000",
  42768=>"000000011",
  42769=>"111000000",
  42770=>"000001000",
  42771=>"110110110",
  42772=>"000000001",
  42773=>"111011011",
  42774=>"001111111",
  42775=>"111111111",
  42776=>"100110110",
  42777=>"111000000",
  42778=>"111111010",
  42779=>"001011001",
  42780=>"111111111",
  42781=>"000000000",
  42782=>"000000010",
  42783=>"000000001",
  42784=>"110011111",
  42785=>"110110111",
  42786=>"111110010",
  42787=>"000000000",
  42788=>"011001000",
  42789=>"010000000",
  42790=>"100100100",
  42791=>"111110110",
  42792=>"111110000",
  42793=>"111101111",
  42794=>"110100000",
  42795=>"111111111",
  42796=>"111111111",
  42797=>"101100010",
  42798=>"000000000",
  42799=>"000000000",
  42800=>"001001111",
  42801=>"001111111",
  42802=>"000111111",
  42803=>"000011000",
  42804=>"000011111",
  42805=>"111110100",
  42806=>"101101111",
  42807=>"000000000",
  42808=>"000000111",
  42809=>"000000000",
  42810=>"110110010",
  42811=>"111111111",
  42812=>"000000100",
  42813=>"100000000",
  42814=>"110111100",
  42815=>"111111111",
  42816=>"000100110",
  42817=>"101001101",
  42818=>"010010110",
  42819=>"111111000",
  42820=>"000100111",
  42821=>"111111111",
  42822=>"000000001",
  42823=>"111111111",
  42824=>"001010010",
  42825=>"111011011",
  42826=>"111001101",
  42827=>"101101111",
  42828=>"000000000",
  42829=>"110010000",
  42830=>"000000000",
  42831=>"001001011",
  42832=>"110111111",
  42833=>"000010110",
  42834=>"000001111",
  42835=>"000001001",
  42836=>"000000010",
  42837=>"111111111",
  42838=>"111111111",
  42839=>"000000110",
  42840=>"100111111",
  42841=>"000000000",
  42842=>"000010110",
  42843=>"111110110",
  42844=>"011000011",
  42845=>"000000000",
  42846=>"111000000",
  42847=>"110000000",
  42848=>"111100101",
  42849=>"000000000",
  42850=>"111100100",
  42851=>"000000111",
  42852=>"000000110",
  42853=>"000000000",
  42854=>"000110111",
  42855=>"100100000",
  42856=>"111011111",
  42857=>"000000110",
  42858=>"111000100",
  42859=>"100111111",
  42860=>"101111111",
  42861=>"111010011",
  42862=>"011010000",
  42863=>"000010110",
  42864=>"001111111",
  42865=>"000000000",
  42866=>"000111010",
  42867=>"000011000",
  42868=>"111111111",
  42869=>"011011001",
  42870=>"000000010",
  42871=>"000000011",
  42872=>"111100100",
  42873=>"000010000",
  42874=>"000010000",
  42875=>"011011111",
  42876=>"110010000",
  42877=>"111111010",
  42878=>"001111111",
  42879=>"000000000",
  42880=>"000000000",
  42881=>"111101101",
  42882=>"010100110",
  42883=>"000111111",
  42884=>"001111111",
  42885=>"001001011",
  42886=>"000000001",
  42887=>"111011001",
  42888=>"000000000",
  42889=>"111101001",
  42890=>"000110110",
  42891=>"111111111",
  42892=>"111111111",
  42893=>"000000001",
  42894=>"000011000",
  42895=>"000000001",
  42896=>"000000000",
  42897=>"111111011",
  42898=>"111111001",
  42899=>"010110111",
  42900=>"001000000",
  42901=>"000000000",
  42902=>"111110111",
  42903=>"111111111",
  42904=>"111000000",
  42905=>"110110110",
  42906=>"111110110",
  42907=>"001111111",
  42908=>"111101111",
  42909=>"111111100",
  42910=>"001001001",
  42911=>"000000000",
  42912=>"010011111",
  42913=>"111111111",
  42914=>"110010010",
  42915=>"111011011",
  42916=>"111100000",
  42917=>"000000110",
  42918=>"000110111",
  42919=>"111001001",
  42920=>"111111111",
  42921=>"111101111",
  42922=>"111111111",
  42923=>"001001111",
  42924=>"011001001",
  42925=>"000100000",
  42926=>"110110000",
  42927=>"000000000",
  42928=>"000000000",
  42929=>"010010000",
  42930=>"000000000",
  42931=>"101000011",
  42932=>"110000000",
  42933=>"000000000",
  42934=>"000110110",
  42935=>"000100111",
  42936=>"111010110",
  42937=>"010011111",
  42938=>"000000000",
  42939=>"111111101",
  42940=>"001000000",
  42941=>"100100100",
  42942=>"011110110",
  42943=>"111000011",
  42944=>"101111111",
  42945=>"111011000",
  42946=>"101000000",
  42947=>"110000010",
  42948=>"101000000",
  42949=>"001001000",
  42950=>"110100000",
  42951=>"111111111",
  42952=>"111101111",
  42953=>"001011111",
  42954=>"111100100",
  42955=>"000000000",
  42956=>"000110111",
  42957=>"000000110",
  42958=>"110110100",
  42959=>"011000000",
  42960=>"000000000",
  42961=>"111111111",
  42962=>"000100000",
  42963=>"001000000",
  42964=>"111110110",
  42965=>"100000000",
  42966=>"000000000",
  42967=>"011001001",
  42968=>"000000000",
  42969=>"100001001",
  42970=>"001000000",
  42971=>"011101111",
  42972=>"000010011",
  42973=>"111111111",
  42974=>"000000111",
  42975=>"000100110",
  42976=>"011011010",
  42977=>"001000001",
  42978=>"111111100",
  42979=>"000000000",
  42980=>"111001111",
  42981=>"010111110",
  42982=>"001000000",
  42983=>"011011111",
  42984=>"110111000",
  42985=>"000000111",
  42986=>"000000000",
  42987=>"000110111",
  42988=>"111111101",
  42989=>"111110111",
  42990=>"101101101",
  42991=>"011111111",
  42992=>"111001000",
  42993=>"010000000",
  42994=>"111111000",
  42995=>"111110111",
  42996=>"000000000",
  42997=>"101101001",
  42998=>"111011111",
  42999=>"001101101",
  43000=>"000000000",
  43001=>"100000000",
  43002=>"011010000",
  43003=>"111111001",
  43004=>"000111111",
  43005=>"001001000",
  43006=>"111111111",
  43007=>"000000000",
  43008=>"001000000",
  43009=>"000000000",
  43010=>"000000111",
  43011=>"101101001",
  43012=>"000000111",
  43013=>"000001111",
  43014=>"011000111",
  43015=>"100000000",
  43016=>"111111000",
  43017=>"000000001",
  43018=>"000010000",
  43019=>"100111000",
  43020=>"001111010",
  43021=>"001001111",
  43022=>"000000111",
  43023=>"001001101",
  43024=>"111000000",
  43025=>"000111111",
  43026=>"101001001",
  43027=>"000000100",
  43028=>"001000000",
  43029=>"111000000",
  43030=>"111111111",
  43031=>"111001011",
  43032=>"111010000",
  43033=>"001011011",
  43034=>"000000000",
  43035=>"100000000",
  43036=>"100110000",
  43037=>"100100100",
  43038=>"001001111",
  43039=>"000000000",
  43040=>"000000011",
  43041=>"000000111",
  43042=>"001111111",
  43043=>"111000000",
  43044=>"000000110",
  43045=>"111001001",
  43046=>"001000001",
  43047=>"111111111",
  43048=>"111000100",
  43049=>"111111111",
  43050=>"001000111",
  43051=>"000100101",
  43052=>"111111111",
  43053=>"111101000",
  43054=>"000000011",
  43055=>"001000110",
  43056=>"111111111",
  43057=>"010010000",
  43058=>"000000001",
  43059=>"000000011",
  43060=>"000111111",
  43061=>"111011011",
  43062=>"111111101",
  43063=>"001111000",
  43064=>"000000001",
  43065=>"000111111",
  43066=>"111111111",
  43067=>"111111111",
  43068=>"111000110",
  43069=>"100111110",
  43070=>"000001001",
  43071=>"110010111",
  43072=>"111111011",
  43073=>"000000000",
  43074=>"001000000",
  43075=>"000000000",
  43076=>"111001000",
  43077=>"010011011",
  43078=>"010000000",
  43079=>"111100000",
  43080=>"110111110",
  43081=>"100000111",
  43082=>"000000000",
  43083=>"001001111",
  43084=>"111111101",
  43085=>"111111111",
  43086=>"000000000",
  43087=>"111111111",
  43088=>"111111111",
  43089=>"111111110",
  43090=>"000000000",
  43091=>"011000000",
  43092=>"000000011",
  43093=>"000111111",
  43094=>"100000000",
  43095=>"111111111",
  43096=>"000110111",
  43097=>"111111111",
  43098=>"111101011",
  43099=>"100100110",
  43100=>"000000000",
  43101=>"000100001",
  43102=>"101001000",
  43103=>"111111000",
  43104=>"000001000",
  43105=>"111111011",
  43106=>"000000000",
  43107=>"011111000",
  43108=>"000111000",
  43109=>"000010111",
  43110=>"111111111",
  43111=>"110101101",
  43112=>"111101010",
  43113=>"111111000",
  43114=>"000000100",
  43115=>"000111001",
  43116=>"000100000",
  43117=>"000111111",
  43118=>"111111000",
  43119=>"000000000",
  43120=>"000111111",
  43121=>"000111111",
  43122=>"000000000",
  43123=>"000001111",
  43124=>"011011010",
  43125=>"000111111",
  43126=>"000000000",
  43127=>"000000000",
  43128=>"000000000",
  43129=>"111110110",
  43130=>"011000000",
  43131=>"000000000",
  43132=>"111100100",
  43133=>"000000000",
  43134=>"000000000",
  43135=>"011011111",
  43136=>"111111111",
  43137=>"100000000",
  43138=>"111000000",
  43139=>"001000000",
  43140=>"110010111",
  43141=>"000000111",
  43142=>"000101000",
  43143=>"111000100",
  43144=>"111101111",
  43145=>"111100000",
  43146=>"100111000",
  43147=>"111010000",
  43148=>"000000000",
  43149=>"001001111",
  43150=>"000011000",
  43151=>"101111111",
  43152=>"000000000",
  43153=>"111111111",
  43154=>"000000000",
  43155=>"000111111",
  43156=>"011001000",
  43157=>"111111011",
  43158=>"111101001",
  43159=>"111111111",
  43160=>"000000001",
  43161=>"111101100",
  43162=>"001000000",
  43163=>"111100000",
  43164=>"111111111",
  43165=>"000110110",
  43166=>"000000111",
  43167=>"001000000",
  43168=>"100000111",
  43169=>"111000000",
  43170=>"111111111",
  43171=>"100111111",
  43172=>"000000000",
  43173=>"000000000",
  43174=>"101111110",
  43175=>"110111110",
  43176=>"111111111",
  43177=>"000000000",
  43178=>"000000111",
  43179=>"000100111",
  43180=>"000000111",
  43181=>"111111110",
  43182=>"000000000",
  43183=>"110000000",
  43184=>"001000000",
  43185=>"100001000",
  43186=>"111111111",
  43187=>"111001000",
  43188=>"000111111",
  43189=>"101111111",
  43190=>"001000111",
  43191=>"110111111",
  43192=>"101111111",
  43193=>"111111111",
  43194=>"100100001",
  43195=>"000000000",
  43196=>"000000000",
  43197=>"000011011",
  43198=>"000001001",
  43199=>"000000000",
  43200=>"111111111",
  43201=>"000101111",
  43202=>"000011011",
  43203=>"000110000",
  43204=>"000001111",
  43205=>"001111111",
  43206=>"000000101",
  43207=>"000110110",
  43208=>"111110111",
  43209=>"000110000",
  43210=>"100000100",
  43211=>"101101111",
  43212=>"111000100",
  43213=>"000000001",
  43214=>"100100111",
  43215=>"100100000",
  43216=>"000000111",
  43217=>"111110110",
  43218=>"000100011",
  43219=>"001111111",
  43220=>"111000101",
  43221=>"110111010",
  43222=>"100111001",
  43223=>"000110111",
  43224=>"000000100",
  43225=>"000000000",
  43226=>"111111111",
  43227=>"111100101",
  43228=>"111111111",
  43229=>"111110000",
  43230=>"000100111",
  43231=>"101000000",
  43232=>"110000000",
  43233=>"000111010",
  43234=>"100101001",
  43235=>"111111111",
  43236=>"111000000",
  43237=>"000000111",
  43238=>"111001001",
  43239=>"000000111",
  43240=>"000010000",
  43241=>"000000000",
  43242=>"001000100",
  43243=>"000000010",
  43244=>"111111000",
  43245=>"000000110",
  43246=>"000000000",
  43247=>"111001111",
  43248=>"000000000",
  43249=>"110100000",
  43250=>"000010000",
  43251=>"111111001",
  43252=>"000000111",
  43253=>"111111011",
  43254=>"000000000",
  43255=>"110000000",
  43256=>"011111111",
  43257=>"000000000",
  43258=>"000000000",
  43259=>"000001001",
  43260=>"000100100",
  43261=>"110110000",
  43262=>"110100100",
  43263=>"111101111",
  43264=>"000000000",
  43265=>"000000110",
  43266=>"000000000",
  43267=>"000000000",
  43268=>"000000000",
  43269=>"001000001",
  43270=>"000001111",
  43271=>"000000100",
  43272=>"000000000",
  43273=>"000010000",
  43274=>"111000100",
  43275=>"111111000",
  43276=>"100000101",
  43277=>"110100111",
  43278=>"111111111",
  43279=>"000000000",
  43280=>"101000000",
  43281=>"000000000",
  43282=>"111011000",
  43283=>"000000000",
  43284=>"000000000",
  43285=>"000111111",
  43286=>"111111111",
  43287=>"111111100",
  43288=>"000000000",
  43289=>"000100111",
  43290=>"000100000",
  43291=>"001011111",
  43292=>"011111111",
  43293=>"000000000",
  43294=>"001000000",
  43295=>"101000000",
  43296=>"111011000",
  43297=>"111111111",
  43298=>"111111000",
  43299=>"111000001",
  43300=>"111000000",
  43301=>"000000000",
  43302=>"100100110",
  43303=>"111011000",
  43304=>"000000000",
  43305=>"000000000",
  43306=>"111111010",
  43307=>"100101000",
  43308=>"111110000",
  43309=>"011111010",
  43310=>"111110111",
  43311=>"000000100",
  43312=>"110111000",
  43313=>"111111111",
  43314=>"111000000",
  43315=>"000000000",
  43316=>"110000001",
  43317=>"111000000",
  43318=>"100100111",
  43319=>"111000000",
  43320=>"001000000",
  43321=>"111111101",
  43322=>"000000000",
  43323=>"000100111",
  43324=>"001001111",
  43325=>"000000000",
  43326=>"111111011",
  43327=>"101000000",
  43328=>"011011011",
  43329=>"000000000",
  43330=>"010111111",
  43331=>"100100000",
  43332=>"111000000",
  43333=>"101111111",
  43334=>"100111110",
  43335=>"011000000",
  43336=>"000000001",
  43337=>"111111000",
  43338=>"001111010",
  43339=>"000100110",
  43340=>"000111111",
  43341=>"110000111",
  43342=>"001000000",
  43343=>"000111011",
  43344=>"000000111",
  43345=>"111111111",
  43346=>"000111111",
  43347=>"000000000",
  43348=>"000000000",
  43349=>"011001011",
  43350=>"110111111",
  43351=>"100000110",
  43352=>"101011000",
  43353=>"111111110",
  43354=>"110110000",
  43355=>"100000110",
  43356=>"111000000",
  43357=>"001011111",
  43358=>"110110101",
  43359=>"011011010",
  43360=>"110011001",
  43361=>"001011111",
  43362=>"000111111",
  43363=>"111111111",
  43364=>"011000000",
  43365=>"000000000",
  43366=>"111111111",
  43367=>"111111110",
  43368=>"001000000",
  43369=>"000111000",
  43370=>"000011011",
  43371=>"001110010",
  43372=>"111111111",
  43373=>"111111111",
  43374=>"111111000",
  43375=>"110000000",
  43376=>"011011000",
  43377=>"111111111",
  43378=>"111111111",
  43379=>"000000000",
  43380=>"000000000",
  43381=>"000011000",
  43382=>"010111110",
  43383=>"011000000",
  43384=>"000111111",
  43385=>"000000000",
  43386=>"111111000",
  43387=>"100000001",
  43388=>"000000111",
  43389=>"001001111",
  43390=>"100000000",
  43391=>"000000100",
  43392=>"000110111",
  43393=>"111111111",
  43394=>"011001000",
  43395=>"000000110",
  43396=>"111111111",
  43397=>"110000000",
  43398=>"100000110",
  43399=>"001011000",
  43400=>"001000001",
  43401=>"000000010",
  43402=>"000111111",
  43403=>"111111000",
  43404=>"111100000",
  43405=>"000111110",
  43406=>"111111111",
  43407=>"111111000",
  43408=>"000000000",
  43409=>"111111101",
  43410=>"111111111",
  43411=>"000110000",
  43412=>"111011001",
  43413=>"010111000",
  43414=>"010110110",
  43415=>"111010000",
  43416=>"000011111",
  43417=>"111101000",
  43418=>"111111111",
  43419=>"000000000",
  43420=>"101000100",
  43421=>"000000110",
  43422=>"000000101",
  43423=>"000000111",
  43424=>"111101111",
  43425=>"111111110",
  43426=>"110001000",
  43427=>"111001101",
  43428=>"000111111",
  43429=>"111111100",
  43430=>"110000000",
  43431=>"111111001",
  43432=>"000000110",
  43433=>"001001100",
  43434=>"100000000",
  43435=>"100001000",
  43436=>"000111010",
  43437=>"111001000",
  43438=>"111111111",
  43439=>"111000000",
  43440=>"110100000",
  43441=>"110000000",
  43442=>"001101111",
  43443=>"110000000",
  43444=>"100111111",
  43445=>"000000000",
  43446=>"000000000",
  43447=>"000000100",
  43448=>"111110000",
  43449=>"000001001",
  43450=>"000100000",
  43451=>"111111111",
  43452=>"011000000",
  43453=>"111000001",
  43454=>"101000000",
  43455=>"100001111",
  43456=>"000000110",
  43457=>"000000000",
  43458=>"111110000",
  43459=>"000000000",
  43460=>"100111111",
  43461=>"100110111",
  43462=>"000000000",
  43463=>"111111111",
  43464=>"000000001",
  43465=>"000000000",
  43466=>"000000000",
  43467=>"000000000",
  43468=>"111111000",
  43469=>"111111011",
  43470=>"111011000",
  43471=>"111000000",
  43472=>"000000001",
  43473=>"000000000",
  43474=>"000000000",
  43475=>"000000000",
  43476=>"000000000",
  43477=>"111111111",
  43478=>"111111001",
  43479=>"110111110",
  43480=>"111111111",
  43481=>"111111111",
  43482=>"111111000",
  43483=>"000010000",
  43484=>"000000000",
  43485=>"101101000",
  43486=>"000011001",
  43487=>"000000100",
  43488=>"000000000",
  43489=>"000000000",
  43490=>"000000100",
  43491=>"111111011",
  43492=>"110010011",
  43493=>"011000000",
  43494=>"000111000",
  43495=>"111100000",
  43496=>"000000111",
  43497=>"111111111",
  43498=>"110111001",
  43499=>"011111000",
  43500=>"110000000",
  43501=>"111111011",
  43502=>"000000000",
  43503=>"000100110",
  43504=>"100100000",
  43505=>"000000110",
  43506=>"100110010",
  43507=>"000000000",
  43508=>"111111110",
  43509=>"001111111",
  43510=>"000000000",
  43511=>"010000000",
  43512=>"000100100",
  43513=>"000100111",
  43514=>"000010010",
  43515=>"111000011",
  43516=>"011000000",
  43517=>"101111111",
  43518=>"011011111",
  43519=>"000000000",
  43520=>"001001001",
  43521=>"000010000",
  43522=>"110111111",
  43523=>"111111100",
  43524=>"001011111",
  43525=>"000100100",
  43526=>"111011111",
  43527=>"000111111",
  43528=>"000000100",
  43529=>"111111111",
  43530=>"000000000",
  43531=>"000000000",
  43532=>"000100000",
  43533=>"111011001",
  43534=>"111111011",
  43535=>"111111111",
  43536=>"100000111",
  43537=>"000000000",
  43538=>"000000001",
  43539=>"110100011",
  43540=>"000000000",
  43541=>"000000000",
  43542=>"010010100",
  43543=>"111111011",
  43544=>"001000000",
  43545=>"110110111",
  43546=>"100000000",
  43547=>"011111001",
  43548=>"000111111",
  43549=>"111111111",
  43550=>"011111011",
  43551=>"111011001",
  43552=>"000010011",
  43553=>"111111000",
  43554=>"011111111",
  43555=>"000001001",
  43556=>"000010111",
  43557=>"000000000",
  43558=>"010111111",
  43559=>"001001000",
  43560=>"000111111",
  43561=>"000010000",
  43562=>"111111101",
  43563=>"111011111",
  43564=>"000011011",
  43565=>"000000110",
  43566=>"000000001",
  43567=>"000110110",
  43568=>"110000000",
  43569=>"001000000",
  43570=>"100100110",
  43571=>"000110111",
  43572=>"100110000",
  43573=>"000000000",
  43574=>"001111100",
  43575=>"001000110",
  43576=>"001100000",
  43577=>"110100000",
  43578=>"101000000",
  43579=>"000010111",
  43580=>"111100000",
  43581=>"100000000",
  43582=>"101110110",
  43583=>"100000000",
  43584=>"011011111",
  43585=>"111101000",
  43586=>"111000111",
  43587=>"111111000",
  43588=>"111100101",
  43589=>"001000111",
  43590=>"111110000",
  43591=>"000000000",
  43592=>"111111111",
  43593=>"111000000",
  43594=>"011111111",
  43595=>"111000000",
  43596=>"000101010",
  43597=>"000000000",
  43598=>"010111111",
  43599=>"011001011",
  43600=>"011111111",
  43601=>"000000000",
  43602=>"001111110",
  43603=>"010111000",
  43604=>"111111000",
  43605=>"001111111",
  43606=>"000000011",
  43607=>"111000000",
  43608=>"111101000",
  43609=>"000000000",
  43610=>"110111000",
  43611=>"110001111",
  43612=>"000000000",
  43613=>"000000001",
  43614=>"111111000",
  43615=>"001000000",
  43616=>"000001000",
  43617=>"111110111",
  43618=>"011000000",
  43619=>"000000000",
  43620=>"001001111",
  43621=>"000000101",
  43622=>"000000111",
  43623=>"001001011",
  43624=>"100100000",
  43625=>"111000011",
  43626=>"111000000",
  43627=>"000100111",
  43628=>"001001100",
  43629=>"001000111",
  43630=>"111111000",
  43631=>"111111000",
  43632=>"011011000",
  43633=>"000000111",
  43634=>"111111100",
  43635=>"000000000",
  43636=>"111000000",
  43637=>"011000011",
  43638=>"000000000",
  43639=>"000001001",
  43640=>"111011001",
  43641=>"111000100",
  43642=>"011000011",
  43643=>"000000000",
  43644=>"100111111",
  43645=>"011000111",
  43646=>"111000000",
  43647=>"110110111",
  43648=>"111111000",
  43649=>"011000110",
  43650=>"111111100",
  43651=>"000000010",
  43652=>"111111111",
  43653=>"111111111",
  43654=>"111011000",
  43655=>"010011011",
  43656=>"110111111",
  43657=>"111000000",
  43658=>"000100000",
  43659=>"100111110",
  43660=>"111011000",
  43661=>"111100111",
  43662=>"100000000",
  43663=>"111111111",
  43664=>"110000000",
  43665=>"011000000",
  43666=>"001111111",
  43667=>"111111111",
  43668=>"111100000",
  43669=>"111111000",
  43670=>"000000000",
  43671=>"111100000",
  43672=>"111111110",
  43673=>"000000111",
  43674=>"010000000",
  43675=>"101011111",
  43676=>"000000000",
  43677=>"001101001",
  43678=>"000000111",
  43679=>"110100111",
  43680=>"111111001",
  43681=>"111111000",
  43682=>"001111111",
  43683=>"001011111",
  43684=>"000001011",
  43685=>"000001111",
  43686=>"000110111",
  43687=>"001011001",
  43688=>"000000000",
  43689=>"110000000",
  43690=>"111000000",
  43691=>"100111111",
  43692=>"001011111",
  43693=>"100100000",
  43694=>"000000011",
  43695=>"111111011",
  43696=>"100000000",
  43697=>"111111100",
  43698=>"000010010",
  43699=>"111111001",
  43700=>"000000111",
  43701=>"111101111",
  43702=>"111111111",
  43703=>"100000000",
  43704=>"100101111",
  43705=>"111111111",
  43706=>"000000000",
  43707=>"111111000",
  43708=>"001111111",
  43709=>"000000000",
  43710=>"111111101",
  43711=>"111111111",
  43712=>"000000000",
  43713=>"011111111",
  43714=>"111000010",
  43715=>"110111000",
  43716=>"111111111",
  43717=>"000000000",
  43718=>"100000000",
  43719=>"000100100",
  43720=>"000000100",
  43721=>"100000000",
  43722=>"100100101",
  43723=>"001001011",
  43724=>"100100101",
  43725=>"000000000",
  43726=>"111111011",
  43727=>"000001111",
  43728=>"110110000",
  43729=>"010000000",
  43730=>"000100110",
  43731=>"111011111",
  43732=>"000101111",
  43733=>"110110111",
  43734=>"000000000",
  43735=>"000111111",
  43736=>"101000000",
  43737=>"000000000",
  43738=>"000000000",
  43739=>"000000111",
  43740=>"111001101",
  43741=>"100100110",
  43742=>"011011000",
  43743=>"011111111",
  43744=>"101111000",
  43745=>"100011000",
  43746=>"000000000",
  43747=>"000000000",
  43748=>"011010011",
  43749=>"111111100",
  43750=>"111000000",
  43751=>"111010000",
  43752=>"000000000",
  43753=>"111111111",
  43754=>"111111001",
  43755=>"011011001",
  43756=>"110111111",
  43757=>"000000000",
  43758=>"000011111",
  43759=>"111101111",
  43760=>"110100000",
  43761=>"111111110",
  43762=>"111001111",
  43763=>"000000101",
  43764=>"111111000",
  43765=>"000000000",
  43766=>"011111111",
  43767=>"000100100",
  43768=>"101100111",
  43769=>"000000000",
  43770=>"111000011",
  43771=>"000011000",
  43772=>"101100010",
  43773=>"011000111",
  43774=>"000000000",
  43775=>"001001001",
  43776=>"110000000",
  43777=>"111111111",
  43778=>"000000010",
  43779=>"111101101",
  43780=>"000000000",
  43781=>"111000000",
  43782=>"000000111",
  43783=>"111111001",
  43784=>"111111000",
  43785=>"110001000",
  43786=>"111000000",
  43787=>"111111111",
  43788=>"110100000",
  43789=>"001000000",
  43790=>"001011111",
  43791=>"100110000",
  43792=>"111000000",
  43793=>"111111001",
  43794=>"000000111",
  43795=>"111111001",
  43796=>"111111011",
  43797=>"011000000",
  43798=>"111001110",
  43799=>"111111010",
  43800=>"100101101",
  43801=>"010111001",
  43802=>"111111110",
  43803=>"111111011",
  43804=>"000001111",
  43805=>"001101111",
  43806=>"001001000",
  43807=>"000000111",
  43808=>"100111111",
  43809=>"011000011",
  43810=>"111111010",
  43811=>"111111111",
  43812=>"100100000",
  43813=>"000000100",
  43814=>"111111000",
  43815=>"000000001",
  43816=>"000000000",
  43817=>"111111001",
  43818=>"000000000",
  43819=>"111111111",
  43820=>"111100100",
  43821=>"101111111",
  43822=>"000000111",
  43823=>"111000100",
  43824=>"000000111",
  43825=>"111111111",
  43826=>"111010000",
  43827=>"010111111",
  43828=>"000000000",
  43829=>"111100110",
  43830=>"000000000",
  43831=>"111111110",
  43832=>"000011000",
  43833=>"111100111",
  43834=>"110000000",
  43835=>"000111111",
  43836=>"001000100",
  43837=>"101100111",
  43838=>"011111110",
  43839=>"111111001",
  43840=>"111111111",
  43841=>"000000101",
  43842=>"100000110",
  43843=>"111000000",
  43844=>"111111000",
  43845=>"110101011",
  43846=>"111001000",
  43847=>"111111111",
  43848=>"000110111",
  43849=>"000000000",
  43850=>"000000000",
  43851=>"001000100",
  43852=>"111011111",
  43853=>"111111000",
  43854=>"000001011",
  43855=>"100100100",
  43856=>"011011100",
  43857=>"100011111",
  43858=>"101000110",
  43859=>"111111111",
  43860=>"000000000",
  43861=>"001011000",
  43862=>"011000000",
  43863=>"000011111",
  43864=>"000100000",
  43865=>"000000000",
  43866=>"110111111",
  43867=>"000000111",
  43868=>"000000001",
  43869=>"100001111",
  43870=>"000000000",
  43871=>"000001010",
  43872=>"110111000",
  43873=>"111111111",
  43874=>"000110000",
  43875=>"000000001",
  43876=>"110100110",
  43877=>"000100001",
  43878=>"000111111",
  43879=>"000001111",
  43880=>"110110110",
  43881=>"000110111",
  43882=>"110110111",
  43883=>"111111100",
  43884=>"000111111",
  43885=>"000000100",
  43886=>"000000000",
  43887=>"000000111",
  43888=>"010011111",
  43889=>"111111111",
  43890=>"100111111",
  43891=>"000100110",
  43892=>"111000000",
  43893=>"111001000",
  43894=>"101111111",
  43895=>"000000100",
  43896=>"111111111",
  43897=>"000000111",
  43898=>"111111111",
  43899=>"000000000",
  43900=>"111110000",
  43901=>"000000111",
  43902=>"111111000",
  43903=>"000000000",
  43904=>"000100111",
  43905=>"011011101",
  43906=>"001000000",
  43907=>"000000000",
  43908=>"000111011",
  43909=>"011011011",
  43910=>"111111001",
  43911=>"100000000",
  43912=>"000000000",
  43913=>"100000110",
  43914=>"000010000",
  43915=>"111110010",
  43916=>"111111111",
  43917=>"000000101",
  43918=>"000000010",
  43919=>"000110111",
  43920=>"111111000",
  43921=>"001001001",
  43922=>"000111111",
  43923=>"100000001",
  43924=>"111111111",
  43925=>"000000000",
  43926=>"000000000",
  43927=>"000000100",
  43928=>"000000000",
  43929=>"001001111",
  43930=>"111111000",
  43931=>"000000100",
  43932=>"101000000",
  43933=>"000000011",
  43934=>"001001011",
  43935=>"000000000",
  43936=>"011011001",
  43937=>"001011000",
  43938=>"000000110",
  43939=>"000000011",
  43940=>"110100000",
  43941=>"000010010",
  43942=>"000000000",
  43943=>"011111011",
  43944=>"000000011",
  43945=>"111011011",
  43946=>"111111111",
  43947=>"111101000",
  43948=>"110100000",
  43949=>"000000000",
  43950=>"100100111",
  43951=>"110110111",
  43952=>"011111111",
  43953=>"000111111",
  43954=>"000000101",
  43955=>"001001011",
  43956=>"100011011",
  43957=>"111111111",
  43958=>"101111011",
  43959=>"100000000",
  43960=>"000000111",
  43961=>"100111111",
  43962=>"000111111",
  43963=>"001000111",
  43964=>"000000000",
  43965=>"101000110",
  43966=>"000100110",
  43967=>"101100100",
  43968=>"100101000",
  43969=>"111110010",
  43970=>"111111111",
  43971=>"000000000",
  43972=>"000000111",
  43973=>"111110000",
  43974=>"010000011",
  43975=>"101000000",
  43976=>"110011111",
  43977=>"110110000",
  43978=>"100000000",
  43979=>"011111111",
  43980=>"111001010",
  43981=>"111111001",
  43982=>"000000010",
  43983=>"000010011",
  43984=>"000000011",
  43985=>"111111000",
  43986=>"111100111",
  43987=>"111111111",
  43988=>"100100100",
  43989=>"010011000",
  43990=>"111111000",
  43991=>"000000101",
  43992=>"110111110",
  43993=>"011101111",
  43994=>"100111111",
  43995=>"011001000",
  43996=>"100100000",
  43997=>"000000111",
  43998=>"010011111",
  43999=>"011001001",
  44000=>"111000000",
  44001=>"001000000",
  44002=>"010000000",
  44003=>"011011111",
  44004=>"000111111",
  44005=>"111111111",
  44006=>"111111111",
  44007=>"000000000",
  44008=>"000000001",
  44009=>"000000111",
  44010=>"000100110",
  44011=>"000100111",
  44012=>"000100101",
  44013=>"000000000",
  44014=>"111010000",
  44015=>"110111000",
  44016=>"001001111",
  44017=>"111111111",
  44018=>"101111110",
  44019=>"000000010",
  44020=>"111111111",
  44021=>"011011001",
  44022=>"000111101",
  44023=>"000100111",
  44024=>"001001111",
  44025=>"000000000",
  44026=>"111000000",
  44027=>"111101000",
  44028=>"000100000",
  44029=>"111011001",
  44030=>"011000000",
  44031=>"101000001",
  44032=>"111011111",
  44033=>"111111111",
  44034=>"000001111",
  44035=>"111111111",
  44036=>"001000001",
  44037=>"001000010",
  44038=>"000000000",
  44039=>"101000000",
  44040=>"111111000",
  44041=>"100000000",
  44042=>"000000000",
  44043=>"000000001",
  44044=>"000000000",
  44045=>"000000011",
  44046=>"000000100",
  44047=>"111111111",
  44048=>"011111111",
  44049=>"000000000",
  44050=>"000000000",
  44051=>"000000000",
  44052=>"111111111",
  44053=>"110110111",
  44054=>"000000000",
  44055=>"111111111",
  44056=>"110110110",
  44057=>"100110000",
  44058=>"101000011",
  44059=>"110110100",
  44060=>"000000000",
  44061=>"000000000",
  44062=>"011011110",
  44063=>"111111111",
  44064=>"000000010",
  44065=>"111111111",
  44066=>"111100000",
  44067=>"100000111",
  44068=>"001001000",
  44069=>"010001001",
  44070=>"111111110",
  44071=>"111111000",
  44072=>"011011000",
  44073=>"111101000",
  44074=>"000000000",
  44075=>"110110110",
  44076=>"111101011",
  44077=>"110111111",
  44078=>"001001000",
  44079=>"111111111",
  44080=>"000000111",
  44081=>"000000000",
  44082=>"000100001",
  44083=>"000000000",
  44084=>"110110000",
  44085=>"101011011",
  44086=>"000111111",
  44087=>"011010111",
  44088=>"111111111",
  44089=>"111101111",
  44090=>"000000000",
  44091=>"111111011",
  44092=>"111100000",
  44093=>"000111111",
  44094=>"011011111",
  44095=>"111111111",
  44096=>"000001111",
  44097=>"111110111",
  44098=>"111000000",
  44099=>"101000000",
  44100=>"111111111",
  44101=>"111110110",
  44102=>"111001000",
  44103=>"000000010",
  44104=>"111111111",
  44105=>"000000110",
  44106=>"101000000",
  44107=>"001001001",
  44108=>"000111000",
  44109=>"000000001",
  44110=>"111111110",
  44111=>"000000101",
  44112=>"000000000",
  44113=>"000000110",
  44114=>"000000000",
  44115=>"000000110",
  44116=>"001001011",
  44117=>"000111101",
  44118=>"000000100",
  44119=>"000000000",
  44120=>"111111111",
  44121=>"100000111",
  44122=>"001111111",
  44123=>"110100101",
  44124=>"111111111",
  44125=>"000001000",
  44126=>"100000000",
  44127=>"000111111",
  44128=>"111111110",
  44129=>"111000100",
  44130=>"111111111",
  44131=>"010000000",
  44132=>"101100111",
  44133=>"111100100",
  44134=>"010000111",
  44135=>"000000000",
  44136=>"111111111",
  44137=>"110111111",
  44138=>"111001111",
  44139=>"000000000",
  44140=>"111111111",
  44141=>"000000000",
  44142=>"001001000",
  44143=>"001111000",
  44144=>"000000111",
  44145=>"111011001",
  44146=>"010010011",
  44147=>"111111111",
  44148=>"111100000",
  44149=>"000001011",
  44150=>"111111111",
  44151=>"001001101",
  44152=>"111111010",
  44153=>"000000000",
  44154=>"001001111",
  44155=>"111111111",
  44156=>"010000000",
  44157=>"010000000",
  44158=>"010001001",
  44159=>"111111110",
  44160=>"000000000",
  44161=>"000111111",
  44162=>"000001111",
  44163=>"000000000",
  44164=>"111101000",
  44165=>"000000000",
  44166=>"000100000",
  44167=>"000001011",
  44168=>"100000000",
  44169=>"000000000",
  44170=>"000000000",
  44171=>"000000000",
  44172=>"111111111",
  44173=>"110110000",
  44174=>"110111101",
  44175=>"111111111",
  44176=>"111111111",
  44177=>"111111111",
  44178=>"000111111",
  44179=>"001000000",
  44180=>"111111011",
  44181=>"111111111",
  44182=>"111111111",
  44183=>"111111111",
  44184=>"001000001",
  44185=>"111111111",
  44186=>"111111111",
  44187=>"111001000",
  44188=>"000000000",
  44189=>"100000000",
  44190=>"110111111",
  44191=>"110110100",
  44192=>"000000000",
  44193=>"101101101",
  44194=>"111111111",
  44195=>"111111110",
  44196=>"110111111",
  44197=>"110000000",
  44198=>"111111111",
  44199=>"100100000",
  44200=>"000000000",
  44201=>"000000000",
  44202=>"000000000",
  44203=>"000000000",
  44204=>"111111111",
  44205=>"000000001",
  44206=>"000000000",
  44207=>"011011001",
  44208=>"000000100",
  44209=>"000000000",
  44210=>"110111111",
  44211=>"111111000",
  44212=>"001001111",
  44213=>"011111111",
  44214=>"111001111",
  44215=>"111101001",
  44216=>"000111111",
  44217=>"010000100",
  44218=>"001011111",
  44219=>"011000000",
  44220=>"000000000",
  44221=>"111101000",
  44222=>"111111111",
  44223=>"000000000",
  44224=>"000000100",
  44225=>"000000000",
  44226=>"000000111",
  44227=>"111111111",
  44228=>"000100000",
  44229=>"111111111",
  44230=>"011001111",
  44231=>"000000011",
  44232=>"111111111",
  44233=>"000000000",
  44234=>"011000100",
  44235=>"011011000",
  44236=>"001000111",
  44237=>"000000000",
  44238=>"111111111",
  44239=>"001001111",
  44240=>"001000100",
  44241=>"001101101",
  44242=>"011011111",
  44243=>"000000001",
  44244=>"000000010",
  44245=>"111111111",
  44246=>"111111111",
  44247=>"111000100",
  44248=>"111111111",
  44249=>"011001001",
  44250=>"000000000",
  44251=>"000000000",
  44252=>"111111111",
  44253=>"111111111",
  44254=>"000000000",
  44255=>"001011001",
  44256=>"111111000",
  44257=>"111111111",
  44258=>"000000000",
  44259=>"111111111",
  44260=>"111111111",
  44261=>"110111111",
  44262=>"010000000",
  44263=>"111111000",
  44264=>"111111111",
  44265=>"111011111",
  44266=>"111111111",
  44267=>"000000000",
  44268=>"111000000",
  44269=>"000000000",
  44270=>"111111000",
  44271=>"000011000",
  44272=>"000000011",
  44273=>"000000000",
  44274=>"011000001",
  44275=>"000000000",
  44276=>"000111111",
  44277=>"000001111",
  44278=>"111110000",
  44279=>"001000000",
  44280=>"011000010",
  44281=>"000000000",
  44282=>"011000000",
  44283=>"111111111",
  44284=>"111111100",
  44285=>"111111111",
  44286=>"000000111",
  44287=>"100111111",
  44288=>"111111111",
  44289=>"110110100",
  44290=>"110000111",
  44291=>"011000000",
  44292=>"111111111",
  44293=>"000000100",
  44294=>"001101111",
  44295=>"111111111",
  44296=>"111011111",
  44297=>"001111111",
  44298=>"000100100",
  44299=>"111111110",
  44300=>"111111100",
  44301=>"010111111",
  44302=>"000000000",
  44303=>"001011000",
  44304=>"111011001",
  44305=>"100100010",
  44306=>"111111111",
  44307=>"100000000",
  44308=>"111111011",
  44309=>"000000011",
  44310=>"011011011",
  44311=>"100000001",
  44312=>"000000001",
  44313=>"111111111",
  44314=>"111111111",
  44315=>"000000110",
  44316=>"111110111",
  44317=>"000000000",
  44318=>"111001000",
  44319=>"110111111",
  44320=>"000000000",
  44321=>"001001000",
  44322=>"111000100",
  44323=>"010000000",
  44324=>"001001001",
  44325=>"111000100",
  44326=>"000011111",
  44327=>"110000000",
  44328=>"001101101",
  44329=>"110111111",
  44330=>"000000010",
  44331=>"010010011",
  44332=>"111111000",
  44333=>"111111110",
  44334=>"000000000",
  44335=>"110000000",
  44336=>"001001001",
  44337=>"111111111",
  44338=>"000001111",
  44339=>"111000101",
  44340=>"000000000",
  44341=>"111111000",
  44342=>"000001001",
  44343=>"111111111",
  44344=>"111111111",
  44345=>"000000000",
  44346=>"111111111",
  44347=>"001000000",
  44348=>"000000000",
  44349=>"001011000",
  44350=>"000001001",
  44351=>"111111001",
  44352=>"111100000",
  44353=>"000000011",
  44354=>"000110111",
  44355=>"111111111",
  44356=>"001000111",
  44357=>"110010100",
  44358=>"111111111",
  44359=>"111011011",
  44360=>"100000100",
  44361=>"111111110",
  44362=>"000011111",
  44363=>"000000011",
  44364=>"000000000",
  44365=>"000000111",
  44366=>"000000001",
  44367=>"011001001",
  44368=>"110011000",
  44369=>"000000000",
  44370=>"000000000",
  44371=>"000000001",
  44372=>"000000111",
  44373=>"000100000",
  44374=>"001001001",
  44375=>"111000000",
  44376=>"111000000",
  44377=>"000000100",
  44378=>"010010001",
  44379=>"001000000",
  44380=>"100000000",
  44381=>"000000000",
  44382=>"000000000",
  44383=>"001001001",
  44384=>"111111111",
  44385=>"000000000",
  44386=>"100110111",
  44387=>"000000000",
  44388=>"111111111",
  44389=>"000011011",
  44390=>"000000000",
  44391=>"111111111",
  44392=>"110110111",
  44393=>"001000000",
  44394=>"000110010",
  44395=>"111111111",
  44396=>"111011001",
  44397=>"001000111",
  44398=>"000000000",
  44399=>"111111111",
  44400=>"001001111",
  44401=>"111111001",
  44402=>"111111111",
  44403=>"000000000",
  44404=>"000000000",
  44405=>"111111111",
  44406=>"111111111",
  44407=>"111111111",
  44408=>"100110100",
  44409=>"000000000",
  44410=>"111111111",
  44411=>"011100000",
  44412=>"000000100",
  44413=>"111111111",
  44414=>"001000000",
  44415=>"111111111",
  44416=>"000000000",
  44417=>"001000001",
  44418=>"101101000",
  44419=>"000000000",
  44420=>"000000000",
  44421=>"111000011",
  44422=>"001000100",
  44423=>"100000000",
  44424=>"111111111",
  44425=>"111111111",
  44426=>"111111111",
  44427=>"011000000",
  44428=>"000110000",
  44429=>"111111111",
  44430=>"111111111",
  44431=>"111111111",
  44432=>"011001010",
  44433=>"110010000",
  44434=>"111111111",
  44435=>"000111111",
  44436=>"111111111",
  44437=>"111111111",
  44438=>"000000000",
  44439=>"111010010",
  44440=>"001000000",
  44441=>"101111100",
  44442=>"111111111",
  44443=>"000000000",
  44444=>"111111110",
  44445=>"000000001",
  44446=>"000000000",
  44447=>"111111111",
  44448=>"111111110",
  44449=>"110000000",
  44450=>"111111101",
  44451=>"000000100",
  44452=>"100111111",
  44453=>"111111111",
  44454=>"111111111",
  44455=>"000000000",
  44456=>"100111001",
  44457=>"000000110",
  44458=>"011111111",
  44459=>"111111111",
  44460=>"111111101",
  44461=>"000000000",
  44462=>"001000001",
  44463=>"111111111",
  44464=>"010000110",
  44465=>"001000001",
  44466=>"111000000",
  44467=>"110000000",
  44468=>"010000000",
  44469=>"000000111",
  44470=>"110111111",
  44471=>"011110000",
  44472=>"100110100",
  44473=>"011011111",
  44474=>"011111111",
  44475=>"111000111",
  44476=>"011111001",
  44477=>"111111111",
  44478=>"111000000",
  44479=>"001101000",
  44480=>"111110000",
  44481=>"000000000",
  44482=>"000000000",
  44483=>"111111011",
  44484=>"000100111",
  44485=>"001000001",
  44486=>"000000000",
  44487=>"111111111",
  44488=>"011011001",
  44489=>"110100100",
  44490=>"001000000",
  44491=>"000000111",
  44492=>"000000110",
  44493=>"000000001",
  44494=>"000000000",
  44495=>"111111000",
  44496=>"111100000",
  44497=>"011100000",
  44498=>"101001001",
  44499=>"000000001",
  44500=>"011111111",
  44501=>"001001111",
  44502=>"111111000",
  44503=>"000000111",
  44504=>"111111110",
  44505=>"111000000",
  44506=>"000001000",
  44507=>"001001001",
  44508=>"001000000",
  44509=>"111111101",
  44510=>"000111000",
  44511=>"110100100",
  44512=>"111111000",
  44513=>"111110000",
  44514=>"111111111",
  44515=>"111010010",
  44516=>"111111111",
  44517=>"111111011",
  44518=>"111111111",
  44519=>"000000011",
  44520=>"000000100",
  44521=>"000000101",
  44522=>"000000000",
  44523=>"111111000",
  44524=>"000011000",
  44525=>"111000000",
  44526=>"010000000",
  44527=>"111001001",
  44528=>"000000000",
  44529=>"000000000",
  44530=>"111111111",
  44531=>"111111100",
  44532=>"000000000",
  44533=>"111111110",
  44534=>"111111111",
  44535=>"111011001",
  44536=>"111010010",
  44537=>"000000000",
  44538=>"111011111",
  44539=>"100111111",
  44540=>"000111001",
  44541=>"000000000",
  44542=>"000000000",
  44543=>"111111000",
  44544=>"110111111",
  44545=>"000001001",
  44546=>"000000110",
  44547=>"111111111",
  44548=>"111110000",
  44549=>"000000000",
  44550=>"000111111",
  44551=>"111111111",
  44552=>"111000000",
  44553=>"111001111",
  44554=>"000000000",
  44555=>"110110000",
  44556=>"100110100",
  44557=>"111000100",
  44558=>"001111111",
  44559=>"100100100",
  44560=>"000000100",
  44561=>"110111100",
  44562=>"010111000",
  44563=>"111111100",
  44564=>"000000000",
  44565=>"111000000",
  44566=>"000000001",
  44567=>"111111110",
  44568=>"100000000",
  44569=>"111111111",
  44570=>"111010000",
  44571=>"000001111",
  44572=>"111111110",
  44573=>"000110110",
  44574=>"000011111",
  44575=>"000000111",
  44576=>"110110111",
  44577=>"111100001",
  44578=>"110110111",
  44579=>"111011001",
  44580=>"000001111",
  44581=>"110111000",
  44582=>"001001001",
  44583=>"101001111",
  44584=>"000010010",
  44585=>"111111000",
  44586=>"000000000",
  44587=>"000000111",
  44588=>"001111100",
  44589=>"110110000",
  44590=>"101101000",
  44591=>"010011111",
  44592=>"000000101",
  44593=>"111111110",
  44594=>"010000011",
  44595=>"001001100",
  44596=>"110111111",
  44597=>"111111110",
  44598=>"000000011",
  44599=>"001011000",
  44600=>"111111111",
  44601=>"100000001",
  44602=>"110010110",
  44603=>"011000001",
  44604=>"101100100",
  44605=>"111010000",
  44606=>"010011111",
  44607=>"111111011",
  44608=>"000100111",
  44609=>"001111111",
  44610=>"001001001",
  44611=>"010000101",
  44612=>"110100100",
  44613=>"000000001",
  44614=>"000000000",
  44615=>"101001101",
  44616=>"000010111",
  44617=>"111111111",
  44618=>"111000000",
  44619=>"111111111",
  44620=>"111111000",
  44621=>"110111000",
  44622=>"001001000",
  44623=>"111000101",
  44624=>"000001111",
  44625=>"000001111",
  44626=>"111101000",
  44627=>"100010000",
  44628=>"111111010",
  44629=>"111110000",
  44630=>"111110010",
  44631=>"001001000",
  44632=>"111110111",
  44633=>"111001101",
  44634=>"110001001",
  44635=>"000000100",
  44636=>"000000000",
  44637=>"001000111",
  44638=>"011001001",
  44639=>"000010000",
  44640=>"001111110",
  44641=>"000001101",
  44642=>"000101000",
  44643=>"111011011",
  44644=>"110010000",
  44645=>"111000111",
  44646=>"000000010",
  44647=>"111111111",
  44648=>"111011011",
  44649=>"001000101",
  44650=>"001000000",
  44651=>"110111000",
  44652=>"001011111",
  44653=>"000101111",
  44654=>"111100000",
  44655=>"111110110",
  44656=>"101001000",
  44657=>"000001010",
  44658=>"000010111",
  44659=>"001001111",
  44660=>"001111111",
  44661=>"010110111",
  44662=>"011111111",
  44663=>"101000110",
  44664=>"100000001",
  44665=>"011000000",
  44666=>"101000000",
  44667=>"111111011",
  44668=>"000111111",
  44669=>"001000000",
  44670=>"000000101",
  44671=>"101101001",
  44672=>"000001011",
  44673=>"111000000",
  44674=>"000111100",
  44675=>"111110110",
  44676=>"000001111",
  44677=>"111111000",
  44678=>"111111110",
  44679=>"011011001",
  44680=>"111001001",
  44681=>"100000001",
  44682=>"000000100",
  44683=>"111011111",
  44684=>"000000110",
  44685=>"110000100",
  44686=>"111011000",
  44687=>"000111111",
  44688=>"001101111",
  44689=>"100001001",
  44690=>"100110000",
  44691=>"001000000",
  44692=>"111111111",
  44693=>"110100000",
  44694=>"101000000",
  44695=>"111101101",
  44696=>"001001101",
  44697=>"000000000",
  44698=>"110111111",
  44699=>"000000011",
  44700=>"001000011",
  44701=>"110111011",
  44702=>"111101000",
  44703=>"000111111",
  44704=>"010000000",
  44705=>"100000000",
  44706=>"111111010",
  44707=>"000111111",
  44708=>"101000000",
  44709=>"000000110",
  44710=>"111000011",
  44711=>"111010100",
  44712=>"001000000",
  44713=>"000001001",
  44714=>"111101111",
  44715=>"101001111",
  44716=>"111111111",
  44717=>"101101111",
  44718=>"000000110",
  44719=>"111000100",
  44720=>"111110000",
  44721=>"100000111",
  44722=>"111110000",
  44723=>"000000000",
  44724=>"000000011",
  44725=>"001001111",
  44726=>"000010011",
  44727=>"111111111",
  44728=>"001111111",
  44729=>"111111111",
  44730=>"111000000",
  44731=>"111000000",
  44732=>"001111111",
  44733=>"100000111",
  44734=>"111111111",
  44735=>"111111110",
  44736=>"100000100",
  44737=>"000000001",
  44738=>"110010000",
  44739=>"110110010",
  44740=>"000000110",
  44741=>"001001000",
  44742=>"101001000",
  44743=>"111010000",
  44744=>"001000100",
  44745=>"101000000",
  44746=>"000000000",
  44747=>"101101111",
  44748=>"111111110",
  44749=>"100110110",
  44750=>"000001100",
  44751=>"110000000",
  44752=>"000000011",
  44753=>"000001000",
  44754=>"000000011",
  44755=>"110100101",
  44756=>"100010010",
  44757=>"111111111",
  44758=>"111100111",
  44759=>"001001111",
  44760=>"111000000",
  44761=>"001000001",
  44762=>"111111111",
  44763=>"111110100",
  44764=>"111000001",
  44765=>"000000011",
  44766=>"000000111",
  44767=>"000000001",
  44768=>"111111111",
  44769=>"001000000",
  44770=>"000000000",
  44771=>"101001111",
  44772=>"000110111",
  44773=>"000000001",
  44774=>"110110000",
  44775=>"111111110",
  44776=>"001000111",
  44777=>"111111111",
  44778=>"111111111",
  44779=>"001101001",
  44780=>"100000000",
  44781=>"110111110",
  44782=>"111111111",
  44783=>"100000000",
  44784=>"111110111",
  44785=>"011001000",
  44786=>"111111111",
  44787=>"000000100",
  44788=>"001000110",
  44789=>"000001011",
  44790=>"111110110",
  44791=>"000100100",
  44792=>"011000010",
  44793=>"000111111",
  44794=>"111000001",
  44795=>"111001000",
  44796=>"111111111",
  44797=>"001001101",
  44798=>"001000000",
  44799=>"110111111",
  44800=>"111000110",
  44801=>"100000001",
  44802=>"000010011",
  44803=>"000001011",
  44804=>"001001001",
  44805=>"000000000",
  44806=>"000000000",
  44807=>"110110000",
  44808=>"111111111",
  44809=>"000000000",
  44810=>"110111111",
  44811=>"110111111",
  44812=>"001001001",
  44813=>"100100111",
  44814=>"110110000",
  44815=>"011011011",
  44816=>"010100000",
  44817=>"000000000",
  44818=>"101001000",
  44819=>"100000001",
  44820=>"000000010",
  44821=>"000000000",
  44822=>"001111111",
  44823=>"110111111",
  44824=>"110000010",
  44825=>"111111001",
  44826=>"000000001",
  44827=>"111101011",
  44828=>"111100100",
  44829=>"111000000",
  44830=>"010100111",
  44831=>"100001001",
  44832=>"010000000",
  44833=>"101000001",
  44834=>"000011111",
  44835=>"111111111",
  44836=>"000000010",
  44837=>"111001000",
  44838=>"111111100",
  44839=>"001000110",
  44840=>"000000001",
  44841=>"110111110",
  44842=>"000000000",
  44843=>"000000011",
  44844=>"000000111",
  44845=>"111110110",
  44846=>"000000000",
  44847=>"100001111",
  44848=>"001000000",
  44849=>"110111000",
  44850=>"110111000",
  44851=>"001111111",
  44852=>"001001000",
  44853=>"111100011",
  44854=>"000000000",
  44855=>"000000100",
  44856=>"000001111",
  44857=>"000001001",
  44858=>"000000101",
  44859=>"111111111",
  44860=>"000000011",
  44861=>"111001001",
  44862=>"100101111",
  44863=>"000000000",
  44864=>"001101111",
  44865=>"000000000",
  44866=>"001000000",
  44867=>"001000000",
  44868=>"001001000",
  44869=>"101100111",
  44870=>"111111111",
  44871=>"111111111",
  44872=>"111000001",
  44873=>"000000000",
  44874=>"111001001",
  44875=>"101000000",
  44876=>"000000000",
  44877=>"111111111",
  44878=>"110000011",
  44879=>"010010100",
  44880=>"000110111",
  44881=>"100100000",
  44882=>"000011111",
  44883=>"111111111",
  44884=>"000000000",
  44885=>"001011111",
  44886=>"111101101",
  44887=>"000000000",
  44888=>"000000011",
  44889=>"100000010",
  44890=>"111111101",
  44891=>"000000000",
  44892=>"111011100",
  44893=>"000001000",
  44894=>"000001101",
  44895=>"000010000",
  44896=>"000000110",
  44897=>"001001001",
  44898=>"011010000",
  44899=>"000100000",
  44900=>"110110110",
  44901=>"101111111",
  44902=>"000101000",
  44903=>"110111111",
  44904=>"001000000",
  44905=>"010001101",
  44906=>"111111000",
  44907=>"101000001",
  44908=>"100010111",
  44909=>"000000000",
  44910=>"110111000",
  44911=>"100000000",
  44912=>"001001000",
  44913=>"001000000",
  44914=>"000000111",
  44915=>"110010000",
  44916=>"011011111",
  44917=>"011011111",
  44918=>"100100000",
  44919=>"001001101",
  44920=>"000000000",
  44921=>"111101000",
  44922=>"000000001",
  44923=>"100111111",
  44924=>"100000000",
  44925=>"000000000",
  44926=>"100000111",
  44927=>"000001001",
  44928=>"110100111",
  44929=>"001101101",
  44930=>"100000100",
  44931=>"001000001",
  44932=>"010111000",
  44933=>"000000000",
  44934=>"000000001",
  44935=>"111111000",
  44936=>"000000000",
  44937=>"010000000",
  44938=>"110110010",
  44939=>"000110110",
  44940=>"111101000",
  44941=>"111110000",
  44942=>"100111111",
  44943=>"000111000",
  44944=>"111111111",
  44945=>"110110111",
  44946=>"000110110",
  44947=>"000000110",
  44948=>"001001101",
  44949=>"000000000",
  44950=>"111110110",
  44951=>"011111111",
  44952=>"000001111",
  44953=>"000000001",
  44954=>"000000000",
  44955=>"110111111",
  44956=>"111111010",
  44957=>"111111111",
  44958=>"101100111",
  44959=>"111011000",
  44960=>"100001111",
  44961=>"111000011",
  44962=>"111001101",
  44963=>"001001111",
  44964=>"001001111",
  44965=>"010011000",
  44966=>"000000000",
  44967=>"001000001",
  44968=>"100101111",
  44969=>"111111000",
  44970=>"111111111",
  44971=>"000001001",
  44972=>"000000010",
  44973=>"000000110",
  44974=>"101001001",
  44975=>"111000000",
  44976=>"111101100",
  44977=>"111111110",
  44978=>"101001111",
  44979=>"000000001",
  44980=>"000000000",
  44981=>"001000000",
  44982=>"111101000",
  44983=>"000000110",
  44984=>"000000111",
  44985=>"111100100",
  44986=>"001111101",
  44987=>"000001000",
  44988=>"000000000",
  44989=>"000000000",
  44990=>"101001001",
  44991=>"001001111",
  44992=>"011000001",
  44993=>"101001101",
  44994=>"000001000",
  44995=>"111010000",
  44996=>"110110000",
  44997=>"101001000",
  44998=>"111001000",
  44999=>"011111110",
  45000=>"001000000",
  45001=>"000000000",
  45002=>"001001101",
  45003=>"000000000",
  45004=>"111111110",
  45005=>"001111011",
  45006=>"111100100",
  45007=>"111101101",
  45008=>"111111111",
  45009=>"111000000",
  45010=>"111111111",
  45011=>"101110111",
  45012=>"011001011",
  45013=>"111111000",
  45014=>"111111000",
  45015=>"011011010",
  45016=>"111000000",
  45017=>"000000000",
  45018=>"000001000",
  45019=>"111100000",
  45020=>"101100100",
  45021=>"000000000",
  45022=>"101111011",
  45023=>"101111110",
  45024=>"001101000",
  45025=>"000111111",
  45026=>"100100111",
  45027=>"111111111",
  45028=>"001111101",
  45029=>"000000000",
  45030=>"000000001",
  45031=>"111000000",
  45032=>"100111011",
  45033=>"111111000",
  45034=>"001001101",
  45035=>"111100101",
  45036=>"001001101",
  45037=>"000111111",
  45038=>"101001001",
  45039=>"111101001",
  45040=>"100000000",
  45041=>"110110000",
  45042=>"011000000",
  45043=>"001001001",
  45044=>"100000000",
  45045=>"111111011",
  45046=>"111111000",
  45047=>"100011011",
  45048=>"010000100",
  45049=>"000011001",
  45050=>"010110111",
  45051=>"001001100",
  45052=>"111000111",
  45053=>"111001000",
  45054=>"101101101",
  45055=>"000000000",
  45056=>"110111000",
  45057=>"111111111",
  45058=>"111101001",
  45059=>"111110001",
  45060=>"001000110",
  45061=>"101000000",
  45062=>"111111111",
  45063=>"101001001",
  45064=>"000000111",
  45065=>"011010000",
  45066=>"000000001",
  45067=>"011111100",
  45068=>"000110100",
  45069=>"000000100",
  45070=>"111111000",
  45071=>"000000111",
  45072=>"111101000",
  45073=>"111111111",
  45074=>"000000000",
  45075=>"111010000",
  45076=>"101000101",
  45077=>"111111111",
  45078=>"000001111",
  45079=>"000000111",
  45080=>"001001001",
  45081=>"111111111",
  45082=>"101111000",
  45083=>"001110000",
  45084=>"000000000",
  45085=>"001001001",
  45086=>"000111111",
  45087=>"100110111",
  45088=>"000000000",
  45089=>"000111111",
  45090=>"111111000",
  45091=>"011010000",
  45092=>"100000000",
  45093=>"010110000",
  45094=>"001001000",
  45095=>"111111111",
  45096=>"000000001",
  45097=>"111111111",
  45098=>"111011011",
  45099=>"111000010",
  45100=>"001001111",
  45101=>"000000000",
  45102=>"000100001",
  45103=>"111001001",
  45104=>"000000000",
  45105=>"000000111",
  45106=>"100100100",
  45107=>"111111101",
  45108=>"000111011",
  45109=>"100110100",
  45110=>"111111111",
  45111=>"000000100",
  45112=>"111111000",
  45113=>"001011111",
  45114=>"000111110",
  45115=>"000000111",
  45116=>"101000111",
  45117=>"111000001",
  45118=>"111111011",
  45119=>"001001100",
  45120=>"000000101",
  45121=>"110110111",
  45122=>"000000111",
  45123=>"011000000",
  45124=>"000001001",
  45125=>"010011011",
  45126=>"000000001",
  45127=>"111111111",
  45128=>"100111001",
  45129=>"111111111",
  45130=>"111111111",
  45131=>"011000110",
  45132=>"001001001",
  45133=>"111000100",
  45134=>"101001001",
  45135=>"000000010",
  45136=>"000000110",
  45137=>"000000000",
  45138=>"011011000",
  45139=>"000000000",
  45140=>"110110110",
  45141=>"000000100",
  45142=>"101110111",
  45143=>"000000111",
  45144=>"011001000",
  45145=>"111100111",
  45146=>"000001010",
  45147=>"110000100",
  45148=>"001001111",
  45149=>"101100111",
  45150=>"001000100",
  45151=>"101001000",
  45152=>"001001011",
  45153=>"110111000",
  45154=>"000000100",
  45155=>"000001001",
  45156=>"011010001",
  45157=>"111100000",
  45158=>"000011000",
  45159=>"111111111",
  45160=>"100110110",
  45161=>"000000010",
  45162=>"100000000",
  45163=>"000110111",
  45164=>"111111000",
  45165=>"111111100",
  45166=>"110000000",
  45167=>"011011001",
  45168=>"100111111",
  45169=>"011000000",
  45170=>"000000000",
  45171=>"001000000",
  45172=>"111111111",
  45173=>"111000001",
  45174=>"000000000",
  45175=>"111111110",
  45176=>"000000011",
  45177=>"000000000",
  45178=>"000110111",
  45179=>"000000001",
  45180=>"100100100",
  45181=>"000111111",
  45182=>"000111111",
  45183=>"100111101",
  45184=>"000000111",
  45185=>"111110010",
  45186=>"000110000",
  45187=>"001000001",
  45188=>"000000100",
  45189=>"111101000",
  45190=>"001000001",
  45191=>"000000111",
  45192=>"111001000",
  45193=>"110100111",
  45194=>"000000110",
  45195=>"000101110",
  45196=>"111001000",
  45197=>"111111000",
  45198=>"000111100",
  45199=>"000000000",
  45200=>"101101001",
  45201=>"000100111",
  45202=>"000010001",
  45203=>"000100100",
  45204=>"000000000",
  45205=>"101100111",
  45206=>"111100110",
  45207=>"001001011",
  45208=>"101000000",
  45209=>"000000100",
  45210=>"100100110",
  45211=>"000000101",
  45212=>"100000101",
  45213=>"011110100",
  45214=>"001000111",
  45215=>"000101111",
  45216=>"000011111",
  45217=>"011111111",
  45218=>"111111101",
  45219=>"000110110",
  45220=>"000111111",
  45221=>"111111100",
  45222=>"111111111",
  45223=>"000000000",
  45224=>"100100110",
  45225=>"111111111",
  45226=>"000110111",
  45227=>"111001000",
  45228=>"001001011",
  45229=>"000110011",
  45230=>"111101110",
  45231=>"011001001",
  45232=>"111111111",
  45233=>"100100111",
  45234=>"111111111",
  45235=>"000000000",
  45236=>"110111111",
  45237=>"111111111",
  45238=>"000001001",
  45239=>"000100111",
  45240=>"000000000",
  45241=>"000001111",
  45242=>"000000000",
  45243=>"101010110",
  45244=>"001000001",
  45245=>"001000111",
  45246=>"111111111",
  45247=>"000111111",
  45248=>"000000000",
  45249=>"111111101",
  45250=>"100111111",
  45251=>"111011000",
  45252=>"001001001",
  45253=>"000000000",
  45254=>"011011010",
  45255=>"001111101",
  45256=>"010110110",
  45257=>"001001100",
  45258=>"011111110",
  45259=>"000000000",
  45260=>"000000111",
  45261=>"000000000",
  45262=>"110110000",
  45263=>"000110111",
  45264=>"111111110",
  45265=>"101101000",
  45266=>"011011011",
  45267=>"111111111",
  45268=>"001101111",
  45269=>"110110110",
  45270=>"000000001",
  45271=>"000000101",
  45272=>"000000000",
  45273=>"101110100",
  45274=>"000000101",
  45275=>"000111111",
  45276=>"000000000",
  45277=>"001000000",
  45278=>"111111000",
  45279=>"000000000",
  45280=>"000000000",
  45281=>"010000000",
  45282=>"010011011",
  45283=>"111100011",
  45284=>"000111111",
  45285=>"111001111",
  45286=>"000000000",
  45287=>"111111000",
  45288=>"111111111",
  45289=>"000000101",
  45290=>"000000100",
  45291=>"111111000",
  45292=>"000001011",
  45293=>"100100000",
  45294=>"000000000",
  45295=>"000000000",
  45296=>"000000100",
  45297=>"011011111",
  45298=>"000011111",
  45299=>"010011011",
  45300=>"110000110",
  45301=>"111111100",
  45302=>"000011001",
  45303=>"000001011",
  45304=>"111011110",
  45305=>"000000111",
  45306=>"111101111",
  45307=>"101101000",
  45308=>"010110111",
  45309=>"111111111",
  45310=>"100010010",
  45311=>"000000111",
  45312=>"110111110",
  45313=>"001001001",
  45314=>"111111111",
  45315=>"110111111",
  45316=>"111111110",
  45317=>"110111111",
  45318=>"000000000",
  45319=>"111100000",
  45320=>"111111011",
  45321=>"000001001",
  45322=>"000111111",
  45323=>"000000001",
  45324=>"001001000",
  45325=>"000000000",
  45326=>"000000100",
  45327=>"000000011",
  45328=>"000000110",
  45329=>"011110000",
  45330=>"111101111",
  45331=>"010111111",
  45332=>"010111111",
  45333=>"011011000",
  45334=>"001100100",
  45335=>"111111100",
  45336=>"000111001",
  45337=>"101000001",
  45338=>"101111000",
  45339=>"000000110",
  45340=>"111111000",
  45341=>"111100000",
  45342=>"000000111",
  45343=>"000001001",
  45344=>"111111000",
  45345=>"111111111",
  45346=>"100100000",
  45347=>"111111011",
  45348=>"111111001",
  45349=>"000000111",
  45350=>"111111010",
  45351=>"001001001",
  45352=>"000000011",
  45353=>"111111010",
  45354=>"011011101",
  45355=>"100000000",
  45356=>"110110111",
  45357=>"000000001",
  45358=>"001000000",
  45359=>"111100010",
  45360=>"000111001",
  45361=>"111111000",
  45362=>"000000110",
  45363=>"000000000",
  45364=>"000000000",
  45365=>"111111111",
  45366=>"101011111",
  45367=>"000000000",
  45368=>"000001000",
  45369=>"101101101",
  45370=>"000000111",
  45371=>"011010000",
  45372=>"000101111",
  45373=>"111111001",
  45374=>"001111111",
  45375=>"111011100",
  45376=>"001001001",
  45377=>"111111010",
  45378=>"001001111",
  45379=>"001001111",
  45380=>"111110000",
  45381=>"110000000",
  45382=>"000000111",
  45383=>"001001111",
  45384=>"111111111",
  45385=>"111111000",
  45386=>"111111001",
  45387=>"110100000",
  45388=>"010010010",
  45389=>"000000101",
  45390=>"111111111",
  45391=>"000000111",
  45392=>"001000011",
  45393=>"001000111",
  45394=>"110000001",
  45395=>"111000000",
  45396=>"000001111",
  45397=>"011011011",
  45398=>"111111001",
  45399=>"100100000",
  45400=>"001001000",
  45401=>"111001000",
  45402=>"011000111",
  45403=>"100111000",
  45404=>"111111111",
  45405=>"000000111",
  45406=>"111111101",
  45407=>"111001000",
  45408=>"100011001",
  45409=>"111111111",
  45410=>"000111111",
  45411=>"111001000",
  45412=>"100111110",
  45413=>"000000000",
  45414=>"000011000",
  45415=>"111111100",
  45416=>"001000001",
  45417=>"111111111",
  45418=>"000000000",
  45419=>"111111000",
  45420=>"000011111",
  45421=>"011000000",
  45422=>"111110110",
  45423=>"000000001",
  45424=>"000000000",
  45425=>"000000111",
  45426=>"000000101",
  45427=>"111011011",
  45428=>"111110110",
  45429=>"101111111",
  45430=>"111101000",
  45431=>"000100101",
  45432=>"000000000",
  45433=>"111110000",
  45434=>"000000110",
  45435=>"011011011",
  45436=>"000000000",
  45437=>"111101000",
  45438=>"000000010",
  45439=>"111111111",
  45440=>"110000100",
  45441=>"000111111",
  45442=>"100110110",
  45443=>"101000000",
  45444=>"100100100",
  45445=>"111111111",
  45446=>"111001001",
  45447=>"101100111",
  45448=>"101001111",
  45449=>"000000000",
  45450=>"111111111",
  45451=>"000000000",
  45452=>"101001100",
  45453=>"001000000",
  45454=>"001001000",
  45455=>"000001011",
  45456=>"000011001",
  45457=>"111101000",
  45458=>"000111000",
  45459=>"011011111",
  45460=>"000000000",
  45461=>"010110010",
  45462=>"010111000",
  45463=>"110111100",
  45464=>"010000000",
  45465=>"000001111",
  45466=>"000000101",
  45467=>"011111111",
  45468=>"000000111",
  45469=>"000000101",
  45470=>"000000000",
  45471=>"000100000",
  45472=>"110110111",
  45473=>"111000000",
  45474=>"111111110",
  45475=>"111100100",
  45476=>"111111111",
  45477=>"000000111",
  45478=>"111111111",
  45479=>"011000000",
  45480=>"111111011",
  45481=>"101000111",
  45482=>"000000001",
  45483=>"000000000",
  45484=>"000000001",
  45485=>"100000101",
  45486=>"110000000",
  45487=>"111111111",
  45488=>"100000100",
  45489=>"010010111",
  45490=>"111110110",
  45491=>"000000111",
  45492=>"000000000",
  45493=>"100001111",
  45494=>"111111000",
  45495=>"000000101",
  45496=>"000000000",
  45497=>"000000000",
  45498=>"111110000",
  45499=>"000111111",
  45500=>"000100111",
  45501=>"111111111",
  45502=>"100100000",
  45503=>"000000100",
  45504=>"111111110",
  45505=>"011011011",
  45506=>"000001111",
  45507=>"111111111",
  45508=>"111111000",
  45509=>"000000000",
  45510=>"000100100",
  45511=>"111000001",
  45512=>"111000111",
  45513=>"100101111",
  45514=>"000101111",
  45515=>"100000000",
  45516=>"010011011",
  45517=>"001111000",
  45518=>"000001001",
  45519=>"000111111",
  45520=>"111001000",
  45521=>"011001111",
  45522=>"001001000",
  45523=>"000001011",
  45524=>"011000001",
  45525=>"000100111",
  45526=>"100111111",
  45527=>"001111111",
  45528=>"111101111",
  45529=>"000000110",
  45530=>"001000000",
  45531=>"111111111",
  45532=>"111111111",
  45533=>"000000101",
  45534=>"111111111",
  45535=>"011001001",
  45536=>"000001001",
  45537=>"000111111",
  45538=>"000000111",
  45539=>"111011111",
  45540=>"111111111",
  45541=>"111110100",
  45542=>"111101100",
  45543=>"100000100",
  45544=>"000001001",
  45545=>"111011010",
  45546=>"100000000",
  45547=>"000000000",
  45548=>"111001000",
  45549=>"000110110",
  45550=>"000000000",
  45551=>"011011001",
  45552=>"000000111",
  45553=>"000000100",
  45554=>"111111111",
  45555=>"111111111",
  45556=>"000001111",
  45557=>"100111011",
  45558=>"111111011",
  45559=>"100101011",
  45560=>"111111000",
  45561=>"001000010",
  45562=>"111001000",
  45563=>"000001001",
  45564=>"001000000",
  45565=>"111111111",
  45566=>"110111000",
  45567=>"111101111",
  45568=>"001001111",
  45569=>"111000000",
  45570=>"000000000",
  45571=>"000000111",
  45572=>"001111001",
  45573=>"101000000",
  45574=>"000010110",
  45575=>"000000000",
  45576=>"001111000",
  45577=>"110110110",
  45578=>"001001000",
  45579=>"111111111",
  45580=>"000110111",
  45581=>"100100111",
  45582=>"000100110",
  45583=>"000000000",
  45584=>"011011011",
  45585=>"000010001",
  45586=>"000000000",
  45587=>"111111111",
  45588=>"111000000",
  45589=>"111111111",
  45590=>"000000000",
  45591=>"111101100",
  45592=>"000000000",
  45593=>"000000000",
  45594=>"001001001",
  45595=>"110110111",
  45596=>"000000000",
  45597=>"111011011",
  45598=>"011011011",
  45599=>"111010111",
  45600=>"000000011",
  45601=>"111111111",
  45602=>"000000000",
  45603=>"011111111",
  45604=>"111111111",
  45605=>"001001001",
  45606=>"011111111",
  45607=>"111111110",
  45608=>"000000000",
  45609=>"001000000",
  45610=>"001111111",
  45611=>"110110111",
  45612=>"110111000",
  45613=>"111111101",
  45614=>"001000000",
  45615=>"000000000",
  45616=>"000000000",
  45617=>"000011011",
  45618=>"000110100",
  45619=>"100100000",
  45620=>"000000110",
  45621=>"111111111",
  45622=>"011000110",
  45623=>"000001001",
  45624=>"111111110",
  45625=>"000000000",
  45626=>"111111111",
  45627=>"000010000",
  45628=>"001001111",
  45629=>"101100000",
  45630=>"001100010",
  45631=>"000000010",
  45632=>"000000111",
  45633=>"100110100",
  45634=>"111111111",
  45635=>"000110111",
  45636=>"000111001",
  45637=>"111111111",
  45638=>"001000001",
  45639=>"111111111",
  45640=>"001011011",
  45641=>"011010000",
  45642=>"110000000",
  45643=>"000000000",
  45644=>"011000001",
  45645=>"110110000",
  45646=>"111000000",
  45647=>"111111111",
  45648=>"100000000",
  45649=>"000000000",
  45650=>"000000111",
  45651=>"111111111",
  45652=>"000000000",
  45653=>"111110000",
  45654=>"000011010",
  45655=>"000111111",
  45656=>"000000101",
  45657=>"000000000",
  45658=>"100000000",
  45659=>"001011001",
  45660=>"000000000",
  45661=>"000111011",
  45662=>"000010000",
  45663=>"100100100",
  45664=>"001000001",
  45665=>"001001111",
  45666=>"001110000",
  45667=>"000000000",
  45668=>"000000000",
  45669=>"000000100",
  45670=>"000010000",
  45671=>"000000000",
  45672=>"000000110",
  45673=>"111111111",
  45674=>"110110110",
  45675=>"000000000",
  45676=>"110111111",
  45677=>"000000000",
  45678=>"001111011",
  45679=>"111011011",
  45680=>"110001001",
  45681=>"000000000",
  45682=>"110110110",
  45683=>"111101110",
  45684=>"000000000",
  45685=>"111111111",
  45686=>"000111111",
  45687=>"010011011",
  45688=>"000000111",
  45689=>"000000000",
  45690=>"000000101",
  45691=>"111111111",
  45692=>"001001011",
  45693=>"110111111",
  45694=>"000000000",
  45695=>"000000000",
  45696=>"000000000",
  45697=>"000111110",
  45698=>"100000000",
  45699=>"111111111",
  45700=>"111101100",
  45701=>"111001001",
  45702=>"001001011",
  45703=>"111111110",
  45704=>"000000000",
  45705=>"010010111",
  45706=>"111110111",
  45707=>"111111111",
  45708=>"000000000",
  45709=>"000000111",
  45710=>"100110110",
  45711=>"011110000",
  45712=>"000000000",
  45713=>"001000000",
  45714=>"000000000",
  45715=>"100000000",
  45716=>"000000111",
  45717=>"001101111",
  45718=>"111110100",
  45719=>"111100000",
  45720=>"000000000",
  45721=>"111111111",
  45722=>"011000111",
  45723=>"000101000",
  45724=>"000110000",
  45725=>"100000000",
  45726=>"110111111",
  45727=>"111111111",
  45728=>"111111111",
  45729=>"111111111",
  45730=>"111111111",
  45731=>"111110110",
  45732=>"000000111",
  45733=>"001011011",
  45734=>"111001000",
  45735=>"011010111",
  45736=>"111111111",
  45737=>"000000000",
  45738=>"000110110",
  45739=>"110000000",
  45740=>"111111001",
  45741=>"000000000",
  45742=>"000100100",
  45743=>"110001000",
  45744=>"000000000",
  45745=>"001000000",
  45746=>"111111110",
  45747=>"000101111",
  45748=>"001001001",
  45749=>"000000001",
  45750=>"000000000",
  45751=>"111111111",
  45752=>"111111111",
  45753=>"000000000",
  45754=>"000000000",
  45755=>"000111111",
  45756=>"001000001",
  45757=>"000000001",
  45758=>"010000001",
  45759=>"111111111",
  45760=>"011001111",
  45761=>"111111111",
  45762=>"000001011",
  45763=>"101101111",
  45764=>"110110000",
  45765=>"001000101",
  45766=>"111111111",
  45767=>"000000000",
  45768=>"000110111",
  45769=>"111111010",
  45770=>"001000001",
  45771=>"000000000",
  45772=>"000000111",
  45773=>"000000001",
  45774=>"111111111",
  45775=>"000000000",
  45776=>"100000000",
  45777=>"111111110",
  45778=>"000000000",
  45779=>"011100000",
  45780=>"000000000",
  45781=>"011111111",
  45782=>"000000000",
  45783=>"111111111",
  45784=>"111101111",
  45785=>"011000000",
  45786=>"111000000",
  45787=>"111111100",
  45788=>"111111111",
  45789=>"000000000",
  45790=>"111011001",
  45791=>"000000000",
  45792=>"111111111",
  45793=>"111111111",
  45794=>"111000000",
  45795=>"111111111",
  45796=>"110111111",
  45797=>"000100100",
  45798=>"000000110",
  45799=>"101101101",
  45800=>"111101111",
  45801=>"111000000",
  45802=>"010111000",
  45803=>"000000100",
  45804=>"000010111",
  45805=>"111111111",
  45806=>"111111111",
  45807=>"000000000",
  45808=>"111111010",
  45809=>"111111111",
  45810=>"111001000",
  45811=>"000110100",
  45812=>"000010110",
  45813=>"111000001",
  45814=>"111100111",
  45815=>"011011111",
  45816=>"000000000",
  45817=>"111111011",
  45818=>"000000000",
  45819=>"000000000",
  45820=>"111100000",
  45821=>"000000000",
  45822=>"101001101",
  45823=>"000000000",
  45824=>"000000000",
  45825=>"100000000",
  45826=>"111111100",
  45827=>"000001001",
  45828=>"011011111",
  45829=>"111111111",
  45830=>"000000000",
  45831=>"111111110",
  45832=>"111111111",
  45833=>"000000000",
  45834=>"000000000",
  45835=>"111100100",
  45836=>"000010010",
  45837=>"101100111",
  45838=>"111111011",
  45839=>"110100000",
  45840=>"111111111",
  45841=>"001100110",
  45842=>"000000000",
  45843=>"000000000",
  45844=>"000000000",
  45845=>"000000100",
  45846=>"111111011",
  45847=>"000001111",
  45848=>"011111111",
  45849=>"111111111",
  45850=>"111111111",
  45851=>"000000000",
  45852=>"000010110",
  45853=>"111111111",
  45854=>"000000000",
  45855=>"011111111",
  45856=>"000000000",
  45857=>"111111100",
  45858=>"001000000",
  45859=>"110101111",
  45860=>"100100000",
  45861=>"000001001",
  45862=>"111111111",
  45863=>"000000000",
  45864=>"110100111",
  45865=>"000000000",
  45866=>"101101000",
  45867=>"000000000",
  45868=>"000000100",
  45869=>"011011111",
  45870=>"000111111",
  45871=>"111111111",
  45872=>"110000001",
  45873=>"111111111",
  45874=>"011000000",
  45875=>"111101000",
  45876=>"000000000",
  45877=>"111111101",
  45878=>"111111111",
  45879=>"111111111",
  45880=>"000000000",
  45881=>"000000000",
  45882=>"000000000",
  45883=>"111111110",
  45884=>"000001001",
  45885=>"000001111",
  45886=>"111111010",
  45887=>"000000101",
  45888=>"000000110",
  45889=>"010000000",
  45890=>"111111000",
  45891=>"000000000",
  45892=>"111111001",
  45893=>"000000000",
  45894=>"000000010",
  45895=>"010111111",
  45896=>"101111011",
  45897=>"000000000",
  45898=>"000000000",
  45899=>"111111111",
  45900=>"110000001",
  45901=>"111000111",
  45902=>"010010100",
  45903=>"011011011",
  45904=>"111101111",
  45905=>"100000111",
  45906=>"000000000",
  45907=>"100110101",
  45908=>"000000001",
  45909=>"011011001",
  45910=>"111111000",
  45911=>"111100111",
  45912=>"111111111",
  45913=>"111111111",
  45914=>"001001011",
  45915=>"010010100",
  45916=>"110111101",
  45917=>"110111111",
  45918=>"000000110",
  45919=>"000011011",
  45920=>"000001111",
  45921=>"111000101",
  45922=>"110100110",
  45923=>"000001001",
  45924=>"000111110",
  45925=>"000000000",
  45926=>"111111111",
  45927=>"000000001",
  45928=>"111011111",
  45929=>"111111010",
  45930=>"000000001",
  45931=>"111001000",
  45932=>"110011001",
  45933=>"110110110",
  45934=>"111001001",
  45935=>"000001000",
  45936=>"000000000",
  45937=>"001000000",
  45938=>"111011011",
  45939=>"111011011",
  45940=>"110110110",
  45941=>"000001101",
  45942=>"000000000",
  45943=>"000000000",
  45944=>"000000000",
  45945=>"111001111",
  45946=>"001000000",
  45947=>"111101101",
  45948=>"000000000",
  45949=>"011111000",
  45950=>"001000110",
  45951=>"000000000",
  45952=>"110001001",
  45953=>"111000000",
  45954=>"111111111",
  45955=>"010010000",
  45956=>"111111111",
  45957=>"000000111",
  45958=>"000000000",
  45959=>"001011111",
  45960=>"000000000",
  45961=>"000000000",
  45962=>"000000000",
  45963=>"000000000",
  45964=>"101111111",
  45965=>"001111011",
  45966=>"111111101",
  45967=>"111110000",
  45968=>"000000001",
  45969=>"111111111",
  45970=>"001001000",
  45971=>"000000000",
  45972=>"111111111",
  45973=>"000000000",
  45974=>"000000000",
  45975=>"110000100",
  45976=>"000000111",
  45977=>"000001001",
  45978=>"111100100",
  45979=>"100110100",
  45980=>"000011011",
  45981=>"000000001",
  45982=>"000110000",
  45983=>"111001001",
  45984=>"111011000",
  45985=>"111110110",
  45986=>"000001111",
  45987=>"100000111",
  45988=>"101111111",
  45989=>"111111111",
  45990=>"110110111",
  45991=>"111011000",
  45992=>"000001000",
  45993=>"000001111",
  45994=>"111111101",
  45995=>"000000000",
  45996=>"000000000",
  45997=>"011000000",
  45998=>"000000001",
  45999=>"000000010",
  46000=>"000111111",
  46001=>"000000001",
  46002=>"111110101",
  46003=>"000000000",
  46004=>"010000000",
  46005=>"010110000",
  46006=>"111111111",
  46007=>"111110110",
  46008=>"100000111",
  46009=>"111111111",
  46010=>"000001011",
  46011=>"000000111",
  46012=>"111111111",
  46013=>"111111111",
  46014=>"000000101",
  46015=>"100100000",
  46016=>"111111010",
  46017=>"000000101",
  46018=>"111000000",
  46019=>"000000000",
  46020=>"111100100",
  46021=>"111011111",
  46022=>"000000101",
  46023=>"000111011",
  46024=>"000111111",
  46025=>"111010111",
  46026=>"111111111",
  46027=>"111110000",
  46028=>"000000000",
  46029=>"101000111",
  46030=>"000000101",
  46031=>"110000000",
  46032=>"000000000",
  46033=>"000000000",
  46034=>"111111111",
  46035=>"111111100",
  46036=>"110110110",
  46037=>"111111111",
  46038=>"101100001",
  46039=>"001111101",
  46040=>"100110000",
  46041=>"110110110",
  46042=>"111111111",
  46043=>"000000111",
  46044=>"111100100",
  46045=>"000000001",
  46046=>"111111111",
  46047=>"111111011",
  46048=>"000001111",
  46049=>"000000000",
  46050=>"111111111",
  46051=>"000000000",
  46052=>"000000010",
  46053=>"000000000",
  46054=>"111111110",
  46055=>"111000111",
  46056=>"111101101",
  46057=>"111111111",
  46058=>"110100100",
  46059=>"000101001",
  46060=>"000000000",
  46061=>"111101100",
  46062=>"000000000",
  46063=>"000000110",
  46064=>"000000000",
  46065=>"111111111",
  46066=>"000101111",
  46067=>"010000000",
  46068=>"111111111",
  46069=>"000000000",
  46070=>"111111111",
  46071=>"000010011",
  46072=>"011011000",
  46073=>"011000000",
  46074=>"000110110",
  46075=>"101001101",
  46076=>"100111111",
  46077=>"100001111",
  46078=>"000000110",
  46079=>"000000000",
  46080=>"111111111",
  46081=>"000001000",
  46082=>"110000000",
  46083=>"111111111",
  46084=>"110100001",
  46085=>"000000000",
  46086=>"010111111",
  46087=>"000000000",
  46088=>"111011111",
  46089=>"111111000",
  46090=>"001000000",
  46091=>"010000000",
  46092=>"111111111",
  46093=>"011111000",
  46094=>"100100000",
  46095=>"111111111",
  46096=>"100110111",
  46097=>"000000000",
  46098=>"010011000",
  46099=>"000000101",
  46100=>"011001111",
  46101=>"000000000",
  46102=>"000111000",
  46103=>"001101100",
  46104=>"110100111",
  46105=>"100000000",
  46106=>"000000000",
  46107=>"111111101",
  46108=>"010111111",
  46109=>"111000000",
  46110=>"110100000",
  46111=>"111111111",
  46112=>"100001101",
  46113=>"000110011",
  46114=>"100001000",
  46115=>"100101000",
  46116=>"111111000",
  46117=>"110110111",
  46118=>"111111001",
  46119=>"010000000",
  46120=>"111110111",
  46121=>"010011010",
  46122=>"100111111",
  46123=>"000000001",
  46124=>"000000111",
  46125=>"001111111",
  46126=>"000100111",
  46127=>"000010111",
  46128=>"000100111",
  46129=>"000000000",
  46130=>"111110100",
  46131=>"101001001",
  46132=>"111101001",
  46133=>"111011011",
  46134=>"111001001",
  46135=>"111000000",
  46136=>"001000111",
  46137=>"010011111",
  46138=>"000100100",
  46139=>"110111111",
  46140=>"111111101",
  46141=>"111101110",
  46142=>"001111111",
  46143=>"000000000",
  46144=>"011000110",
  46145=>"000101111",
  46146=>"111000000",
  46147=>"011000110",
  46148=>"011001000",
  46149=>"000110000",
  46150=>"000000000",
  46151=>"111111111",
  46152=>"000010111",
  46153=>"000000000",
  46154=>"000000000",
  46155=>"111111111",
  46156=>"001001001",
  46157=>"111111111",
  46158=>"000000000",
  46159=>"111000111",
  46160=>"111100000",
  46161=>"111111111",
  46162=>"111111100",
  46163=>"111111000",
  46164=>"000110000",
  46165=>"000000000",
  46166=>"111100110",
  46167=>"000000000",
  46168=>"111110100",
  46169=>"000000000",
  46170=>"000011111",
  46171=>"110110011",
  46172=>"111111101",
  46173=>"000111111",
  46174=>"001000100",
  46175=>"010110111",
  46176=>"000000000",
  46177=>"000000000",
  46178=>"000000111",
  46179=>"111000000",
  46180=>"101100000",
  46181=>"000100111",
  46182=>"111111111",
  46183=>"000110000",
  46184=>"101111111",
  46185=>"111111111",
  46186=>"011000000",
  46187=>"100000111",
  46188=>"111101111",
  46189=>"111000000",
  46190=>"000000000",
  46191=>"000001000",
  46192=>"000000111",
  46193=>"101100111",
  46194=>"100100000",
  46195=>"111111111",
  46196=>"000011111",
  46197=>"001000100",
  46198=>"000111111",
  46199=>"000000000",
  46200=>"001111001",
  46201=>"000000000",
  46202=>"000100111",
  46203=>"000110000",
  46204=>"111000000",
  46205=>"010010000",
  46206=>"000000111",
  46207=>"000000000",
  46208=>"111111111",
  46209=>"000000000",
  46210=>"110000100",
  46211=>"100110010",
  46212=>"000000000",
  46213=>"010000100",
  46214=>"001011001",
  46215=>"111111000",
  46216=>"000000000",
  46217=>"011011011",
  46218=>"111100000",
  46219=>"000110111",
  46220=>"000000000",
  46221=>"000111111",
  46222=>"000011111",
  46223=>"111111110",
  46224=>"000111111",
  46225=>"111111001",
  46226=>"000001111",
  46227=>"000111111",
  46228=>"111011111",
  46229=>"100000111",
  46230=>"000000000",
  46231=>"001000000",
  46232=>"111111111",
  46233=>"000111100",
  46234=>"000110111",
  46235=>"000000111",
  46236=>"010000000",
  46237=>"000000101",
  46238=>"000000000",
  46239=>"000000111",
  46240=>"000111111",
  46241=>"111110000",
  46242=>"111111111",
  46243=>"111111111",
  46244=>"111001111",
  46245=>"000010111",
  46246=>"000000000",
  46247=>"110110000",
  46248=>"111111111",
  46249=>"100000000",
  46250=>"111000000",
  46251=>"000100000",
  46252=>"000000000",
  46253=>"110011001",
  46254=>"110111001",
  46255=>"000001001",
  46256=>"111111111",
  46257=>"000000000",
  46258=>"111111000",
  46259=>"111111000",
  46260=>"001000000",
  46261=>"010010000",
  46262=>"111001000",
  46263=>"111011000",
  46264=>"100000000",
  46265=>"000000000",
  46266=>"111001001",
  46267=>"111000011",
  46268=>"010010111",
  46269=>"111011000",
  46270=>"000001111",
  46271=>"001111111",
  46272=>"111100000",
  46273=>"111000000",
  46274=>"000000111",
  46275=>"000000000",
  46276=>"111111011",
  46277=>"000000000",
  46278=>"000000000",
  46279=>"011011001",
  46280=>"001011011",
  46281=>"000000010",
  46282=>"111100111",
  46283=>"011011000",
  46284=>"000010000",
  46285=>"101000001",
  46286=>"000111111",
  46287=>"000000100",
  46288=>"000000000",
  46289=>"000011001",
  46290=>"111111111",
  46291=>"011011010",
  46292=>"111101000",
  46293=>"111111111",
  46294=>"010000000",
  46295=>"111101000",
  46296=>"111000000",
  46297=>"111111111",
  46298=>"000000000",
  46299=>"000000000",
  46300=>"000000000",
  46301=>"111000001",
  46302=>"001111111",
  46303=>"111000001",
  46304=>"101111111",
  46305=>"000000111",
  46306=>"111000110",
  46307=>"111111111",
  46308=>"001001000",
  46309=>"011001100",
  46310=>"111001000",
  46311=>"000000000",
  46312=>"111111111",
  46313=>"011000001",
  46314=>"111100000",
  46315=>"111111100",
  46316=>"101111101",
  46317=>"100000001",
  46318=>"111111001",
  46319=>"111011000",
  46320=>"011111111",
  46321=>"110011011",
  46322=>"111111000",
  46323=>"111001101",
  46324=>"010010110",
  46325=>"000000110",
  46326=>"000000000",
  46327=>"111110000",
  46328=>"100101111",
  46329=>"000000110",
  46330=>"001000110",
  46331=>"000000000",
  46332=>"000010111",
  46333=>"001001111",
  46334=>"000000000",
  46335=>"001111111",
  46336=>"100000000",
  46337=>"100111000",
  46338=>"100000001",
  46339=>"000000000",
  46340=>"100100100",
  46341=>"001000000",
  46342=>"000000001",
  46343=>"101000000",
  46344=>"000111111",
  46345=>"111111000",
  46346=>"111111111",
  46347=>"001111000",
  46348=>"111001001",
  46349=>"000001111",
  46350=>"000100000",
  46351=>"000000000",
  46352=>"010111111",
  46353=>"111111000",
  46354=>"111000001",
  46355=>"010000000",
  46356=>"111111000",
  46357=>"111011111",
  46358=>"000100011",
  46359=>"100000100",
  46360=>"100111100",
  46361=>"000000000",
  46362=>"000000000",
  46363=>"111111000",
  46364=>"100111001",
  46365=>"000000000",
  46366=>"000000000",
  46367=>"111101000",
  46368=>"111111000",
  46369=>"111000001",
  46370=>"000000000",
  46371=>"101111111",
  46372=>"111111111",
  46373=>"111111101",
  46374=>"111001001",
  46375=>"111100100",
  46376=>"111000000",
  46377=>"000000100",
  46378=>"111111111",
  46379=>"111011011",
  46380=>"110010000",
  46381=>"111111111",
  46382=>"000000000",
  46383=>"011000000",
  46384=>"000110110",
  46385=>"000000000",
  46386=>"111000000",
  46387=>"110000000",
  46388=>"000000000",
  46389=>"001000000",
  46390=>"000000111",
  46391=>"000111000",
  46392=>"111000000",
  46393=>"000000111",
  46394=>"010000111",
  46395=>"111111111",
  46396=>"101101100",
  46397=>"011010000",
  46398=>"011000110",
  46399=>"000000000",
  46400=>"111111000",
  46401=>"111011011",
  46402=>"001100110",
  46403=>"000101000",
  46404=>"000000000",
  46405=>"111111111",
  46406=>"111000000",
  46407=>"000001111",
  46408=>"000000110",
  46409=>"000111000",
  46410=>"011001000",
  46411=>"001000100",
  46412=>"111000000",
  46413=>"001000000",
  46414=>"111111101",
  46415=>"011110100",
  46416=>"011011110",
  46417=>"000000111",
  46418=>"111111000",
  46419=>"000001000",
  46420=>"000000000",
  46421=>"111111000",
  46422=>"100000011",
  46423=>"101000000",
  46424=>"000000001",
  46425=>"000111111",
  46426=>"000000000",
  46427=>"001001111",
  46428=>"000001111",
  46429=>"111111101",
  46430=>"110000000",
  46431=>"000000111",
  46432=>"110110010",
  46433=>"110100000",
  46434=>"110000000",
  46435=>"000000111",
  46436=>"001001000",
  46437=>"000000000",
  46438=>"111111111",
  46439=>"111111011",
  46440=>"110000001",
  46441=>"111000111",
  46442=>"000000000",
  46443=>"000000001",
  46444=>"011011000",
  46445=>"100000000",
  46446=>"010000000",
  46447=>"000000000",
  46448=>"000001000",
  46449=>"010000000",
  46450=>"000111111",
  46451=>"110110110",
  46452=>"111000111",
  46453=>"100110111",
  46454=>"111100111",
  46455=>"111010000",
  46456=>"000001111",
  46457=>"111110111",
  46458=>"010001000",
  46459=>"000000000",
  46460=>"101001111",
  46461=>"011001000",
  46462=>"100101111",
  46463=>"000000000",
  46464=>"111111111",
  46465=>"001001111",
  46466=>"010111111",
  46467=>"000000001",
  46468=>"000111111",
  46469=>"000000000",
  46470=>"000000000",
  46471=>"000000000",
  46472=>"000000000",
  46473=>"100100100",
  46474=>"000000110",
  46475=>"000000000",
  46476=>"000011110",
  46477=>"110100000",
  46478=>"111111111",
  46479=>"111001001",
  46480=>"000000000",
  46481=>"000001011",
  46482=>"100100000",
  46483=>"000100000",
  46484=>"000111111",
  46485=>"010010010",
  46486=>"111001111",
  46487=>"111001001",
  46488=>"000111111",
  46489=>"000000000",
  46490=>"001011111",
  46491=>"110100000",
  46492=>"010111111",
  46493=>"111111111",
  46494=>"010000000",
  46495=>"111000100",
  46496=>"011000011",
  46497=>"110111111",
  46498=>"111000000",
  46499=>"111111111",
  46500=>"100110111",
  46501=>"000000000",
  46502=>"001000000",
  46503=>"001111001",
  46504=>"000110100",
  46505=>"000000000",
  46506=>"111100111",
  46507=>"111000000",
  46508=>"000000000",
  46509=>"000000000",
  46510=>"111010110",
  46511=>"000000000",
  46512=>"000011111",
  46513=>"000111111",
  46514=>"111111000",
  46515=>"110111111",
  46516=>"000001111",
  46517=>"001001000",
  46518=>"000101111",
  46519=>"000010001",
  46520=>"000000011",
  46521=>"010011111",
  46522=>"111000100",
  46523=>"110110000",
  46524=>"111000011",
  46525=>"011111111",
  46526=>"111111000",
  46527=>"110011111",
  46528=>"111111111",
  46529=>"000101111",
  46530=>"000000000",
  46531=>"000001111",
  46532=>"101101000",
  46533=>"110110100",
  46534=>"001001101",
  46535=>"111111000",
  46536=>"110100111",
  46537=>"000000000",
  46538=>"011011000",
  46539=>"000000100",
  46540=>"011000000",
  46541=>"000000000",
  46542=>"000000000",
  46543=>"000000000",
  46544=>"000111000",
  46545=>"111000110",
  46546=>"000001001",
  46547=>"111000111",
  46548=>"000110110",
  46549=>"000100111",
  46550=>"111111111",
  46551=>"111101110",
  46552=>"111000000",
  46553=>"000111000",
  46554=>"000000000",
  46555=>"011000000",
  46556=>"111111010",
  46557=>"000000101",
  46558=>"111111111",
  46559=>"010001011",
  46560=>"000110000",
  46561=>"111000000",
  46562=>"111111100",
  46563=>"111111000",
  46564=>"111111111",
  46565=>"000000110",
  46566=>"111101111",
  46567=>"010000000",
  46568=>"000111111",
  46569=>"111111110",
  46570=>"000000000",
  46571=>"111111000",
  46572=>"111111111",
  46573=>"110100100",
  46574=>"000000000",
  46575=>"111000001",
  46576=>"010010010",
  46577=>"011000000",
  46578=>"011010111",
  46579=>"111101001",
  46580=>"000000000",
  46581=>"111110000",
  46582=>"100111000",
  46583=>"111110110",
  46584=>"100000000",
  46585=>"011000000",
  46586=>"000001000",
  46587=>"000000000",
  46588=>"110011111",
  46589=>"101110111",
  46590=>"111111101",
  46591=>"110110000",
  46592=>"000000100",
  46593=>"000000000",
  46594=>"000000001",
  46595=>"111111111",
  46596=>"111111111",
  46597=>"001000000",
  46598=>"000000011",
  46599=>"000000000",
  46600=>"000000000",
  46601=>"000100111",
  46602=>"001001111",
  46603=>"000000111",
  46604=>"000000110",
  46605=>"111110011",
  46606=>"000000000",
  46607=>"000011011",
  46608=>"110100100",
  46609=>"010011111",
  46610=>"011000000",
  46611=>"000000000",
  46612=>"001001001",
  46613=>"011111111",
  46614=>"101100000",
  46615=>"000000000",
  46616=>"000000111",
  46617=>"000000101",
  46618=>"111111101",
  46619=>"001000000",
  46620=>"111111111",
  46621=>"111110000",
  46622=>"000011011",
  46623=>"100100000",
  46624=>"000000100",
  46625=>"111000001",
  46626=>"111111111",
  46627=>"001101101",
  46628=>"111111100",
  46629=>"000101111",
  46630=>"000000000",
  46631=>"011001011",
  46632=>"001000001",
  46633=>"101101111",
  46634=>"111111111",
  46635=>"000000111",
  46636=>"111111111",
  46637=>"101100000",
  46638=>"110000000",
  46639=>"000000000",
  46640=>"001001111",
  46641=>"111111111",
  46642=>"111100110",
  46643=>"000000000",
  46644=>"000000011",
  46645=>"000110110",
  46646=>"000000000",
  46647=>"111111111",
  46648=>"111111111",
  46649=>"001111000",
  46650=>"110110111",
  46651=>"111111111",
  46652=>"000000000",
  46653=>"000000111",
  46654=>"000000000",
  46655=>"111001101",
  46656=>"110011001",
  46657=>"000101111",
  46658=>"000000100",
  46659=>"011111101",
  46660=>"000110110",
  46661=>"111110000",
  46662=>"011001000",
  46663=>"000000000",
  46664=>"110011111",
  46665=>"000000001",
  46666=>"010111111",
  46667=>"110110000",
  46668=>"000110111",
  46669=>"000000000",
  46670=>"000011000",
  46671=>"000000000",
  46672=>"110111111",
  46673=>"000000101",
  46674=>"000010011",
  46675=>"000001111",
  46676=>"000000000",
  46677=>"110000010",
  46678=>"001011111",
  46679=>"000000111",
  46680=>"000000000",
  46681=>"111111111",
  46682=>"111111111",
  46683=>"000010000",
  46684=>"000000000",
  46685=>"000000010",
  46686=>"111011111",
  46687=>"000000001",
  46688=>"100101111",
  46689=>"000000000",
  46690=>"111001001",
  46691=>"000101111",
  46692=>"000100111",
  46693=>"001001000",
  46694=>"000110000",
  46695=>"000111111",
  46696=>"001001011",
  46697=>"000000001",
  46698=>"000000111",
  46699=>"111111111",
  46700=>"000000001",
  46701=>"100000000",
  46702=>"010010000",
  46703=>"111111111",
  46704=>"111111111",
  46705=>"111101111",
  46706=>"000000111",
  46707=>"000011001",
  46708=>"111111111",
  46709=>"000001000",
  46710=>"100100000",
  46711=>"000000000",
  46712=>"111011101",
  46713=>"111111111",
  46714=>"111111111",
  46715=>"010000000",
  46716=>"000110111",
  46717=>"000000010",
  46718=>"100100111",
  46719=>"001011011",
  46720=>"001011011",
  46721=>"000000000",
  46722=>"100111110",
  46723=>"000000111",
  46724=>"010010010",
  46725=>"111111111",
  46726=>"001001110",
  46727=>"111111010",
  46728=>"000000000",
  46729=>"000000000",
  46730=>"011011111",
  46731=>"110000000",
  46732=>"111001100",
  46733=>"000000000",
  46734=>"000000100",
  46735=>"000000111",
  46736=>"111111000",
  46737=>"111111111",
  46738=>"100000000",
  46739=>"111110000",
  46740=>"000111111",
  46741=>"110000000",
  46742=>"111111100",
  46743=>"011000000",
  46744=>"000011111",
  46745=>"000000000",
  46746=>"000000010",
  46747=>"000000000",
  46748=>"100000000",
  46749=>"000000001",
  46750=>"000000101",
  46751=>"001111111",
  46752=>"111111111",
  46753=>"111111101",
  46754=>"111111111",
  46755=>"110001011",
  46756=>"001000101",
  46757=>"100100100",
  46758=>"111110001",
  46759=>"001001011",
  46760=>"111111111",
  46761=>"111111111",
  46762=>"000001011",
  46763=>"111111110",
  46764=>"111111111",
  46765=>"010011111",
  46766=>"000000101",
  46767=>"000011000",
  46768=>"110111111",
  46769=>"000000001",
  46770=>"010110010",
  46771=>"111111101",
  46772=>"111111000",
  46773=>"000000000",
  46774=>"011010111",
  46775=>"101001000",
  46776=>"000000000",
  46777=>"001000101",
  46778=>"001001011",
  46779=>"111101000",
  46780=>"110111111",
  46781=>"101001001",
  46782=>"111110111",
  46783=>"101101101",
  46784=>"000011000",
  46785=>"010000100",
  46786=>"000000000",
  46787=>"111011000",
  46788=>"000000000",
  46789=>"111111111",
  46790=>"110110000",
  46791=>"000011000",
  46792=>"001000000",
  46793=>"000000000",
  46794=>"000010110",
  46795=>"010011011",
  46796=>"011011010",
  46797=>"001111111",
  46798=>"010100110",
  46799=>"111111111",
  46800=>"000000100",
  46801=>"000000000",
  46802=>"111000001",
  46803=>"000011000",
  46804=>"111000000",
  46805=>"000000000",
  46806=>"101101000",
  46807=>"000000000",
  46808=>"011011100",
  46809=>"010000100",
  46810=>"000010010",
  46811=>"011111011",
  46812=>"000000111",
  46813=>"111100100",
  46814=>"111111111",
  46815=>"000000111",
  46816=>"111111111",
  46817=>"000111111",
  46818=>"110000111",
  46819=>"111111111",
  46820=>"111111111",
  46821=>"000000000",
  46822=>"000000000",
  46823=>"100100111",
  46824=>"111000000",
  46825=>"100100111",
  46826=>"111011001",
  46827=>"111111000",
  46828=>"000000000",
  46829=>"011000000",
  46830=>"101111111",
  46831=>"000000111",
  46832=>"011111111",
  46833=>"111111111",
  46834=>"001111111",
  46835=>"010000100",
  46836=>"010000011",
  46837=>"000000111",
  46838=>"111111000",
  46839=>"110111010",
  46840=>"000000000",
  46841=>"000000000",
  46842=>"111011001",
  46843=>"101111111",
  46844=>"010010110",
  46845=>"100000001",
  46846=>"000001000",
  46847=>"000001111",
  46848=>"001011001",
  46849=>"110100000",
  46850=>"111111111",
  46851=>"111111111",
  46852=>"000000100",
  46853=>"000000000",
  46854=>"001000000",
  46855=>"111111101",
  46856=>"000000010",
  46857=>"000000000",
  46858=>"111011001",
  46859=>"000110111",
  46860=>"111011000",
  46861=>"110010000",
  46862=>"000000000",
  46863=>"111111111",
  46864=>"111111111",
  46865=>"110000000",
  46866=>"111111111",
  46867=>"111111111",
  46868=>"011000111",
  46869=>"000000000",
  46870=>"100000110",
  46871=>"010010001",
  46872=>"111111111",
  46873=>"110000000",
  46874=>"000000010",
  46875=>"111000100",
  46876=>"000000011",
  46877=>"000000111",
  46878=>"111111111",
  46879=>"011011111",
  46880=>"000000110",
  46881=>"101111111",
  46882=>"111111000",
  46883=>"111010000",
  46884=>"011111111",
  46885=>"011001011",
  46886=>"011010011",
  46887=>"000000000",
  46888=>"000000000",
  46889=>"011111000",
  46890=>"111101101",
  46891=>"111000111",
  46892=>"000000000",
  46893=>"000000100",
  46894=>"111111110",
  46895=>"000011011",
  46896=>"111111101",
  46897=>"111111111",
  46898=>"110110111",
  46899=>"000000000",
  46900=>"000000111",
  46901=>"000000001",
  46902=>"111000000",
  46903=>"000000111",
  46904=>"000100110",
  46905=>"101000000",
  46906=>"111111111",
  46907=>"111111111",
  46908=>"011011111",
  46909=>"010010100",
  46910=>"000000000",
  46911=>"000100111",
  46912=>"111100100",
  46913=>"000000000",
  46914=>"000100000",
  46915=>"111100111",
  46916=>"111111111",
  46917=>"000000000",
  46918=>"110011011",
  46919=>"000000000",
  46920=>"111111010",
  46921=>"010011011",
  46922=>"000000000",
  46923=>"111101101",
  46924=>"111000010",
  46925=>"010000111",
  46926=>"110111100",
  46927=>"001001000",
  46928=>"100110000",
  46929=>"000000111",
  46930=>"111111111",
  46931=>"000000000",
  46932=>"000000011",
  46933=>"001001001",
  46934=>"001000000",
  46935=>"000011001",
  46936=>"111111111",
  46937=>"100100101",
  46938=>"111111111",
  46939=>"000000110",
  46940=>"100111111",
  46941=>"000000111",
  46942=>"000000000",
  46943=>"100000000",
  46944=>"111111111",
  46945=>"111111111",
  46946=>"111111111",
  46947=>"111111111",
  46948=>"000010010",
  46949=>"000000000",
  46950=>"111010000",
  46951=>"000000000",
  46952=>"110101001",
  46953=>"100111111",
  46954=>"000000100",
  46955=>"111001001",
  46956=>"000000000",
  46957=>"001000011",
  46958=>"001001001",
  46959=>"111111110",
  46960=>"000000000",
  46961=>"111111110",
  46962=>"011011000",
  46963=>"111111111",
  46964=>"111111111",
  46965=>"101000100",
  46966=>"100100000",
  46967=>"000000000",
  46968=>"111111111",
  46969=>"111110011",
  46970=>"000111111",
  46971=>"100000111",
  46972=>"000100111",
  46973=>"110000000",
  46974=>"000000111",
  46975=>"111111011",
  46976=>"001001111",
  46977=>"111111101",
  46978=>"000011011",
  46979=>"000100100",
  46980=>"000000000",
  46981=>"001001101",
  46982=>"000100100",
  46983=>"000000000",
  46984=>"000000000",
  46985=>"000000100",
  46986=>"101001001",
  46987=>"111001000",
  46988=>"011000111",
  46989=>"010011000",
  46990=>"011011110",
  46991=>"000000000",
  46992=>"000010000",
  46993=>"111111111",
  46994=>"111111010",
  46995=>"111011011",
  46996=>"000000000",
  46997=>"000000111",
  46998=>"111101011",
  46999=>"000100000",
  47000=>"111111001",
  47001=>"111100101",
  47002=>"100111111",
  47003=>"000000100",
  47004=>"111111111",
  47005=>"111001001",
  47006=>"101001001",
  47007=>"111111111",
  47008=>"011111001",
  47009=>"000100110",
  47010=>"000011001",
  47011=>"001000000",
  47012=>"110110111",
  47013=>"101111111",
  47014=>"111111111",
  47015=>"000000000",
  47016=>"100010001",
  47017=>"000000111",
  47018=>"000000010",
  47019=>"111111111",
  47020=>"000000000",
  47021=>"111111000",
  47022=>"000000000",
  47023=>"000000110",
  47024=>"111000000",
  47025=>"111111111",
  47026=>"001000111",
  47027=>"000111111",
  47028=>"111111111",
  47029=>"000000000",
  47030=>"111111111",
  47031=>"110110000",
  47032=>"111111111",
  47033=>"111110010",
  47034=>"000000000",
  47035=>"011000011",
  47036=>"111111111",
  47037=>"000000100",
  47038=>"111011111",
  47039=>"110000110",
  47040=>"011111100",
  47041=>"000000000",
  47042=>"000000000",
  47043=>"111011010",
  47044=>"111111001",
  47045=>"011110110",
  47046=>"001111000",
  47047=>"000000000",
  47048=>"000000000",
  47049=>"011001110",
  47050=>"000000000",
  47051=>"000000001",
  47052=>"010000000",
  47053=>"000000101",
  47054=>"111111111",
  47055=>"101101000",
  47056=>"111111111",
  47057=>"010000000",
  47058=>"100100001",
  47059=>"111111111",
  47060=>"100100000",
  47061=>"111101000",
  47062=>"000000111",
  47063=>"000100100",
  47064=>"000010111",
  47065=>"100100110",
  47066=>"011100000",
  47067=>"011000000",
  47068=>"000000011",
  47069=>"111101111",
  47070=>"000100100",
  47071=>"000000000",
  47072=>"111111111",
  47073=>"000000000",
  47074=>"111001000",
  47075=>"011011000",
  47076=>"111011111",
  47077=>"001001001",
  47078=>"010011100",
  47079=>"000000000",
  47080=>"011010000",
  47081=>"000000000",
  47082=>"011011111",
  47083=>"001111111",
  47084=>"111111001",
  47085=>"000001011",
  47086=>"111111111",
  47087=>"001011111",
  47088=>"000000011",
  47089=>"111110110",
  47090=>"111111111",
  47091=>"001001001",
  47092=>"000111111",
  47093=>"000000000",
  47094=>"000001001",
  47095=>"010110000",
  47096=>"101000000",
  47097=>"000000111",
  47098=>"110110010",
  47099=>"000000000",
  47100=>"000000001",
  47101=>"110111100",
  47102=>"000011100",
  47103=>"111011001",
  47104=>"111111010",
  47105=>"111110110",
  47106=>"010111111",
  47107=>"000111111",
  47108=>"111111111",
  47109=>"001001000",
  47110=>"001001001",
  47111=>"000000110",
  47112=>"111111111",
  47113=>"100101101",
  47114=>"111111000",
  47115=>"011111111",
  47116=>"000110111",
  47117=>"000010111",
  47118=>"111111111",
  47119=>"111111111",
  47120=>"110100110",
  47121=>"111111111",
  47122=>"000000110",
  47123=>"011001001",
  47124=>"000000111",
  47125=>"000000000",
  47126=>"110111111",
  47127=>"001000100",
  47128=>"110111111",
  47129=>"011011011",
  47130=>"010011111",
  47131=>"111100100",
  47132=>"111101111",
  47133=>"111111111",
  47134=>"111111111",
  47135=>"111111111",
  47136=>"110110010",
  47137=>"100000010",
  47138=>"111111111",
  47139=>"111011011",
  47140=>"001000001",
  47141=>"010111001",
  47142=>"111111111",
  47143=>"000000000",
  47144=>"000000000",
  47145=>"000000110",
  47146=>"100100100",
  47147=>"000000000",
  47148=>"100100000",
  47149=>"000111110",
  47150=>"000000000",
  47151=>"000000000",
  47152=>"000000111",
  47153=>"001111111",
  47154=>"110110111",
  47155=>"010111011",
  47156=>"000000000",
  47157=>"011011111",
  47158=>"000000000",
  47159=>"011110010",
  47160=>"000000100",
  47161=>"010110100",
  47162=>"001000001",
  47163=>"000000000",
  47164=>"110000000",
  47165=>"011000000",
  47166=>"110110000",
  47167=>"000111111",
  47168=>"001111111",
  47169=>"111111011",
  47170=>"001111001",
  47171=>"000011111",
  47172=>"001001001",
  47173=>"000000000",
  47174=>"111111110",
  47175=>"000000000",
  47176=>"000000000",
  47177=>"000000001",
  47178=>"000001001",
  47179=>"111000000",
  47180=>"011011111",
  47181=>"011000001",
  47182=>"111101101",
  47183=>"111111111",
  47184=>"111000000",
  47185=>"000000000",
  47186=>"000001000",
  47187=>"000000011",
  47188=>"000000000",
  47189=>"110111111",
  47190=>"111111011",
  47191=>"000000000",
  47192=>"111111000",
  47193=>"000000000",
  47194=>"110110000",
  47195=>"000000111",
  47196=>"111100000",
  47197=>"000000000",
  47198=>"001011111",
  47199=>"110111001",
  47200=>"000000000",
  47201=>"001001001",
  47202=>"001000000",
  47203=>"010010000",
  47204=>"001000000",
  47205=>"101111111",
  47206=>"110111111",
  47207=>"000000000",
  47208=>"010110000",
  47209=>"000111000",
  47210=>"000000000",
  47211=>"100111111",
  47212=>"000000000",
  47213=>"100100000",
  47214=>"000000000",
  47215=>"100100000",
  47216=>"110110111",
  47217=>"111111111",
  47218=>"101101101",
  47219=>"000000000",
  47220=>"001001000",
  47221=>"000000000",
  47222=>"100100000",
  47223=>"000000000",
  47224=>"110110110",
  47225=>"001001101",
  47226=>"000000000",
  47227=>"111111111",
  47228=>"000010000",
  47229=>"011111111",
  47230=>"111111000",
  47231=>"111111110",
  47232=>"111110100",
  47233=>"010111111",
  47234=>"100110100",
  47235=>"111101001",
  47236=>"110111011",
  47237=>"111111110",
  47238=>"000001110",
  47239=>"111111110",
  47240=>"000000001",
  47241=>"000000000",
  47242=>"111111111",
  47243=>"111111111",
  47244=>"011111111",
  47245=>"000000000",
  47246=>"000001111",
  47247=>"111111111",
  47248=>"000000000",
  47249=>"111111111",
  47250=>"000000000",
  47251=>"011111010",
  47252=>"000010010",
  47253=>"110110111",
  47254=>"000110000",
  47255=>"000000000",
  47256=>"110000011",
  47257=>"000001001",
  47258=>"111000001",
  47259=>"111111111",
  47260=>"111111011",
  47261=>"111111111",
  47262=>"000111111",
  47263=>"000000000",
  47264=>"000000010",
  47265=>"011001000",
  47266=>"011000000",
  47267=>"110111011",
  47268=>"000000000",
  47269=>"011111011",
  47270=>"010110010",
  47271=>"111110110",
  47272=>"000100110",
  47273=>"000100100",
  47274=>"111111111",
  47275=>"000000000",
  47276=>"000000000",
  47277=>"000011111",
  47278=>"110111111",
  47279=>"001011010",
  47280=>"110110100",
  47281=>"111111111",
  47282=>"000000010",
  47283=>"000000000",
  47284=>"111111111",
  47285=>"000110110",
  47286=>"000000111",
  47287=>"011011011",
  47288=>"000000100",
  47289=>"100111111",
  47290=>"000111111",
  47291=>"000000011",
  47292=>"111111111",
  47293=>"111111000",
  47294=>"000110111",
  47295=>"000000101",
  47296=>"111111010",
  47297=>"111110000",
  47298=>"111111111",
  47299=>"000000111",
  47300=>"111111111",
  47301=>"111111111",
  47302=>"000001000",
  47303=>"111111110",
  47304=>"111000100",
  47305=>"101000001",
  47306=>"111011011",
  47307=>"011011011",
  47308=>"010111000",
  47309=>"111110000",
  47310=>"000000001",
  47311=>"000000111",
  47312=>"110111111",
  47313=>"110110111",
  47314=>"111011000",
  47315=>"101001111",
  47316=>"000000000",
  47317=>"000000000",
  47318=>"000000000",
  47319=>"000000000",
  47320=>"000000000",
  47321=>"110111011",
  47322=>"000000000",
  47323=>"111110011",
  47324=>"010111111",
  47325=>"000111111",
  47326=>"111111111",
  47327=>"110000110",
  47328=>"000000000",
  47329=>"000000000",
  47330=>"000100110",
  47331=>"000000000",
  47332=>"111011111",
  47333=>"111110111",
  47334=>"000000011",
  47335=>"100111111",
  47336=>"100100000",
  47337=>"001001000",
  47338=>"000010011",
  47339=>"111111111",
  47340=>"111101100",
  47341=>"000000000",
  47342=>"000000000",
  47343=>"110110000",
  47344=>"111110100",
  47345=>"011010000",
  47346=>"111111111",
  47347=>"101000001",
  47348=>"000111111",
  47349=>"100000000",
  47350=>"100100110",
  47351=>"100111000",
  47352=>"010110011",
  47353=>"110111101",
  47354=>"011111001",
  47355=>"110100000",
  47356=>"100110111",
  47357=>"000000000",
  47358=>"111111100",
  47359=>"111111111",
  47360=>"011011011",
  47361=>"100100100",
  47362=>"000000000",
  47363=>"010100100",
  47364=>"110100100",
  47365=>"100100111",
  47366=>"111111010",
  47367=>"110000001",
  47368=>"000000000",
  47369=>"000000111",
  47370=>"111011000",
  47371=>"111111100",
  47372=>"110110110",
  47373=>"000100100",
  47374=>"100010000",
  47375=>"000100100",
  47376=>"000010010",
  47377=>"000011011",
  47378=>"011000000",
  47379=>"000100000",
  47380=>"011001011",
  47381=>"000100100",
  47382=>"000100000",
  47383=>"100111111",
  47384=>"110010010",
  47385=>"000000001",
  47386=>"111111111",
  47387=>"111111111",
  47388=>"001001111",
  47389=>"000000111",
  47390=>"110111111",
  47391=>"111111111",
  47392=>"000000000",
  47393=>"000000110",
  47394=>"000000110",
  47395=>"000011111",
  47396=>"000000110",
  47397=>"100000001",
  47398=>"110111100",
  47399=>"000000000",
  47400=>"111111100",
  47401=>"000000001",
  47402=>"111111111",
  47403=>"000101101",
  47404=>"100000111",
  47405=>"000011111",
  47406=>"110110111",
  47407=>"000000100",
  47408=>"000011111",
  47409=>"111111000",
  47410=>"111111111",
  47411=>"010110111",
  47412=>"111111011",
  47413=>"000110111",
  47414=>"011111100",
  47415=>"100110100",
  47416=>"000000110",
  47417=>"000000000",
  47418=>"000000000",
  47419=>"001111111",
  47420=>"110110100",
  47421=>"000000000",
  47422=>"000000000",
  47423=>"010010001",
  47424=>"000000000",
  47425=>"111111111",
  47426=>"111111111",
  47427=>"110010110",
  47428=>"000000110",
  47429=>"111100100",
  47430=>"100000000",
  47431=>"010001011",
  47432=>"111111000",
  47433=>"111000000",
  47434=>"000000100",
  47435=>"000000001",
  47436=>"110111000",
  47437=>"010111111",
  47438=>"111110111",
  47439=>"001001001",
  47440=>"101100000",
  47441=>"000000000",
  47442=>"111101111",
  47443=>"111111111",
  47444=>"000000100",
  47445=>"110111011",
  47446=>"011111111",
  47447=>"111101001",
  47448=>"111111111",
  47449=>"111111011",
  47450=>"001000100",
  47451=>"000000000",
  47452=>"010010011",
  47453=>"000000000",
  47454=>"000000011",
  47455=>"001001001",
  47456=>"111111010",
  47457=>"000000000",
  47458=>"111111111",
  47459=>"110100111",
  47460=>"000000011",
  47461=>"000000000",
  47462=>"101111000",
  47463=>"111011001",
  47464=>"000100100",
  47465=>"100100100",
  47466=>"110110110",
  47467=>"111111111",
  47468=>"000000000",
  47469=>"000001001",
  47470=>"001111111",
  47471=>"111110000",
  47472=>"111101110",
  47473=>"000000000",
  47474=>"111111111",
  47475=>"011111111",
  47476=>"101001001",
  47477=>"111111111",
  47478=>"000111110",
  47479=>"000000000",
  47480=>"111000000",
  47481=>"000000110",
  47482=>"011001011",
  47483=>"011111111",
  47484=>"000000000",
  47485=>"000000111",
  47486=>"011011011",
  47487=>"000000000",
  47488=>"100100101",
  47489=>"000000010",
  47490=>"000000000",
  47491=>"111001011",
  47492=>"111111111",
  47493=>"011010000",
  47494=>"000000110",
  47495=>"000100001",
  47496=>"000000000",
  47497=>"011011111",
  47498=>"111111111",
  47499=>"000001001",
  47500=>"111111111",
  47501=>"000000000",
  47502=>"000110010",
  47503=>"111111100",
  47504=>"110110000",
  47505=>"110111111",
  47506=>"001011000",
  47507=>"111110110",
  47508=>"000000000",
  47509=>"000010010",
  47510=>"000011001",
  47511=>"000000000",
  47512=>"111111111",
  47513=>"111000100",
  47514=>"001000000",
  47515=>"000000110",
  47516=>"000100111",
  47517=>"111111111",
  47518=>"000010010",
  47519=>"000000000",
  47520=>"111011011",
  47521=>"111110110",
  47522=>"001011011",
  47523=>"111111111",
  47524=>"011111111",
  47525=>"111011111",
  47526=>"000000001",
  47527=>"111100111",
  47528=>"000000000",
  47529=>"000000000",
  47530=>"000110111",
  47531=>"000000000",
  47532=>"111111111",
  47533=>"100100100",
  47534=>"011000111",
  47535=>"000000000",
  47536=>"000000000",
  47537=>"000000000",
  47538=>"011001001",
  47539=>"111111111",
  47540=>"000000000",
  47541=>"000000000",
  47542=>"000000100",
  47543=>"000000111",
  47544=>"111111111",
  47545=>"111111111",
  47546=>"000000000",
  47547=>"000000000",
  47548=>"000000000",
  47549=>"111111111",
  47550=>"001000000",
  47551=>"000000000",
  47552=>"000000000",
  47553=>"111110111",
  47554=>"111111111",
  47555=>"001111111",
  47556=>"000000000",
  47557=>"001000110",
  47558=>"000010110",
  47559=>"000000000",
  47560=>"000000000",
  47561=>"000000000",
  47562=>"000000001",
  47563=>"000000111",
  47564=>"010110110",
  47565=>"111111000",
  47566=>"100111110",
  47567=>"111111111",
  47568=>"000000000",
  47569=>"000001000",
  47570=>"111011111",
  47571=>"111111110",
  47572=>"110111111",
  47573=>"110110000",
  47574=>"011111111",
  47575=>"100000011",
  47576=>"000000111",
  47577=>"111001011",
  47578=>"000000111",
  47579=>"000000010",
  47580=>"011111110",
  47581=>"011011011",
  47582=>"111111111",
  47583=>"111011000",
  47584=>"000000000",
  47585=>"111111101",
  47586=>"001001001",
  47587=>"000000000",
  47588=>"110110010",
  47589=>"110110110",
  47590=>"000000000",
  47591=>"000000000",
  47592=>"000000000",
  47593=>"111111111",
  47594=>"111111111",
  47595=>"000001101",
  47596=>"000000001",
  47597=>"000000000",
  47598=>"111111111",
  47599=>"111111111",
  47600=>"000000000",
  47601=>"000111111",
  47602=>"110111000",
  47603=>"000000000",
  47604=>"000000000",
  47605=>"111110000",
  47606=>"110110000",
  47607=>"111111111",
  47608=>"100100000",
  47609=>"000000000",
  47610=>"110000000",
  47611=>"000000000",
  47612=>"000000000",
  47613=>"111110101",
  47614=>"111111111",
  47615=>"010111111",
  47616=>"101111000",
  47617=>"111100111",
  47618=>"101000111",
  47619=>"111111111",
  47620=>"101101000",
  47621=>"111100001",
  47622=>"000000100",
  47623=>"000000000",
  47624=>"000101100",
  47625=>"001111111",
  47626=>"111000000",
  47627=>"000001011",
  47628=>"000100100",
  47629=>"000000000",
  47630=>"000000111",
  47631=>"010001101",
  47632=>"111111011",
  47633=>"000000000",
  47634=>"000101000",
  47635=>"000000000",
  47636=>"001001000",
  47637=>"111111111",
  47638=>"100111000",
  47639=>"000100111",
  47640=>"111111111",
  47641=>"110111111",
  47642=>"101101001",
  47643=>"000000000",
  47644=>"111111111",
  47645=>"111111000",
  47646=>"000011111",
  47647=>"000000100",
  47648=>"000000001",
  47649=>"000000101",
  47650=>"000000000",
  47651=>"000000110",
  47652=>"000000111",
  47653=>"000000000",
  47654=>"111111111",
  47655=>"011010011",
  47656=>"111111111",
  47657=>"000000100",
  47658=>"110111111",
  47659=>"111000000",
  47660=>"000000111",
  47661=>"111111010",
  47662=>"000000000",
  47663=>"011111111",
  47664=>"000001001",
  47665=>"000110111",
  47666=>"011000011",
  47667=>"000000000",
  47668=>"111111111",
  47669=>"000000111",
  47670=>"010110010",
  47671=>"000011011",
  47672=>"100000111",
  47673=>"011110111",
  47674=>"110111011",
  47675=>"000000000",
  47676=>"000000000",
  47677=>"011011010",
  47678=>"111111111",
  47679=>"101000001",
  47680=>"111111111",
  47681=>"111111111",
  47682=>"010011111",
  47683=>"100000110",
  47684=>"111100000",
  47685=>"000111111",
  47686=>"001001001",
  47687=>"111110111",
  47688=>"110110000",
  47689=>"010111110",
  47690=>"111111011",
  47691=>"111001001",
  47692=>"000000000",
  47693=>"111111111",
  47694=>"000000000",
  47695=>"111100100",
  47696=>"000000000",
  47697=>"111111100",
  47698=>"110110110",
  47699=>"110111011",
  47700=>"001001001",
  47701=>"011011000",
  47702=>"111111101",
  47703=>"000000000",
  47704=>"000001101",
  47705=>"101000001",
  47706=>"001101111",
  47707=>"000001001",
  47708=>"001011010",
  47709=>"111001111",
  47710=>"000000000",
  47711=>"111111111",
  47712=>"110110111",
  47713=>"001000000",
  47714=>"100000000",
  47715=>"000000000",
  47716=>"000000110",
  47717=>"111111111",
  47718=>"001111000",
  47719=>"111111111",
  47720=>"100000101",
  47721=>"000000001",
  47722=>"000000000",
  47723=>"000000011",
  47724=>"101001111",
  47725=>"111000000",
  47726=>"111111111",
  47727=>"000110110",
  47728=>"111111011",
  47729=>"110110111",
  47730=>"000000001",
  47731=>"010000000",
  47732=>"000000000",
  47733=>"000000000",
  47734=>"001001000",
  47735=>"111000111",
  47736=>"100100111",
  47737=>"000001001",
  47738=>"101100100",
  47739=>"000000000",
  47740=>"111110110",
  47741=>"001000000",
  47742=>"111111111",
  47743=>"111111010",
  47744=>"000000100",
  47745=>"000000000",
  47746=>"000000011",
  47747=>"011000000",
  47748=>"000000101",
  47749=>"111111111",
  47750=>"111111111",
  47751=>"001000000",
  47752=>"000000000",
  47753=>"000000100",
  47754=>"000000100",
  47755=>"000000100",
  47756=>"111111111",
  47757=>"100000100",
  47758=>"000101111",
  47759=>"000000000",
  47760=>"011111011",
  47761=>"000000000",
  47762=>"111111110",
  47763=>"110110111",
  47764=>"000100000",
  47765=>"000000000",
  47766=>"011000000",
  47767=>"000000000",
  47768=>"000000000",
  47769=>"000000001",
  47770=>"110110111",
  47771=>"111110000",
  47772=>"000001000",
  47773=>"000000000",
  47774=>"000001011",
  47775=>"000001111",
  47776=>"011110111",
  47777=>"111011001",
  47778=>"001001000",
  47779=>"000010011",
  47780=>"001100000",
  47781=>"010111111",
  47782=>"000000000",
  47783=>"111111111",
  47784=>"001000000",
  47785=>"011111111",
  47786=>"000000000",
  47787=>"111111110",
  47788=>"111111111",
  47789=>"000011000",
  47790=>"001100100",
  47791=>"111111111",
  47792=>"010010011",
  47793=>"111111000",
  47794=>"111111111",
  47795=>"100000000",
  47796=>"110110110",
  47797=>"111111100",
  47798=>"111111000",
  47799=>"001001000",
  47800=>"111111111",
  47801=>"111111111",
  47802=>"001111111",
  47803=>"111111111",
  47804=>"111000000",
  47805=>"000001111",
  47806=>"111111111",
  47807=>"001001111",
  47808=>"100000000",
  47809=>"000010110",
  47810=>"000000111",
  47811=>"000000000",
  47812=>"110111110",
  47813=>"000000011",
  47814=>"011001000",
  47815=>"110110000",
  47816=>"000000000",
  47817=>"010000000",
  47818=>"111111011",
  47819=>"100100100",
  47820=>"001111111",
  47821=>"111100000",
  47822=>"000000010",
  47823=>"110010000",
  47824=>"110000000",
  47825=>"000000000",
  47826=>"111111111",
  47827=>"000000000",
  47828=>"001001111",
  47829=>"111111111",
  47830=>"111000100",
  47831=>"111011011",
  47832=>"101000000",
  47833=>"000110111",
  47834=>"000111010",
  47835=>"111111110",
  47836=>"010000000",
  47837=>"000001001",
  47838=>"011000011",
  47839=>"000000000",
  47840=>"001001001",
  47841=>"111111111",
  47842=>"110111011",
  47843=>"111111011",
  47844=>"000000100",
  47845=>"000000110",
  47846=>"111111111",
  47847=>"111111111",
  47848=>"000000000",
  47849=>"000000001",
  47850=>"010010010",
  47851=>"110110111",
  47852=>"111111000",
  47853=>"001000111",
  47854=>"111111111",
  47855=>"111111111",
  47856=>"111111111",
  47857=>"111111111",
  47858=>"000000001",
  47859=>"000000000",
  47860=>"110000000",
  47861=>"111111111",
  47862=>"011011001",
  47863=>"110110000",
  47864=>"110100100",
  47865=>"011000000",
  47866=>"111011111",
  47867=>"000000110",
  47868=>"000010111",
  47869=>"111000000",
  47870=>"000111100",
  47871=>"111111111",
  47872=>"000000000",
  47873=>"011111111",
  47874=>"100100000",
  47875=>"100000000",
  47876=>"000000000",
  47877=>"111000011",
  47878=>"000000000",
  47879=>"111111111",
  47880=>"111111000",
  47881=>"111111111",
  47882=>"000000010",
  47883=>"000011111",
  47884=>"111111111",
  47885=>"111111000",
  47886=>"111101111",
  47887=>"000000000",
  47888=>"101101110",
  47889=>"000000000",
  47890=>"111111000",
  47891=>"111111111",
  47892=>"000000000",
  47893=>"000000000",
  47894=>"000001001",
  47895=>"000000101",
  47896=>"000011011",
  47897=>"111011110",
  47898=>"100000000",
  47899=>"000001001",
  47900=>"001001011",
  47901=>"011111111",
  47902=>"000000000",
  47903=>"000110000",
  47904=>"110111000",
  47905=>"000000000",
  47906=>"011100000",
  47907=>"111111011",
  47908=>"101101111",
  47909=>"111001111",
  47910=>"000000000",
  47911=>"010000001",
  47912=>"000000001",
  47913=>"000010010",
  47914=>"111111011",
  47915=>"111100000",
  47916=>"111111111",
  47917=>"000001111",
  47918=>"000000001",
  47919=>"111111111",
  47920=>"100100110",
  47921=>"111111000",
  47922=>"000001000",
  47923=>"000000000",
  47924=>"000000000",
  47925=>"000000101",
  47926=>"011111101",
  47927=>"001011000",
  47928=>"000000000",
  47929=>"111111000",
  47930=>"001001100",
  47931=>"000000000",
  47932=>"000000000",
  47933=>"011011000",
  47934=>"000111111",
  47935=>"111111111",
  47936=>"101000101",
  47937=>"001111001",
  47938=>"000000000",
  47939=>"001000000",
  47940=>"111111011",
  47941=>"000000101",
  47942=>"000000000",
  47943=>"000000000",
  47944=>"000000111",
  47945=>"000000000",
  47946=>"110111010",
  47947=>"001101001",
  47948=>"000000000",
  47949=>"000000100",
  47950=>"011010011",
  47951=>"100100110",
  47952=>"111011111",
  47953=>"110110100",
  47954=>"000000000",
  47955=>"111000011",
  47956=>"111111111",
  47957=>"111111111",
  47958=>"000000001",
  47959=>"000011111",
  47960=>"111010001",
  47961=>"110111010",
  47962=>"111111111",
  47963=>"111111111",
  47964=>"000000000",
  47965=>"001001111",
  47966=>"111010000",
  47967=>"110101111",
  47968=>"000000000",
  47969=>"001001011",
  47970=>"000010011",
  47971=>"111111000",
  47972=>"000000000",
  47973=>"000000000",
  47974=>"001001111",
  47975=>"110000001",
  47976=>"010010010",
  47977=>"111110110",
  47978=>"100000000",
  47979=>"111111000",
  47980=>"100000110",
  47981=>"000001111",
  47982=>"000000000",
  47983=>"001110101",
  47984=>"000000000",
  47985=>"000000101",
  47986=>"000110110",
  47987=>"100111111",
  47988=>"111111010",
  47989=>"111111111",
  47990=>"000000001",
  47991=>"110000000",
  47992=>"100000100",
  47993=>"111110100",
  47994=>"111000000",
  47995=>"000010000",
  47996=>"100111110",
  47997=>"111100000",
  47998=>"000010111",
  47999=>"100100100",
  48000=>"000011011",
  48001=>"011010111",
  48002=>"000111111",
  48003=>"101101111",
  48004=>"101000100",
  48005=>"111111110",
  48006=>"111111000",
  48007=>"111110011",
  48008=>"000000000",
  48009=>"000100100",
  48010=>"110010010",
  48011=>"001000100",
  48012=>"001001111",
  48013=>"000011111",
  48014=>"000000111",
  48015=>"000000100",
  48016=>"000000000",
  48017=>"111011000",
  48018=>"110110010",
  48019=>"001001001",
  48020=>"110000000",
  48021=>"000001000",
  48022=>"111101100",
  48023=>"100000000",
  48024=>"100000000",
  48025=>"111110110",
  48026=>"000000000",
  48027=>"001111111",
  48028=>"111110000",
  48029=>"000000001",
  48030=>"000000000",
  48031=>"001000111",
  48032=>"111111111",
  48033=>"000010011",
  48034=>"111111111",
  48035=>"111101111",
  48036=>"001000100",
  48037=>"000000000",
  48038=>"111111111",
  48039=>"001001000",
  48040=>"000000000",
  48041=>"000001111",
  48042=>"010110110",
  48043=>"111001000",
  48044=>"000000110",
  48045=>"000000000",
  48046=>"101100000",
  48047=>"111111000",
  48048=>"111111111",
  48049=>"110111111",
  48050=>"010000000",
  48051=>"000000000",
  48052=>"111111111",
  48053=>"001111111",
  48054=>"011111110",
  48055=>"111111111",
  48056=>"110011000",
  48057=>"011111000",
  48058=>"000110110",
  48059=>"000000000",
  48060=>"000000000",
  48061=>"001100100",
  48062=>"111000000",
  48063=>"011010010",
  48064=>"000000000",
  48065=>"000000000",
  48066=>"000000000",
  48067=>"000000000",
  48068=>"000000001",
  48069=>"110111111",
  48070=>"000100000",
  48071=>"001111111",
  48072=>"000000000",
  48073=>"000000111",
  48074=>"011000011",
  48075=>"000000001",
  48076=>"000000111",
  48077=>"111111111",
  48078=>"001000000",
  48079=>"000000000",
  48080=>"000000000",
  48081=>"000000000",
  48082=>"000000010",
  48083=>"000000101",
  48084=>"111100100",
  48085=>"000111111",
  48086=>"001000000",
  48087=>"000011101",
  48088=>"000000010",
  48089=>"111111111",
  48090=>"000111111",
  48091=>"110000000",
  48092=>"110111111",
  48093=>"111111001",
  48094=>"001001001",
  48095=>"001111111",
  48096=>"000000000",
  48097=>"110110110",
  48098=>"000000111",
  48099=>"000000111",
  48100=>"111111111",
  48101=>"111111111",
  48102=>"011000011",
  48103=>"111000000",
  48104=>"010000011",
  48105=>"000000000",
  48106=>"110111111",
  48107=>"110100101",
  48108=>"011010010",
  48109=>"000010000",
  48110=>"111111111",
  48111=>"111111101",
  48112=>"100100111",
  48113=>"011001111",
  48114=>"011001011",
  48115=>"001000000",
  48116=>"011111011",
  48117=>"111000001",
  48118=>"111110110",
  48119=>"110100110",
  48120=>"110111110",
  48121=>"000000011",
  48122=>"100000000",
  48123=>"111111111",
  48124=>"000000000",
  48125=>"010111111",
  48126=>"111011011",
  48127=>"000000111",
  48128=>"111111111",
  48129=>"101000000",
  48130=>"111111111",
  48131=>"111111110",
  48132=>"100110111",
  48133=>"000000111",
  48134=>"000000000",
  48135=>"111101000",
  48136=>"000000010",
  48137=>"000000111",
  48138=>"111111111",
  48139=>"111111111",
  48140=>"111111110",
  48141=>"111111111",
  48142=>"000000001",
  48143=>"000000000",
  48144=>"101000000",
  48145=>"100111111",
  48146=>"011110100",
  48147=>"000000000",
  48148=>"111011111",
  48149=>"000000000",
  48150=>"000001000",
  48151=>"111111000",
  48152=>"111111000",
  48153=>"100100110",
  48154=>"000000011",
  48155=>"111100000",
  48156=>"000000001",
  48157=>"100010111",
  48158=>"000010011",
  48159=>"111111000",
  48160=>"000001001",
  48161=>"000000000",
  48162=>"111001000",
  48163=>"000000011",
  48164=>"000000111",
  48165=>"000000111",
  48166=>"111111011",
  48167=>"000000001",
  48168=>"111111111",
  48169=>"000000000",
  48170=>"111011011",
  48171=>"111000111",
  48172=>"100000000",
  48173=>"111110011",
  48174=>"000000011",
  48175=>"111111000",
  48176=>"000000111",
  48177=>"000000111",
  48178=>"000000000",
  48179=>"000000000",
  48180=>"111111100",
  48181=>"100100111",
  48182=>"001000000",
  48183=>"111111111",
  48184=>"111111111",
  48185=>"111000011",
  48186=>"000111111",
  48187=>"000011111",
  48188=>"100000111",
  48189=>"111111011",
  48190=>"101000001",
  48191=>"000000000",
  48192=>"000000000",
  48193=>"011011000",
  48194=>"000000111",
  48195=>"000000000",
  48196=>"100110111",
  48197=>"011001000",
  48198=>"110110000",
  48199=>"000000000",
  48200=>"111111001",
  48201=>"111111000",
  48202=>"000000111",
  48203=>"111110111",
  48204=>"000000111",
  48205=>"001001001",
  48206=>"000000000",
  48207=>"111000000",
  48208=>"111111000",
  48209=>"000000111",
  48210=>"000000000",
  48211=>"011111000",
  48212=>"000000001",
  48213=>"000001111",
  48214=>"111011011",
  48215=>"000000000",
  48216=>"111111111",
  48217=>"101101101",
  48218=>"000000000",
  48219=>"001000000",
  48220=>"111111111",
  48221=>"000000000",
  48222=>"000111111",
  48223=>"011010011",
  48224=>"111111111",
  48225=>"000000000",
  48226=>"000011001",
  48227=>"000000000",
  48228=>"000001111",
  48229=>"111101111",
  48230=>"000001111",
  48231=>"000000110",
  48232=>"000000000",
  48233=>"000000000",
  48234=>"011111111",
  48235=>"000010010",
  48236=>"110110001",
  48237=>"111111111",
  48238=>"111111111",
  48239=>"001101000",
  48240=>"111011000",
  48241=>"111000000",
  48242=>"011011111",
  48243=>"100100111",
  48244=>"111111001",
  48245=>"110110110",
  48246=>"000000010",
  48247=>"000001000",
  48248=>"000000111",
  48249=>"000111011",
  48250=>"111011000",
  48251=>"000000111",
  48252=>"110110100",
  48253=>"111111110",
  48254=>"111011000",
  48255=>"011000000",
  48256=>"111010111",
  48257=>"111000000",
  48258=>"111000000",
  48259=>"000000001",
  48260=>"100110000",
  48261=>"001001101",
  48262=>"100001111",
  48263=>"111111111",
  48264=>"110111000",
  48265=>"111000000",
  48266=>"000000000",
  48267=>"111001100",
  48268=>"011111000",
  48269=>"000000000",
  48270=>"000000100",
  48271=>"000011110",
  48272=>"010111000",
  48273=>"110110111",
  48274=>"000000000",
  48275=>"110111111",
  48276=>"111111010",
  48277=>"000010111",
  48278=>"111111000",
  48279=>"000000000",
  48280=>"000000111",
  48281=>"000000000",
  48282=>"111111010",
  48283=>"111001000",
  48284=>"100110110",
  48285=>"000000000",
  48286=>"111111000",
  48287=>"000000111",
  48288=>"001001000",
  48289=>"111111111",
  48290=>"111111110",
  48291=>"111111000",
  48292=>"001000000",
  48293=>"000001001",
  48294=>"111111111",
  48295=>"001111111",
  48296=>"111111000",
  48297=>"000011010",
  48298=>"100100000",
  48299=>"000000111",
  48300=>"111011011",
  48301=>"111011111",
  48302=>"000000111",
  48303=>"000000000",
  48304=>"001001000",
  48305=>"011011101",
  48306=>"110111111",
  48307=>"111111111",
  48308=>"111001100",
  48309=>"011000001",
  48310=>"000111111",
  48311=>"000000000",
  48312=>"111111001",
  48313=>"000001000",
  48314=>"000000000",
  48315=>"000001001",
  48316=>"000000000",
  48317=>"000110101",
  48318=>"111111000",
  48319=>"100111111",
  48320=>"000000000",
  48321=>"001111010",
  48322=>"111111111",
  48323=>"100111111",
  48324=>"000110100",
  48325=>"000111111",
  48326=>"010110111",
  48327=>"000000000",
  48328=>"000111111",
  48329=>"000000000",
  48330=>"000000100",
  48331=>"000000010",
  48332=>"110110000",
  48333=>"000111111",
  48334=>"000100000",
  48335=>"111101000",
  48336=>"111100110",
  48337=>"001000000",
  48338=>"110100000",
  48339=>"111001000",
  48340=>"111111111",
  48341=>"010111100",
  48342=>"000000010",
  48343=>"110111111",
  48344=>"000010100",
  48345=>"000000000",
  48346=>"111111111",
  48347=>"000000111",
  48348=>"110111100",
  48349=>"111111000",
  48350=>"000000000",
  48351=>"000000000",
  48352=>"111111011",
  48353=>"111111111",
  48354=>"000111001",
  48355=>"011000000",
  48356=>"100100000",
  48357=>"100110111",
  48358=>"000011111",
  48359=>"001000000",
  48360=>"111110111",
  48361=>"001000000",
  48362=>"000000101",
  48363=>"110110000",
  48364=>"111111111",
  48365=>"110110111",
  48366=>"000100111",
  48367=>"111111111",
  48368=>"000111111",
  48369=>"000000000",
  48370=>"001000000",
  48371=>"001001000",
  48372=>"111111111",
  48373=>"011110100",
  48374=>"111001001",
  48375=>"000000011",
  48376=>"111111111",
  48377=>"111111111",
  48378=>"000000111",
  48379=>"110110110",
  48380=>"000000000",
  48381=>"101111110",
  48382=>"000000000",
  48383=>"000000001",
  48384=>"000000000",
  48385=>"111011011",
  48386=>"000000111",
  48387=>"111111000",
  48388=>"000000000",
  48389=>"000010111",
  48390=>"000000000",
  48391=>"111111001",
  48392=>"111111000",
  48393=>"000000000",
  48394=>"000000000",
  48395=>"000000011",
  48396=>"111111111",
  48397=>"000000010",
  48398=>"000000110",
  48399=>"011111111",
  48400=>"010100100",
  48401=>"110111111",
  48402=>"111101111",
  48403=>"000000001",
  48404=>"111111111",
  48405=>"000000000",
  48406=>"100111100",
  48407=>"000000000",
  48408=>"000000111",
  48409=>"110000000",
  48410=>"111111100",
  48411=>"111111111",
  48412=>"111111111",
  48413=>"000000010",
  48414=>"111000000",
  48415=>"111111111",
  48416=>"111001011",
  48417=>"111111111",
  48418=>"111111001",
  48419=>"000110111",
  48420=>"101001000",
  48421=>"000100000",
  48422=>"111111111",
  48423=>"000000001",
  48424=>"000000000",
  48425=>"000010111",
  48426=>"011111000",
  48427=>"111111000",
  48428=>"111111111",
  48429=>"001001111",
  48430=>"110000000",
  48431=>"000000111",
  48432=>"111111111",
  48433=>"111111111",
  48434=>"111111111",
  48435=>"000010011",
  48436=>"111101010",
  48437=>"000000000",
  48438=>"100111000",
  48439=>"001001000",
  48440=>"111010000",
  48441=>"000010111",
  48442=>"111111110",
  48443=>"110111111",
  48444=>"011011000",
  48445=>"011111011",
  48446=>"000000000",
  48447=>"111010110",
  48448=>"011000000",
  48449=>"000000000",
  48450=>"111111111",
  48451=>"000001000",
  48452=>"000000111",
  48453=>"111111000",
  48454=>"010000000",
  48455=>"000000111",
  48456=>"111111000",
  48457=>"111111000",
  48458=>"001000000",
  48459=>"111111111",
  48460=>"000000010",
  48461=>"100000111",
  48462=>"001100000",
  48463=>"101100110",
  48464=>"111111001",
  48465=>"111110100",
  48466=>"100000000",
  48467=>"001111011",
  48468=>"111000001",
  48469=>"000001001",
  48470=>"111001000",
  48471=>"111111001",
  48472=>"011111111",
  48473=>"111111000",
  48474=>"000000011",
  48475=>"111111000",
  48476=>"000000111",
  48477=>"000100110",
  48478=>"011111101",
  48479=>"110111111",
  48480=>"100111101",
  48481=>"000000100",
  48482=>"000000100",
  48483=>"000001011",
  48484=>"100100111",
  48485=>"000000010",
  48486=>"100000001",
  48487=>"001001001",
  48488=>"111111110",
  48489=>"100110001",
  48490=>"101111111",
  48491=>"111011000",
  48492=>"001100000",
  48493=>"000000000",
  48494=>"000111110",
  48495=>"001010000",
  48496=>"110000110",
  48497=>"011010000",
  48498=>"000000000",
  48499=>"000000000",
  48500=>"000000010",
  48501=>"000000000",
  48502=>"000000000",
  48503=>"000000111",
  48504=>"101100111",
  48505=>"111111000",
  48506=>"111111000",
  48507=>"110100000",
  48508=>"111100111",
  48509=>"111111000",
  48510=>"000000000",
  48511=>"000000111",
  48512=>"111111101",
  48513=>"101111111",
  48514=>"111111000",
  48515=>"111111111",
  48516=>"111111110",
  48517=>"011111011",
  48518=>"000111111",
  48519=>"100000000",
  48520=>"110100110",
  48521=>"001001001",
  48522=>"000111111",
  48523=>"111111011",
  48524=>"011011001",
  48525=>"000111111",
  48526=>"111111111",
  48527=>"000000000",
  48528=>"000000000",
  48529=>"000000001",
  48530=>"011011111",
  48531=>"110100100",
  48532=>"111111110",
  48533=>"000011001",
  48534=>"101001111",
  48535=>"000000000",
  48536=>"111111111",
  48537=>"000000000",
  48538=>"000001111",
  48539=>"101100100",
  48540=>"101000000",
  48541=>"111110000",
  48542=>"000000000",
  48543=>"001011000",
  48544=>"000101111",
  48545=>"000000011",
  48546=>"001000000",
  48547=>"000000111",
  48548=>"000000100",
  48549=>"110010000",
  48550=>"000000000",
  48551=>"111000000",
  48552=>"000000010",
  48553=>"000000001",
  48554=>"101000111",
  48555=>"000000100",
  48556=>"001000000",
  48557=>"001111111",
  48558=>"000000000",
  48559=>"000011011",
  48560=>"000000000",
  48561=>"000000000",
  48562=>"111000001",
  48563=>"111111111",
  48564=>"000000111",
  48565=>"000001000",
  48566=>"011011011",
  48567=>"111000000",
  48568=>"000000111",
  48569=>"111111111",
  48570=>"000000100",
  48571=>"111111111",
  48572=>"111100110",
  48573=>"000111111",
  48574=>"000000000",
  48575=>"110110000",
  48576=>"111111011",
  48577=>"000000111",
  48578=>"111111100",
  48579=>"110111111",
  48580=>"000000100",
  48581=>"110110110",
  48582=>"000000000",
  48583=>"110000110",
  48584=>"111000000",
  48585=>"111111111",
  48586=>"001000111",
  48587=>"000000000",
  48588=>"000011111",
  48589=>"100000001",
  48590=>"110000000",
  48591=>"000000000",
  48592=>"110110010",
  48593=>"000000000",
  48594=>"000000110",
  48595=>"000000000",
  48596=>"000000111",
  48597=>"000100111",
  48598=>"001111111",
  48599=>"001001001",
  48600=>"000000000",
  48601=>"001111001",
  48602=>"111111111",
  48603=>"111111111",
  48604=>"000000000",
  48605=>"000000000",
  48606=>"111110011",
  48607=>"000111001",
  48608=>"000000000",
  48609=>"100000000",
  48610=>"011111110",
  48611=>"110111111",
  48612=>"010010000",
  48613=>"100100111",
  48614=>"111111111",
  48615=>"011000111",
  48616=>"111111000",
  48617=>"000000111",
  48618=>"000100110",
  48619=>"101111000",
  48620=>"111111111",
  48621=>"001001000",
  48622=>"000000000",
  48623=>"000000000",
  48624=>"000000000",
  48625=>"000000000",
  48626=>"000000000",
  48627=>"111111111",
  48628=>"111111111",
  48629=>"000000000",
  48630=>"000010000",
  48631=>"110110111",
  48632=>"000001111",
  48633=>"110111010",
  48634=>"111111000",
  48635=>"111111000",
  48636=>"110000011",
  48637=>"000000000",
  48638=>"000100000",
  48639=>"001110111",
  48640=>"111000000",
  48641=>"111111111",
  48642=>"111001000",
  48643=>"110111111",
  48644=>"000000011",
  48645=>"111011000",
  48646=>"111111111",
  48647=>"000001111",
  48648=>"111111111",
  48649=>"111111100",
  48650=>"000000000",
  48651=>"111100000",
  48652=>"111111000",
  48653=>"000110010",
  48654=>"111100000",
  48655=>"000000111",
  48656=>"000000001",
  48657=>"111111000",
  48658=>"111111111",
  48659=>"111000000",
  48660=>"000000000",
  48661=>"000010010",
  48662=>"000110111",
  48663=>"000000000",
  48664=>"001111111",
  48665=>"111111111",
  48666=>"111111111",
  48667=>"111000000",
  48668=>"101000011",
  48669=>"100011111",
  48670=>"001011011",
  48671=>"000000111",
  48672=>"000011000",
  48673=>"000111111",
  48674=>"001110100",
  48675=>"000000001",
  48676=>"111000100",
  48677=>"000000100",
  48678=>"001000000",
  48679=>"011010000",
  48680=>"000100111",
  48681=>"111111000",
  48682=>"111111111",
  48683=>"000000001",
  48684=>"000000111",
  48685=>"110110111",
  48686=>"000100111",
  48687=>"011000000",
  48688=>"111111010",
  48689=>"110101111",
  48690=>"011011011",
  48691=>"000110000",
  48692=>"000000000",
  48693=>"111111000",
  48694=>"000001000",
  48695=>"000110111",
  48696=>"000000000",
  48697=>"111111000",
  48698=>"000000000",
  48699=>"111111000",
  48700=>"111010111",
  48701=>"000011000",
  48702=>"010111111",
  48703=>"111111111",
  48704=>"011001000",
  48705=>"111000000",
  48706=>"000000000",
  48707=>"000000111",
  48708=>"000000000",
  48709=>"000000000",
  48710=>"101011001",
  48711=>"111111011",
  48712=>"011011000",
  48713=>"111001111",
  48714=>"000001000",
  48715=>"110000000",
  48716=>"100100000",
  48717=>"000000001",
  48718=>"111000000",
  48719=>"001000001",
  48720=>"000000000",
  48721=>"100111111",
  48722=>"111111001",
  48723=>"111101000",
  48724=>"000000000",
  48725=>"000000000",
  48726=>"111101000",
  48727=>"000000000",
  48728=>"110110111",
  48729=>"111001000",
  48730=>"010111000",
  48731=>"000010011",
  48732=>"111111000",
  48733=>"111111000",
  48734=>"111111001",
  48735=>"001001000",
  48736=>"000110110",
  48737=>"011111111",
  48738=>"101100001",
  48739=>"101101111",
  48740=>"100000000",
  48741=>"001001000",
  48742=>"111111011",
  48743=>"000000111",
  48744=>"000000111",
  48745=>"111111111",
  48746=>"111111000",
  48747=>"000000100",
  48748=>"111111111",
  48749=>"111111111",
  48750=>"101101111",
  48751=>"000000000",
  48752=>"000111111",
  48753=>"111111000",
  48754=>"000000011",
  48755=>"111111111",
  48756=>"111111110",
  48757=>"101001001",
  48758=>"111101000",
  48759=>"101100001",
  48760=>"110001000",
  48761=>"001111111",
  48762=>"101001000",
  48763=>"000001000",
  48764=>"011001001",
  48765=>"000000110",
  48766=>"111111000",
  48767=>"000000000",
  48768=>"000000011",
  48769=>"111101000",
  48770=>"000111111",
  48771=>"111111111",
  48772=>"000000111",
  48773=>"111111000",
  48774=>"111111001",
  48775=>"000000001",
  48776=>"000000000",
  48777=>"000111000",
  48778=>"101000000",
  48779=>"001011001",
  48780=>"111111101",
  48781=>"000000000",
  48782=>"110000000",
  48783=>"000000001",
  48784=>"111000000",
  48785=>"111000000",
  48786=>"000000111",
  48787=>"000000110",
  48788=>"111111111",
  48789=>"011111111",
  48790=>"110111111",
  48791=>"111000000",
  48792=>"000000000",
  48793=>"111100100",
  48794=>"101111111",
  48795=>"000000000",
  48796=>"111100100",
  48797=>"000111111",
  48798=>"111111110",
  48799=>"000000111",
  48800=>"000000000",
  48801=>"000100011",
  48802=>"000111111",
  48803=>"111111111",
  48804=>"001001001",
  48805=>"111111111",
  48806=>"111111011",
  48807=>"001011000",
  48808=>"000111111",
  48809=>"111111111",
  48810=>"101111110",
  48811=>"000000111",
  48812=>"011000000",
  48813=>"110110000",
  48814=>"110111011",
  48815=>"000001111",
  48816=>"000111000",
  48817=>"111001111",
  48818=>"111001011",
  48819=>"111111000",
  48820=>"000001111",
  48821=>"111111111",
  48822=>"111111010",
  48823=>"000111100",
  48824=>"110100111",
  48825=>"011111111",
  48826=>"000000001",
  48827=>"000000000",
  48828=>"111000000",
  48829=>"100000100",
  48830=>"000000010",
  48831=>"111111011",
  48832=>"111101000",
  48833=>"001111011",
  48834=>"000000100",
  48835=>"000000111",
  48836=>"100000000",
  48837=>"000001000",
  48838=>"000000100",
  48839=>"001111000",
  48840=>"111111111",
  48841=>"001000101",
  48842=>"111101110",
  48843=>"111111111",
  48844=>"111000000",
  48845=>"000000000",
  48846=>"000010001",
  48847=>"000000111",
  48848=>"000011000",
  48849=>"111111010",
  48850=>"111011000",
  48851=>"000010010",
  48852=>"100111111",
  48853=>"011111001",
  48854=>"111011010",
  48855=>"111111100",
  48856=>"000000011",
  48857=>"001000000",
  48858=>"000000000",
  48859=>"000000110",
  48860=>"111111101",
  48861=>"000011111",
  48862=>"000000000",
  48863=>"000110000",
  48864=>"000000001",
  48865=>"011001000",
  48866=>"111111111",
  48867=>"000111010",
  48868=>"111111111",
  48869=>"000000110",
  48870=>"111111111",
  48871=>"000000111",
  48872=>"111101110",
  48873=>"111111111",
  48874=>"111111111",
  48875=>"000100000",
  48876=>"111101101",
  48877=>"011011000",
  48878=>"000001000",
  48879=>"011001000",
  48880=>"000111101",
  48881=>"000111111",
  48882=>"111001000",
  48883=>"000011000",
  48884=>"111111111",
  48885=>"000000000",
  48886=>"100100000",
  48887=>"111111111",
  48888=>"111111111",
  48889=>"011001000",
  48890=>"011111111",
  48891=>"000000000",
  48892=>"011010110",
  48893=>"111001001",
  48894=>"000000000",
  48895=>"111111011",
  48896=>"111111000",
  48897=>"111111110",
  48898=>"111111000",
  48899=>"111111111",
  48900=>"000000000",
  48901=>"100100000",
  48902=>"111101100",
  48903=>"011111000",
  48904=>"001011001",
  48905=>"111000000",
  48906=>"111110111",
  48907=>"000000110",
  48908=>"110110111",
  48909=>"010111110",
  48910=>"000000000",
  48911=>"111111000",
  48912=>"011111111",
  48913=>"000000111",
  48914=>"000000000",
  48915=>"011111101",
  48916=>"111001000",
  48917=>"000000000",
  48918=>"011010111",
  48919=>"001000000",
  48920=>"000000011",
  48921=>"101101000",
  48922=>"000000000",
  48923=>"000000001",
  48924=>"100111100",
  48925=>"000000000",
  48926=>"000000111",
  48927=>"001001011",
  48928=>"011010000",
  48929=>"000000111",
  48930=>"011110000",
  48931=>"000000000",
  48932=>"001000000",
  48933=>"101110111",
  48934=>"110001000",
  48935=>"000000110",
  48936=>"001110100",
  48937=>"101100110",
  48938=>"000000111",
  48939=>"011011011",
  48940=>"000000110",
  48941=>"000000000",
  48942=>"001001001",
  48943=>"000000101",
  48944=>"000000000",
  48945=>"111111000",
  48946=>"111111011",
  48947=>"110111111",
  48948=>"111111001",
  48949=>"111111111",
  48950=>"101110000",
  48951=>"001000111",
  48952=>"000000000",
  48953=>"111111000",
  48954=>"001001111",
  48955=>"111000000",
  48956=>"111111011",
  48957=>"000111011",
  48958=>"010110111",
  48959=>"111111011",
  48960=>"000000000",
  48961=>"001001011",
  48962=>"111101000",
  48963=>"001000111",
  48964=>"111111111",
  48965=>"000111111",
  48966=>"000000000",
  48967=>"111111000",
  48968=>"000000000",
  48969=>"101001001",
  48970=>"000100111",
  48971=>"100100100",
  48972=>"000000000",
  48973=>"111111111",
  48974=>"000000000",
  48975=>"011011111",
  48976=>"000001011",
  48977=>"110110000",
  48978=>"111111111",
  48979=>"000000000",
  48980=>"101101101",
  48981=>"111001001",
  48982=>"111111001",
  48983=>"111111000",
  48984=>"111111111",
  48985=>"000000010",
  48986=>"000000111",
  48987=>"000000001",
  48988=>"000000010",
  48989=>"000001000",
  48990=>"111111000",
  48991=>"000000100",
  48992=>"001001111",
  48993=>"000000011",
  48994=>"111101000",
  48995=>"111111111",
  48996=>"010010111",
  48997=>"000000000",
  48998=>"001001111",
  48999=>"001000000",
  49000=>"000001001",
  49001=>"000111111",
  49002=>"111111100",
  49003=>"000100000",
  49004=>"111111001",
  49005=>"000000000",
  49006=>"000111111",
  49007=>"000000000",
  49008=>"000000000",
  49009=>"110111110",
  49010=>"000111011",
  49011=>"011111111",
  49012=>"111111111",
  49013=>"011100100",
  49014=>"000100111",
  49015=>"000000000",
  49016=>"000001111",
  49017=>"101111111",
  49018=>"000000000",
  49019=>"000110010",
  49020=>"000000001",
  49021=>"000111011",
  49022=>"000100000",
  49023=>"111111111",
  49024=>"000000111",
  49025=>"001000000",
  49026=>"100100110",
  49027=>"111100111",
  49028=>"011010000",
  49029=>"011011111",
  49030=>"000000111",
  49031=>"000011111",
  49032=>"000000000",
  49033=>"011000000",
  49034=>"001000001",
  49035=>"001001001",
  49036=>"011001000",
  49037=>"101001111",
  49038=>"000000000",
  49039=>"000010111",
  49040=>"010111011",
  49041=>"111101000",
  49042=>"110000000",
  49043=>"111111110",
  49044=>"000000000",
  49045=>"111110010",
  49046=>"111111101",
  49047=>"111000000",
  49048=>"000111111",
  49049=>"000000000",
  49050=>"000000101",
  49051=>"011001011",
  49052=>"111000000",
  49053=>"100110000",
  49054=>"000000011",
  49055=>"000000111",
  49056=>"001001000",
  49057=>"111111001",
  49058=>"011111101",
  49059=>"000101111",
  49060=>"001000100",
  49061=>"010000001",
  49062=>"000111000",
  49063=>"111111101",
  49064=>"110110000",
  49065=>"000000000",
  49066=>"011011111",
  49067=>"000111111",
  49068=>"000000000",
  49069=>"111111101",
  49070=>"000000000",
  49071=>"111111111",
  49072=>"000000111",
  49073=>"100000000",
  49074=>"000000000",
  49075=>"000000010",
  49076=>"101001000",
  49077=>"000110111",
  49078=>"001000111",
  49079=>"000110111",
  49080=>"000000111",
  49081=>"111100100",
  49082=>"111101100",
  49083=>"000100000",
  49084=>"000100000",
  49085=>"111001000",
  49086=>"000000000",
  49087=>"001000001",
  49088=>"010110000",
  49089=>"000001000",
  49090=>"111111111",
  49091=>"000000000",
  49092=>"000000111",
  49093=>"111111000",
  49094=>"111111000",
  49095=>"000000000",
  49096=>"111111000",
  49097=>"111111000",
  49098=>"111111000",
  49099=>"111001100",
  49100=>"000000000",
  49101=>"111111111",
  49102=>"111111110",
  49103=>"100110111",
  49104=>"111001000",
  49105=>"000001111",
  49106=>"111111110",
  49107=>"111111111",
  49108=>"111111111",
  49109=>"000100000",
  49110=>"000000110",
  49111=>"110000001",
  49112=>"111110100",
  49113=>"000000000",
  49114=>"111010010",
  49115=>"111111110",
  49116=>"000011111",
  49117=>"011011010",
  49118=>"101000000",
  49119=>"110110111",
  49120=>"000000001",
  49121=>"111111100",
  49122=>"111111111",
  49123=>"111111000",
  49124=>"000000000",
  49125=>"100000110",
  49126=>"111010000",
  49127=>"001111011",
  49128=>"111111111",
  49129=>"000000110",
  49130=>"000111111",
  49131=>"111111100",
  49132=>"000000000",
  49133=>"011000000",
  49134=>"110111010",
  49135=>"000001111",
  49136=>"000000001",
  49137=>"000111000",
  49138=>"001000101",
  49139=>"100000111",
  49140=>"111111011",
  49141=>"000010111",
  49142=>"011000000",
  49143=>"111111100",
  49144=>"011011001",
  49145=>"000000010",
  49146=>"001111111",
  49147=>"111000000",
  49148=>"001001000",
  49149=>"110110000",
  49150=>"010111000",
  49151=>"000111111",
  49152=>"001101001",
  49153=>"000000110",
  49154=>"001000001",
  49155=>"000000111",
  49156=>"010110110",
  49157=>"000000000",
  49158=>"000110001",
  49159=>"111111011",
  49160=>"010001101",
  49161=>"000000000",
  49162=>"000010010",
  49163=>"111111111",
  49164=>"000001000",
  49165=>"111111111",
  49166=>"100111110",
  49167=>"000111010",
  49168=>"101110110",
  49169=>"000111111",
  49170=>"000000001",
  49171=>"000000000",
  49172=>"000000001",
  49173=>"001001001",
  49174=>"000001001",
  49175=>"000100110",
  49176=>"110110100",
  49177=>"011000110",
  49178=>"000000000",
  49179=>"110110110",
  49180=>"000000000",
  49181=>"100110111",
  49182=>"001001001",
  49183=>"111111111",
  49184=>"110110000",
  49185=>"100000000",
  49186=>"001000111",
  49187=>"100100110",
  49188=>"000000001",
  49189=>"001001001",
  49190=>"011001111",
  49191=>"111011011",
  49192=>"011001000",
  49193=>"000000100",
  49194=>"001000001",
  49195=>"111010111",
  49196=>"000001001",
  49197=>"001001101",
  49198=>"000000000",
  49199=>"110110111",
  49200=>"110110010",
  49201=>"000000101",
  49202=>"001001111",
  49203=>"111111000",
  49204=>"000010000",
  49205=>"101100100",
  49206=>"000010000",
  49207=>"111110011",
  49208=>"000100000",
  49209=>"111110000",
  49210=>"111111000",
  49211=>"000000000",
  49212=>"111111110",
  49213=>"010111001",
  49214=>"010010010",
  49215=>"111001100",
  49216=>"000010000",
  49217=>"111111110",
  49218=>"111011000",
  49219=>"111111111",
  49220=>"100100000",
  49221=>"011011010",
  49222=>"101101111",
  49223=>"111111111",
  49224=>"011011101",
  49225=>"001001001",
  49226=>"111111111",
  49227=>"111110000",
  49228=>"000011001",
  49229=>"111111111",
  49230=>"101101011",
  49231=>"001001000",
  49232=>"000101101",
  49233=>"101101001",
  49234=>"000000000",
  49235=>"111100000",
  49236=>"000111111",
  49237=>"000000111",
  49238=>"001011011",
  49239=>"110110110",
  49240=>"000100100",
  49241=>"111100100",
  49242=>"001001011",
  49243=>"000110110",
  49244=>"111111111",
  49245=>"111111111",
  49246=>"111011001",
  49247=>"110000000",
  49248=>"000010110",
  49249=>"100110110",
  49250=>"000000000",
  49251=>"000001000",
  49252=>"010000001",
  49253=>"100000000",
  49254=>"101101101",
  49255=>"000000110",
  49256=>"011010011",
  49257=>"000000000",
  49258=>"111010000",
  49259=>"111111001",
  49260=>"111111111",
  49261=>"110110110",
  49262=>"101001001",
  49263=>"100111111",
  49264=>"001000000",
  49265=>"111100000",
  49266=>"111111000",
  49267=>"001001001",
  49268=>"000001101",
  49269=>"111011001",
  49270=>"111001001",
  49271=>"011011000",
  49272=>"000000110",
  49273=>"100010111",
  49274=>"001001000",
  49275=>"101101101",
  49276=>"100110000",
  49277=>"000001111",
  49278=>"110110110",
  49279=>"000001001",
  49280=>"001000000",
  49281=>"000010011",
  49282=>"011011111",
  49283=>"110000000",
  49284=>"100110110",
  49285=>"100000000",
  49286=>"110000000",
  49287=>"000011110",
  49288=>"000000000",
  49289=>"111000000",
  49290=>"111100100",
  49291=>"000000000",
  49292=>"110110011",
  49293=>"010000010",
  49294=>"110110000",
  49295=>"111111111",
  49296=>"101001001",
  49297=>"000001101",
  49298=>"000000000",
  49299=>"011001001",
  49300=>"111110111",
  49301=>"011001111",
  49302=>"000100111",
  49303=>"001001101",
  49304=>"001001000",
  49305=>"000000001",
  49306=>"010110111",
  49307=>"010111011",
  49308=>"110010000",
  49309=>"000010010",
  49310=>"111111111",
  49311=>"111111111",
  49312=>"001111101",
  49313=>"000111111",
  49314=>"110110100",
  49315=>"111101101",
  49316=>"101111101",
  49317=>"111111111",
  49318=>"101111000",
  49319=>"010010000",
  49320=>"111000011",
  49321=>"010110110",
  49322=>"011001001",
  49323=>"111111111",
  49324=>"000001001",
  49325=>"111101101",
  49326=>"100100111",
  49327=>"010010110",
  49328=>"111111111",
  49329=>"100110100",
  49330=>"111111111",
  49331=>"110111111",
  49332=>"010110000",
  49333=>"001001101",
  49334=>"000000000",
  49335=>"111101100",
  49336=>"011011010",
  49337=>"101101101",
  49338=>"001001001",
  49339=>"001010010",
  49340=>"000000000",
  49341=>"111000000",
  49342=>"111111111",
  49343=>"110111011",
  49344=>"001000100",
  49345=>"000010110",
  49346=>"011000000",
  49347=>"000000111",
  49348=>"000000110",
  49349=>"000000000",
  49350=>"111111101",
  49351=>"111111110",
  49352=>"110110110",
  49353=>"010110111",
  49354=>"000110000",
  49355=>"000000001",
  49356=>"111111100",
  49357=>"010110110",
  49358=>"001001111",
  49359=>"001000001",
  49360=>"111010111",
  49361=>"000000010",
  49362=>"001111111",
  49363=>"100000101",
  49364=>"111111111",
  49365=>"010000111",
  49366=>"000000010",
  49367=>"110000101",
  49368=>"110000000",
  49369=>"110010111",
  49370=>"100000001",
  49371=>"100000110",
  49372=>"001001101",
  49373=>"111101101",
  49374=>"000000000",
  49375=>"001001011",
  49376=>"011011000",
  49377=>"000110000",
  49378=>"101101110",
  49379=>"111011011",
  49380=>"000000001",
  49381=>"111111111",
  49382=>"111010000",
  49383=>"000110110",
  49384=>"111010111",
  49385=>"100000000",
  49386=>"000000000",
  49387=>"000110111",
  49388=>"000000100",
  49389=>"100100111",
  49390=>"110010000",
  49391=>"000000101",
  49392=>"110000000",
  49393=>"000000001",
  49394=>"111001001",
  49395=>"001001001",
  49396=>"001000001",
  49397=>"000000100",
  49398=>"000100100",
  49399=>"000110111",
  49400=>"111111111",
  49401=>"000010010",
  49402=>"111111111",
  49403=>"000010111",
  49404=>"000001001",
  49405=>"111010000",
  49406=>"101101111",
  49407=>"000000001",
  49408=>"111111111",
  49409=>"101101101",
  49410=>"001000100",
  49411=>"000000100",
  49412=>"001000100",
  49413=>"000111111",
  49414=>"001001101",
  49415=>"001010000",
  49416=>"111111111",
  49417=>"101101111",
  49418=>"111101000",
  49419=>"000000000",
  49420=>"001001001",
  49421=>"111111111",
  49422=>"000000100",
  49423=>"000000000",
  49424=>"001001001",
  49425=>"010000011",
  49426=>"101000000",
  49427=>"110000100",
  49428=>"011011011",
  49429=>"000000110",
  49430=>"001100101",
  49431=>"110110110",
  49432=>"110110001",
  49433=>"111001001",
  49434=>"110011001",
  49435=>"010000000",
  49436=>"100111111",
  49437=>"010000000",
  49438=>"111111111",
  49439=>"001001011",
  49440=>"000100100",
  49441=>"001010011",
  49442=>"111110111",
  49443=>"110111111",
  49444=>"111111111",
  49445=>"000000000",
  49446=>"000000000",
  49447=>"110010000",
  49448=>"000111111",
  49449=>"000000000",
  49450=>"000110111",
  49451=>"001111111",
  49452=>"001001000",
  49453=>"001001011",
  49454=>"111111111",
  49455=>"111000111",
  49456=>"100100101",
  49457=>"000011001",
  49458=>"111110111",
  49459=>"111111111",
  49460=>"110111110",
  49461=>"101011111",
  49462=>"001001111",
  49463=>"000000000",
  49464=>"011001000",
  49465=>"111111111",
  49466=>"001000000",
  49467=>"001000111",
  49468=>"100000011",
  49469=>"110110001",
  49470=>"000010110",
  49471=>"110110111",
  49472=>"000001001",
  49473=>"000000111",
  49474=>"001000001",
  49475=>"101101101",
  49476=>"110110010",
  49477=>"001000011",
  49478=>"000000100",
  49479=>"100000001",
  49480=>"010100100",
  49481=>"000000010",
  49482=>"111111110",
  49483=>"100100110",
  49484=>"000000110",
  49485=>"111000000",
  49486=>"110110010",
  49487=>"110011001",
  49488=>"000111111",
  49489=>"001001111",
  49490=>"111111111",
  49491=>"010110111",
  49492=>"000000000",
  49493=>"110010010",
  49494=>"000110110",
  49495=>"000001001",
  49496=>"000001000",
  49497=>"110110110",
  49498=>"111111111",
  49499=>"001001101",
  49500=>"000110111",
  49501=>"010000000",
  49502=>"000001101",
  49503=>"110110111",
  49504=>"001111111",
  49505=>"000000001",
  49506=>"100000000",
  49507=>"000100111",
  49508=>"010011111",
  49509=>"001001000",
  49510=>"011000001",
  49511=>"000000001",
  49512=>"001001001",
  49513=>"000000000",
  49514=>"001011111",
  49515=>"000010110",
  49516=>"111011011",
  49517=>"000001110",
  49518=>"000000000",
  49519=>"110011111",
  49520=>"000100110",
  49521=>"100010000",
  49522=>"000001000",
  49523=>"111111001",
  49524=>"011000000",
  49525=>"000001110",
  49526=>"111100011",
  49527=>"000000000",
  49528=>"000000111",
  49529=>"111011001",
  49530=>"000000100",
  49531=>"000000000",
  49532=>"111011000",
  49533=>"111010000",
  49534=>"110000000",
  49535=>"101000000",
  49536=>"001000100",
  49537=>"111111000",
  49538=>"110110110",
  49539=>"000000000",
  49540=>"110111100",
  49541=>"001001001",
  49542=>"000000000",
  49543=>"001101001",
  49544=>"001000001",
  49545=>"110111111",
  49546=>"000000000",
  49547=>"000000111",
  49548=>"000000000",
  49549=>"000000000",
  49550=>"011011111",
  49551=>"000000000",
  49552=>"000001001",
  49553=>"110110110",
  49554=>"011010111",
  49555=>"011001111",
  49556=>"010100111",
  49557=>"000000000",
  49558=>"111110110",
  49559=>"111001001",
  49560=>"000000001",
  49561=>"011111111",
  49562=>"010011011",
  49563=>"000001001",
  49564=>"011111111",
  49565=>"101111111",
  49566=>"001001001",
  49567=>"000111111",
  49568=>"000001001",
  49569=>"110000000",
  49570=>"011010010",
  49571=>"111000000",
  49572=>"000010000",
  49573=>"000111010",
  49574=>"000000000",
  49575=>"111111111",
  49576=>"000111111",
  49577=>"001011001",
  49578=>"000000000",
  49579=>"001011111",
  49580=>"000000000",
  49581=>"001001000",
  49582=>"001001111",
  49583=>"111011000",
  49584=>"101101111",
  49585=>"000000000",
  49586=>"000001001",
  49587=>"111111111",
  49588=>"000110111",
  49589=>"101000000",
  49590=>"000000100",
  49591=>"000010111",
  49592=>"111111001",
  49593=>"110110111",
  49594=>"000001001",
  49595=>"001001101",
  49596=>"000000000",
  49597=>"110010111",
  49598=>"000001111",
  49599=>"001000100",
  49600=>"101001000",
  49601=>"011011001",
  49602=>"000000000",
  49603=>"000000000",
  49604=>"001011001",
  49605=>"000000100",
  49606=>"100110110",
  49607=>"001011111",
  49608=>"111001101",
  49609=>"101000000",
  49610=>"001001001",
  49611=>"000000011",
  49612=>"111111001",
  49613=>"110110010",
  49614=>"010000000",
  49615=>"101100000",
  49616=>"100000111",
  49617=>"000000001",
  49618=>"000010110",
  49619=>"001001001",
  49620=>"001011111",
  49621=>"000001001",
  49622=>"000000000",
  49623=>"111111100",
  49624=>"000001111",
  49625=>"010010101",
  49626=>"001001111",
  49627=>"100101101",
  49628=>"110110110",
  49629=>"000000001",
  49630=>"110000110",
  49631=>"001101001",
  49632=>"111101000",
  49633=>"111001001",
  49634=>"000000000",
  49635=>"101001111",
  49636=>"100101101",
  49637=>"101110110",
  49638=>"000000100",
  49639=>"000000001",
  49640=>"000000000",
  49641=>"001000000",
  49642=>"000001101",
  49643=>"111111000",
  49644=>"100000000",
  49645=>"100111101",
  49646=>"001000001",
  49647=>"111110110",
  49648=>"001001101",
  49649=>"000000000",
  49650=>"111110111",
  49651=>"111111011",
  49652=>"111001000",
  49653=>"000000000",
  49654=>"110111111",
  49655=>"100100100",
  49656=>"111101101",
  49657=>"000001101",
  49658=>"000001111",
  49659=>"101001001",
  49660=>"011111111",
  49661=>"010110110",
  49662=>"111110100",
  49663=>"101001101",
  49664=>"111111111",
  49665=>"000000000",
  49666=>"000000000",
  49667=>"000000000",
  49668=>"111111111",
  49669=>"111001000",
  49670=>"001111111",
  49671=>"111111111",
  49672=>"100110011",
  49673=>"101111001",
  49674=>"111100000",
  49675=>"000011111",
  49676=>"000000001",
  49677=>"001111111",
  49678=>"100101101",
  49679=>"111111111",
  49680=>"110110111",
  49681=>"000000000",
  49682=>"000111111",
  49683=>"100000000",
  49684=>"111111111",
  49685=>"111111000",
  49686=>"001000010",
  49687=>"000000011",
  49688=>"000000000",
  49689=>"111111111",
  49690=>"000000111",
  49691=>"111110100",
  49692=>"000000000",
  49693=>"111111111",
  49694=>"111110111",
  49695=>"111111000",
  49696=>"100101001",
  49697=>"110110110",
  49698=>"110100110",
  49699=>"111000011",
  49700=>"000000000",
  49701=>"000000000",
  49702=>"011000001",
  49703=>"111111111",
  49704=>"100111111",
  49705=>"100000000",
  49706=>"111111111",
  49707=>"111000000",
  49708=>"000000000",
  49709=>"000000000",
  49710=>"111111111",
  49711=>"001001111",
  49712=>"000000000",
  49713=>"000000000",
  49714=>"000100110",
  49715=>"000000000",
  49716=>"000001000",
  49717=>"011001000",
  49718=>"111111000",
  49719=>"110100000",
  49720=>"000100111",
  49721=>"111111111",
  49722=>"111111111",
  49723=>"111000000",
  49724=>"000000000",
  49725=>"100100000",
  49726=>"000000000",
  49727=>"110100111",
  49728=>"111111100",
  49729=>"111100111",
  49730=>"111111111",
  49731=>"001101001",
  49732=>"000000000",
  49733=>"000111011",
  49734=>"000000000",
  49735=>"101001000",
  49736=>"011000011",
  49737=>"001000001",
  49738=>"111111111",
  49739=>"110111110",
  49740=>"000100111",
  49741=>"100011001",
  49742=>"111111111",
  49743=>"000000100",
  49744=>"111111111",
  49745=>"111111111",
  49746=>"000110111",
  49747=>"001001011",
  49748=>"000111010",
  49749=>"000110010",
  49750=>"001000100",
  49751=>"000000000",
  49752=>"000100001",
  49753=>"000000000",
  49754=>"000010010",
  49755=>"100011011",
  49756=>"000000110",
  49757=>"111111001",
  49758=>"111001111",
  49759=>"100101100",
  49760=>"111110111",
  49761=>"111000000",
  49762=>"000100100",
  49763=>"111111111",
  49764=>"111111111",
  49765=>"000000000",
  49766=>"111111111",
  49767=>"111111001",
  49768=>"000111110",
  49769=>"111111111",
  49770=>"000000000",
  49771=>"111111111",
  49772=>"010010100",
  49773=>"111111101",
  49774=>"111111111",
  49775=>"111111111",
  49776=>"000000101",
  49777=>"101111111",
  49778=>"111111101",
  49779=>"001001111",
  49780=>"000000000",
  49781=>"111110001",
  49782=>"111010010",
  49783=>"000100100",
  49784=>"000001001",
  49785=>"111111111",
  49786=>"000100100",
  49787=>"111111111",
  49788=>"110110110",
  49789=>"000010010",
  49790=>"000010110",
  49791=>"111111111",
  49792=>"011111111",
  49793=>"000000000",
  49794=>"000000111",
  49795=>"110000011",
  49796=>"111111110",
  49797=>"111111111",
  49798=>"101111110",
  49799=>"000011111",
  49800=>"111111101",
  49801=>"000000000",
  49802=>"000100000",
  49803=>"111111111",
  49804=>"111111111",
  49805=>"100000000",
  49806=>"000000000",
  49807=>"111111111",
  49808=>"110111111",
  49809=>"001000000",
  49810=>"111111100",
  49811=>"000100000",
  49812=>"111011000",
  49813=>"100101011",
  49814=>"111111111",
  49815=>"111111000",
  49816=>"101100111",
  49817=>"111101111",
  49818=>"110111010",
  49819=>"000000000",
  49820=>"000000000",
  49821=>"000000100",
  49822=>"111111111",
  49823=>"000000000",
  49824=>"000000000",
  49825=>"000100000",
  49826=>"111111111",
  49827=>"110111111",
  49828=>"000000000",
  49829=>"111000101",
  49830=>"000000111",
  49831=>"110111011",
  49832=>"011111111",
  49833=>"111111111",
  49834=>"111110111",
  49835=>"111000001",
  49836=>"011111110",
  49837=>"110000000",
  49838=>"100100110",
  49839=>"011100000",
  49840=>"111000000",
  49841=>"110010011",
  49842=>"111111010",
  49843=>"000000000",
  49844=>"111111001",
  49845=>"000000000",
  49846=>"000000000",
  49847=>"101111111",
  49848=>"101000000",
  49849=>"000000000",
  49850=>"000000000",
  49851=>"111100111",
  49852=>"111111111",
  49853=>"000000000",
  49854=>"001000111",
  49855=>"111111111",
  49856=>"000000000",
  49857=>"001001000",
  49858=>"111111111",
  49859=>"000000000",
  49860=>"111000001",
  49861=>"000000000",
  49862=>"011011011",
  49863=>"100110100",
  49864=>"000000011",
  49865=>"111000100",
  49866=>"101101101",
  49867=>"011011000",
  49868=>"100101111",
  49869=>"000001111",
  49870=>"000000000",
  49871=>"000000000",
  49872=>"000001111",
  49873=>"000000110",
  49874=>"000000111",
  49875=>"111000000",
  49876=>"000111111",
  49877=>"110110110",
  49878=>"000000000",
  49879=>"000000110",
  49880=>"001100000",
  49881=>"000000000",
  49882=>"001000000",
  49883=>"000000111",
  49884=>"000110100",
  49885=>"000000000",
  49886=>"001111110",
  49887=>"001011011",
  49888=>"111111110",
  49889=>"000100111",
  49890=>"000000111",
  49891=>"111101000",
  49892=>"101001001",
  49893=>"111111111",
  49894=>"000000000",
  49895=>"100111111",
  49896=>"111111111",
  49897=>"000001000",
  49898=>"000000000",
  49899=>"001000000",
  49900=>"011011111",
  49901=>"000000011",
  49902=>"000000111",
  49903=>"000000000",
  49904=>"110010000",
  49905=>"111110111",
  49906=>"111000000",
  49907=>"000000000",
  49908=>"011011111",
  49909=>"111000000",
  49910=>"111011111",
  49911=>"111111111",
  49912=>"001000000",
  49913=>"110111111",
  49914=>"111001000",
  49915=>"000111111",
  49916=>"000110111",
  49917=>"111001001",
  49918=>"111110111",
  49919=>"000111111",
  49920=>"000000100",
  49921=>"000000000",
  49922=>"000000000",
  49923=>"111111111",
  49924=>"001001001",
  49925=>"111111111",
  49926=>"111110110",
  49927=>"101111111",
  49928=>"000100100",
  49929=>"000000000",
  49930=>"000000000",
  49931=>"100100001",
  49932=>"001001011",
  49933=>"001011011",
  49934=>"110110100",
  49935=>"100001111",
  49936=>"110110000",
  49937=>"111111111",
  49938=>"000000001",
  49939=>"000000001",
  49940=>"000000000",
  49941=>"111111111",
  49942=>"000001001",
  49943=>"110111111",
  49944=>"000000000",
  49945=>"000110000",
  49946=>"011001000",
  49947=>"111101111",
  49948=>"111111111",
  49949=>"111111111",
  49950=>"000000000",
  49951=>"000000100",
  49952=>"111111011",
  49953=>"101111000",
  49954=>"111111111",
  49955=>"000000000",
  49956=>"010000000",
  49957=>"000001101",
  49958=>"110110110",
  49959=>"011000000",
  49960=>"111111111",
  49961=>"111000000",
  49962=>"111101111",
  49963=>"000000010",
  49964=>"111111110",
  49965=>"110111111",
  49966=>"000000000",
  49967=>"000000000",
  49968=>"111111111",
  49969=>"111111001",
  49970=>"000000110",
  49971=>"100100110",
  49972=>"111111111",
  49973=>"000000100",
  49974=>"111111000",
  49975=>"111100001",
  49976=>"000000000",
  49977=>"000000000",
  49978=>"111011000",
  49979=>"111011000",
  49980=>"000000000",
  49981=>"000000011",
  49982=>"010001000",
  49983=>"111111000",
  49984=>"111111111",
  49985=>"000000000",
  49986=>"111000000",
  49987=>"100000000",
  49988=>"100000000",
  49989=>"111000000",
  49990=>"000001000",
  49991=>"111111111",
  49992=>"111000000",
  49993=>"000000001",
  49994=>"111100101",
  49995=>"110111110",
  49996=>"000000000",
  49997=>"001001000",
  49998=>"000100100",
  49999=>"000000000",
  50000=>"000001100",
  50001=>"001001111",
  50002=>"001000000",
  50003=>"000000000",
  50004=>"000000110",
  50005=>"011011011",
  50006=>"111111111",
  50007=>"111111111",
  50008=>"111111111",
  50009=>"000000000",
  50010=>"000000001",
  50011=>"000000010",
  50012=>"000000000",
  50013=>"000000000",
  50014=>"000000000",
  50015=>"001011111",
  50016=>"000100110",
  50017=>"000000000",
  50018=>"101101100",
  50019=>"111111111",
  50020=>"000000000",
  50021=>"000000000",
  50022=>"111000000",
  50023=>"000000000",
  50024=>"001000001",
  50025=>"011111000",
  50026=>"000000000",
  50027=>"111111110",
  50028=>"011011111",
  50029=>"111111111",
  50030=>"011111111",
  50031=>"111011000",
  50032=>"000010110",
  50033=>"100100111",
  50034=>"000000100",
  50035=>"000000000",
  50036=>"000101001",
  50037=>"100100100",
  50038=>"000000101",
  50039=>"111111111",
  50040=>"011001000",
  50041=>"111111111",
  50042=>"000000010",
  50043=>"110000000",
  50044=>"000011111",
  50045=>"000000000",
  50046=>"000000001",
  50047=>"111111111",
  50048=>"000000000",
  50049=>"111100000",
  50050=>"011011011",
  50051=>"111111111",
  50052=>"000111111",
  50053=>"000100111",
  50054=>"110010000",
  50055=>"000100100",
  50056=>"000001000",
  50057=>"111000000",
  50058=>"111111111",
  50059=>"100111111",
  50060=>"001000111",
  50061=>"110110110",
  50062=>"100110111",
  50063=>"000000000",
  50064=>"000001000",
  50065=>"111111111",
  50066=>"111011111",
  50067=>"000000000",
  50068=>"111010000",
  50069=>"000000000",
  50070=>"000000000",
  50071=>"111001000",
  50072=>"111111100",
  50073=>"111111111",
  50074=>"111111111",
  50075=>"000000000",
  50076=>"000000000",
  50077=>"111110111",
  50078=>"001001001",
  50079=>"000000000",
  50080=>"000001011",
  50081=>"000000000",
  50082=>"100000111",
  50083=>"111011111",
  50084=>"000100110",
  50085=>"000000000",
  50086=>"111111111",
  50087=>"111111111",
  50088=>"000000000",
  50089=>"011111111",
  50090=>"011011000",
  50091=>"111111101",
  50092=>"111111000",
  50093=>"000000000",
  50094=>"111000100",
  50095=>"100100101",
  50096=>"111110111",
  50097=>"111111111",
  50098=>"111111111",
  50099=>"011011111",
  50100=>"000100100",
  50101=>"110100111",
  50102=>"111101011",
  50103=>"100101111",
  50104=>"011110111",
  50105=>"111011000",
  50106=>"000000000",
  50107=>"101111110",
  50108=>"110110010",
  50109=>"000001011",
  50110=>"000101111",
  50111=>"000000010",
  50112=>"100111111",
  50113=>"000000000",
  50114=>"111111111",
  50115=>"011111111",
  50116=>"001001101",
  50117=>"000000000",
  50118=>"000000111",
  50119=>"000010111",
  50120=>"111111010",
  50121=>"110110000",
  50122=>"101100111",
  50123=>"000000000",
  50124=>"000000000",
  50125=>"000000000",
  50126=>"011001000",
  50127=>"111111001",
  50128=>"111111111",
  50129=>"000000000",
  50130=>"111111111",
  50131=>"111000000",
  50132=>"110010111",
  50133=>"000000000",
  50134=>"000100001",
  50135=>"000100100",
  50136=>"111100111",
  50137=>"000000001",
  50138=>"000001000",
  50139=>"100000000",
  50140=>"000000000",
  50141=>"000100111",
  50142=>"000010000",
  50143=>"100100001",
  50144=>"111100000",
  50145=>"111100100",
  50146=>"111111001",
  50147=>"111111111",
  50148=>"111000000",
  50149=>"010000000",
  50150=>"001101111",
  50151=>"111111000",
  50152=>"111111011",
  50153=>"111111001",
  50154=>"111111110",
  50155=>"111111111",
  50156=>"111111010",
  50157=>"100100100",
  50158=>"000000000",
  50159=>"011000000",
  50160=>"000000000",
  50161=>"000000011",
  50162=>"000000000",
  50163=>"001001001",
  50164=>"111111111",
  50165=>"000011011",
  50166=>"011010000",
  50167=>"011011010",
  50168=>"001000001",
  50169=>"001011111",
  50170=>"110110000",
  50171=>"000000000",
  50172=>"100111111",
  50173=>"111101100",
  50174=>"111111010",
  50175=>"111110110",
  50176=>"001001001",
  50177=>"000000000",
  50178=>"001111111",
  50179=>"000000000",
  50180=>"001001011",
  50181=>"000010000",
  50182=>"000001000",
  50183=>"101000101",
  50184=>"011011000",
  50185=>"100110111",
  50186=>"000000000",
  50187=>"000000011",
  50188=>"011011000",
  50189=>"110000001",
  50190=>"001011000",
  50191=>"000000000",
  50192=>"111011111",
  50193=>"000000001",
  50194=>"100100000",
  50195=>"111110110",
  50196=>"111000000",
  50197=>"000000000",
  50198=>"001000000",
  50199=>"011111111",
  50200=>"000000000",
  50201=>"001011000",
  50202=>"111111111",
  50203=>"111011000",
  50204=>"011011011",
  50205=>"000000000",
  50206=>"111001000",
  50207=>"111111111",
  50208=>"011110110",
  50209=>"111001001",
  50210=>"001000000",
  50211=>"000000001",
  50212=>"110011000",
  50213=>"000000111",
  50214=>"110110111",
  50215=>"000000001",
  50216=>"000001011",
  50217=>"010110010",
  50218=>"000000000",
  50219=>"011000000",
  50220=>"111111111",
  50221=>"000100000",
  50222=>"111111001",
  50223=>"000000000",
  50224=>"110110110",
  50225=>"000000000",
  50226=>"000001000",
  50227=>"000000000",
  50228=>"000111111",
  50229=>"011011000",
  50230=>"000001100",
  50231=>"111111111",
  50232=>"010010001",
  50233=>"000010111",
  50234=>"000000000",
  50235=>"111000000",
  50236=>"111101111",
  50237=>"001011011",
  50238=>"100100111",
  50239=>"000000000",
  50240=>"000001011",
  50241=>"110010000",
  50242=>"000011111",
  50243=>"011011111",
  50244=>"111111111",
  50245=>"000000001",
  50246=>"111111000",
  50247=>"001111111",
  50248=>"111001000",
  50249=>"000000001",
  50250=>"000010111",
  50251=>"111111111",
  50252=>"001111110",
  50253=>"010111111",
  50254=>"100100100",
  50255=>"000000000",
  50256=>"101100000",
  50257=>"111110111",
  50258=>"000001001",
  50259=>"111011011",
  50260=>"100100000",
  50261=>"100001000",
  50262=>"101100000",
  50263=>"001001111",
  50264=>"000000000",
  50265=>"000000011",
  50266=>"111000000",
  50267=>"111111010",
  50268=>"000000000",
  50269=>"111000000",
  50270=>"000000110",
  50271=>"100100000",
  50272=>"000000000",
  50273=>"000000000",
  50274=>"111010011",
  50275=>"110110100",
  50276=>"111100000",
  50277=>"111111110",
  50278=>"111111111",
  50279=>"111111011",
  50280=>"000000000",
  50281=>"111111111",
  50282=>"011000011",
  50283=>"000000001",
  50284=>"001111110",
  50285=>"111111111",
  50286=>"000000110",
  50287=>"000000110",
  50288=>"001000000",
  50289=>"001111111",
  50290=>"000000001",
  50291=>"011000000",
  50292=>"111111011",
  50293=>"000000000",
  50294=>"111111111",
  50295=>"000000000",
  50296=>"000000000",
  50297=>"111111001",
  50298=>"000111000",
  50299=>"010000010",
  50300=>"110110110",
  50301=>"000111111",
  50302=>"001001001",
  50303=>"010011011",
  50304=>"000000110",
  50305=>"001000000",
  50306=>"000000110",
  50307=>"111110111",
  50308=>"111011011",
  50309=>"111111111",
  50310=>"111111010",
  50311=>"111011000",
  50312=>"111000000",
  50313=>"001111111",
  50314=>"000000000",
  50315=>"111111111",
  50316=>"000100001",
  50317=>"000000000",
  50318=>"010010110",
  50319=>"111001111",
  50320=>"000000000",
  50321=>"111100100",
  50322=>"000110111",
  50323=>"000000000",
  50324=>"000010010",
  50325=>"110110100",
  50326=>"000000000",
  50327=>"011000000",
  50328=>"011111111",
  50329=>"110011011",
  50330=>"000000000",
  50331=>"000000000",
  50332=>"111111110",
  50333=>"000001000",
  50334=>"111111111",
  50335=>"000000001",
  50336=>"000000000",
  50337=>"000000000",
  50338=>"000000000",
  50339=>"111010000",
  50340=>"001101011",
  50341=>"001001111",
  50342=>"111111111",
  50343=>"000111111",
  50344=>"111111111",
  50345=>"000001000",
  50346=>"000000111",
  50347=>"111011011",
  50348=>"100000000",
  50349=>"011111110",
  50350=>"111111111",
  50351=>"000001001",
  50352=>"111111100",
  50353=>"000000000",
  50354=>"011111011",
  50355=>"000000000",
  50356=>"000000000",
  50357=>"111111111",
  50358=>"000100100",
  50359=>"000000000",
  50360=>"001000001",
  50361=>"111001001",
  50362=>"000100111",
  50363=>"111111111",
  50364=>"000000100",
  50365=>"001000000",
  50366=>"000111110",
  50367=>"000000000",
  50368=>"000000100",
  50369=>"111110100",
  50370=>"111111111",
  50371=>"111111111",
  50372=>"000110001",
  50373=>"111011000",
  50374=>"000000001",
  50375=>"110110111",
  50376=>"000001111",
  50377=>"111111111",
  50378=>"111110000",
  50379=>"000000110",
  50380=>"110111000",
  50381=>"110010000",
  50382=>"110111111",
  50383=>"000000000",
  50384=>"011101111",
  50385=>"010110110",
  50386=>"111111001",
  50387=>"001000010",
  50388=>"000000110",
  50389=>"100000000",
  50390=>"111011111",
  50391=>"010010110",
  50392=>"011010000",
  50393=>"011111111",
  50394=>"000000000",
  50395=>"111111111",
  50396=>"000000000",
  50397=>"111111111",
  50398=>"111111111",
  50399=>"111111111",
  50400=>"101000000",
  50401=>"011001111",
  50402=>"000011011",
  50403=>"111110000",
  50404=>"000000000",
  50405=>"110110000",
  50406=>"111110110",
  50407=>"111111111",
  50408=>"011011000",
  50409=>"111111110",
  50410=>"101001101",
  50411=>"000000000",
  50412=>"000101000",
  50413=>"111111111",
  50414=>"111111111",
  50415=>"000000000",
  50416=>"100000000",
  50417=>"000110110",
  50418=>"011111111",
  50419=>"111111111",
  50420=>"000000000",
  50421=>"011001001",
  50422=>"011011011",
  50423=>"111111111",
  50424=>"000000000",
  50425=>"111111111",
  50426=>"111001001",
  50427=>"001011111",
  50428=>"000000000",
  50429=>"001111001",
  50430=>"111010010",
  50431=>"000000000",
  50432=>"011111111",
  50433=>"011111001",
  50434=>"000001110",
  50435=>"111111111",
  50436=>"111111001",
  50437=>"000001101",
  50438=>"100000000",
  50439=>"110111111",
  50440=>"000000101",
  50441=>"111001000",
  50442=>"000000000",
  50443=>"000000000",
  50444=>"011111111",
  50445=>"111111110",
  50446=>"110000000",
  50447=>"111101000",
  50448=>"000110011",
  50449=>"000000101",
  50450=>"000000111",
  50451=>"111111111",
  50452=>"111110000",
  50453=>"000001001",
  50454=>"111111111",
  50455=>"011011111",
  50456=>"111001001",
  50457=>"010000000",
  50458=>"000000000",
  50459=>"111101111",
  50460=>"000000001",
  50461=>"100100111",
  50462=>"000000111",
  50463=>"111101101",
  50464=>"111111111",
  50465=>"001000000",
  50466=>"111111000",
  50467=>"111001001",
  50468=>"001000000",
  50469=>"111111111",
  50470=>"110100111",
  50471=>"000100000",
  50472=>"110000000",
  50473=>"000000000",
  50474=>"111110000",
  50475=>"100000000",
  50476=>"001000001",
  50477=>"111111111",
  50478=>"000000000",
  50479=>"000000000",
  50480=>"111111111",
  50481=>"100111010",
  50482=>"001001000",
  50483=>"111000000",
  50484=>"111100000",
  50485=>"111111001",
  50486=>"000010000",
  50487=>"111111111",
  50488=>"000000111",
  50489=>"000000001",
  50490=>"000000000",
  50491=>"111111110",
  50492=>"110110111",
  50493=>"110110111",
  50494=>"000000000",
  50495=>"001000000",
  50496=>"011011101",
  50497=>"100100100",
  50498=>"011001000",
  50499=>"000000111",
  50500=>"000000110",
  50501=>"110000110",
  50502=>"000000000",
  50503=>"110111111",
  50504=>"000000000",
  50505=>"000000000",
  50506=>"001000000",
  50507=>"111111111",
  50508=>"100000110",
  50509=>"101011001",
  50510=>"000000000",
  50511=>"111111111",
  50512=>"100111111",
  50513=>"000000011",
  50514=>"101111111",
  50515=>"011011010",
  50516=>"000000000",
  50517=>"011011001",
  50518=>"111111111",
  50519=>"000000000",
  50520=>"000000000",
  50521=>"111111111",
  50522=>"001001000",
  50523=>"000001111",
  50524=>"000000000",
  50525=>"000000100",
  50526=>"001001101",
  50527=>"100000001",
  50528=>"000101111",
  50529=>"111111111",
  50530=>"111100000",
  50531=>"100100111",
  50532=>"011001000",
  50533=>"000000000",
  50534=>"111111111",
  50535=>"111010010",
  50536=>"111111111",
  50537=>"010010010",
  50538=>"010111111",
  50539=>"000000010",
  50540=>"111001010",
  50541=>"101111111",
  50542=>"111111111",
  50543=>"111101101",
  50544=>"011000000",
  50545=>"111111111",
  50546=>"111111111",
  50547=>"100110010",
  50548=>"000011000",
  50549=>"111011000",
  50550=>"111111000",
  50551=>"111111000",
  50552=>"010000000",
  50553=>"011111111",
  50554=>"011111001",
  50555=>"000000110",
  50556=>"010010011",
  50557=>"001111011",
  50558=>"010110111",
  50559=>"000111110",
  50560=>"111111111",
  50561=>"101000010",
  50562=>"000000000",
  50563=>"000000000",
  50564=>"000000000",
  50565=>"000000000",
  50566=>"100100000",
  50567=>"000100000",
  50568=>"000000000",
  50569=>"000000000",
  50570=>"111111111",
  50571=>"110011000",
  50572=>"000000101",
  50573=>"111101100",
  50574=>"111111111",
  50575=>"111111000",
  50576=>"111111111",
  50577=>"011011111",
  50578=>"111111111",
  50579=>"001000100",
  50580=>"111000000",
  50581=>"000000000",
  50582=>"111101001",
  50583=>"011011111",
  50584=>"011011111",
  50585=>"000000000",
  50586=>"000000000",
  50587=>"000000000",
  50588=>"000001001",
  50589=>"111011011",
  50590=>"001001100",
  50591=>"101011111",
  50592=>"111100110",
  50593=>"000000000",
  50594=>"001111111",
  50595=>"011011011",
  50596=>"111111111",
  50597=>"111111111",
  50598=>"111000001",
  50599=>"011000011",
  50600=>"010000000",
  50601=>"000000001",
  50602=>"111111110",
  50603=>"111001001",
  50604=>"000000000",
  50605=>"111111111",
  50606=>"000100111",
  50607=>"110000010",
  50608=>"000000000",
  50609=>"110111111",
  50610=>"111101111",
  50611=>"000000000",
  50612=>"000101100",
  50613=>"001001111",
  50614=>"111111111",
  50615=>"110000000",
  50616=>"011111111",
  50617=>"111111110",
  50618=>"010000000",
  50619=>"000101111",
  50620=>"000000000",
  50621=>"111110100",
  50622=>"110111000",
  50623=>"001101000",
  50624=>"111010000",
  50625=>"111011011",
  50626=>"000000000",
  50627=>"011111111",
  50628=>"111101000",
  50629=>"100111110",
  50630=>"011011011",
  50631=>"000000000",
  50632=>"111111111",
  50633=>"000110010",
  50634=>"000000000",
  50635=>"101111111",
  50636=>"010000110",
  50637=>"111111010",
  50638=>"000000000",
  50639=>"110110111",
  50640=>"111111001",
  50641=>"000000000",
  50642=>"111111111",
  50643=>"111111110",
  50644=>"111111110",
  50645=>"000001111",
  50646=>"000000111",
  50647=>"000011000",
  50648=>"111110111",
  50649=>"111111111",
  50650=>"111111111",
  50651=>"000000000",
  50652=>"101001000",
  50653=>"111111110",
  50654=>"010010000",
  50655=>"001001011",
  50656=>"000111111",
  50657=>"000000000",
  50658=>"000000000",
  50659=>"111110000",
  50660=>"001001000",
  50661=>"111111111",
  50662=>"000000101",
  50663=>"110110110",
  50664=>"111111011",
  50665=>"000000000",
  50666=>"000000010",
  50667=>"000001001",
  50668=>"001001000",
  50669=>"100100110",
  50670=>"000000000",
  50671=>"001101111",
  50672=>"000000011",
  50673=>"000000110",
  50674=>"111111011",
  50675=>"000000000",
  50676=>"001001000",
  50677=>"110100100",
  50678=>"000000000",
  50679=>"000000001",
  50680=>"111111111",
  50681=>"000000001",
  50682=>"011011000",
  50683=>"111111111",
  50684=>"111111110",
  50685=>"000000000",
  50686=>"111001111",
  50687=>"000000000",
  50688=>"111110111",
  50689=>"000011111",
  50690=>"111111010",
  50691=>"000000001",
  50692=>"100000000",
  50693=>"101100100",
  50694=>"111111111",
  50695=>"101101100",
  50696=>"001100000",
  50697=>"111110100",
  50698=>"111100000",
  50699=>"001111111",
  50700=>"000000000",
  50701=>"000000000",
  50702=>"001000111",
  50703=>"000000111",
  50704=>"000110111",
  50705=>"110110111",
  50706=>"100110111",
  50707=>"000000000",
  50708=>"111111111",
  50709=>"000000000",
  50710=>"000000001",
  50711=>"000000000",
  50712=>"111011011",
  50713=>"011001001",
  50714=>"110110100",
  50715=>"010011011",
  50716=>"010010000",
  50717=>"000000100",
  50718=>"000000000",
  50719=>"000111111",
  50720=>"111111011",
  50721=>"110110111",
  50722=>"111111100",
  50723=>"110111110",
  50724=>"011001011",
  50725=>"000100000",
  50726=>"111111101",
  50727=>"111101001",
  50728=>"111111000",
  50729=>"110110100",
  50730=>"101000000",
  50731=>"000110000",
  50732=>"000010111",
  50733=>"000000100",
  50734=>"101111111",
  50735=>"000100011",
  50736=>"111111111",
  50737=>"111111111",
  50738=>"001001001",
  50739=>"111111111",
  50740=>"111111101",
  50741=>"001011011",
  50742=>"000000000",
  50743=>"111111100",
  50744=>"000000001",
  50745=>"000000010",
  50746=>"111111100",
  50747=>"110110000",
  50748=>"001000111",
  50749=>"111111001",
  50750=>"110110111",
  50751=>"111000001",
  50752=>"111101111",
  50753=>"000000000",
  50754=>"111111111",
  50755=>"110000110",
  50756=>"000001000",
  50757=>"001111111",
  50758=>"000000000",
  50759=>"110111111",
  50760=>"111100100",
  50761=>"111010010",
  50762=>"000000001",
  50763=>"111111111",
  50764=>"001000000",
  50765=>"100000000",
  50766=>"000001101",
  50767=>"000111011",
  50768=>"101111001",
  50769=>"100100110",
  50770=>"111011011",
  50771=>"010010000",
  50772=>"111100000",
  50773=>"111111111",
  50774=>"000000000",
  50775=>"001001001",
  50776=>"000100111",
  50777=>"110110110",
  50778=>"000000000",
  50779=>"000000000",
  50780=>"111111111",
  50781=>"110011001",
  50782=>"000000000",
  50783=>"011111011",
  50784=>"111000000",
  50785=>"000000101",
  50786=>"111000000",
  50787=>"110000111",
  50788=>"111000100",
  50789=>"000000000",
  50790=>"100100100",
  50791=>"111100111",
  50792=>"000000011",
  50793=>"111111111",
  50794=>"011011000",
  50795=>"000010000",
  50796=>"011111111",
  50797=>"000000000",
  50798=>"000011111",
  50799=>"111111111",
  50800=>"000111111",
  50801=>"001111110",
  50802=>"100100101",
  50803=>"111001000",
  50804=>"000000000",
  50805=>"000110110",
  50806=>"000000000",
  50807=>"101101100",
  50808=>"000001111",
  50809=>"111001000",
  50810=>"100111111",
  50811=>"000000000",
  50812=>"111111111",
  50813=>"000000000",
  50814=>"011111000",
  50815=>"111101000",
  50816=>"111101001",
  50817=>"100110111",
  50818=>"111111111",
  50819=>"111000111",
  50820=>"000000001",
  50821=>"100011001",
  50822=>"001111111",
  50823=>"000000000",
  50824=>"111111010",
  50825=>"111100100",
  50826=>"111111111",
  50827=>"000000001",
  50828=>"111111111",
  50829=>"000000001",
  50830=>"111111011",
  50831=>"000000000",
  50832=>"000101000",
  50833=>"001000000",
  50834=>"000000001",
  50835=>"111111001",
  50836=>"110101110",
  50837=>"111111111",
  50838=>"000000000",
  50839=>"100111000",
  50840=>"111110100",
  50841=>"101100000",
  50842=>"000110000",
  50843=>"111111111",
  50844=>"011000000",
  50845=>"111011001",
  50846=>"101110111",
  50847=>"001111101",
  50848=>"100111111",
  50849=>"011000000",
  50850=>"001000000",
  50851=>"000000000",
  50852=>"000000010",
  50853=>"000000110",
  50854=>"000000000",
  50855=>"000000100",
  50856=>"000000011",
  50857=>"000000000",
  50858=>"011000000",
  50859=>"111111111",
  50860=>"111111000",
  50861=>"000000000",
  50862=>"100110000",
  50863=>"000000101",
  50864=>"100111110",
  50865=>"001001100",
  50866=>"100100100",
  50867=>"010110111",
  50868=>"000011111",
  50869=>"110111011",
  50870=>"000000000",
  50871=>"001000000",
  50872=>"111101100",
  50873=>"000000100",
  50874=>"100100101",
  50875=>"111111011",
  50876=>"011110000",
  50877=>"000001111",
  50878=>"000000000",
  50879=>"100000011",
  50880=>"111111111",
  50881=>"000000000",
  50882=>"000000000",
  50883=>"111100000",
  50884=>"111111111",
  50885=>"000000000",
  50886=>"111111111",
  50887=>"111111111",
  50888=>"000000000",
  50889=>"000000001",
  50890=>"000000001",
  50891=>"111111111",
  50892=>"000110110",
  50893=>"100110110",
  50894=>"011111000",
  50895=>"101111111",
  50896=>"000000000",
  50897=>"001001111",
  50898=>"000000000",
  50899=>"000000000",
  50900=>"100110000",
  50901=>"000011011",
  50902=>"000000110",
  50903=>"000000000",
  50904=>"011011000",
  50905=>"100100000",
  50906=>"000000000",
  50907=>"000010111",
  50908=>"000011111",
  50909=>"000111110",
  50910=>"111001000",
  50911=>"111111111",
  50912=>"011011000",
  50913=>"000011011",
  50914=>"111111100",
  50915=>"111000000",
  50916=>"111010011",
  50917=>"000000000",
  50918=>"011111111",
  50919=>"000000000",
  50920=>"111011001",
  50921=>"000000000",
  50922=>"010110111",
  50923=>"001001011",
  50924=>"000010111",
  50925=>"000000010",
  50926=>"100101111",
  50927=>"010111000",
  50928=>"000000101",
  50929=>"000000000",
  50930=>"001011001",
  50931=>"100100011",
  50932=>"111111111",
  50933=>"011011001",
  50934=>"001011111",
  50935=>"111111110",
  50936=>"111111111",
  50937=>"000000000",
  50938=>"000000000",
  50939=>"000100110",
  50940=>"000000000",
  50941=>"000000110",
  50942=>"000000000",
  50943=>"000000000",
  50944=>"110111011",
  50945=>"111111110",
  50946=>"000000000",
  50947=>"000001111",
  50948=>"111111111",
  50949=>"111111001",
  50950=>"111000000",
  50951=>"111111111",
  50952=>"111011000",
  50953=>"001001111",
  50954=>"000010000",
  50955=>"111111111",
  50956=>"100000000",
  50957=>"000001111",
  50958=>"111111100",
  50959=>"000000100",
  50960=>"011011111",
  50961=>"111110100",
  50962=>"100100000",
  50963=>"101000000",
  50964=>"000000000",
  50965=>"000000001",
  50966=>"001011011",
  50967=>"011001001",
  50968=>"000000000",
  50969=>"111000000",
  50970=>"000000100",
  50971=>"010000000",
  50972=>"101000111",
  50973=>"111111111",
  50974=>"000000000",
  50975=>"110110010",
  50976=>"000000010",
  50977=>"000000000",
  50978=>"111111001",
  50979=>"000010000",
  50980=>"111111101",
  50981=>"111111111",
  50982=>"010010011",
  50983=>"100100110",
  50984=>"000010110",
  50985=>"100111111",
  50986=>"100111111",
  50987=>"111111111",
  50988=>"011010000",
  50989=>"110110000",
  50990=>"110000000",
  50991=>"111111111",
  50992=>"111111111",
  50993=>"111111111",
  50994=>"111111111",
  50995=>"001000001",
  50996=>"010010110",
  50997=>"110111111",
  50998=>"000000111",
  50999=>"101100000",
  51000=>"000000000",
  51001=>"010000000",
  51002=>"000000010",
  51003=>"000000111",
  51004=>"111111111",
  51005=>"100110111",
  51006=>"011111111",
  51007=>"101111010",
  51008=>"000110000",
  51009=>"000000000",
  51010=>"000001001",
  51011=>"111111111",
  51012=>"000000100",
  51013=>"000000000",
  51014=>"000100111",
  51015=>"000000000",
  51016=>"110111111",
  51017=>"111111111",
  51018=>"000001000",
  51019=>"011111001",
  51020=>"100100100",
  51021=>"111111101",
  51022=>"100000001",
  51023=>"100000001",
  51024=>"011010011",
  51025=>"001000011",
  51026=>"000000000",
  51027=>"011000000",
  51028=>"001110110",
  51029=>"001011011",
  51030=>"110111111",
  51031=>"111111111",
  51032=>"010011011",
  51033=>"001000000",
  51034=>"111111111",
  51035=>"111011000",
  51036=>"000000100",
  51037=>"111111101",
  51038=>"000000000",
  51039=>"000000000",
  51040=>"111001111",
  51041=>"100000000",
  51042=>"000011011",
  51043=>"110110111",
  51044=>"111010011",
  51045=>"101111111",
  51046=>"110110001",
  51047=>"001000000",
  51048=>"000101111",
  51049=>"111111111",
  51050=>"111111111",
  51051=>"011111111",
  51052=>"000011000",
  51053=>"100000000",
  51054=>"011000000",
  51055=>"111111101",
  51056=>"000001111",
  51057=>"111111111",
  51058=>"000101111",
  51059=>"110100100",
  51060=>"000000000",
  51061=>"001000000",
  51062=>"111111111",
  51063=>"000010110",
  51064=>"000001101",
  51065=>"000011110",
  51066=>"000000010",
  51067=>"111111101",
  51068=>"011111000",
  51069=>"111110100",
  51070=>"111111111",
  51071=>"111111111",
  51072=>"111011011",
  51073=>"000000111",
  51074=>"001001011",
  51075=>"111110000",
  51076=>"000000010",
  51077=>"100000000",
  51078=>"111110111",
  51079=>"000101001",
  51080=>"000000000",
  51081=>"111111111",
  51082=>"111111111",
  51083=>"000010000",
  51084=>"111111111",
  51085=>"111111111",
  51086=>"111111111",
  51087=>"000001000",
  51088=>"100111111",
  51089=>"001001000",
  51090=>"000000000",
  51091=>"101001000",
  51092=>"111111100",
  51093=>"001010111",
  51094=>"000000000",
  51095=>"000011110",
  51096=>"000001011",
  51097=>"001001011",
  51098=>"011111011",
  51099=>"111111111",
  51100=>"111111111",
  51101=>"111111111",
  51102=>"100100000",
  51103=>"000000000",
  51104=>"000000011",
  51105=>"110110010",
  51106=>"111111110",
  51107=>"100111111",
  51108=>"101101101",
  51109=>"000000000",
  51110=>"001000000",
  51111=>"111111111",
  51112=>"111111111",
  51113=>"100110110",
  51114=>"000000000",
  51115=>"100000000",
  51116=>"001000000",
  51117=>"101101111",
  51118=>"111111001",
  51119=>"001001011",
  51120=>"111111111",
  51121=>"111011011",
  51122=>"110010000",
  51123=>"000000000",
  51124=>"111000000",
  51125=>"000000001",
  51126=>"100101001",
  51127=>"111011011",
  51128=>"000111111",
  51129=>"110111111",
  51130=>"100100111",
  51131=>"111111100",
  51132=>"000000000",
  51133=>"000111111",
  51134=>"000000010",
  51135=>"110001111",
  51136=>"000000001",
  51137=>"000000000",
  51138=>"000000000",
  51139=>"000100100",
  51140=>"000000000",
  51141=>"000011001",
  51142=>"111111110",
  51143=>"000000000",
  51144=>"110010010",
  51145=>"111011111",
  51146=>"111111111",
  51147=>"000000000",
  51148=>"000000000",
  51149=>"111111110",
  51150=>"000000000",
  51151=>"000000000",
  51152=>"000000000",
  51153=>"100001000",
  51154=>"111110100",
  51155=>"100110101",
  51156=>"110110110",
  51157=>"110110010",
  51158=>"000000000",
  51159=>"001001011",
  51160=>"000000001",
  51161=>"000100100",
  51162=>"101101111",
  51163=>"111111111",
  51164=>"001000000",
  51165=>"111111111",
  51166=>"111111000",
  51167=>"001000010",
  51168=>"000000000",
  51169=>"000000000",
  51170=>"111001111",
  51171=>"101000000",
  51172=>"000000011",
  51173=>"100110011",
  51174=>"000001000",
  51175=>"001001001",
  51176=>"000111001",
  51177=>"111110111",
  51178=>"111000101",
  51179=>"111101111",
  51180=>"011111111",
  51181=>"110010000",
  51182=>"100110100",
  51183=>"010010010",
  51184=>"000000000",
  51185=>"111111111",
  51186=>"001000001",
  51187=>"111111111",
  51188=>"111111001",
  51189=>"000110000",
  51190=>"011011111",
  51191=>"001011111",
  51192=>"000000000",
  51193=>"110110011",
  51194=>"111111111",
  51195=>"110111111",
  51196=>"000000000",
  51197=>"111111100",
  51198=>"100000001",
  51199=>"100000001",
  51200=>"011011111",
  51201=>"111111111",
  51202=>"111000000",
  51203=>"000011011",
  51204=>"111111111",
  51205=>"001000001",
  51206=>"111000000",
  51207=>"000000011",
  51208=>"100000001",
  51209=>"010000000",
  51210=>"111111111",
  51211=>"111011000",
  51212=>"000000110",
  51213=>"001000000",
  51214=>"011111110",
  51215=>"111111111",
  51216=>"000011011",
  51217=>"111111111",
  51218=>"111001001",
  51219=>"111111111",
  51220=>"000000110",
  51221=>"000111111",
  51222=>"000000001",
  51223=>"001001000",
  51224=>"000000000",
  51225=>"000100111",
  51226=>"111100000",
  51227=>"110000100",
  51228=>"000000111",
  51229=>"000000111",
  51230=>"111011010",
  51231=>"000011111",
  51232=>"110000011",
  51233=>"100100111",
  51234=>"111000000",
  51235=>"000000010",
  51236=>"111001000",
  51237=>"100111100",
  51238=>"111110000",
  51239=>"000111111",
  51240=>"111000000",
  51241=>"111111111",
  51242=>"000000111",
  51243=>"000000000",
  51244=>"000101001",
  51245=>"111111000",
  51246=>"111100110",
  51247=>"111111000",
  51248=>"001111010",
  51249=>"111111011",
  51250=>"111111000",
  51251=>"111000000",
  51252=>"101111100",
  51253=>"101100100",
  51254=>"111101000",
  51255=>"000000000",
  51256=>"111010010",
  51257=>"111111111",
  51258=>"111101111",
  51259=>"111111000",
  51260=>"001000000",
  51261=>"111111111",
  51262=>"111111111",
  51263=>"101000000",
  51264=>"000111111",
  51265=>"100110110",
  51266=>"000000000",
  51267=>"010111000",
  51268=>"001000011",
  51269=>"000111111",
  51270=>"001111111",
  51271=>"110000000",
  51272=>"000000001",
  51273=>"000000111",
  51274=>"000000001",
  51275=>"000111010",
  51276=>"000100010",
  51277=>"111001111",
  51278=>"111000111",
  51279=>"110111111",
  51280=>"000111111",
  51281=>"000111111",
  51282=>"110000001",
  51283=>"001001000",
  51284=>"111101001",
  51285=>"111000011",
  51286=>"111100000",
  51287=>"011111111",
  51288=>"001101111",
  51289=>"000000111",
  51290=>"100000100",
  51291=>"111111110",
  51292=>"000000111",
  51293=>"000000000",
  51294=>"000000111",
  51295=>"111111011",
  51296=>"000110111",
  51297=>"000000000",
  51298=>"101000101",
  51299=>"111111111",
  51300=>"000000111",
  51301=>"000000000",
  51302=>"111111010",
  51303=>"111001101",
  51304=>"000000000",
  51305=>"000001011",
  51306=>"100110111",
  51307=>"111111111",
  51308=>"111111110",
  51309=>"111111110",
  51310=>"101000000",
  51311=>"111101101",
  51312=>"111111000",
  51313=>"000010000",
  51314=>"110110000",
  51315=>"001011110",
  51316=>"110111111",
  51317=>"111111000",
  51318=>"000000100",
  51319=>"111111111",
  51320=>"011000000",
  51321=>"010101111",
  51322=>"000000000",
  51323=>"111011000",
  51324=>"000000000",
  51325=>"000111111",
  51326=>"111110000",
  51327=>"111111111",
  51328=>"111111111",
  51329=>"111111000",
  51330=>"111101111",
  51331=>"000111001",
  51332=>"111101001",
  51333=>"000000000",
  51334=>"110110110",
  51335=>"111000000",
  51336=>"001001000",
  51337=>"000000000",
  51338=>"000000000",
  51339=>"111111111",
  51340=>"000100111",
  51341=>"111111111",
  51342=>"011110000",
  51343=>"111000000",
  51344=>"000000000",
  51345=>"111111111",
  51346=>"000101101",
  51347=>"111111111",
  51348=>"110111011",
  51349=>"111101111",
  51350=>"000000001",
  51351=>"011001001",
  51352=>"001001011",
  51353=>"001011001",
  51354=>"111110000",
  51355=>"110000000",
  51356=>"010000111",
  51357=>"111111111",
  51358=>"110010000",
  51359=>"000101111",
  51360=>"111111110",
  51361=>"111100111",
  51362=>"100111100",
  51363=>"111100101",
  51364=>"000100000",
  51365=>"000111111",
  51366=>"000000000",
  51367=>"111011011",
  51368=>"000000011",
  51369=>"111001000",
  51370=>"000000001",
  51371=>"111001111",
  51372=>"010010110",
  51373=>"111011000",
  51374=>"111000111",
  51375=>"100100111",
  51376=>"000000111",
  51377=>"111111111",
  51378=>"000000000",
  51379=>"000000000",
  51380=>"000000010",
  51381=>"000000000",
  51382=>"111101111",
  51383=>"111010111",
  51384=>"000000000",
  51385=>"000010111",
  51386=>"000000000",
  51387=>"000010010",
  51388=>"111001001",
  51389=>"111111111",
  51390=>"000011000",
  51391=>"100000000",
  51392=>"011000110",
  51393=>"111111000",
  51394=>"000111111",
  51395=>"011001010",
  51396=>"111001101",
  51397=>"011011000",
  51398=>"011011011",
  51399=>"101111111",
  51400=>"000000000",
  51401=>"001100100",
  51402=>"000001001",
  51403=>"111000001",
  51404=>"000000000",
  51405=>"001101111",
  51406=>"011011011",
  51407=>"110011000",
  51408=>"111111111",
  51409=>"111000111",
  51410=>"101111111",
  51411=>"000111111",
  51412=>"001100111",
  51413=>"000100000",
  51414=>"111111111",
  51415=>"110010000",
  51416=>"111111101",
  51417=>"000000010",
  51418=>"000001000",
  51419=>"001001100",
  51420=>"110010010",
  51421=>"010000000",
  51422=>"000100111",
  51423=>"111101000",
  51424=>"100000101",
  51425=>"100100110",
  51426=>"000000100",
  51427=>"001000000",
  51428=>"000000000",
  51429=>"101101101",
  51430=>"000110010",
  51431=>"000000010",
  51432=>"000001111",
  51433=>"111011000",
  51434=>"011111111",
  51435=>"111111000",
  51436=>"011001000",
  51437=>"111111101",
  51438=>"011000101",
  51439=>"000000000",
  51440=>"000000000",
  51441=>"011011111",
  51442=>"111000000",
  51443=>"111110010",
  51444=>"000000000",
  51445=>"011011111",
  51446=>"110110111",
  51447=>"111111111",
  51448=>"111000000",
  51449=>"111101011",
  51450=>"000000001",
  51451=>"111101001",
  51452=>"111110000",
  51453=>"110110100",
  51454=>"001001001",
  51455=>"111000000",
  51456=>"010111111",
  51457=>"010011010",
  51458=>"000000000",
  51459=>"000000001",
  51460=>"111000000",
  51461=>"111111111",
  51462=>"011111011",
  51463=>"000000000",
  51464=>"100111111",
  51465=>"000010010",
  51466=>"111101101",
  51467=>"000000000",
  51468=>"000000000",
  51469=>"111111111",
  51470=>"111111111",
  51471=>"000111111",
  51472=>"111001000",
  51473=>"000000000",
  51474=>"000000000",
  51475=>"001111100",
  51476=>"101001111",
  51477=>"111111111",
  51478=>"110110000",
  51479=>"111111111",
  51480=>"000000110",
  51481=>"000000000",
  51482=>"111111001",
  51483=>"111111111",
  51484=>"111011000",
  51485=>"000000000",
  51486=>"000101111",
  51487=>"100100111",
  51488=>"000110111",
  51489=>"100000111",
  51490=>"001111111",
  51491=>"111011111",
  51492=>"000000100",
  51493=>"000000110",
  51494=>"001101011",
  51495=>"000000110",
  51496=>"111111100",
  51497=>"001111111",
  51498=>"000111111",
  51499=>"000000000",
  51500=>"110110010",
  51501=>"011111111",
  51502=>"000000111",
  51503=>"011011011",
  51504=>"011001011",
  51505=>"111001000",
  51506=>"000000000",
  51507=>"111111111",
  51508=>"000000000",
  51509=>"011111111",
  51510=>"000111111",
  51511=>"010111111",
  51512=>"111111010",
  51513=>"111000000",
  51514=>"001000000",
  51515=>"111111111",
  51516=>"011011011",
  51517=>"000000000",
  51518=>"000001111",
  51519=>"000000000",
  51520=>"010011000",
  51521=>"000110000",
  51522=>"000110111",
  51523=>"000000000",
  51524=>"000000001",
  51525=>"110000000",
  51526=>"001111111",
  51527=>"111111111",
  51528=>"111111111",
  51529=>"111000110",
  51530=>"001000000",
  51531=>"000100001",
  51532=>"000000110",
  51533=>"101110111",
  51534=>"011111011",
  51535=>"101100100",
  51536=>"001001111",
  51537=>"000111010",
  51538=>"011110000",
  51539=>"000000000",
  51540=>"111011000",
  51541=>"111110111",
  51542=>"110111011",
  51543=>"000111111",
  51544=>"111110000",
  51545=>"000000000",
  51546=>"111111011",
  51547=>"000001111",
  51548=>"011111110",
  51549=>"100100110",
  51550=>"111000101",
  51551=>"110111110",
  51552=>"100010000",
  51553=>"001000000",
  51554=>"100110110",
  51555=>"000000000",
  51556=>"111111111",
  51557=>"001001111",
  51558=>"101101111",
  51559=>"111111111",
  51560=>"010010000",
  51561=>"111110000",
  51562=>"111000000",
  51563=>"100110101",
  51564=>"011001001",
  51565=>"000011000",
  51566=>"110111001",
  51567=>"000000000",
  51568=>"111111111",
  51569=>"000000100",
  51570=>"010111111",
  51571=>"011011001",
  51572=>"111110110",
  51573=>"100100000",
  51574=>"000111111",
  51575=>"000110111",
  51576=>"101001000",
  51577=>"111001101",
  51578=>"001101111",
  51579=>"000101111",
  51580=>"111101001",
  51581=>"011000000",
  51582=>"001001010",
  51583=>"111111111",
  51584=>"001000001",
  51585=>"111111001",
  51586=>"000011111",
  51587=>"000000000",
  51588=>"111101101",
  51589=>"000000000",
  51590=>"010110110",
  51591=>"111000000",
  51592=>"011000000",
  51593=>"111111111",
  51594=>"001001001",
  51595=>"000000000",
  51596=>"000000111",
  51597=>"011011100",
  51598=>"111111110",
  51599=>"100010010",
  51600=>"111000000",
  51601=>"000000001",
  51602=>"100000111",
  51603=>"111111111",
  51604=>"000000001",
  51605=>"111111100",
  51606=>"000010111",
  51607=>"111111111",
  51608=>"110100000",
  51609=>"011001001",
  51610=>"000000000",
  51611=>"100101000",
  51612=>"000000001",
  51613=>"111001100",
  51614=>"111001010",
  51615=>"000000010",
  51616=>"111111111",
  51617=>"010010000",
  51618=>"000111110",
  51619=>"111111000",
  51620=>"000010010",
  51621=>"000000001",
  51622=>"000100000",
  51623=>"111111111",
  51624=>"001000000",
  51625=>"110111111",
  51626=>"111000000",
  51627=>"011100111",
  51628=>"000111111",
  51629=>"000101111",
  51630=>"000000100",
  51631=>"000000000",
  51632=>"000111110",
  51633=>"001000000",
  51634=>"111111111",
  51635=>"111111101",
  51636=>"000000000",
  51637=>"000000010",
  51638=>"111110000",
  51639=>"100111111",
  51640=>"000000000",
  51641=>"001001000",
  51642=>"001001101",
  51643=>"000100101",
  51644=>"100000000",
  51645=>"000010010",
  51646=>"000000000",
  51647=>"010010010",
  51648=>"001000000",
  51649=>"000000000",
  51650=>"000000000",
  51651=>"000000000",
  51652=>"110000010",
  51653=>"000100000",
  51654=>"111111000",
  51655=>"111111100",
  51656=>"000000000",
  51657=>"000110000",
  51658=>"000111111",
  51659=>"000000000",
  51660=>"001011011",
  51661=>"000010110",
  51662=>"111100101",
  51663=>"101100100",
  51664=>"101100000",
  51665=>"000110111",
  51666=>"001111011",
  51667=>"011111111",
  51668=>"000000000",
  51669=>"011010111",
  51670=>"111101000",
  51671=>"100100101",
  51672=>"010111001",
  51673=>"111110111",
  51674=>"100100101",
  51675=>"011000001",
  51676=>"010000000",
  51677=>"110111111",
  51678=>"000000100",
  51679=>"000000011",
  51680=>"111100000",
  51681=>"111111111",
  51682=>"000000011",
  51683=>"111011010",
  51684=>"100000000",
  51685=>"000000111",
  51686=>"000000111",
  51687=>"111111111",
  51688=>"111111111",
  51689=>"001111111",
  51690=>"001111111",
  51691=>"111000001",
  51692=>"000111111",
  51693=>"111111001",
  51694=>"001011111",
  51695=>"111011011",
  51696=>"000000000",
  51697=>"111111000",
  51698=>"000111111",
  51699=>"000000000",
  51700=>"000010011",
  51701=>"101111111",
  51702=>"111111110",
  51703=>"011011011",
  51704=>"000000000",
  51705=>"001001001",
  51706=>"111100100",
  51707=>"011011000",
  51708=>"111111101",
  51709=>"111001000",
  51710=>"011111111",
  51711=>"000000000",
  51712=>"000000100",
  51713=>"000001000",
  51714=>"111111010",
  51715=>"000100111",
  51716=>"000000100",
  51717=>"001111111",
  51718=>"111111000",
  51719=>"111000000",
  51720=>"000000000",
  51721=>"111111111",
  51722=>"001000100",
  51723=>"111111111",
  51724=>"110110100",
  51725=>"111111111",
  51726=>"100111011",
  51727=>"000001011",
  51728=>"111101111",
  51729=>"000011000",
  51730=>"000000100",
  51731=>"011111011",
  51732=>"101101111",
  51733=>"111111111",
  51734=>"001111111",
  51735=>"111111100",
  51736=>"001000001",
  51737=>"110110111",
  51738=>"001000111",
  51739=>"111011000",
  51740=>"000000000",
  51741=>"111111000",
  51742=>"000011011",
  51743=>"100000000",
  51744=>"111111000",
  51745=>"100110111",
  51746=>"001001001",
  51747=>"001001001",
  51748=>"111111111",
  51749=>"111111111",
  51750=>"000000000",
  51751=>"000001111",
  51752=>"000000000",
  51753=>"111111111",
  51754=>"001000000",
  51755=>"111100101",
  51756=>"000000000",
  51757=>"000110000",
  51758=>"000000000",
  51759=>"100001111",
  51760=>"111000001",
  51761=>"101101000",
  51762=>"001001000",
  51763=>"111111011",
  51764=>"101001001",
  51765=>"010000000",
  51766=>"001000000",
  51767=>"111111111",
  51768=>"000000000",
  51769=>"000000011",
  51770=>"111000101",
  51771=>"000000000",
  51772=>"101000000",
  51773=>"000000000",
  51774=>"111111111",
  51775=>"000000111",
  51776=>"000010000",
  51777=>"110110110",
  51778=>"111111111",
  51779=>"000101111",
  51780=>"110100000",
  51781=>"111110000",
  51782=>"010110000",
  51783=>"000000000",
  51784=>"111111011",
  51785=>"111000000",
  51786=>"111111111",
  51787=>"001000111",
  51788=>"000001111",
  51789=>"110110000",
  51790=>"001100100",
  51791=>"111111111",
  51792=>"111111111",
  51793=>"001000111",
  51794=>"000000000",
  51795=>"100100000",
  51796=>"111000000",
  51797=>"101001110",
  51798=>"000011111",
  51799=>"001001111",
  51800=>"010001000",
  51801=>"111001011",
  51802=>"000011111",
  51803=>"111100111",
  51804=>"000000010",
  51805=>"000000000",
  51806=>"111110011",
  51807=>"000011011",
  51808=>"110010000",
  51809=>"111100111",
  51810=>"011111100",
  51811=>"000101111",
  51812=>"100100110",
  51813=>"111111011",
  51814=>"001000101",
  51815=>"000000000",
  51816=>"000100000",
  51817=>"111111011",
  51818=>"110001111",
  51819=>"000000000",
  51820=>"001111100",
  51821=>"001000001",
  51822=>"000000001",
  51823=>"000000000",
  51824=>"000001000",
  51825=>"010010111",
  51826=>"000000000",
  51827=>"000000000",
  51828=>"000000000",
  51829=>"000100110",
  51830=>"111111111",
  51831=>"001000000",
  51832=>"011111110",
  51833=>"000000111",
  51834=>"000001001",
  51835=>"101000000",
  51836=>"100110100",
  51837=>"111101111",
  51838=>"000000000",
  51839=>"111000000",
  51840=>"000001111",
  51841=>"111111111",
  51842=>"010000000",
  51843=>"011011001",
  51844=>"000000001",
  51845=>"000000000",
  51846=>"111100100",
  51847=>"010000000",
  51848=>"101000000",
  51849=>"110000111",
  51850=>"110010000",
  51851=>"000000000",
  51852=>"000000101",
  51853=>"001000000",
  51854=>"000010011",
  51855=>"000111111",
  51856=>"111011000",
  51857=>"000000000",
  51858=>"001110111",
  51859=>"110110100",
  51860=>"110110000",
  51861=>"111000110",
  51862=>"110111111",
  51863=>"001111111",
  51864=>"000000000",
  51865=>"111111111",
  51866=>"101001000",
  51867=>"000011011",
  51868=>"101001111",
  51869=>"111101000",
  51870=>"000000111",
  51871=>"000000111",
  51872=>"111111111",
  51873=>"010100000",
  51874=>"111111000",
  51875=>"111111000",
  51876=>"000100000",
  51877=>"111111111",
  51878=>"000100111",
  51879=>"001001111",
  51880=>"110101000",
  51881=>"000111111",
  51882=>"000000000",
  51883=>"111111111",
  51884=>"000001111",
  51885=>"001001011",
  51886=>"000000000",
  51887=>"110000000",
  51888=>"010111010",
  51889=>"111110010",
  51890=>"111111011",
  51891=>"001000111",
  51892=>"111111111",
  51893=>"001111111",
  51894=>"111111111",
  51895=>"100101011",
  51896=>"000001000",
  51897=>"000010000",
  51898=>"000000000",
  51899=>"000000011",
  51900=>"101111111",
  51901=>"111111110",
  51902=>"111101000",
  51903=>"001111111",
  51904=>"111110010",
  51905=>"000000000",
  51906=>"111111111",
  51907=>"000000000",
  51908=>"111111111",
  51909=>"001001001",
  51910=>"111000011",
  51911=>"000000000",
  51912=>"000111111",
  51913=>"001000000",
  51914=>"000000000",
  51915=>"000000010",
  51916=>"111111001",
  51917=>"111111000",
  51918=>"111101111",
  51919=>"111110111",
  51920=>"000011111",
  51921=>"000000000",
  51922=>"000000000",
  51923=>"101000000",
  51924=>"000100100",
  51925=>"111111011",
  51926=>"000000000",
  51927=>"111111101",
  51928=>"001000001",
  51929=>"111110111",
  51930=>"111111111",
  51931=>"111111101",
  51932=>"110111111",
  51933=>"111111111",
  51934=>"000111111",
  51935=>"000000001",
  51936=>"000000011",
  51937=>"010111110",
  51938=>"001111111",
  51939=>"000011001",
  51940=>"000010011",
  51941=>"111100110",
  51942=>"111110111",
  51943=>"111110000",
  51944=>"000000000",
  51945=>"000000000",
  51946=>"111000000",
  51947=>"101111001",
  51948=>"001001111",
  51949=>"101001000",
  51950=>"000010011",
  51951=>"011001000",
  51952=>"111101111",
  51953=>"111101101",
  51954=>"000011011",
  51955=>"001111111",
  51956=>"100000000",
  51957=>"100110100",
  51958=>"001001001",
  51959=>"111111001",
  51960=>"111111111",
  51961=>"001000000",
  51962=>"000000100",
  51963=>"111111000",
  51964=>"011100110",
  51965=>"000000100",
  51966=>"000000011",
  51967=>"101000111",
  51968=>"111111100",
  51969=>"101100000",
  51970=>"111111001",
  51971=>"000000000",
  51972=>"111111010",
  51973=>"000000110",
  51974=>"100111011",
  51975=>"111111100",
  51976=>"000010000",
  51977=>"000000000",
  51978=>"111111111",
  51979=>"010010000",
  51980=>"111010000",
  51981=>"000000000",
  51982=>"111111111",
  51983=>"000000111",
  51984=>"111101111",
  51985=>"111111001",
  51986=>"101100111",
  51987=>"001111111",
  51988=>"111111111",
  51989=>"000000000",
  51990=>"001001001",
  51991=>"000000001",
  51992=>"010010101",
  51993=>"000101111",
  51994=>"101100101",
  51995=>"000000111",
  51996=>"110111111",
  51997=>"110111000",
  51998=>"000000000",
  51999=>"000000000",
  52000=>"000001001",
  52001=>"000000000",
  52002=>"111010010",
  52003=>"001001001",
  52004=>"000100100",
  52005=>"111111111",
  52006=>"101111011",
  52007=>"110100101",
  52008=>"000000100",
  52009=>"111111111",
  52010=>"110000000",
  52011=>"111111011",
  52012=>"111110111",
  52013=>"101101011",
  52014=>"000000000",
  52015=>"111100000",
  52016=>"001111111",
  52017=>"111000000",
  52018=>"001001000",
  52019=>"000000111",
  52020=>"101100100",
  52021=>"011111111",
  52022=>"011010111",
  52023=>"001001001",
  52024=>"000010000",
  52025=>"001001000",
  52026=>"011011111",
  52027=>"000000000",
  52028=>"000000000",
  52029=>"111111000",
  52030=>"000000010",
  52031=>"000100111",
  52032=>"000010000",
  52033=>"111111111",
  52034=>"000000000",
  52035=>"001011111",
  52036=>"110110000",
  52037=>"000111111",
  52038=>"001000000",
  52039=>"000000000",
  52040=>"000000101",
  52041=>"000000000",
  52042=>"001001001",
  52043=>"001111011",
  52044=>"110100111",
  52045=>"000010110",
  52046=>"111111111",
  52047=>"000100100",
  52048=>"011011011",
  52049=>"000000001",
  52050=>"111000000",
  52051=>"000000000",
  52052=>"111111000",
  52053=>"001001001",
  52054=>"000000101",
  52055=>"000111111",
  52056=>"000001000",
  52057=>"011111001",
  52058=>"000001011",
  52059=>"111111010",
  52060=>"010111111",
  52061=>"000110111",
  52062=>"110100111",
  52063=>"101000000",
  52064=>"001111111",
  52065=>"101100100",
  52066=>"000110111",
  52067=>"001110110",
  52068=>"000000000",
  52069=>"000000100",
  52070=>"000001111",
  52071=>"100000000",
  52072=>"100110110",
  52073=>"110110011",
  52074=>"011010000",
  52075=>"000111111",
  52076=>"111110110",
  52077=>"000000000",
  52078=>"100100101",
  52079=>"000000000",
  52080=>"000000000",
  52081=>"111111010",
  52082=>"111000001",
  52083=>"010111000",
  52084=>"000000000",
  52085=>"000000000",
  52086=>"000000000",
  52087=>"011001001",
  52088=>"000100100",
  52089=>"000100110",
  52090=>"101000111",
  52091=>"111111111",
  52092=>"111000000",
  52093=>"111101111",
  52094=>"011000101",
  52095=>"000000001",
  52096=>"110110000",
  52097=>"000000000",
  52098=>"111111111",
  52099=>"111101101",
  52100=>"111000111",
  52101=>"011111111",
  52102=>"101101000",
  52103=>"111111111",
  52104=>"111101111",
  52105=>"100000010",
  52106=>"000000101",
  52107=>"111111011",
  52108=>"000000111",
  52109=>"001111001",
  52110=>"101111111",
  52111=>"111101000",
  52112=>"000000000",
  52113=>"111111100",
  52114=>"000000000",
  52115=>"100100100",
  52116=>"010010000",
  52117=>"000010110",
  52118=>"000000000",
  52119=>"000100110",
  52120=>"111111000",
  52121=>"001011000",
  52122=>"000000000",
  52123=>"111111111",
  52124=>"000000001",
  52125=>"000000000",
  52126=>"111111000",
  52127=>"111111001",
  52128=>"111111011",
  52129=>"000000011",
  52130=>"111000000",
  52131=>"000110000",
  52132=>"111010000",
  52133=>"010111110",
  52134=>"001001001",
  52135=>"000111101",
  52136=>"000000000",
  52137=>"000101111",
  52138=>"111111111",
  52139=>"000000000",
  52140=>"101101111",
  52141=>"111011001",
  52142=>"000000000",
  52143=>"000000000",
  52144=>"100100100",
  52145=>"111111011",
  52146=>"000000000",
  52147=>"000000011",
  52148=>"000000111",
  52149=>"111000100",
  52150=>"000101000",
  52151=>"101100101",
  52152=>"000000111",
  52153=>"001111011",
  52154=>"110000000",
  52155=>"111101101",
  52156=>"110111111",
  52157=>"111111111",
  52158=>"111000000",
  52159=>"000100000",
  52160=>"000000100",
  52161=>"111111111",
  52162=>"000000000",
  52163=>"111011010",
  52164=>"000111101",
  52165=>"000000000",
  52166=>"000001111",
  52167=>"010110000",
  52168=>"011000000",
  52169=>"000000000",
  52170=>"101100101",
  52171=>"111001111",
  52172=>"000000111",
  52173=>"000111111",
  52174=>"101000001",
  52175=>"000000001",
  52176=>"100110111",
  52177=>"111101011",
  52178=>"000100110",
  52179=>"000000000",
  52180=>"101101001",
  52181=>"110111100",
  52182=>"000000111",
  52183=>"001011001",
  52184=>"101011011",
  52185=>"000000111",
  52186=>"001001101",
  52187=>"000010000",
  52188=>"111111011",
  52189=>"000000000",
  52190=>"111110100",
  52191=>"110110010",
  52192=>"100000000",
  52193=>"111111111",
  52194=>"000000000",
  52195=>"000000111",
  52196=>"111011011",
  52197=>"111011000",
  52198=>"100000000",
  52199=>"000000101",
  52200=>"111111101",
  52201=>"111111111",
  52202=>"111000000",
  52203=>"111111000",
  52204=>"011001000",
  52205=>"000000100",
  52206=>"000000111",
  52207=>"001100101",
  52208=>"111111110",
  52209=>"111111111",
  52210=>"111011001",
  52211=>"111111011",
  52212=>"101000011",
  52213=>"110100000",
  52214=>"001000101",
  52215=>"000000000",
  52216=>"011111110",
  52217=>"001001000",
  52218=>"111000000",
  52219=>"111111111",
  52220=>"011011111",
  52221=>"111111111",
  52222=>"111011000",
  52223=>"111111111",
  52224=>"000000111",
  52225=>"011001000",
  52226=>"001000000",
  52227=>"011111111",
  52228=>"100000111",
  52229=>"110101111",
  52230=>"000000000",
  52231=>"111001111",
  52232=>"100100000",
  52233=>"111010000",
  52234=>"000000000",
  52235=>"001000000",
  52236=>"001000000",
  52237=>"100111111",
  52238=>"011011000",
  52239=>"000000000",
  52240=>"000110111",
  52241=>"000100000",
  52242=>"111111111",
  52243=>"001000100",
  52244=>"111111111",
  52245=>"000000000",
  52246=>"000000000",
  52247=>"111111101",
  52248=>"110111111",
  52249=>"001001000",
  52250=>"001000000",
  52251=>"000000001",
  52252=>"111111111",
  52253=>"001000000",
  52254=>"000000000",
  52255=>"100100000",
  52256=>"000000001",
  52257=>"111111011",
  52258=>"000000000",
  52259=>"000000000",
  52260=>"000000000",
  52261=>"111111000",
  52262=>"111111111",
  52263=>"000000000",
  52264=>"001000011",
  52265=>"011111111",
  52266=>"000000111",
  52267=>"111000001",
  52268=>"000000000",
  52269=>"000000100",
  52270=>"111111101",
  52271=>"001000001",
  52272=>"000111110",
  52273=>"000000111",
  52274=>"000000000",
  52275=>"001110100",
  52276=>"000001101",
  52277=>"000000000",
  52278=>"000000000",
  52279=>"000000000",
  52280=>"000000111",
  52281=>"111111110",
  52282=>"111111111",
  52283=>"000101111",
  52284=>"111011000",
  52285=>"000000000",
  52286=>"000010000",
  52287=>"111000000",
  52288=>"111111111",
  52289=>"101111001",
  52290=>"101000000",
  52291=>"111110011",
  52292=>"000100110",
  52293=>"001001110",
  52294=>"111111111",
  52295=>"000000000",
  52296=>"111010000",
  52297=>"111111111",
  52298=>"111000000",
  52299=>"111010111",
  52300=>"011000000",
  52301=>"111111111",
  52302=>"000011111",
  52303=>"111111110",
  52304=>"000000110",
  52305=>"101000000",
  52306=>"001001101",
  52307=>"001001011",
  52308=>"000100111",
  52309=>"110110111",
  52310=>"000000000",
  52311=>"111111111",
  52312=>"111111111",
  52313=>"100111010",
  52314=>"111111000",
  52315=>"100100000",
  52316=>"000000000",
  52317=>"011000000",
  52318=>"111000000",
  52319=>"000000000",
  52320=>"000001000",
  52321=>"000110110",
  52322=>"111000000",
  52323=>"000000000",
  52324=>"000000000",
  52325=>"000000000",
  52326=>"001000000",
  52327=>"111111100",
  52328=>"000111111",
  52329=>"000000000",
  52330=>"101000101",
  52331=>"001000000",
  52332=>"000100111",
  52333=>"111111111",
  52334=>"111111000",
  52335=>"110100000",
  52336=>"000000000",
  52337=>"000000111",
  52338=>"111111101",
  52339=>"000011010",
  52340=>"000000111",
  52341=>"000000000",
  52342=>"100100011",
  52343=>"000000000",
  52344=>"111111111",
  52345=>"110100000",
  52346=>"000000110",
  52347=>"111111111",
  52348=>"100000100",
  52349=>"001001111",
  52350=>"111000000",
  52351=>"111111111",
  52352=>"000000000",
  52353=>"111111111",
  52354=>"111111110",
  52355=>"110100110",
  52356=>"000110110",
  52357=>"000000111",
  52358=>"111011000",
  52359=>"000000000",
  52360=>"111111111",
  52361=>"000000000",
  52362=>"110111000",
  52363=>"000000000",
  52364=>"000000000",
  52365=>"111111111",
  52366=>"111111111",
  52367=>"000000000",
  52368=>"000000111",
  52369=>"000100001",
  52370=>"000000110",
  52371=>"011011001",
  52372=>"100111111",
  52373=>"110100100",
  52374=>"111111111",
  52375=>"111000000",
  52376=>"000001101",
  52377=>"111001100",
  52378=>"001000000",
  52379=>"000011111",
  52380=>"100110111",
  52381=>"000011111",
  52382=>"111111111",
  52383=>"111111111",
  52384=>"111101001",
  52385=>"000110110",
  52386=>"000000010",
  52387=>"111111111",
  52388=>"011001101",
  52389=>"111111000",
  52390=>"100000000",
  52391=>"000110110",
  52392=>"000000111",
  52393=>"111111000",
  52394=>"111000110",
  52395=>"000000000",
  52396=>"000011011",
  52397=>"000000000",
  52398=>"001000001",
  52399=>"000000001",
  52400=>"111111111",
  52401=>"111101100",
  52402=>"111011010",
  52403=>"000000000",
  52404=>"000000000",
  52405=>"100111111",
  52406=>"001101111",
  52407=>"111111111",
  52408=>"100111100",
  52409=>"000000111",
  52410=>"000000111",
  52411=>"000000000",
  52412=>"000000111",
  52413=>"100100000",
  52414=>"000100111",
  52415=>"000000000",
  52416=>"001000001",
  52417=>"010000000",
  52418=>"011000001",
  52419=>"101111111",
  52420=>"111111111",
  52421=>"001000111",
  52422=>"100111111",
  52423=>"000011111",
  52424=>"000110111",
  52425=>"111100100",
  52426=>"000000000",
  52427=>"000000000",
  52428=>"001111110",
  52429=>"000000000",
  52430=>"111111000",
  52431=>"111001001",
  52432=>"000000011",
  52433=>"000000000",
  52434=>"000000000",
  52435=>"111001111",
  52436=>"111000000",
  52437=>"000000101",
  52438=>"000000010",
  52439=>"010011011",
  52440=>"111111111",
  52441=>"100111100",
  52442=>"110010000",
  52443=>"000000111",
  52444=>"011011111",
  52445=>"010010000",
  52446=>"000011111",
  52447=>"000110111",
  52448=>"000000000",
  52449=>"000100111",
  52450=>"111010001",
  52451=>"100100100",
  52452=>"100111000",
  52453=>"001000100",
  52454=>"111111111",
  52455=>"000001111",
  52456=>"011011000",
  52457=>"110010000",
  52458=>"110110111",
  52459=>"000111111",
  52460=>"000110100",
  52461=>"000100111",
  52462=>"000000000",
  52463=>"000000000",
  52464=>"111111011",
  52465=>"111111000",
  52466=>"111111111",
  52467=>"001001111",
  52468=>"000100100",
  52469=>"001000000",
  52470=>"010111111",
  52471=>"111111111",
  52472=>"001001000",
  52473=>"000000000",
  52474=>"111111111",
  52475=>"111111110",
  52476=>"000100111",
  52477=>"000011111",
  52478=>"000110001",
  52479=>"111111111",
  52480=>"011001001",
  52481=>"011010010",
  52482=>"000000111",
  52483=>"000000000",
  52484=>"000111111",
  52485=>"110100000",
  52486=>"000000000",
  52487=>"000000000",
  52488=>"110111111",
  52489=>"110000000",
  52490=>"111011001",
  52491=>"000100000",
  52492=>"111111111",
  52493=>"000000000",
  52494=>"111110000",
  52495=>"000000110",
  52496=>"111111111",
  52497=>"000000000",
  52498=>"111100111",
  52499=>"111010110",
  52500=>"111001011",
  52501=>"110111011",
  52502=>"000111111",
  52503=>"111111111",
  52504=>"000000001",
  52505=>"111101001",
  52506=>"010000000",
  52507=>"000100011",
  52508=>"111111010",
  52509=>"100100111",
  52510=>"000000000",
  52511=>"111111000",
  52512=>"000111000",
  52513=>"100101001",
  52514=>"111001111",
  52515=>"001001101",
  52516=>"000000000",
  52517=>"110111111",
  52518=>"001111111",
  52519=>"100111111",
  52520=>"010111010",
  52521=>"101001001",
  52522=>"000110000",
  52523=>"100111111",
  52524=>"000000111",
  52525=>"110111111",
  52526=>"000111111",
  52527=>"001111111",
  52528=>"110111111",
  52529=>"000000111",
  52530=>"100000000",
  52531=>"110111111",
  52532=>"101000000",
  52533=>"111111111",
  52534=>"111111001",
  52535=>"111000000",
  52536=>"000000111",
  52537=>"111111111",
  52538=>"000100111",
  52539=>"111111111",
  52540=>"010010000",
  52541=>"111111001",
  52542=>"111111111",
  52543=>"000100100",
  52544=>"010000000",
  52545=>"001000001",
  52546=>"000000000",
  52547=>"111000111",
  52548=>"110111011",
  52549=>"000101101",
  52550=>"000000000",
  52551=>"111101111",
  52552=>"000000010",
  52553=>"000000000",
  52554=>"111111000",
  52555=>"000111111",
  52556=>"000000111",
  52557=>"000111000",
  52558=>"111111111",
  52559=>"100100000",
  52560=>"111111011",
  52561=>"111111000",
  52562=>"111111011",
  52563=>"000000110",
  52564=>"000000000",
  52565=>"001000000",
  52566=>"111111111",
  52567=>"000000000",
  52568=>"000000000",
  52569=>"000000000",
  52570=>"111111011",
  52571=>"111111111",
  52572=>"111111100",
  52573=>"111111011",
  52574=>"111011111",
  52575=>"111111111",
  52576=>"000111001",
  52577=>"111111001",
  52578=>"011001000",
  52579=>"000000000",
  52580=>"000100100",
  52581=>"111111111",
  52582=>"000000000",
  52583=>"000000110",
  52584=>"000001000",
  52585=>"000000010",
  52586=>"111111100",
  52587=>"000000001",
  52588=>"110010000",
  52589=>"111001111",
  52590=>"001011001",
  52591=>"110000000",
  52592=>"010000000",
  52593=>"000110100",
  52594=>"011111111",
  52595=>"000000011",
  52596=>"011111111",
  52597=>"001001001",
  52598=>"110110100",
  52599=>"000111111",
  52600=>"111111001",
  52601=>"000111111",
  52602=>"000000001",
  52603=>"011111000",
  52604=>"111110000",
  52605=>"111100000",
  52606=>"111010000",
  52607=>"111111001",
  52608=>"001011000",
  52609=>"110011011",
  52610=>"000000000",
  52611=>"111111000",
  52612=>"000000111",
  52613=>"111101101",
  52614=>"111110000",
  52615=>"000010110",
  52616=>"010000000",
  52617=>"000000000",
  52618=>"010100100",
  52619=>"110111111",
  52620=>"111111111",
  52621=>"111011000",
  52622=>"000100111",
  52623=>"011000000",
  52624=>"000000111",
  52625=>"111111111",
  52626=>"110110111",
  52627=>"100000000",
  52628=>"011111000",
  52629=>"010111111",
  52630=>"111110111",
  52631=>"000000000",
  52632=>"000000001",
  52633=>"010010010",
  52634=>"111111111",
  52635=>"100010111",
  52636=>"000000111",
  52637=>"001000011",
  52638=>"100000101",
  52639=>"000000000",
  52640=>"000111111",
  52641=>"011001000",
  52642=>"000000000",
  52643=>"100100000",
  52644=>"111100100",
  52645=>"000111111",
  52646=>"100000000",
  52647=>"000000000",
  52648=>"000000000",
  52649=>"000100110",
  52650=>"000001000",
  52651=>"111111111",
  52652=>"000000000",
  52653=>"111111100",
  52654=>"000100111",
  52655=>"111111000",
  52656=>"000110000",
  52657=>"000000111",
  52658=>"100111100",
  52659=>"111111111",
  52660=>"000000011",
  52661=>"001111111",
  52662=>"111111101",
  52663=>"111111000",
  52664=>"000110000",
  52665=>"111111010",
  52666=>"111111111",
  52667=>"111101111",
  52668=>"111111111",
  52669=>"111000100",
  52670=>"100111111",
  52671=>"000000000",
  52672=>"000000000",
  52673=>"111110000",
  52674=>"000000111",
  52675=>"111111111",
  52676=>"000000000",
  52677=>"000000000",
  52678=>"100000111",
  52679=>"111111111",
  52680=>"111111111",
  52681=>"111110111",
  52682=>"101101101",
  52683=>"111111000",
  52684=>"111111000",
  52685=>"101000000",
  52686=>"000000010",
  52687=>"100000010",
  52688=>"000111111",
  52689=>"000100111",
  52690=>"111110000",
  52691=>"010010000",
  52692=>"100100110",
  52693=>"111111011",
  52694=>"000000111",
  52695=>"100000000",
  52696=>"100000001",
  52697=>"000000101",
  52698=>"000010111",
  52699=>"100000000",
  52700=>"010111111",
  52701=>"000000011",
  52702=>"110100110",
  52703=>"000010000",
  52704=>"000000000",
  52705=>"000000000",
  52706=>"000010000",
  52707=>"101111111",
  52708=>"000010011",
  52709=>"000000000",
  52710=>"000000100",
  52711=>"110110111",
  52712=>"111010000",
  52713=>"000000110",
  52714=>"111111111",
  52715=>"001000000",
  52716=>"100001000",
  52717=>"100000000",
  52718=>"000000100",
  52719=>"100100111",
  52720=>"000000111",
  52721=>"111111000",
  52722=>"011000111",
  52723=>"100111111",
  52724=>"111111111",
  52725=>"111100111",
  52726=>"000000000",
  52727=>"000000000",
  52728=>"000100000",
  52729=>"000001011",
  52730=>"111110111",
  52731=>"000010111",
  52732=>"011111111",
  52733=>"000000110",
  52734=>"111111000",
  52735=>"100000000",
  52736=>"000000001",
  52737=>"010000000",
  52738=>"101101101",
  52739=>"111111111",
  52740=>"000000010",
  52741=>"000000111",
  52742=>"000000000",
  52743=>"000000111",
  52744=>"111111000",
  52745=>"011011111",
  52746=>"000000101",
  52747=>"111111111",
  52748=>"010110111",
  52749=>"000000000",
  52750=>"100100111",
  52751=>"000000000",
  52752=>"110111110",
  52753=>"000000000",
  52754=>"011001000",
  52755=>"000000111",
  52756=>"001100000",
  52757=>"000110111",
  52758=>"001111111",
  52759=>"011011011",
  52760=>"100100111",
  52761=>"111000000",
  52762=>"111111110",
  52763=>"100100001",
  52764=>"111000000",
  52765=>"000110111",
  52766=>"111111111",
  52767=>"110110100",
  52768=>"100000000",
  52769=>"101111111",
  52770=>"000000000",
  52771=>"001000111",
  52772=>"000000000",
  52773=>"010010000",
  52774=>"110000000",
  52775=>"110110100",
  52776=>"001000000",
  52777=>"000000000",
  52778=>"000000000",
  52779=>"000000100",
  52780=>"000000000",
  52781=>"110000000",
  52782=>"011011011",
  52783=>"111111111",
  52784=>"010111000",
  52785=>"001101000",
  52786=>"000110010",
  52787=>"000111100",
  52788=>"000000000",
  52789=>"100000101",
  52790=>"001001111",
  52791=>"111111100",
  52792=>"100000000",
  52793=>"110100110",
  52794=>"000000000",
  52795=>"000010000",
  52796=>"001000000",
  52797=>"110110111",
  52798=>"101111111",
  52799=>"000001011",
  52800=>"111111111",
  52801=>"111011011",
  52802=>"000110000",
  52803=>"000001011",
  52804=>"000001001",
  52805=>"001000000",
  52806=>"110110100",
  52807=>"111111111",
  52808=>"111111000",
  52809=>"111111111",
  52810=>"000111010",
  52811=>"101101001",
  52812=>"010110000",
  52813=>"111111111",
  52814=>"011111111",
  52815=>"000000000",
  52816=>"111111111",
  52817=>"011011011",
  52818=>"110111000",
  52819=>"001000000",
  52820=>"000000111",
  52821=>"110111110",
  52822=>"101101000",
  52823=>"111111111",
  52824=>"000000000",
  52825=>"111001111",
  52826=>"000111111",
  52827=>"110111111",
  52828=>"100000000",
  52829=>"000000000",
  52830=>"000010111",
  52831=>"111111010",
  52832=>"000000111",
  52833=>"011111111",
  52834=>"111111111",
  52835=>"111111111",
  52836=>"001001000",
  52837=>"011000111",
  52838=>"000100111",
  52839=>"010000000",
  52840=>"111111001",
  52841=>"000000000",
  52842=>"000000000",
  52843=>"011111111",
  52844=>"101001011",
  52845=>"000000000",
  52846=>"111111000",
  52847=>"111111000",
  52848=>"000111111",
  52849=>"110000000",
  52850=>"111111111",
  52851=>"111111000",
  52852=>"111111100",
  52853=>"000000000",
  52854=>"011111000",
  52855=>"001001111",
  52856=>"000000000",
  52857=>"000000001",
  52858=>"101101100",
  52859=>"000001001",
  52860=>"011001100",
  52861=>"000010000",
  52862=>"111111010",
  52863=>"101000000",
  52864=>"111111111",
  52865=>"010111111",
  52866=>"000000100",
  52867=>"000000000",
  52868=>"001000000",
  52869=>"000000000",
  52870=>"110110000",
  52871=>"000000000",
  52872=>"111100000",
  52873=>"011110111",
  52874=>"111111110",
  52875=>"111111001",
  52876=>"110111111",
  52877=>"111111111",
  52878=>"111111111",
  52879=>"110111111",
  52880=>"000000000",
  52881=>"100010110",
  52882=>"111111110",
  52883=>"111111011",
  52884=>"010001000",
  52885=>"111100100",
  52886=>"111111111",
  52887=>"001000000",
  52888=>"000000000",
  52889=>"000000000",
  52890=>"011000000",
  52891=>"010000000",
  52892=>"000000000",
  52893=>"001000101",
  52894=>"111111111",
  52895=>"000000001",
  52896=>"001000110",
  52897=>"000001100",
  52898=>"000000000",
  52899=>"000000101",
  52900=>"111111101",
  52901=>"100110110",
  52902=>"000000111",
  52903=>"011011011",
  52904=>"111111011",
  52905=>"001111111",
  52906=>"000000000",
  52907=>"000001111",
  52908=>"000000000",
  52909=>"111100101",
  52910=>"000010000",
  52911=>"100110100",
  52912=>"000000000",
  52913=>"000000000",
  52914=>"011111011",
  52915=>"111111111",
  52916=>"110111111",
  52917=>"110111110",
  52918=>"111111111",
  52919=>"111111111",
  52920=>"000000110",
  52921=>"000000000",
  52922=>"111111101",
  52923=>"100100111",
  52924=>"001000001",
  52925=>"000000000",
  52926=>"001011111",
  52927=>"111011000",
  52928=>"111100111",
  52929=>"000000000",
  52930=>"100100100",
  52931=>"000000000",
  52932=>"011011111",
  52933=>"000010010",
  52934=>"000000100",
  52935=>"101100001",
  52936=>"111111111",
  52937=>"101111111",
  52938=>"000011001",
  52939=>"000000000",
  52940=>"110110111",
  52941=>"111111110",
  52942=>"000000010",
  52943=>"000000000",
  52944=>"000001100",
  52945=>"011011011",
  52946=>"010111111",
  52947=>"000000001",
  52948=>"000110100",
  52949=>"000000000",
  52950=>"111011011",
  52951=>"000000000",
  52952=>"111101111",
  52953=>"100100100",
  52954=>"000000101",
  52955=>"111111110",
  52956=>"111111101",
  52957=>"000111111",
  52958=>"000000111",
  52959=>"011110111",
  52960=>"000000000",
  52961=>"000000010",
  52962=>"000000000",
  52963=>"111110000",
  52964=>"011011100",
  52965=>"111101101",
  52966=>"111111011",
  52967=>"111111101",
  52968=>"001001000",
  52969=>"000000001",
  52970=>"001101111",
  52971=>"000000111",
  52972=>"010110110",
  52973=>"000110110",
  52974=>"010001111",
  52975=>"001000100",
  52976=>"000000100",
  52977=>"011011011",
  52978=>"000000000",
  52979=>"011010110",
  52980=>"000000000",
  52981=>"111111111",
  52982=>"101111111",
  52983=>"000000000",
  52984=>"111111111",
  52985=>"101100100",
  52986=>"110100000",
  52987=>"000001011",
  52988=>"110101111",
  52989=>"001111111",
  52990=>"000000111",
  52991=>"111111111",
  52992=>"000000000",
  52993=>"111011101",
  52994=>"010111010",
  52995=>"011011000",
  52996=>"000110100",
  52997=>"111101100",
  52998=>"111111111",
  52999=>"111111111",
  53000=>"111110111",
  53001=>"000000000",
  53002=>"000000000",
  53003=>"011000000",
  53004=>"111111111",
  53005=>"100000000",
  53006=>"111010100",
  53007=>"000111111",
  53008=>"110110101",
  53009=>"100100100",
  53010=>"111111110",
  53011=>"111101100",
  53012=>"111011000",
  53013=>"111111111",
  53014=>"100100110",
  53015=>"111111011",
  53016=>"011111010",
  53017=>"111110000",
  53018=>"111111111",
  53019=>"000000000",
  53020=>"011111110",
  53021=>"110111010",
  53022=>"111111111",
  53023=>"110110110",
  53024=>"110110000",
  53025=>"101100000",
  53026=>"100110111",
  53027=>"001000000",
  53028=>"111111111",
  53029=>"011000000",
  53030=>"010011011",
  53031=>"110110010",
  53032=>"111100000",
  53033=>"000000000",
  53034=>"010110110",
  53035=>"011011001",
  53036=>"100101111",
  53037=>"100100100",
  53038=>"111111111",
  53039=>"100000000",
  53040=>"001111111",
  53041=>"101101111",
  53042=>"011111111",
  53043=>"000110111",
  53044=>"111101100",
  53045=>"111110010",
  53046=>"111111101",
  53047=>"111111111",
  53048=>"111111111",
  53049=>"011000000",
  53050=>"111000000",
  53051=>"000000111",
  53052=>"100000000",
  53053=>"101111110",
  53054=>"111101001",
  53055=>"100001111",
  53056=>"000000111",
  53057=>"100010000",
  53058=>"000100000",
  53059=>"010110111",
  53060=>"111111000",
  53061=>"011010000",
  53062=>"000000000",
  53063=>"111111000",
  53064=>"111111111",
  53065=>"011101000",
  53066=>"001110100",
  53067=>"111111111",
  53068=>"000000000",
  53069=>"100000000",
  53070=>"110110111",
  53071=>"111111100",
  53072=>"111101100",
  53073=>"110000000",
  53074=>"000000000",
  53075=>"111111111",
  53076=>"111101001",
  53077=>"001000000",
  53078=>"000000000",
  53079=>"111111111",
  53080=>"000111110",
  53081=>"111111111",
  53082=>"000000111",
  53083=>"001111010",
  53084=>"001000100",
  53085=>"000000000",
  53086=>"111111110",
  53087=>"000000000",
  53088=>"111111110",
  53089=>"111101111",
  53090=>"111111111",
  53091=>"001000000",
  53092=>"011101111",
  53093=>"100100110",
  53094=>"000000000",
  53095=>"011000001",
  53096=>"111110110",
  53097=>"011010000",
  53098=>"000000110",
  53099=>"111111111",
  53100=>"111011001",
  53101=>"001001000",
  53102=>"110100001",
  53103=>"111111000",
  53104=>"011111111",
  53105=>"000001000",
  53106=>"011001001",
  53107=>"000110011",
  53108=>"011111011",
  53109=>"110111111",
  53110=>"001001011",
  53111=>"000000010",
  53112=>"001001111",
  53113=>"000111010",
  53114=>"000000000",
  53115=>"010110000",
  53116=>"000000000",
  53117=>"011011111",
  53118=>"111000111",
  53119=>"101000000",
  53120=>"001001011",
  53121=>"111110111",
  53122=>"100110111",
  53123=>"000111111",
  53124=>"010011011",
  53125=>"000000010",
  53126=>"011110110",
  53127=>"011010011",
  53128=>"001000100",
  53129=>"111111111",
  53130=>"111010011",
  53131=>"011011111",
  53132=>"111111111",
  53133=>"111110100",
  53134=>"100000001",
  53135=>"010111010",
  53136=>"001001101",
  53137=>"000000000",
  53138=>"001111110",
  53139=>"000000000",
  53140=>"000000001",
  53141=>"000010010",
  53142=>"000000000",
  53143=>"001001111",
  53144=>"000101000",
  53145=>"011111111",
  53146=>"111001001",
  53147=>"101111111",
  53148=>"111111111",
  53149=>"110110000",
  53150=>"000000100",
  53151=>"110000000",
  53152=>"000000000",
  53153=>"111111111",
  53154=>"111111111",
  53155=>"001101111",
  53156=>"000001011",
  53157=>"111111010",
  53158=>"000000111",
  53159=>"000000100",
  53160=>"101111110",
  53161=>"111100000",
  53162=>"001011011",
  53163=>"000100100",
  53164=>"111111111",
  53165=>"111111111",
  53166=>"111111110",
  53167=>"001000000",
  53168=>"110111111",
  53169=>"000001111",
  53170=>"100100000",
  53171=>"000100000",
  53172=>"000000000",
  53173=>"111110110",
  53174=>"010011111",
  53175=>"000000001",
  53176=>"100100100",
  53177=>"011001000",
  53178=>"111100100",
  53179=>"110110110",
  53180=>"000000000",
  53181=>"000001001",
  53182=>"111111110",
  53183=>"101111011",
  53184=>"000000000",
  53185=>"111111111",
  53186=>"111111111",
  53187=>"111111110",
  53188=>"000000001",
  53189=>"101001111",
  53190=>"111111111",
  53191=>"100101100",
  53192=>"111111111",
  53193=>"111111111",
  53194=>"001100000",
  53195=>"011110000",
  53196=>"111111101",
  53197=>"111000101",
  53198=>"111111110",
  53199=>"000000111",
  53200=>"011111111",
  53201=>"000111111",
  53202=>"101000000",
  53203=>"111111110",
  53204=>"000100010",
  53205=>"111111111",
  53206=>"111111111",
  53207=>"001000000",
  53208=>"000000000",
  53209=>"011010000",
  53210=>"111111000",
  53211=>"111111111",
  53212=>"000000001",
  53213=>"111111111",
  53214=>"000000000",
  53215=>"100011011",
  53216=>"001000111",
  53217=>"000000000",
  53218=>"110110000",
  53219=>"111111100",
  53220=>"000000000",
  53221=>"111111110",
  53222=>"100100110",
  53223=>"111111001",
  53224=>"100110110",
  53225=>"000100100",
  53226=>"111111111",
  53227=>"001000001",
  53228=>"000110111",
  53229=>"101111011",
  53230=>"111111111",
  53231=>"000011111",
  53232=>"000000100",
  53233=>"000111111",
  53234=>"000000000",
  53235=>"000110110",
  53236=>"001111111",
  53237=>"000000000",
  53238=>"000000000",
  53239=>"111111111",
  53240=>"111111111",
  53241=>"011111110",
  53242=>"011111111",
  53243=>"001000110",
  53244=>"011000000",
  53245=>"100000000",
  53246=>"010010110",
  53247=>"000000101",
  53248=>"111111001",
  53249=>"001111011",
  53250=>"111011000",
  53251=>"111111111",
  53252=>"000000001",
  53253=>"011000000",
  53254=>"111001111",
  53255=>"110000101",
  53256=>"001111111",
  53257=>"100000000",
  53258=>"000000001",
  53259=>"000000001",
  53260=>"111001001",
  53261=>"000000111",
  53262=>"011011011",
  53263=>"000000000",
  53264=>"000000110",
  53265=>"111111000",
  53266=>"000000000",
  53267=>"111011111",
  53268=>"110111000",
  53269=>"000000100",
  53270=>"100100111",
  53271=>"111011111",
  53272=>"111000000",
  53273=>"101001001",
  53274=>"111111111",
  53275=>"000000001",
  53276=>"010011111",
  53277=>"000000000",
  53278=>"111011111",
  53279=>"100000000",
  53280=>"111111001",
  53281=>"100111111",
  53282=>"000011111",
  53283=>"111100000",
  53284=>"110000101",
  53285=>"111001111",
  53286=>"110100100",
  53287=>"010000000",
  53288=>"000000000",
  53289=>"100000000",
  53290=>"000000101",
  53291=>"110100100",
  53292=>"000000000",
  53293=>"111011111",
  53294=>"111111001",
  53295=>"000000000",
  53296=>"100111111",
  53297=>"111111111",
  53298=>"011011111",
  53299=>"100100110",
  53300=>"011111000",
  53301=>"111001000",
  53302=>"000111101",
  53303=>"001100111",
  53304=>"000000101",
  53305=>"110100111",
  53306=>"000000001",
  53307=>"001000011",
  53308=>"100000100",
  53309=>"000011001",
  53310=>"110110100",
  53311=>"000000000",
  53312=>"111111111",
  53313=>"111000000",
  53314=>"110000000",
  53315=>"000000000",
  53316=>"111111011",
  53317=>"000000000",
  53318=>"000001000",
  53319=>"111111111",
  53320=>"011010010",
  53321=>"111000000",
  53322=>"111111010",
  53323=>"001111111",
  53324=>"100100001",
  53325=>"110110110",
  53326=>"000000000",
  53327=>"111111111",
  53328=>"000000000",
  53329=>"110100111",
  53330=>"000000000",
  53331=>"011011110",
  53332=>"000000000",
  53333=>"000000000",
  53334=>"000000110",
  53335=>"111110111",
  53336=>"000000010",
  53337=>"000000000",
  53338=>"110110011",
  53339=>"001011111",
  53340=>"111110110",
  53341=>"100111111",
  53342=>"100100110",
  53343=>"000100000",
  53344=>"100100111",
  53345=>"001001111",
  53346=>"001011010",
  53347=>"111011001",
  53348=>"001001111",
  53349=>"111000000",
  53350=>"010111000",
  53351=>"111111000",
  53352=>"000000111",
  53353=>"000000000",
  53354=>"110111111",
  53355=>"111011000",
  53356=>"011000000",
  53357=>"000111000",
  53358=>"000000111",
  53359=>"000000110",
  53360=>"111111111",
  53361=>"100001000",
  53362=>"111111111",
  53363=>"110111111",
  53364=>"001111011",
  53365=>"111111111",
  53366=>"001000000",
  53367=>"111111000",
  53368=>"100000000",
  53369=>"100100000",
  53370=>"110000000",
  53371=>"001000000",
  53372=>"111011011",
  53373=>"100000100",
  53374=>"100000001",
  53375=>"111111111",
  53376=>"000000000",
  53377=>"001001100",
  53378=>"111110110",
  53379=>"000101111",
  53380=>"000000111",
  53381=>"000000000",
  53382=>"000011001",
  53383=>"100100111",
  53384=>"111111111",
  53385=>"000000100",
  53386=>"110000001",
  53387=>"000111111",
  53388=>"001001000",
  53389=>"000000000",
  53390=>"000000111",
  53391=>"100101111",
  53392=>"111111111",
  53393=>"011100011",
  53394=>"111111111",
  53395=>"111111111",
  53396=>"111101011",
  53397=>"111111110",
  53398=>"111111111",
  53399=>"001000111",
  53400=>"111110110",
  53401=>"111111111",
  53402=>"000000110",
  53403=>"111001001",
  53404=>"100100000",
  53405=>"111111111",
  53406=>"111101000",
  53407=>"111000000",
  53408=>"100000000",
  53409=>"111000000",
  53410=>"001111111",
  53411=>"111100100",
  53412=>"111100001",
  53413=>"111111111",
  53414=>"111110111",
  53415=>"101110110",
  53416=>"111111000",
  53417=>"000001111",
  53418=>"111111111",
  53419=>"111100111",
  53420=>"100000100",
  53421=>"011011000",
  53422=>"111111111",
  53423=>"011001111",
  53424=>"000000000",
  53425=>"111000001",
  53426=>"111111111",
  53427=>"111000111",
  53428=>"000010000",
  53429=>"000000000",
  53430=>"111111000",
  53431=>"101000000",
  53432=>"110111100",
  53433=>"000000000",
  53434=>"100010000",
  53435=>"111000100",
  53436=>"010110010",
  53437=>"110111100",
  53438=>"000000000",
  53439=>"010111111",
  53440=>"111101111",
  53441=>"000000000",
  53442=>"000000000",
  53443=>"000000111",
  53444=>"111111001",
  53445=>"000000001",
  53446=>"111001000",
  53447=>"000000000",
  53448=>"000000100",
  53449=>"011001000",
  53450=>"000110110",
  53451=>"000000000",
  53452=>"000000100",
  53453=>"000000000",
  53454=>"000001101",
  53455=>"001000000",
  53456=>"001000000",
  53457=>"111111111",
  53458=>"011111000",
  53459=>"111111111",
  53460=>"001101111",
  53461=>"101001001",
  53462=>"000000000",
  53463=>"010111110",
  53464=>"101101001",
  53465=>"000110111",
  53466=>"000000000",
  53467=>"000111111",
  53468=>"000000100",
  53469=>"111111111",
  53470=>"001100111",
  53471=>"000001110",
  53472=>"011001111",
  53473=>"111111110",
  53474=>"111111000",
  53475=>"110110110",
  53476=>"111111110",
  53477=>"111100111",
  53478=>"110110111",
  53479=>"110000111",
  53480=>"111111111",
  53481=>"100111111",
  53482=>"110011110",
  53483=>"000000001",
  53484=>"111111111",
  53485=>"000111000",
  53486=>"111011000",
  53487=>"111111001",
  53488=>"110110010",
  53489=>"111111111",
  53490=>"111111111",
  53491=>"110110000",
  53492=>"110101111",
  53493=>"001000000",
  53494=>"111111001",
  53495=>"111111111",
  53496=>"100000001",
  53497=>"100000000",
  53498=>"000000011",
  53499=>"000000000",
  53500=>"000100000",
  53501=>"010011011",
  53502=>"111111111",
  53503=>"000000010",
  53504=>"110000000",
  53505=>"111101101",
  53506=>"000000000",
  53507=>"001100100",
  53508=>"010011111",
  53509=>"001001000",
  53510=>"111000111",
  53511=>"111111111",
  53512=>"110011000",
  53513=>"000000000",
  53514=>"011001111",
  53515=>"000000111",
  53516=>"011111111",
  53517=>"000111111",
  53518=>"110101101",
  53519=>"000011001",
  53520=>"110111110",
  53521=>"100100111",
  53522=>"000000000",
  53523=>"001001000",
  53524=>"111111100",
  53525=>"111001011",
  53526=>"001011001",
  53527=>"001000000",
  53528=>"011001111",
  53529=>"101100111",
  53530=>"001000000",
  53531=>"000000000",
  53532=>"111111101",
  53533=>"111111111",
  53534=>"000000110",
  53535=>"111111111",
  53536=>"001111111",
  53537=>"100101001",
  53538=>"001101000",
  53539=>"011111011",
  53540=>"000101111",
  53541=>"000000001",
  53542=>"111111111",
  53543=>"111001101",
  53544=>"111111111",
  53545=>"110010111",
  53546=>"000001111",
  53547=>"011010000",
  53548=>"111110000",
  53549=>"111101111",
  53550=>"111010010",
  53551=>"000000001",
  53552=>"000000110",
  53553=>"110110100",
  53554=>"101000001",
  53555=>"111110010",
  53556=>"000000000",
  53557=>"111111111",
  53558=>"000010010",
  53559=>"111101001",
  53560=>"000000011",
  53561=>"101011111",
  53562=>"100110111",
  53563=>"011010111",
  53564=>"110110110",
  53565=>"000110111",
  53566=>"111101101",
  53567=>"100001001",
  53568=>"111101000",
  53569=>"111111111",
  53570=>"001000001",
  53571=>"000000000",
  53572=>"000000000",
  53573=>"000110101",
  53574=>"001000000",
  53575=>"111111110",
  53576=>"000100100",
  53577=>"111000000",
  53578=>"001011111",
  53579=>"110000000",
  53580=>"001101111",
  53581=>"000100111",
  53582=>"110111111",
  53583=>"000011011",
  53584=>"111110110",
  53585=>"110111110",
  53586=>"111111111",
  53587=>"000000000",
  53588=>"110011111",
  53589=>"111110010",
  53590=>"111111111",
  53591=>"111111111",
  53592=>"111111111",
  53593=>"000000001",
  53594=>"001000000",
  53595=>"000000100",
  53596=>"000000110",
  53597=>"101000000",
  53598=>"111001000",
  53599=>"110110111",
  53600=>"001001000",
  53601=>"011111110",
  53602=>"111100110",
  53603=>"100111111",
  53604=>"000101111",
  53605=>"000000000",
  53606=>"000111011",
  53607=>"001011100",
  53608=>"101101011",
  53609=>"111111111",
  53610=>"111101101",
  53611=>"100010010",
  53612=>"000011000",
  53613=>"111111110",
  53614=>"000000000",
  53615=>"111001101",
  53616=>"000000100",
  53617=>"111111000",
  53618=>"000001000",
  53619=>"111111101",
  53620=>"111001111",
  53621=>"110110111",
  53622=>"011011011",
  53623=>"000111111",
  53624=>"111111110",
  53625=>"001101101",
  53626=>"000000000",
  53627=>"110110110",
  53628=>"010000001",
  53629=>"110110000",
  53630=>"000010010",
  53631=>"111001001",
  53632=>"001011111",
  53633=>"000001001",
  53634=>"010010000",
  53635=>"110111011",
  53636=>"010010000",
  53637=>"000000000",
  53638=>"000001111",
  53639=>"000000001",
  53640=>"111000001",
  53641=>"110000111",
  53642=>"011000000",
  53643=>"000000001",
  53644=>"101000111",
  53645=>"101101111",
  53646=>"000000000",
  53647=>"110110100",
  53648=>"111111111",
  53649=>"111000000",
  53650=>"111111001",
  53651=>"001011011",
  53652=>"111001100",
  53653=>"000110111",
  53654=>"111111111",
  53655=>"011001001",
  53656=>"111110000",
  53657=>"000000100",
  53658=>"000110111",
  53659=>"001000101",
  53660=>"111111101",
  53661=>"000000000",
  53662=>"001000000",
  53663=>"000000000",
  53664=>"000010000",
  53665=>"111111111",
  53666=>"000000100",
  53667=>"000011111",
  53668=>"111110000",
  53669=>"100000000",
  53670=>"101001001",
  53671=>"011000000",
  53672=>"000000000",
  53673=>"001000000",
  53674=>"111011010",
  53675=>"000000000",
  53676=>"000010000",
  53677=>"000000111",
  53678=>"111111101",
  53679=>"010100111",
  53680=>"111101101",
  53681=>"111111111",
  53682=>"111000111",
  53683=>"000000000",
  53684=>"000101111",
  53685=>"001111101",
  53686=>"111011111",
  53687=>"111001000",
  53688=>"000000000",
  53689=>"000000111",
  53690=>"000000001",
  53691=>"111110110",
  53692=>"000000101",
  53693=>"000111110",
  53694=>"000000000",
  53695=>"111111111",
  53696=>"000100100",
  53697=>"100001111",
  53698=>"000000100",
  53699=>"110000000",
  53700=>"111100110",
  53701=>"111111111",
  53702=>"111101101",
  53703=>"000000000",
  53704=>"111010110",
  53705=>"000000111",
  53706=>"000101110",
  53707=>"000000000",
  53708=>"111110010",
  53709=>"000000001",
  53710=>"001000000",
  53711=>"000000000",
  53712=>"000000000",
  53713=>"111111111",
  53714=>"110111111",
  53715=>"000000111",
  53716=>"000000000",
  53717=>"011000000",
  53718=>"010000000",
  53719=>"110000111",
  53720=>"111101001",
  53721=>"000000100",
  53722=>"000011111",
  53723=>"011111111",
  53724=>"110000101",
  53725=>"111111111",
  53726=>"000011111",
  53727=>"111001110",
  53728=>"011111111",
  53729=>"001000100",
  53730=>"111111111",
  53731=>"000000100",
  53732=>"000000110",
  53733=>"000000000",
  53734=>"111111111",
  53735=>"000000111",
  53736=>"111001001",
  53737=>"000110111",
  53738=>"100111111",
  53739=>"111111100",
  53740=>"011000000",
  53741=>"100100000",
  53742=>"000000000",
  53743=>"101000000",
  53744=>"100111111",
  53745=>"011000000",
  53746=>"111000000",
  53747=>"100000000",
  53748=>"111111111",
  53749=>"000000000",
  53750=>"111110111",
  53751=>"111110110",
  53752=>"011000111",
  53753=>"111100110",
  53754=>"000011011",
  53755=>"000000000",
  53756=>"000000000",
  53757=>"001000000",
  53758=>"000000100",
  53759=>"011000000",
  53760=>"111100001",
  53761=>"000000011",
  53762=>"100100100",
  53763=>"000000111",
  53764=>"011011111",
  53765=>"111111011",
  53766=>"111111111",
  53767=>"000100110",
  53768=>"000111111",
  53769=>"000000000",
  53770=>"100000000",
  53771=>"000001001",
  53772=>"111101101",
  53773=>"000100111",
  53774=>"010000100",
  53775=>"111001000",
  53776=>"100100110",
  53777=>"000000000",
  53778=>"111000000",
  53779=>"100000000",
  53780=>"000000000",
  53781=>"111111110",
  53782=>"001111111",
  53783=>"111111111",
  53784=>"100011111",
  53785=>"011001101",
  53786=>"111000000",
  53787=>"000000000",
  53788=>"000010000",
  53789=>"111111111",
  53790=>"000000111",
  53791=>"011100110",
  53792=>"000000111",
  53793=>"110100101",
  53794=>"111111111",
  53795=>"111011011",
  53796=>"000000000",
  53797=>"000000110",
  53798=>"000000011",
  53799=>"111111111",
  53800=>"001111111",
  53801=>"000000010",
  53802=>"001000101",
  53803=>"111100000",
  53804=>"000000000",
  53805=>"111110100",
  53806=>"100000011",
  53807=>"000000000",
  53808=>"000000111",
  53809=>"001001111",
  53810=>"111111111",
  53811=>"111111001",
  53812=>"000001111",
  53813=>"111110100",
  53814=>"000000000",
  53815=>"010110110",
  53816=>"111111111",
  53817=>"011111110",
  53818=>"001001001",
  53819=>"000000000",
  53820=>"000100111",
  53821=>"000000000",
  53822=>"110101001",
  53823=>"111111101",
  53824=>"111100100",
  53825=>"011000100",
  53826=>"000000100",
  53827=>"001100100",
  53828=>"111111111",
  53829=>"000000001",
  53830=>"111111000",
  53831=>"111111111",
  53832=>"011001001",
  53833=>"000000000",
  53834=>"000000000",
  53835=>"111101101",
  53836=>"000000000",
  53837=>"000000000",
  53838=>"100011011",
  53839=>"001000111",
  53840=>"000110110",
  53841=>"100000000",
  53842=>"111111111",
  53843=>"110110010",
  53844=>"000000000",
  53845=>"010111111",
  53846=>"001101101",
  53847=>"000000000",
  53848=>"100110101",
  53849=>"000000111",
  53850=>"000110111",
  53851=>"100100111",
  53852=>"000000000",
  53853=>"100000001",
  53854=>"001001001",
  53855=>"000000100",
  53856=>"111001001",
  53857=>"000000111",
  53858=>"111111011",
  53859=>"010000010",
  53860=>"000000000",
  53861=>"001011011",
  53862=>"011000000",
  53863=>"000001111",
  53864=>"000000001",
  53865=>"110000000",
  53866=>"001000000",
  53867=>"000000000",
  53868=>"111111111",
  53869=>"111111111",
  53870=>"000000000",
  53871=>"111111111",
  53872=>"010011110",
  53873=>"111000000",
  53874=>"000000000",
  53875=>"011000100",
  53876=>"110100100",
  53877=>"111101111",
  53878=>"111111111",
  53879=>"111010000",
  53880=>"000000000",
  53881=>"001001000",
  53882=>"111111101",
  53883=>"110110110",
  53884=>"110110110",
  53885=>"111110111",
  53886=>"001001101",
  53887=>"100111111",
  53888=>"111111111",
  53889=>"001001000",
  53890=>"000000000",
  53891=>"000100010",
  53892=>"000000000",
  53893=>"000000000",
  53894=>"001111111",
  53895=>"111110100",
  53896=>"001001001",
  53897=>"000000110",
  53898=>"001111111",
  53899=>"100111000",
  53900=>"000000011",
  53901=>"000000000",
  53902=>"111110110",
  53903=>"000100000",
  53904=>"100100100",
  53905=>"000100110",
  53906=>"000000000",
  53907=>"100111111",
  53908=>"011001001",
  53909=>"000100100",
  53910=>"000100100",
  53911=>"111111111",
  53912=>"000000101",
  53913=>"111111111",
  53914=>"111110111",
  53915=>"110000000",
  53916=>"000100100",
  53917=>"100001111",
  53918=>"111111111",
  53919=>"000000000",
  53920=>"011111101",
  53921=>"000000110",
  53922=>"111111111",
  53923=>"000000000",
  53924=>"011011011",
  53925=>"001000000",
  53926=>"111111111",
  53927=>"001011111",
  53928=>"000000000",
  53929=>"111011111",
  53930=>"000000000",
  53931=>"001001111",
  53932=>"001111100",
  53933=>"011011111",
  53934=>"111111111",
  53935=>"000000000",
  53936=>"000000000",
  53937=>"000000000",
  53938=>"111111111",
  53939=>"111111111",
  53940=>"001011000",
  53941=>"110110111",
  53942=>"110000000",
  53943=>"000000010",
  53944=>"000000000",
  53945=>"001000000",
  53946=>"001001001",
  53947=>"000000111",
  53948=>"000100100",
  53949=>"000110111",
  53950=>"111111001",
  53951=>"111111111",
  53952=>"010011111",
  53953=>"100000000",
  53954=>"101100100",
  53955=>"111110000",
  53956=>"000000000",
  53957=>"110111000",
  53958=>"011111000",
  53959=>"100000000",
  53960=>"000000100",
  53961=>"101100001",
  53962=>"000000101",
  53963=>"001000001",
  53964=>"111000111",
  53965=>"000111110",
  53966=>"000000000",
  53967=>"001000101",
  53968=>"111111000",
  53969=>"000000001",
  53970=>"100101001",
  53971=>"111000001",
  53972=>"110010111",
  53973=>"001001111",
  53974=>"001001001",
  53975=>"110000000",
  53976=>"111111100",
  53977=>"000110000",
  53978=>"111000000",
  53979=>"000110111",
  53980=>"011111111",
  53981=>"100111111",
  53982=>"111111111",
  53983=>"110111111",
  53984=>"000000001",
  53985=>"111111110",
  53986=>"000000000",
  53987=>"100111111",
  53988=>"111111111",
  53989=>"000001001",
  53990=>"000000000",
  53991=>"000000000",
  53992=>"000111011",
  53993=>"000000101",
  53994=>"000111111",
  53995=>"000000000",
  53996=>"111111110",
  53997=>"110110111",
  53998=>"011000000",
  53999=>"000000000",
  54000=>"100100000",
  54001=>"111111111",
  54002=>"111011011",
  54003=>"101010111",
  54004=>"100110110",
  54005=>"001001000",
  54006=>"111111111",
  54007=>"000111111",
  54008=>"001000000",
  54009=>"000000000",
  54010=>"000000000",
  54011=>"000000000",
  54012=>"011001000",
  54013=>"000000000",
  54014=>"011111000",
  54015=>"000011111",
  54016=>"111001111",
  54017=>"110111111",
  54018=>"101111111",
  54019=>"111110111",
  54020=>"011011010",
  54021=>"000000000",
  54022=>"111101111",
  54023=>"111111111",
  54024=>"110110111",
  54025=>"001000000",
  54026=>"111111111",
  54027=>"111110000",
  54028=>"000000100",
  54029=>"110111111",
  54030=>"000100001",
  54031=>"100000000",
  54032=>"000111111",
  54033=>"100110110",
  54034=>"000000000",
  54035=>"100011011",
  54036=>"000100111",
  54037=>"000000000",
  54038=>"111111000",
  54039=>"000000110",
  54040=>"111011111",
  54041=>"000000011",
  54042=>"000000010",
  54043=>"011010000",
  54044=>"011000000",
  54045=>"110110111",
  54046=>"001111111",
  54047=>"111011111",
  54048=>"011001111",
  54049=>"000011011",
  54050=>"111111111",
  54051=>"000000000",
  54052=>"110110010",
  54053=>"100000100",
  54054=>"010111111",
  54055=>"110010000",
  54056=>"101001111",
  54057=>"000000000",
  54058=>"011111111",
  54059=>"110000000",
  54060=>"110110000",
  54061=>"000011111",
  54062=>"101101101",
  54063=>"000000111",
  54064=>"110000000",
  54065=>"100000000",
  54066=>"111001001",
  54067=>"000000000",
  54068=>"110100100",
  54069=>"111111111",
  54070=>"000001111",
  54071=>"111000100",
  54072=>"001011111",
  54073=>"001000000",
  54074=>"000001001",
  54075=>"111111111",
  54076=>"111100100",
  54077=>"000000001",
  54078=>"011001111",
  54079=>"011111110",
  54080=>"111111100",
  54081=>"111111100",
  54082=>"111111111",
  54083=>"111111111",
  54084=>"000000000",
  54085=>"000000101",
  54086=>"011111100",
  54087=>"001111111",
  54088=>"000000100",
  54089=>"111100000",
  54090=>"000000110",
  54091=>"111111100",
  54092=>"100100100",
  54093=>"000000100",
  54094=>"000100000",
  54095=>"111111011",
  54096=>"100100100",
  54097=>"000000010",
  54098=>"111100101",
  54099=>"000000000",
  54100=>"000000001",
  54101=>"011011011",
  54102=>"110100100",
  54103=>"011111010",
  54104=>"010111111",
  54105=>"000000000",
  54106=>"000000100",
  54107=>"110111000",
  54108=>"010110111",
  54109=>"111111111",
  54110=>"111011001",
  54111=>"110001111",
  54112=>"111111111",
  54113=>"111111111",
  54114=>"011011111",
  54115=>"101111111",
  54116=>"111110110",
  54117=>"000011001",
  54118=>"111110110",
  54119=>"000000000",
  54120=>"001001101",
  54121=>"111111000",
  54122=>"111111110",
  54123=>"100101001",
  54124=>"000000000",
  54125=>"111111111",
  54126=>"111111000",
  54127=>"000000001",
  54128=>"010010010",
  54129=>"000100000",
  54130=>"000111111",
  54131=>"111111111",
  54132=>"111111110",
  54133=>"001111111",
  54134=>"000100110",
  54135=>"110110110",
  54136=>"100000000",
  54137=>"000000000",
  54138=>"000000000",
  54139=>"000000000",
  54140=>"111111111",
  54141=>"101100000",
  54142=>"000001011",
  54143=>"011001000",
  54144=>"000000100",
  54145=>"001001011",
  54146=>"111011111",
  54147=>"000100110",
  54148=>"000000000",
  54149=>"100000011",
  54150=>"000100100",
  54151=>"000001111",
  54152=>"000101101",
  54153=>"000000001",
  54154=>"000000000",
  54155=>"111011000",
  54156=>"000000101",
  54157=>"010000000",
  54158=>"000111111",
  54159=>"101111111",
  54160=>"000000000",
  54161=>"111000000",
  54162=>"000000000",
  54163=>"001011011",
  54164=>"111111100",
  54165=>"000010000",
  54166=>"001111111",
  54167=>"000000011",
  54168=>"111000111",
  54169=>"111111111",
  54170=>"111111111",
  54171=>"111111111",
  54172=>"111111111",
  54173=>"101101000",
  54174=>"101001000",
  54175=>"110100000",
  54176=>"000111011",
  54177=>"111111111",
  54178=>"001001011",
  54179=>"000000111",
  54180=>"000100100",
  54181=>"111111101",
  54182=>"100100101",
  54183=>"000000000",
  54184=>"000000000",
  54185=>"101100000",
  54186=>"000010111",
  54187=>"001010000",
  54188=>"111111000",
  54189=>"011111100",
  54190=>"000000111",
  54191=>"000001000",
  54192=>"110110111",
  54193=>"110111111",
  54194=>"000000111",
  54195=>"010111111",
  54196=>"001011110",
  54197=>"111011000",
  54198=>"100100110",
  54199=>"111111100",
  54200=>"111001011",
  54201=>"100110100",
  54202=>"000001001",
  54203=>"110100110",
  54204=>"000000000",
  54205=>"000110100",
  54206=>"000000000",
  54207=>"100100100",
  54208=>"111010000",
  54209=>"111111000",
  54210=>"000000001",
  54211=>"000000000",
  54212=>"001011101",
  54213=>"000001011",
  54214=>"000000000",
  54215=>"000000000",
  54216=>"101111111",
  54217=>"000000000",
  54218=>"000000000",
  54219=>"000000111",
  54220=>"000000100",
  54221=>"011010000",
  54222=>"011000000",
  54223=>"110110110",
  54224=>"000001011",
  54225=>"000111111",
  54226=>"111111111",
  54227=>"101000000",
  54228=>"111111100",
  54229=>"001111110",
  54230=>"000000000",
  54231=>"111011011",
  54232=>"010010010",
  54233=>"000101100",
  54234=>"111111111",
  54235=>"001011011",
  54236=>"000001111",
  54237=>"100111111",
  54238=>"101101000",
  54239=>"000001011",
  54240=>"111111111",
  54241=>"000100110",
  54242=>"000001001",
  54243=>"000000100",
  54244=>"001000001",
  54245=>"000000101",
  54246=>"000000000",
  54247=>"000000000",
  54248=>"111011011",
  54249=>"000111011",
  54250=>"000000100",
  54251=>"001011111",
  54252=>"111111000",
  54253=>"100110111",
  54254=>"110111011",
  54255=>"000000001",
  54256=>"100100111",
  54257=>"001000000",
  54258=>"001000111",
  54259=>"110100000",
  54260=>"000000000",
  54261=>"010000110",
  54262=>"111111111",
  54263=>"010011001",
  54264=>"111111111",
  54265=>"111111001",
  54266=>"011101001",
  54267=>"100110111",
  54268=>"000000000",
  54269=>"111111111",
  54270=>"000000001",
  54271=>"001001001",
  54272=>"001001001",
  54273=>"100111100",
  54274=>"111111000",
  54275=>"000000000",
  54276=>"111001001",
  54277=>"011110011",
  54278=>"000000111",
  54279=>"100111111",
  54280=>"110111110",
  54281=>"100000000",
  54282=>"111000000",
  54283=>"000000000",
  54284=>"100000000",
  54285=>"101000010",
  54286=>"000101101",
  54287=>"010000000",
  54288=>"000000000",
  54289=>"000010000",
  54290=>"111000000",
  54291=>"111111111",
  54292=>"111111000",
  54293=>"000000001",
  54294=>"111111111",
  54295=>"100100100",
  54296=>"100100110",
  54297=>"110110110",
  54298=>"111111111",
  54299=>"011011011",
  54300=>"111111100",
  54301=>"011111011",
  54302=>"100000011",
  54303=>"000000111",
  54304=>"111110100",
  54305=>"011001001",
  54306=>"111111111",
  54307=>"000000111",
  54308=>"000000000",
  54309=>"000011111",
  54310=>"010000111",
  54311=>"111111111",
  54312=>"000000000",
  54313=>"010111000",
  54314=>"000000001",
  54315=>"100100000",
  54316=>"011111111",
  54317=>"000000000",
  54318=>"011011011",
  54319=>"111101111",
  54320=>"000000111",
  54321=>"010010111",
  54322=>"111011001",
  54323=>"000000000",
  54324=>"010000000",
  54325=>"100000000",
  54326=>"000000001",
  54327=>"000000000",
  54328=>"111111101",
  54329=>"000011111",
  54330=>"100000000",
  54331=>"000000000",
  54332=>"100100111",
  54333=>"111111111",
  54334=>"111000011",
  54335=>"000000000",
  54336=>"100100110",
  54337=>"010010000",
  54338=>"100110111",
  54339=>"000000111",
  54340=>"110110110",
  54341=>"111001100",
  54342=>"111111110",
  54343=>"111100000",
  54344=>"000000000",
  54345=>"110111111",
  54346=>"000000000",
  54347=>"111000000",
  54348=>"111111111",
  54349=>"000000000",
  54350=>"111110110",
  54351=>"000111111",
  54352=>"000000011",
  54353=>"111111111",
  54354=>"101000001",
  54355=>"000000000",
  54356=>"111111111",
  54357=>"011001001",
  54358=>"111011100",
  54359=>"000000000",
  54360=>"100000000",
  54361=>"111111111",
  54362=>"111111110",
  54363=>"000110010",
  54364=>"111111111",
  54365=>"111111111",
  54366=>"011001111",
  54367=>"000001000",
  54368=>"000000111",
  54369=>"010010000",
  54370=>"010101111",
  54371=>"000000110",
  54372=>"011000001",
  54373=>"111100100",
  54374=>"111111111",
  54375=>"000000000",
  54376=>"111011011",
  54377=>"000000111",
  54378=>"000111111",
  54379=>"111111000",
  54380=>"111111001",
  54381=>"111111111",
  54382=>"000000100",
  54383=>"111111111",
  54384=>"111110000",
  54385=>"001101111",
  54386=>"110111011",
  54387=>"011000000",
  54388=>"111111011",
  54389=>"111111111",
  54390=>"010000000",
  54391=>"111111111",
  54392=>"010001000",
  54393=>"110111111",
  54394=>"000000010",
  54395=>"000000000",
  54396=>"000000000",
  54397=>"000011011",
  54398=>"111111111",
  54399=>"000000000",
  54400=>"111111111",
  54401=>"000000000",
  54402=>"000000000",
  54403=>"000000000",
  54404=>"000000110",
  54405=>"101000000",
  54406=>"100100000",
  54407=>"000011001",
  54408=>"000000110",
  54409=>"111110100",
  54410=>"000000111",
  54411=>"110000000",
  54412=>"011111111",
  54413=>"111110000",
  54414=>"111111110",
  54415=>"000000000",
  54416=>"101101000",
  54417=>"000000001",
  54418=>"001100100",
  54419=>"100000000",
  54420=>"011011111",
  54421=>"000000100",
  54422=>"000000000",
  54423=>"000000000",
  54424=>"111100101",
  54425=>"000000100",
  54426=>"110110111",
  54427=>"000001011",
  54428=>"111111111",
  54429=>"111111101",
  54430=>"101001001",
  54431=>"000010000",
  54432=>"111111000",
  54433=>"001111111",
  54434=>"000000000",
  54435=>"000000000",
  54436=>"111111111",
  54437=>"110111111",
  54438=>"000000000",
  54439=>"011110110",
  54440=>"000000100",
  54441=>"111000000",
  54442=>"000000000",
  54443=>"110111111",
  54444=>"001001001",
  54445=>"000101000",
  54446=>"011001101",
  54447=>"000000100",
  54448=>"011111111",
  54449=>"111111111",
  54450=>"111111011",
  54451=>"000111000",
  54452=>"100000000",
  54453=>"111111111",
  54454=>"000000000",
  54455=>"000000000",
  54456=>"111011001",
  54457=>"111111111",
  54458=>"100110100",
  54459=>"011011001",
  54460=>"100100111",
  54461=>"111111111",
  54462=>"111000111",
  54463=>"000000000",
  54464=>"101000000",
  54465=>"111001001",
  54466=>"000000000",
  54467=>"111111111",
  54468=>"111111100",
  54469=>"111111111",
  54470=>"111011011",
  54471=>"000000000",
  54472=>"100111111",
  54473=>"000110000",
  54474=>"011000000",
  54475=>"000100111",
  54476=>"000000000",
  54477=>"000010010",
  54478=>"000000110",
  54479=>"010000000",
  54480=>"001111111",
  54481=>"001010111",
  54482=>"111000000",
  54483=>"001001011",
  54484=>"111100000",
  54485=>"000001000",
  54486=>"100000000",
  54487=>"111111111",
  54488=>"000000000",
  54489=>"000000000",
  54490=>"111111011",
  54491=>"010010000",
  54492=>"110100101",
  54493=>"000000000",
  54494=>"111111111",
  54495=>"100111011",
  54496=>"001011111",
  54497=>"000001010",
  54498=>"000111111",
  54499=>"110110110",
  54500=>"000000001",
  54501=>"110011000",
  54502=>"000000000",
  54503=>"100110100",
  54504=>"000000000",
  54505=>"001001100",
  54506=>"111111111",
  54507=>"011001011",
  54508=>"000000100",
  54509=>"001001101",
  54510=>"000000000",
  54511=>"000100111",
  54512=>"110000110",
  54513=>"100100110",
  54514=>"000000000",
  54515=>"101111001",
  54516=>"000000000",
  54517=>"000100000",
  54518=>"100100100",
  54519=>"001000000",
  54520=>"000000000",
  54521=>"000000000",
  54522=>"111001000",
  54523=>"011000110",
  54524=>"001101111",
  54525=>"111111001",
  54526=>"000001000",
  54527=>"001001000",
  54528=>"100001111",
  54529=>"110100101",
  54530=>"000000000",
  54531=>"000000000",
  54532=>"001001001",
  54533=>"111111111",
  54534=>"111111111",
  54535=>"111111101",
  54536=>"010011011",
  54537=>"111111111",
  54538=>"111111111",
  54539=>"100000011",
  54540=>"111111111",
  54541=>"111111011",
  54542=>"111111011",
  54543=>"000100000",
  54544=>"000100000",
  54545=>"000000000",
  54546=>"000000010",
  54547=>"111111111",
  54548=>"000101111",
  54549=>"111100110",
  54550=>"011011011",
  54551=>"000000000",
  54552=>"011111111",
  54553=>"100111001",
  54554=>"000111111",
  54555=>"011010010",
  54556=>"100100000",
  54557=>"101101111",
  54558=>"000000000",
  54559=>"011110000",
  54560=>"111110111",
  54561=>"000010000",
  54562=>"110100100",
  54563=>"111110000",
  54564=>"110100100",
  54565=>"111111110",
  54566=>"000000001",
  54567=>"011110110",
  54568=>"111111111",
  54569=>"000000001",
  54570=>"000111111",
  54571=>"001011011",
  54572=>"000000000",
  54573=>"100000000",
  54574=>"111111111",
  54575=>"100000101",
  54576=>"000011111",
  54577=>"000000010",
  54578=>"111111111",
  54579=>"000100000",
  54580=>"000000000",
  54581=>"001101101",
  54582=>"111000000",
  54583=>"111111101",
  54584=>"000000000",
  54585=>"111111000",
  54586=>"000000000",
  54587=>"000000111",
  54588=>"111000111",
  54589=>"111110011",
  54590=>"000000000",
  54591=>"100000001",
  54592=>"101100100",
  54593=>"100101101",
  54594=>"000000000",
  54595=>"000000000",
  54596=>"000000000",
  54597=>"111001111",
  54598=>"110110110",
  54599=>"000000000",
  54600=>"000000000",
  54601=>"000000000",
  54602=>"000000000",
  54603=>"001000000",
  54604=>"111111111",
  54605=>"000111111",
  54606=>"000000100",
  54607=>"000110100",
  54608=>"100101100",
  54609=>"000000000",
  54610=>"001011000",
  54611=>"111111111",
  54612=>"000000000",
  54613=>"001001001",
  54614=>"000000000",
  54615=>"111111000",
  54616=>"001000000",
  54617=>"000000000",
  54618=>"111111111",
  54619=>"000011111",
  54620=>"000111110",
  54621=>"000000000",
  54622=>"000000000",
  54623=>"111111111",
  54624=>"000000100",
  54625=>"111000000",
  54626=>"111100000",
  54627=>"111111111",
  54628=>"111111100",
  54629=>"000000000",
  54630=>"010010010",
  54631=>"011000001",
  54632=>"100000011",
  54633=>"111000000",
  54634=>"000000000",
  54635=>"011111111",
  54636=>"110100111",
  54637=>"000000000",
  54638=>"111111111",
  54639=>"101110111",
  54640=>"000000000",
  54641=>"000000110",
  54642=>"011000000",
  54643=>"111111111",
  54644=>"110110001",
  54645=>"100001001",
  54646=>"111001000",
  54647=>"011011001",
  54648=>"010000000",
  54649=>"001000000",
  54650=>"111111111",
  54651=>"000000111",
  54652=>"110111110",
  54653=>"000000000",
  54654=>"000000000",
  54655=>"111111111",
  54656=>"111111011",
  54657=>"110110000",
  54658=>"101101001",
  54659=>"000111111",
  54660=>"011111111",
  54661=>"000000000",
  54662=>"000110000",
  54663=>"001111111",
  54664=>"111111111",
  54665=>"111111111",
  54666=>"111011011",
  54667=>"000000000",
  54668=>"111111111",
  54669=>"111100001",
  54670=>"111111111",
  54671=>"000000000",
  54672=>"000000000",
  54673=>"001011011",
  54674=>"011110110",
  54675=>"101100101",
  54676=>"110000000",
  54677=>"000000000",
  54678=>"000010000",
  54679=>"001000000",
  54680=>"100000000",
  54681=>"111111111",
  54682=>"000000011",
  54683=>"010000000",
  54684=>"000000000",
  54685=>"111000000",
  54686=>"111011111",
  54687=>"011000000",
  54688=>"111111111",
  54689=>"001000010",
  54690=>"110010101",
  54691=>"111111111",
  54692=>"000000000",
  54693=>"000000000",
  54694=>"111111111",
  54695=>"001111111",
  54696=>"111111111",
  54697=>"000000000",
  54698=>"111111111",
  54699=>"111111111",
  54700=>"000000000",
  54701=>"000000000",
  54702=>"000001000",
  54703=>"000110111",
  54704=>"111111100",
  54705=>"111001101",
  54706=>"000000000",
  54707=>"111111000",
  54708=>"011000000",
  54709=>"000000000",
  54710=>"111111111",
  54711=>"110000000",
  54712=>"000000111",
  54713=>"000010110",
  54714=>"000000000",
  54715=>"100110111",
  54716=>"111111111",
  54717=>"111111111",
  54718=>"111111111",
  54719=>"110111111",
  54720=>"000000001",
  54721=>"000000000",
  54722=>"111111110",
  54723=>"010110110",
  54724=>"111100100",
  54725=>"000100100",
  54726=>"000000000",
  54727=>"001000000",
  54728=>"000000000",
  54729=>"000100111",
  54730=>"000001001",
  54731=>"111111111",
  54732=>"000001001",
  54733=>"000110110",
  54734=>"110010110",
  54735=>"000000000",
  54736=>"111110110",
  54737=>"111101000",
  54738=>"111001001",
  54739=>"110110111",
  54740=>"101111011",
  54741=>"011010000",
  54742=>"111111000",
  54743=>"111000000",
  54744=>"110011011",
  54745=>"000010111",
  54746=>"111111111",
  54747=>"111000000",
  54748=>"000110010",
  54749=>"000000111",
  54750=>"000000000",
  54751=>"000000000",
  54752=>"011111010",
  54753=>"101111111",
  54754=>"000111111",
  54755=>"111111000",
  54756=>"111110110",
  54757=>"001001001",
  54758=>"000000110",
  54759=>"000000000",
  54760=>"111000000",
  54761=>"110100000",
  54762=>"000000000",
  54763=>"110110111",
  54764=>"111111111",
  54765=>"011011111",
  54766=>"100100100",
  54767=>"100110110",
  54768=>"000000000",
  54769=>"111111111",
  54770=>"111111000",
  54771=>"001111111",
  54772=>"000000000",
  54773=>"110100110",
  54774=>"011001001",
  54775=>"111001001",
  54776=>"110111110",
  54777=>"000111110",
  54778=>"111111111",
  54779=>"000000100",
  54780=>"111000000",
  54781=>"111011001",
  54782=>"000000100",
  54783=>"000001011",
  54784=>"001101001",
  54785=>"001111001",
  54786=>"000111010",
  54787=>"110111110",
  54788=>"001001001",
  54789=>"000000000",
  54790=>"000000001",
  54791=>"000000000",
  54792=>"100111100",
  54793=>"111111000",
  54794=>"011000011",
  54795=>"110111111",
  54796=>"111001000",
  54797=>"111111111",
  54798=>"000001000",
  54799=>"000000000",
  54800=>"111111111",
  54801=>"111111101",
  54802=>"010111111",
  54803=>"111111011",
  54804=>"111111001",
  54805=>"000000101",
  54806=>"110000011",
  54807=>"110110110",
  54808=>"001011001",
  54809=>"101001101",
  54810=>"000000000",
  54811=>"111000000",
  54812=>"000000000",
  54813=>"100110111",
  54814=>"000000011",
  54815=>"111111111",
  54816=>"001011000",
  54817=>"001001111",
  54818=>"111011001",
  54819=>"000000011",
  54820=>"001111111",
  54821=>"100000000",
  54822=>"100000110",
  54823=>"001111000",
  54824=>"000001000",
  54825=>"000000000",
  54826=>"111111011",
  54827=>"110111010",
  54828=>"111111011",
  54829=>"111111000",
  54830=>"111111100",
  54831=>"010100111",
  54832=>"000100110",
  54833=>"000100101",
  54834=>"110110100",
  54835=>"000000011",
  54836=>"111111111",
  54837=>"111011100",
  54838=>"001110110",
  54839=>"001000000",
  54840=>"000111111",
  54841=>"001001111",
  54842=>"000000000",
  54843=>"000000000",
  54844=>"000000000",
  54845=>"000010111",
  54846=>"000000000",
  54847=>"000100111",
  54848=>"001001001",
  54849=>"110111101",
  54850=>"000000000",
  54851=>"000000000",
  54852=>"000000000",
  54853=>"000100000",
  54854=>"000000000",
  54855=>"000000100",
  54856=>"110100100",
  54857=>"000000000",
  54858=>"111111000",
  54859=>"000000010",
  54860=>"101101001",
  54861=>"111101101",
  54862=>"000111000",
  54863=>"111000111",
  54864=>"000000011",
  54865=>"111111001",
  54866=>"111111111",
  54867=>"000111111",
  54868=>"111111111",
  54869=>"101001000",
  54870=>"000111111",
  54871=>"111100111",
  54872=>"000000000",
  54873=>"111000000",
  54874=>"000000000",
  54875=>"110100111",
  54876=>"010100000",
  54877=>"100000100",
  54878=>"000011111",
  54879=>"111111001",
  54880=>"001000000",
  54881=>"000000000",
  54882=>"000111111",
  54883=>"000000000",
  54884=>"001001000",
  54885=>"000111001",
  54886=>"111111111",
  54887=>"001111111",
  54888=>"000000000",
  54889=>"000111111",
  54890=>"000000001",
  54891=>"000000101",
  54892=>"100001111",
  54893=>"111111111",
  54894=>"101111110",
  54895=>"000000000",
  54896=>"001111011",
  54897=>"011000000",
  54898=>"100100000",
  54899=>"001000100",
  54900=>"101111111",
  54901=>"000100000",
  54902=>"111000000",
  54903=>"000000000",
  54904=>"000101111",
  54905=>"001111111",
  54906=>"000010011",
  54907=>"111111111",
  54908=>"111111111",
  54909=>"111000000",
  54910=>"110111111",
  54911=>"000000000",
  54912=>"000000000",
  54913=>"000100100",
  54914=>"111111111",
  54915=>"000000111",
  54916=>"001000000",
  54917=>"001000101",
  54918=>"000000000",
  54919=>"011000001",
  54920=>"000000000",
  54921=>"000000000",
  54922=>"000000001",
  54923=>"000100111",
  54924=>"000110111",
  54925=>"000111111",
  54926=>"111111111",
  54927=>"001101101",
  54928=>"111111000",
  54929=>"111111100",
  54930=>"011111001",
  54931=>"011111111",
  54932=>"001001001",
  54933=>"100100000",
  54934=>"110111111",
  54935=>"111111001",
  54936=>"011001001",
  54937=>"000110110",
  54938=>"111000010",
  54939=>"000000000",
  54940=>"000000111",
  54941=>"001111000",
  54942=>"000101111",
  54943=>"111111111",
  54944=>"000000111",
  54945=>"000000011",
  54946=>"000000000",
  54947=>"000100000",
  54948=>"110110100",
  54949=>"000111111",
  54950=>"001011111",
  54951=>"111101111",
  54952=>"000000100",
  54953=>"000000001",
  54954=>"000000000",
  54955=>"000000000",
  54956=>"000000010",
  54957=>"100000011",
  54958=>"111101011",
  54959=>"111111011",
  54960=>"000000001",
  54961=>"111111101",
  54962=>"110100000",
  54963=>"000000000",
  54964=>"111111111",
  54965=>"111111111",
  54966=>"110001001",
  54967=>"111111101",
  54968=>"010111001",
  54969=>"111111110",
  54970=>"111110100",
  54971=>"111111011",
  54972=>"011111111",
  54973=>"100101101",
  54974=>"000110111",
  54975=>"111111000",
  54976=>"110111111",
  54977=>"011000001",
  54978=>"000000001",
  54979=>"000000111",
  54980=>"000000000",
  54981=>"111111011",
  54982=>"000111101",
  54983=>"111101001",
  54984=>"000111011",
  54985=>"000000111",
  54986=>"110110111",
  54987=>"111111111",
  54988=>"110111111",
  54989=>"000011011",
  54990=>"000110100",
  54991=>"000111111",
  54992=>"001000000",
  54993=>"111111000",
  54994=>"000101000",
  54995=>"001000000",
  54996=>"000000111",
  54997=>"111011111",
  54998=>"000000000",
  54999=>"000100011",
  55000=>"000101000",
  55001=>"000111011",
  55002=>"000000110",
  55003=>"000101111",
  55004=>"111111111",
  55005=>"010111111",
  55006=>"011111000",
  55007=>"000000111",
  55008=>"001000000",
  55009=>"011111111",
  55010=>"111111101",
  55011=>"000000000",
  55012=>"100000100",
  55013=>"110110100",
  55014=>"000000110",
  55015=>"111111101",
  55016=>"000001000",
  55017=>"000101111",
  55018=>"000000000",
  55019=>"011111111",
  55020=>"111000000",
  55021=>"010000000",
  55022=>"000110111",
  55023=>"000011000",
  55024=>"000100111",
  55025=>"010000000",
  55026=>"000000111",
  55027=>"001001010",
  55028=>"111111111",
  55029=>"111110100",
  55030=>"110110100",
  55031=>"100000000",
  55032=>"000000000",
  55033=>"000000101",
  55034=>"001011111",
  55035=>"111111000",
  55036=>"111110111",
  55037=>"001001011",
  55038=>"000000100",
  55039=>"100100000",
  55040=>"111001001",
  55041=>"111011011",
  55042=>"111101000",
  55043=>"000011011",
  55044=>"000000000",
  55045=>"011010000",
  55046=>"000100110",
  55047=>"111110000",
  55048=>"000000011",
  55049=>"001011010",
  55050=>"110000011",
  55051=>"011111111",
  55052=>"100000111",
  55053=>"000000110",
  55054=>"110000000",
  55055=>"100000000",
  55056=>"001110110",
  55057=>"001001001",
  55058=>"100110100",
  55059=>"000000100",
  55060=>"111111111",
  55061=>"111111011",
  55062=>"111111100",
  55063=>"111110110",
  55064=>"111111111",
  55065=>"000000000",
  55066=>"111111111",
  55067=>"001000000",
  55068=>"000001111",
  55069=>"001001000",
  55070=>"000001011",
  55071=>"000000001",
  55072=>"100111101",
  55073=>"001000101",
  55074=>"000111111",
  55075=>"111111111",
  55076=>"001111111",
  55077=>"000011011",
  55078=>"111111000",
  55079=>"111110011",
  55080=>"011111010",
  55081=>"111111111",
  55082=>"101101101",
  55083=>"000111111",
  55084=>"101101111",
  55085=>"000001001",
  55086=>"000111000",
  55087=>"000010000",
  55088=>"000011111",
  55089=>"111100111",
  55090=>"000111111",
  55091=>"111111111",
  55092=>"000000000",
  55093=>"000100000",
  55094=>"000000000",
  55095=>"110000000",
  55096=>"000111001",
  55097=>"000000000",
  55098=>"000100110",
  55099=>"000000000",
  55100=>"111101111",
  55101=>"000000001",
  55102=>"000000000",
  55103=>"001110111",
  55104=>"000000011",
  55105=>"111111110",
  55106=>"100100001",
  55107=>"000000000",
  55108=>"111111111",
  55109=>"000000000",
  55110=>"000100101",
  55111=>"111111111",
  55112=>"000000010",
  55113=>"001000000",
  55114=>"001001011",
  55115=>"111011011",
  55116=>"110110000",
  55117=>"000011011",
  55118=>"000000001",
  55119=>"001000010",
  55120=>"000000001",
  55121=>"111101111",
  55122=>"000000000",
  55123=>"000000111",
  55124=>"111000000",
  55125=>"101101101",
  55126=>"000000010",
  55127=>"000100111",
  55128=>"000100110",
  55129=>"111100000",
  55130=>"001111110",
  55131=>"000001000",
  55132=>"010111010",
  55133=>"000000000",
  55134=>"000011000",
  55135=>"001001000",
  55136=>"111111011",
  55137=>"000000111",
  55138=>"100110000",
  55139=>"000000000",
  55140=>"110000000",
  55141=>"000011011",
  55142=>"000001101",
  55143=>"000100100",
  55144=>"111011001",
  55145=>"000100011",
  55146=>"000111011",
  55147=>"100000000",
  55148=>"011110111",
  55149=>"111111111",
  55150=>"101111000",
  55151=>"000001010",
  55152=>"000000000",
  55153=>"000000110",
  55154=>"111110010",
  55155=>"001111111",
  55156=>"101111111",
  55157=>"111111111",
  55158=>"000011001",
  55159=>"111000000",
  55160=>"011000001",
  55161=>"001111001",
  55162=>"111101001",
  55163=>"010110111",
  55164=>"111111101",
  55165=>"111110111",
  55166=>"000111111",
  55167=>"000111111",
  55168=>"100000101",
  55169=>"000000110",
  55170=>"000000111",
  55171=>"111111111",
  55172=>"000111111",
  55173=>"100000100",
  55174=>"001000111",
  55175=>"001001010",
  55176=>"000000000",
  55177=>"101001000",
  55178=>"001010000",
  55179=>"111001000",
  55180=>"111111111",
  55181=>"010000000",
  55182=>"010011111",
  55183=>"011101111",
  55184=>"111111111",
  55185=>"111001101",
  55186=>"111111110",
  55187=>"111111110",
  55188=>"101000000",
  55189=>"000000100",
  55190=>"000000111",
  55191=>"100101100",
  55192=>"110111001",
  55193=>"011100110",
  55194=>"111111111",
  55195=>"100111110",
  55196=>"111100110",
  55197=>"000001000",
  55198=>"110000110",
  55199=>"110100000",
  55200=>"110000100",
  55201=>"011110000",
  55202=>"000000100",
  55203=>"110011000",
  55204=>"110100100",
  55205=>"000000000",
  55206=>"000111000",
  55207=>"000000000",
  55208=>"000000000",
  55209=>"010000000",
  55210=>"111011000",
  55211=>"111000000",
  55212=>"111000100",
  55213=>"001101011",
  55214=>"000000111",
  55215=>"000000000",
  55216=>"000000000",
  55217=>"111111111",
  55218=>"111001000",
  55219=>"111000111",
  55220=>"100100000",
  55221=>"111110000",
  55222=>"000000000",
  55223=>"111111010",
  55224=>"000000000",
  55225=>"111111111",
  55226=>"111111000",
  55227=>"111110100",
  55228=>"111111111",
  55229=>"111000000",
  55230=>"000000000",
  55231=>"111001001",
  55232=>"000000000",
  55233=>"111111111",
  55234=>"000000000",
  55235=>"000100100",
  55236=>"000101000",
  55237=>"000000100",
  55238=>"000100111",
  55239=>"011111111",
  55240=>"111000000",
  55241=>"111111111",
  55242=>"000000101",
  55243=>"110111000",
  55244=>"111111111",
  55245=>"000000000",
  55246=>"001001001",
  55247=>"111111111",
  55248=>"000000000",
  55249=>"000000000",
  55250=>"111111111",
  55251=>"000000111",
  55252=>"001001001",
  55253=>"000111111",
  55254=>"000000000",
  55255=>"011000011",
  55256=>"000000000",
  55257=>"100000110",
  55258=>"111111000",
  55259=>"100111111",
  55260=>"000101000",
  55261=>"000000000",
  55262=>"110110000",
  55263=>"010100110",
  55264=>"111111111",
  55265=>"001001010",
  55266=>"111111010",
  55267=>"010000000",
  55268=>"111111111",
  55269=>"111111111",
  55270=>"011101100",
  55271=>"011001001",
  55272=>"111111111",
  55273=>"111111100",
  55274=>"111110000",
  55275=>"000010010",
  55276=>"000000000",
  55277=>"110010011",
  55278=>"000000000",
  55279=>"111111111",
  55280=>"110111111",
  55281=>"000001001",
  55282=>"000000000",
  55283=>"000111000",
  55284=>"110000110",
  55285=>"111100000",
  55286=>"001011011",
  55287=>"100111111",
  55288=>"000000001",
  55289=>"000000001",
  55290=>"000000000",
  55291=>"111111111",
  55292=>"111111011",
  55293=>"000000000",
  55294=>"111111111",
  55295=>"000000000",
  55296=>"111111111",
  55297=>"000110000",
  55298=>"000000000",
  55299=>"000000000",
  55300=>"111111111",
  55301=>"100010000",
  55302=>"100100111",
  55303=>"000000111",
  55304=>"111111111",
  55305=>"000000000",
  55306=>"101001111",
  55307=>"000000000",
  55308=>"111111111",
  55309=>"111111001",
  55310=>"000000000",
  55311=>"000110000",
  55312=>"100111111",
  55313=>"111000110",
  55314=>"111111111",
  55315=>"000110111",
  55316=>"111111111",
  55317=>"111000000",
  55318=>"000000111",
  55319=>"011111110",
  55320=>"111111100",
  55321=>"111111100",
  55322=>"000000011",
  55323=>"110000001",
  55324=>"000000000",
  55325=>"011011001",
  55326=>"111011111",
  55327=>"111101111",
  55328=>"101000000",
  55329=>"000000000",
  55330=>"111111101",
  55331=>"100000000",
  55332=>"001111111",
  55333=>"000011111",
  55334=>"111111101",
  55335=>"011110100",
  55336=>"011000011",
  55337=>"000000011",
  55338=>"010000011",
  55339=>"000000001",
  55340=>"000000110",
  55341=>"011000100",
  55342=>"000110111",
  55343=>"111111111",
  55344=>"111100100",
  55345=>"000000000",
  55346=>"011000000",
  55347=>"000111000",
  55348=>"011111111",
  55349=>"101100110",
  55350=>"000000000",
  55351=>"000000000",
  55352=>"000000000",
  55353=>"011011111",
  55354=>"000000011",
  55355=>"111111111",
  55356=>"000000111",
  55357=>"110000000",
  55358=>"111111111",
  55359=>"000000100",
  55360=>"011011111",
  55361=>"000000000",
  55362=>"111111111",
  55363=>"010000110",
  55364=>"000000000",
  55365=>"000000111",
  55366=>"011000010",
  55367=>"111111111",
  55368=>"111111111",
  55369=>"000000000",
  55370=>"110111111",
  55371=>"000000100",
  55372=>"000000000",
  55373=>"011000110",
  55374=>"110110000",
  55375=>"111000100",
  55376=>"000000000",
  55377=>"100101111",
  55378=>"000000000",
  55379=>"100000000",
  55380=>"000000011",
  55381=>"001011111",
  55382=>"000111111",
  55383=>"000000000",
  55384=>"011000000",
  55385=>"000000000",
  55386=>"111111111",
  55387=>"110110111",
  55388=>"111111111",
  55389=>"111111100",
  55390=>"000000000",
  55391=>"001111000",
  55392=>"000000000",
  55393=>"000010010",
  55394=>"000111111",
  55395=>"100110110",
  55396=>"000101000",
  55397=>"111111111",
  55398=>"000000111",
  55399=>"001000111",
  55400=>"000111111",
  55401=>"001111111",
  55402=>"000010000",
  55403=>"000111111",
  55404=>"100000000",
  55405=>"000000000",
  55406=>"000001111",
  55407=>"000000000",
  55408=>"000001111",
  55409=>"000000111",
  55410=>"111111001",
  55411=>"001011011",
  55412=>"000000000",
  55413=>"001000001",
  55414=>"001000000",
  55415=>"111111111",
  55416=>"001000000",
  55417=>"001001111",
  55418=>"000001001",
  55419=>"000000001",
  55420=>"111100110",
  55421=>"000000000",
  55422=>"001111000",
  55423=>"000000111",
  55424=>"000000000",
  55425=>"111111111",
  55426=>"000000000",
  55427=>"000110111",
  55428=>"000000000",
  55429=>"001101111",
  55430=>"110100000",
  55431=>"111011011",
  55432=>"000110111",
  55433=>"111100000",
  55434=>"111111000",
  55435=>"000000000",
  55436=>"000010000",
  55437=>"000000000",
  55438=>"110111110",
  55439=>"100100000",
  55440=>"011011111",
  55441=>"110110000",
  55442=>"000000100",
  55443=>"000100000",
  55444=>"011010111",
  55445=>"000000100",
  55446=>"000000000",
  55447=>"000000000",
  55448=>"111111100",
  55449=>"111111000",
  55450=>"111011011",
  55451=>"010010000",
  55452=>"000000000",
  55453=>"000000011",
  55454=>"101001000",
  55455=>"111111001",
  55456=>"000010000",
  55457=>"110110011",
  55458=>"010111100",
  55459=>"111011000",
  55460=>"001001110",
  55461=>"100110000",
  55462=>"000111000",
  55463=>"011101111",
  55464=>"000000000",
  55465=>"111110010",
  55466=>"000000001",
  55467=>"010110111",
  55468=>"000111111",
  55469=>"001000001",
  55470=>"111111000",
  55471=>"000111000",
  55472=>"000111111",
  55473=>"111111111",
  55474=>"111111110",
  55475=>"000000000",
  55476=>"001001000",
  55477=>"000011000",
  55478=>"111111111",
  55479=>"000000000",
  55480=>"111111000",
  55481=>"101111111",
  55482=>"111000000",
  55483=>"000000110",
  55484=>"111111111",
  55485=>"001000101",
  55486=>"100111111",
  55487=>"111111001",
  55488=>"111111111",
  55489=>"000111000",
  55490=>"011111001",
  55491=>"000000000",
  55492=>"111111111",
  55493=>"000000000",
  55494=>"011001011",
  55495=>"110011001",
  55496=>"001111111",
  55497=>"100011111",
  55498=>"000000000",
  55499=>"111111111",
  55500=>"110110101",
  55501=>"000000111",
  55502=>"000001001",
  55503=>"000000111",
  55504=>"100110011",
  55505=>"111111000",
  55506=>"000000000",
  55507=>"111111000",
  55508=>"110111000",
  55509=>"111111100",
  55510=>"000001111",
  55511=>"000000000",
  55512=>"000000000",
  55513=>"011111101",
  55514=>"000000010",
  55515=>"000000000",
  55516=>"000000001",
  55517=>"000000000",
  55518=>"000111000",
  55519=>"000000000",
  55520=>"000000000",
  55521=>"001001001",
  55522=>"111011000",
  55523=>"000111111",
  55524=>"000001001",
  55525=>"000000111",
  55526=>"001000000",
  55527=>"000000000",
  55528=>"000000000",
  55529=>"000000111",
  55530=>"111111100",
  55531=>"000000000",
  55532=>"000110111",
  55533=>"001000000",
  55534=>"001011111",
  55535=>"111000001",
  55536=>"000000000",
  55537=>"110111111",
  55538=>"000000010",
  55539=>"111110010",
  55540=>"010000100",
  55541=>"000111101",
  55542=>"000100000",
  55543=>"111001000",
  55544=>"000000000",
  55545=>"001001011",
  55546=>"110111111",
  55547=>"111111111",
  55548=>"001001111",
  55549=>"000110110",
  55550=>"000011111",
  55551=>"001001000",
  55552=>"111111111",
  55553=>"100100111",
  55554=>"000000000",
  55555=>"000000110",
  55556=>"011001000",
  55557=>"000000000",
  55558=>"000000000",
  55559=>"000001000",
  55560=>"000000000",
  55561=>"000000000",
  55562=>"000000000",
  55563=>"000000000",
  55564=>"100000001",
  55565=>"100000000",
  55566=>"010000001",
  55567=>"000000000",
  55568=>"000000000",
  55569=>"000000000",
  55570=>"000000010",
  55571=>"101000000",
  55572=>"000000000",
  55573=>"000000010",
  55574=>"011011011",
  55575=>"111111111",
  55576=>"010011011",
  55577=>"111110000",
  55578=>"000000000",
  55579=>"111110010",
  55580=>"100100111",
  55581=>"000000000",
  55582=>"000000001",
  55583=>"000000110",
  55584=>"110111011",
  55585=>"100111011",
  55586=>"010111111",
  55587=>"010010010",
  55588=>"000000000",
  55589=>"111111001",
  55590=>"110110100",
  55591=>"000000000",
  55592=>"000000000",
  55593=>"000000000",
  55594=>"000110000",
  55595=>"000000000",
  55596=>"110111111",
  55597=>"111010010",
  55598=>"000000000",
  55599=>"000000000",
  55600=>"000011111",
  55601=>"110111001",
  55602=>"111001111",
  55603=>"000000000",
  55604=>"000000000",
  55605=>"111110111",
  55606=>"111001001",
  55607=>"000001001",
  55608=>"000000000",
  55609=>"111111110",
  55610=>"000000111",
  55611=>"111000100",
  55612=>"110101100",
  55613=>"000000000",
  55614=>"000000000",
  55615=>"001000000",
  55616=>"000111111",
  55617=>"000111000",
  55618=>"111111111",
  55619=>"100001001",
  55620=>"110000100",
  55621=>"000000000",
  55622=>"000000111",
  55623=>"000000111",
  55624=>"000000000",
  55625=>"000000000",
  55626=>"000110000",
  55627=>"111101110",
  55628=>"000000001",
  55629=>"000110000",
  55630=>"110000000",
  55631=>"000000000",
  55632=>"001001111",
  55633=>"000000100",
  55634=>"000000011",
  55635=>"111111111",
  55636=>"111011000",
  55637=>"001001001",
  55638=>"001111111",
  55639=>"000011111",
  55640=>"000000101",
  55641=>"111110110",
  55642=>"011011110",
  55643=>"110110000",
  55644=>"000011111",
  55645=>"111111111",
  55646=>"000000000",
  55647=>"000100100",
  55648=>"000000000",
  55649=>"010000100",
  55650=>"110111111",
  55651=>"000111111",
  55652=>"000001001",
  55653=>"000010111",
  55654=>"111000000",
  55655=>"111111111",
  55656=>"111111111",
  55657=>"101101000",
  55658=>"100000000",
  55659=>"000100111",
  55660=>"000000000",
  55661=>"101001111",
  55662=>"000000000",
  55663=>"000010011",
  55664=>"000000000",
  55665=>"000000000",
  55666=>"111111111",
  55667=>"110110110",
  55668=>"000000000",
  55669=>"100000000",
  55670=>"000110110",
  55671=>"111111111",
  55672=>"000000000",
  55673=>"001000010",
  55674=>"111000000",
  55675=>"111111010",
  55676=>"100111111",
  55677=>"101000000",
  55678=>"001011111",
  55679=>"000010111",
  55680=>"111111011",
  55681=>"000000000",
  55682=>"001011000",
  55683=>"000000000",
  55684=>"001111111",
  55685=>"001001001",
  55686=>"000011001",
  55687=>"000110010",
  55688=>"011000000",
  55689=>"111111111",
  55690=>"111111111",
  55691=>"000111111",
  55692=>"111111111",
  55693=>"001011001",
  55694=>"000100000",
  55695=>"001111111",
  55696=>"000000000",
  55697=>"001000000",
  55698=>"001010010",
  55699=>"010111111",
  55700=>"111001000",
  55701=>"001011000",
  55702=>"100110111",
  55703=>"111101111",
  55704=>"010110011",
  55705=>"000011011",
  55706=>"111111111",
  55707=>"000000001",
  55708=>"011111111",
  55709=>"111011111",
  55710=>"111001000",
  55711=>"000000011",
  55712=>"111111111",
  55713=>"000000000",
  55714=>"000011111",
  55715=>"000000010",
  55716=>"100001000",
  55717=>"000011111",
  55718=>"001011111",
  55719=>"111111111",
  55720=>"000111111",
  55721=>"000010000",
  55722=>"001101101",
  55723=>"111110000",
  55724=>"101000000",
  55725=>"111111000",
  55726=>"000000111",
  55727=>"111111000",
  55728=>"011001011",
  55729=>"000001111",
  55730=>"111111001",
  55731=>"000000000",
  55732=>"000000000",
  55733=>"000000000",
  55734=>"000000101",
  55735=>"000111111",
  55736=>"000111111",
  55737=>"111111111",
  55738=>"000000000",
  55739=>"000111111",
  55740=>"000111111",
  55741=>"111111110",
  55742=>"111110100",
  55743=>"000000101",
  55744=>"000111111",
  55745=>"000000010",
  55746=>"111111010",
  55747=>"000000000",
  55748=>"000000101",
  55749=>"000110110",
  55750=>"010000111",
  55751=>"001100100",
  55752=>"111011101",
  55753=>"000000010",
  55754=>"000000000",
  55755=>"100111111",
  55756=>"000000000",
  55757=>"110000100",
  55758=>"100010001",
  55759=>"011111111",
  55760=>"000010000",
  55761=>"000110111",
  55762=>"000011011",
  55763=>"011111111",
  55764=>"000000000",
  55765=>"000000101",
  55766=>"010010111",
  55767=>"111011111",
  55768=>"001001000",
  55769=>"111000101",
  55770=>"000011010",
  55771=>"000010111",
  55772=>"000001111",
  55773=>"000000000",
  55774=>"100000100",
  55775=>"101001101",
  55776=>"000100111",
  55777=>"100000010",
  55778=>"101111100",
  55779=>"000001001",
  55780=>"110110101",
  55781=>"000000111",
  55782=>"111111001",
  55783=>"000000000",
  55784=>"011111111",
  55785=>"111111111",
  55786=>"101100001",
  55787=>"000000000",
  55788=>"111111000",
  55789=>"111100100",
  55790=>"011000000",
  55791=>"110000000",
  55792=>"100000000",
  55793=>"010111111",
  55794=>"000000000",
  55795=>"111110010",
  55796=>"000000000",
  55797=>"000000000",
  55798=>"111111100",
  55799=>"000100110",
  55800=>"101100100",
  55801=>"000000000",
  55802=>"111100110",
  55803=>"001111001",
  55804=>"111111110",
  55805=>"001000000",
  55806=>"000110111",
  55807=>"011011000",
  55808=>"000000100",
  55809=>"000000000",
  55810=>"000000111",
  55811=>"000110000",
  55812=>"000000000",
  55813=>"100000000",
  55814=>"111000000",
  55815=>"110111111",
  55816=>"000010111",
  55817=>"111111111",
  55818=>"000000000",
  55819=>"111111111",
  55820=>"100000000",
  55821=>"000000000",
  55822=>"000100111",
  55823=>"111111011",
  55824=>"111111111",
  55825=>"000000011",
  55826=>"111000011",
  55827=>"000000111",
  55828=>"111111111",
  55829=>"111111111",
  55830=>"010000100",
  55831=>"000000000",
  55832=>"100101100",
  55833=>"100100100",
  55834=>"000000111",
  55835=>"111111010",
  55836=>"111111111",
  55837=>"111111111",
  55838=>"100100100",
  55839=>"000000000",
  55840=>"111111111",
  55841=>"111111111",
  55842=>"000000000",
  55843=>"111000001",
  55844=>"111111111",
  55845=>"110111111",
  55846=>"000000111",
  55847=>"111000000",
  55848=>"000000001",
  55849=>"111111111",
  55850=>"000000111",
  55851=>"110000000",
  55852=>"010000000",
  55853=>"111111001",
  55854=>"001001001",
  55855=>"000100000",
  55856=>"100100000",
  55857=>"111111111",
  55858=>"111111001",
  55859=>"000000000",
  55860=>"000000111",
  55861=>"111101111",
  55862=>"011010000",
  55863=>"111111111",
  55864=>"000001111",
  55865=>"000100110",
  55866=>"111100110",
  55867=>"111111111",
  55868=>"000000000",
  55869=>"000000000",
  55870=>"111000000",
  55871=>"100100111",
  55872=>"000000000",
  55873=>"111111111",
  55874=>"111011011",
  55875=>"000100100",
  55876=>"110011001",
  55877=>"011011000",
  55878=>"000010011",
  55879=>"110110111",
  55880=>"100101001",
  55881=>"111000101",
  55882=>"000000111",
  55883=>"000000011",
  55884=>"011111111",
  55885=>"011000000",
  55886=>"100000000",
  55887=>"111111111",
  55888=>"000000100",
  55889=>"111111111",
  55890=>"111110011",
  55891=>"000101110",
  55892=>"111101111",
  55893=>"101000000",
  55894=>"100100101",
  55895=>"000000000",
  55896=>"000000111",
  55897=>"101000101",
  55898=>"001000111",
  55899=>"001001001",
  55900=>"000001111",
  55901=>"110110111",
  55902=>"000000000",
  55903=>"111111111",
  55904=>"000000000",
  55905=>"000001101",
  55906=>"000000000",
  55907=>"000000000",
  55908=>"000111110",
  55909=>"111000111",
  55910=>"111111111",
  55911=>"111010100",
  55912=>"101000000",
  55913=>"100100111",
  55914=>"000000110",
  55915=>"000110101",
  55916=>"001101000",
  55917=>"000000000",
  55918=>"111111000",
  55919=>"000000000",
  55920=>"100000000",
  55921=>"000000100",
  55922=>"000000111",
  55923=>"000000000",
  55924=>"000000101",
  55925=>"111110000",
  55926=>"000110111",
  55927=>"011111111",
  55928=>"110110000",
  55929=>"000110111",
  55930=>"111001001",
  55931=>"000000000",
  55932=>"110111111",
  55933=>"000100111",
  55934=>"000000000",
  55935=>"111110111",
  55936=>"111111111",
  55937=>"000000101",
  55938=>"000000000",
  55939=>"000001000",
  55940=>"000000111",
  55941=>"000000111",
  55942=>"111111001",
  55943=>"111111111",
  55944=>"000000000",
  55945=>"000111011",
  55946=>"000111111",
  55947=>"000000000",
  55948=>"111111111",
  55949=>"111111111",
  55950=>"000000000",
  55951=>"100000000",
  55952=>"001011111",
  55953=>"000011111",
  55954=>"111110110",
  55955=>"000000011",
  55956=>"000001000",
  55957=>"110110111",
  55958=>"000010110",
  55959=>"000101111",
  55960=>"000000001",
  55961=>"111111100",
  55962=>"110111111",
  55963=>"111111111",
  55964=>"111111111",
  55965=>"111111110",
  55966=>"110100000",
  55967=>"000000000",
  55968=>"110110111",
  55969=>"100000000",
  55970=>"111111010",
  55971=>"000000110",
  55972=>"111011111",
  55973=>"111011011",
  55974=>"000101111",
  55975=>"111111111",
  55976=>"111111110",
  55977=>"000001001",
  55978=>"000000000",
  55979=>"100100111",
  55980=>"111111110",
  55981=>"110111111",
  55982=>"111111111",
  55983=>"111111011",
  55984=>"000010000",
  55985=>"111111100",
  55986=>"111111111",
  55987=>"111101101",
  55988=>"111110110",
  55989=>"111011111",
  55990=>"111111001",
  55991=>"000011000",
  55992=>"000000000",
  55993=>"000000000",
  55994=>"011111011",
  55995=>"111111101",
  55996=>"100000000",
  55997=>"111000000",
  55998=>"000000000",
  55999=>"011011111",
  56000=>"000000000",
  56001=>"000000000",
  56002=>"000000111",
  56003=>"000000001",
  56004=>"110100110",
  56005=>"000000111",
  56006=>"010011000",
  56007=>"111011111",
  56008=>"111111111",
  56009=>"000000111",
  56010=>"100100011",
  56011=>"000000101",
  56012=>"111111111",
  56013=>"111111111",
  56014=>"111111111",
  56015=>"000100100",
  56016=>"000110110",
  56017=>"100100000",
  56018=>"000111000",
  56019=>"010110111",
  56020=>"111000100",
  56021=>"000000001",
  56022=>"000001111",
  56023=>"111000000",
  56024=>"110110100",
  56025=>"110110010",
  56026=>"111000000",
  56027=>"111110110",
  56028=>"111010111",
  56029=>"000001011",
  56030=>"100000000",
  56031=>"000100111",
  56032=>"000000101",
  56033=>"000000110",
  56034=>"000010010",
  56035=>"101010000",
  56036=>"011100000",
  56037=>"100110110",
  56038=>"001101101",
  56039=>"000000111",
  56040=>"000100000",
  56041=>"000000101",
  56042=>"000100111",
  56043=>"100100101",
  56044=>"010011001",
  56045=>"000000011",
  56046=>"000000000",
  56047=>"000111111",
  56048=>"111001000",
  56049=>"111000000",
  56050=>"000000000",
  56051=>"111110111",
  56052=>"111111010",
  56053=>"111111010",
  56054=>"011001111",
  56055=>"111111111",
  56056=>"000000000",
  56057=>"011000001",
  56058=>"100110111",
  56059=>"111111100",
  56060=>"111110000",
  56061=>"000100100",
  56062=>"011111111",
  56063=>"000010111",
  56064=>"111000110",
  56065=>"000000000",
  56066=>"111000000",
  56067=>"000000000",
  56068=>"000001111",
  56069=>"110000000",
  56070=>"111111111",
  56071=>"000000100",
  56072=>"000100111",
  56073=>"000000111",
  56074=>"000011000",
  56075=>"000100111",
  56076=>"111001111",
  56077=>"101100111",
  56078=>"000101101",
  56079=>"111111111",
  56080=>"111110110",
  56081=>"000000110",
  56082=>"000000111",
  56083=>"000000000",
  56084=>"000000000",
  56085=>"001001000",
  56086=>"100001001",
  56087=>"100000001",
  56088=>"000101111",
  56089=>"111111110",
  56090=>"100110111",
  56091=>"000111111",
  56092=>"111111111",
  56093=>"000000110",
  56094=>"000000000",
  56095=>"100000000",
  56096=>"000000011",
  56097=>"000000000",
  56098=>"000000110",
  56099=>"100111111",
  56100=>"111111111",
  56101=>"000000000",
  56102=>"000000000",
  56103=>"000000110",
  56104=>"000100110",
  56105=>"111111111",
  56106=>"111111111",
  56107=>"111101101",
  56108=>"100100001",
  56109=>"000000001",
  56110=>"111111111",
  56111=>"100100110",
  56112=>"000001101",
  56113=>"111111111",
  56114=>"000000000",
  56115=>"000110000",
  56116=>"111000000",
  56117=>"000011011",
  56118=>"000100111",
  56119=>"000000111",
  56120=>"000000000",
  56121=>"000000000",
  56122=>"100100101",
  56123=>"111000000",
  56124=>"000000000",
  56125=>"100000110",
  56126=>"000110110",
  56127=>"000000000",
  56128=>"111001101",
  56129=>"111111110",
  56130=>"100110010",
  56131=>"000000100",
  56132=>"100001110",
  56133=>"000000111",
  56134=>"000000000",
  56135=>"111111111",
  56136=>"000000000",
  56137=>"000000000",
  56138=>"100010000",
  56139=>"000100100",
  56140=>"111110100",
  56141=>"111110000",
  56142=>"100111111",
  56143=>"000000001",
  56144=>"001000100",
  56145=>"111111110",
  56146=>"101000000",
  56147=>"000000000",
  56148=>"111100000",
  56149=>"001011000",
  56150=>"100100000",
  56151=>"110111111",
  56152=>"000001000",
  56153=>"000000111",
  56154=>"111111111",
  56155=>"000111111",
  56156=>"100000010",
  56157=>"000000000",
  56158=>"000000111",
  56159=>"111111111",
  56160=>"000000000",
  56161=>"001000000",
  56162=>"110010111",
  56163=>"000000111",
  56164=>"110100000",
  56165=>"000000000",
  56166=>"000000000",
  56167=>"100111111",
  56168=>"111001001",
  56169=>"111111000",
  56170=>"011001000",
  56171=>"101111010",
  56172=>"000000000",
  56173=>"011011111",
  56174=>"100111000",
  56175=>"000000000",
  56176=>"000000000",
  56177=>"000000000",
  56178=>"100000111",
  56179=>"111111111",
  56180=>"111111011",
  56181=>"110111001",
  56182=>"000000111",
  56183=>"000000001",
  56184=>"110100000",
  56185=>"000000000",
  56186=>"100100111",
  56187=>"000000000",
  56188=>"011011010",
  56189=>"000000001",
  56190=>"111000000",
  56191=>"000000000",
  56192=>"110110110",
  56193=>"000001111",
  56194=>"111111111",
  56195=>"000000000",
  56196=>"000111111",
  56197=>"000000011",
  56198=>"001101111",
  56199=>"110111111",
  56200=>"001001001",
  56201=>"000000000",
  56202=>"100000001",
  56203=>"000011000",
  56204=>"111101111",
  56205=>"111110100",
  56206=>"000000100",
  56207=>"011111001",
  56208=>"000000000",
  56209=>"111111000",
  56210=>"000000000",
  56211=>"000000000",
  56212=>"111111011",
  56213=>"000110011",
  56214=>"111110110",
  56215=>"100100100",
  56216=>"111000000",
  56217=>"111111111",
  56218=>"100100000",
  56219=>"000000000",
  56220=>"000000000",
  56221=>"011000000",
  56222=>"000000000",
  56223=>"111111111",
  56224=>"011000000",
  56225=>"000000100",
  56226=>"111000000",
  56227=>"111111111",
  56228=>"010111110",
  56229=>"000000000",
  56230=>"111111111",
  56231=>"110111111",
  56232=>"111011000",
  56233=>"100100101",
  56234=>"000010000",
  56235=>"111010011",
  56236=>"000000000",
  56237=>"100000000",
  56238=>"001100110",
  56239=>"111111111",
  56240=>"111111100",
  56241=>"000000000",
  56242=>"100111111",
  56243=>"000000101",
  56244=>"011001001",
  56245=>"000000000",
  56246=>"100111111",
  56247=>"100000001",
  56248=>"000000010",
  56249=>"100000100",
  56250=>"011011000",
  56251=>"111000100",
  56252=>"101111111",
  56253=>"111111110",
  56254=>"111111101",
  56255=>"100100100",
  56256=>"111111111",
  56257=>"110111111",
  56258=>"110001000",
  56259=>"010111111",
  56260=>"000000000",
  56261=>"000010000",
  56262=>"000000000",
  56263=>"100100101",
  56264=>"010000011",
  56265=>"000000000",
  56266=>"000000111",
  56267=>"010111001",
  56268=>"000000000",
  56269=>"000000000",
  56270=>"000000000",
  56271=>"111111111",
  56272=>"000110000",
  56273=>"111111111",
  56274=>"110111111",
  56275=>"000000100",
  56276=>"111101111",
  56277=>"010111010",
  56278=>"000000000",
  56279=>"000000000",
  56280=>"111111110",
  56281=>"000100110",
  56282=>"000000000",
  56283=>"111100000",
  56284=>"000000100",
  56285=>"111111111",
  56286=>"000010001",
  56287=>"000000111",
  56288=>"001000000",
  56289=>"000000000",
  56290=>"011111111",
  56291=>"110000000",
  56292=>"110000100",
  56293=>"010010010",
  56294=>"000000010",
  56295=>"000010000",
  56296=>"000000111",
  56297=>"001000000",
  56298=>"110110111",
  56299=>"000000000",
  56300=>"111111000",
  56301=>"011001001",
  56302=>"101100000",
  56303=>"011011111",
  56304=>"001001111",
  56305=>"111111111",
  56306=>"111111111",
  56307=>"000000000",
  56308=>"100001110",
  56309=>"000000000",
  56310=>"111001101",
  56311=>"100100000",
  56312=>"000000111",
  56313=>"001000001",
  56314=>"000000110",
  56315=>"101001001",
  56316=>"000001001",
  56317=>"111000000",
  56318=>"111111010",
  56319=>"000011111",
  56320=>"010111111",
  56321=>"111111111",
  56322=>"011001011",
  56323=>"000001001",
  56324=>"000000000",
  56325=>"000000111",
  56326=>"011001001",
  56327=>"111011001",
  56328=>"110100100",
  56329=>"110000010",
  56330=>"000000000",
  56331=>"000000000",
  56332=>"010010001",
  56333=>"111111111",
  56334=>"001100000",
  56335=>"111111111",
  56336=>"010101001",
  56337=>"111111011",
  56338=>"000000111",
  56339=>"000000000",
  56340=>"000000000",
  56341=>"111011111",
  56342=>"111011111",
  56343=>"011011001",
  56344=>"111110100",
  56345=>"011001010",
  56346=>"100111111",
  56347=>"111110110",
  56348=>"000111110",
  56349=>"110101001",
  56350=>"111110110",
  56351=>"000000111",
  56352=>"000000000",
  56353=>"000000000",
  56354=>"111010111",
  56355=>"111111111",
  56356=>"000000000",
  56357=>"111110000",
  56358=>"111111111",
  56359=>"111111111",
  56360=>"111111111",
  56361=>"000000111",
  56362=>"111111100",
  56363=>"111111000",
  56364=>"111111111",
  56365=>"111111111",
  56366=>"111111111",
  56367=>"001000000",
  56368=>"001100100",
  56369=>"001010111",
  56370=>"111111111",
  56371=>"000000000",
  56372=>"110110000",
  56373=>"000000010",
  56374=>"111111110",
  56375=>"101000000",
  56376=>"000000110",
  56377=>"001111000",
  56378=>"111111111",
  56379=>"101000000",
  56380=>"001001000",
  56381=>"111111111",
  56382=>"000000000",
  56383=>"111111111",
  56384=>"111111111",
  56385=>"111111111",
  56386=>"111111000",
  56387=>"000000111",
  56388=>"011001001",
  56389=>"000000000",
  56390=>"000000111",
  56391=>"011011000",
  56392=>"100110111",
  56393=>"111111111",
  56394=>"111111000",
  56395=>"100101100",
  56396=>"000000000",
  56397=>"101001101",
  56398=>"000000000",
  56399=>"111111111",
  56400=>"111111111",
  56401=>"000000000",
  56402=>"101111101",
  56403=>"011111111",
  56404=>"000000000",
  56405=>"000000101",
  56406=>"111100100",
  56407=>"000000000",
  56408=>"000000000",
  56409=>"000000000",
  56410=>"011001001",
  56411=>"001001001",
  56412=>"001001000",
  56413=>"000100110",
  56414=>"001001111",
  56415=>"000000000",
  56416=>"111111110",
  56417=>"000000011",
  56418=>"111111100",
  56419=>"111111111",
  56420=>"000000000",
  56421=>"111111000",
  56422=>"000000000",
  56423=>"111111111",
  56424=>"111000000",
  56425=>"111101000",
  56426=>"011001000",
  56427=>"000001111",
  56428=>"000000001",
  56429=>"111110010",
  56430=>"111100000",
  56431=>"111111111",
  56432=>"001011111",
  56433=>"000000000",
  56434=>"000000000",
  56435=>"111001000",
  56436=>"000000001",
  56437=>"111111111",
  56438=>"000000000",
  56439=>"000000000",
  56440=>"100110100",
  56441=>"111111111",
  56442=>"001011011",
  56443=>"000000000",
  56444=>"000000000",
  56445=>"011011011",
  56446=>"000000000",
  56447=>"111111111",
  56448=>"110100100",
  56449=>"000100000",
  56450=>"110000000",
  56451=>"110100000",
  56452=>"110111111",
  56453=>"000000111",
  56454=>"000001001",
  56455=>"000000000",
  56456=>"000000000",
  56457=>"000000000",
  56458=>"111101111",
  56459=>"000100000",
  56460=>"100100110",
  56461=>"100100000",
  56462=>"100000000",
  56463=>"011000000",
  56464=>"000000000",
  56465=>"111100111",
  56466=>"101111111",
  56467=>"111111111",
  56468=>"001011011",
  56469=>"100000000",
  56470=>"111111111",
  56471=>"000000000",
  56472=>"111111100",
  56473=>"100100110",
  56474=>"000000000",
  56475=>"111111111",
  56476=>"001000001",
  56477=>"000101111",
  56478=>"100111111",
  56479=>"111000000",
  56480=>"000000110",
  56481=>"111100110",
  56482=>"001011000",
  56483=>"111111111",
  56484=>"011001000",
  56485=>"000000101",
  56486=>"111111000",
  56487=>"010000100",
  56488=>"000000100",
  56489=>"000000000",
  56490=>"000000000",
  56491=>"000000010",
  56492=>"000000000",
  56493=>"111111110",
  56494=>"110100100",
  56495=>"111110100",
  56496=>"000111111",
  56497=>"000110000",
  56498=>"110111111",
  56499=>"111111111",
  56500=>"000000000",
  56501=>"111111100",
  56502=>"010111111",
  56503=>"111111001",
  56504=>"001111111",
  56505=>"111111111",
  56506=>"011001101",
  56507=>"011000000",
  56508=>"111111111",
  56509=>"111110100",
  56510=>"111111011",
  56511=>"000000111",
  56512=>"101111111",
  56513=>"111111111",
  56514=>"000111011",
  56515=>"000000000",
  56516=>"111010100",
  56517=>"011000000",
  56518=>"111111111",
  56519=>"011111111",
  56520=>"010000010",
  56521=>"001000000",
  56522=>"111111111",
  56523=>"001011111",
  56524=>"101111000",
  56525=>"110011000",
  56526=>"000001001",
  56527=>"001000000",
  56528=>"111111111",
  56529=>"101000000",
  56530=>"000000000",
  56531=>"000000000",
  56532=>"000000000",
  56533=>"000000000",
  56534=>"000000000",
  56535=>"111000000",
  56536=>"111111111",
  56537=>"111111000",
  56538=>"111111111",
  56539=>"111110100",
  56540=>"101101000",
  56541=>"000100111",
  56542=>"000000000",
  56543=>"111111111",
  56544=>"111111111",
  56545=>"101001111",
  56546=>"000000010",
  56547=>"001000100",
  56548=>"000000000",
  56549=>"100110000",
  56550=>"111111111",
  56551=>"100000101",
  56552=>"000010111",
  56553=>"100111111",
  56554=>"001000011",
  56555=>"010000000",
  56556=>"111111110",
  56557=>"100110000",
  56558=>"011100000",
  56559=>"111000110",
  56560=>"110111111",
  56561=>"001111000",
  56562=>"000000110",
  56563=>"011111111",
  56564=>"111111000",
  56565=>"000000000",
  56566=>"010000010",
  56567=>"000000000",
  56568=>"111111111",
  56569=>"000000000",
  56570=>"111111111",
  56571=>"000000000",
  56572=>"100100100",
  56573=>"110111111",
  56574=>"111111101",
  56575=>"100000000",
  56576=>"111100100",
  56577=>"111111111",
  56578=>"000111111",
  56579=>"000111111",
  56580=>"111000100",
  56581=>"111111111",
  56582=>"111111111",
  56583=>"000100110",
  56584=>"011011111",
  56585=>"000000001",
  56586=>"111110110",
  56587=>"111111111",
  56588=>"000000000",
  56589=>"000000110",
  56590=>"111111111",
  56591=>"111000101",
  56592=>"010000000",
  56593=>"001110110",
  56594=>"100110000",
  56595=>"000000000",
  56596=>"000000000",
  56597=>"000000000",
  56598=>"000000000",
  56599=>"000111111",
  56600=>"000000000",
  56601=>"000000000",
  56602=>"101111111",
  56603=>"110111111",
  56604=>"011111111",
  56605=>"000110011",
  56606=>"111001111",
  56607=>"111111111",
  56608=>"110011000",
  56609=>"000000100",
  56610=>"111111111",
  56611=>"000000101",
  56612=>"000000000",
  56613=>"000000000",
  56614=>"000000000",
  56615=>"000000000",
  56616=>"111011001",
  56617=>"000100100",
  56618=>"111111100",
  56619=>"000110111",
  56620=>"000000000",
  56621=>"111110110",
  56622=>"111111111",
  56623=>"101111111",
  56624=>"000001111",
  56625=>"111111101",
  56626=>"111111111",
  56627=>"010000000",
  56628=>"111111111",
  56629=>"000000000",
  56630=>"001000001",
  56631=>"000001111",
  56632=>"110000000",
  56633=>"001111100",
  56634=>"111111111",
  56635=>"111111000",
  56636=>"111011111",
  56637=>"000011000",
  56638=>"111111100",
  56639=>"001000000",
  56640=>"000000000",
  56641=>"111001000",
  56642=>"111111100",
  56643=>"000000000",
  56644=>"000000000",
  56645=>"110111111",
  56646=>"000100000",
  56647=>"111111111",
  56648=>"000000000",
  56649=>"111111111",
  56650=>"111100111",
  56651=>"000001001",
  56652=>"111111111",
  56653=>"000000000",
  56654=>"111111111",
  56655=>"110110111",
  56656=>"000001001",
  56657=>"001001011",
  56658=>"000000000",
  56659=>"000000111",
  56660=>"000000010",
  56661=>"111111111",
  56662=>"000110010",
  56663=>"111111111",
  56664=>"000001111",
  56665=>"000000000",
  56666=>"000111111",
  56667=>"111110111",
  56668=>"111111111",
  56669=>"000000000",
  56670=>"000000000",
  56671=>"111111111",
  56672=>"111010000",
  56673=>"111111111",
  56674=>"111001000",
  56675=>"000000010",
  56676=>"010011011",
  56677=>"000000000",
  56678=>"111111111",
  56679=>"001001111",
  56680=>"000000000",
  56681=>"100100000",
  56682=>"000000000",
  56683=>"111101000",
  56684=>"000001111",
  56685=>"011001001",
  56686=>"100100100",
  56687=>"111111101",
  56688=>"000000000",
  56689=>"111111000",
  56690=>"111111111",
  56691=>"000000100",
  56692=>"111000000",
  56693=>"000000000",
  56694=>"000000100",
  56695=>"000011011",
  56696=>"100100111",
  56697=>"111111111",
  56698=>"000000011",
  56699=>"011011111",
  56700=>"011011011",
  56701=>"000000000",
  56702=>"111110100",
  56703=>"000000000",
  56704=>"111111111",
  56705=>"111111111",
  56706=>"000000000",
  56707=>"111000101",
  56708=>"111111111",
  56709=>"011111111",
  56710=>"110111101",
  56711=>"000100100",
  56712=>"111110000",
  56713=>"001000000",
  56714=>"111111111",
  56715=>"111111111",
  56716=>"000000000",
  56717=>"110110110",
  56718=>"000000100",
  56719=>"111101101",
  56720=>"101000000",
  56721=>"111101111",
  56722=>"111111111",
  56723=>"111111111",
  56724=>"011000000",
  56725=>"001001111",
  56726=>"111111111",
  56727=>"000000000",
  56728=>"001000100",
  56729=>"111111111",
  56730=>"011001001",
  56731=>"000101000",
  56732=>"101111111",
  56733=>"100100100",
  56734=>"111111000",
  56735=>"100111111",
  56736=>"101101100",
  56737=>"001001011",
  56738=>"000100110",
  56739=>"111111111",
  56740=>"111100100",
  56741=>"001000001",
  56742=>"100100100",
  56743=>"000110010",
  56744=>"111011111",
  56745=>"011011011",
  56746=>"000000110",
  56747=>"000110110",
  56748=>"000000111",
  56749=>"011001000",
  56750=>"001111111",
  56751=>"000100111",
  56752=>"100110000",
  56753=>"000000000",
  56754=>"111111111",
  56755=>"101111111",
  56756=>"000000000",
  56757=>"000000000",
  56758=>"000000000",
  56759=>"100100000",
  56760=>"111111000",
  56761=>"000100100",
  56762=>"000001000",
  56763=>"110000111",
  56764=>"010010000",
  56765=>"111111111",
  56766=>"101110010",
  56767=>"000000100",
  56768=>"111111111",
  56769=>"000000000",
  56770=>"000000101",
  56771=>"000000000",
  56772=>"001001101",
  56773=>"000000000",
  56774=>"111101000",
  56775=>"000000000",
  56776=>"001000000",
  56777=>"111101101",
  56778=>"001111111",
  56779=>"111111111",
  56780=>"011000001",
  56781=>"000101000",
  56782=>"111001011",
  56783=>"000100110",
  56784=>"000000000",
  56785=>"000001000",
  56786=>"011000000",
  56787=>"111111111",
  56788=>"000000000",
  56789=>"111111001",
  56790=>"000111111",
  56791=>"000110100",
  56792=>"111111111",
  56793=>"110110000",
  56794=>"000000000",
  56795=>"101100100",
  56796=>"001011011",
  56797=>"000000000",
  56798=>"100110110",
  56799=>"001000100",
  56800=>"110111111",
  56801=>"011010110",
  56802=>"111111000",
  56803=>"000000111",
  56804=>"111011001",
  56805=>"000000010",
  56806=>"000101101",
  56807=>"000010000",
  56808=>"000000111",
  56809=>"110000010",
  56810=>"111111111",
  56811=>"001001001",
  56812=>"011100111",
  56813=>"000001001",
  56814=>"100100100",
  56815=>"110111001",
  56816=>"001011000",
  56817=>"111010111",
  56818=>"000000000",
  56819=>"111111111",
  56820=>"111111000",
  56821=>"111111111",
  56822=>"111000000",
  56823=>"000000000",
  56824=>"000000100",
  56825=>"111111111",
  56826=>"000000000",
  56827=>"100000100",
  56828=>"101111111",
  56829=>"111011011",
  56830=>"111110000",
  56831=>"000110010",
  56832=>"111111111",
  56833=>"001001011",
  56834=>"100000000",
  56835=>"001111010",
  56836=>"000000000",
  56837=>"001000100",
  56838=>"110100100",
  56839=>"111111100",
  56840=>"111111111",
  56841=>"000000010",
  56842=>"111011111",
  56843=>"000101000",
  56844=>"100000111",
  56845=>"001011110",
  56846=>"100100101",
  56847=>"010100111",
  56848=>"111111011",
  56849=>"100101111",
  56850=>"000111111",
  56851=>"000100100",
  56852=>"011111011",
  56853=>"111111111",
  56854=>"111000001",
  56855=>"111101110",
  56856=>"010011111",
  56857=>"011011000",
  56858=>"111011111",
  56859=>"011001000",
  56860=>"001000000",
  56861=>"111110100",
  56862=>"001001001",
  56863=>"011110110",
  56864=>"000000000",
  56865=>"110111111",
  56866=>"111111111",
  56867=>"000001000",
  56868=>"000111111",
  56869=>"111110000",
  56870=>"111111111",
  56871=>"011111000",
  56872=>"000000110",
  56873=>"000011111",
  56874=>"000000000",
  56875=>"111111111",
  56876=>"111111111",
  56877=>"000000000",
  56878=>"111111111",
  56879=>"111111111",
  56880=>"111111001",
  56881=>"000000000",
  56882=>"000000100",
  56883=>"000000000",
  56884=>"000000000",
  56885=>"100111111",
  56886=>"000001000",
  56887=>"000000001",
  56888=>"001111111",
  56889=>"001010111",
  56890=>"000010110",
  56891=>"000000101",
  56892=>"100000011",
  56893=>"111011111",
  56894=>"111111111",
  56895=>"111111111",
  56896=>"001001000",
  56897=>"011011011",
  56898=>"111000010",
  56899=>"000000110",
  56900=>"000000101",
  56901=>"010100110",
  56902=>"111000000",
  56903=>"000000000",
  56904=>"111111111",
  56905=>"000000101",
  56906=>"111111100",
  56907=>"111111111",
  56908=>"001000000",
  56909=>"111111111",
  56910=>"000000000",
  56911=>"111111111",
  56912=>"000000100",
  56913=>"110000100",
  56914=>"000000000",
  56915=>"000100000",
  56916=>"100000000",
  56917=>"000000000",
  56918=>"001000000",
  56919=>"000000000",
  56920=>"101011000",
  56921=>"010000000",
  56922=>"011111111",
  56923=>"000010111",
  56924=>"111001111",
  56925=>"000000000",
  56926=>"001000000",
  56927=>"001001110",
  56928=>"000111111",
  56929=>"111111111",
  56930=>"000000000",
  56931=>"101000111",
  56932=>"111111111",
  56933=>"111001000",
  56934=>"001000110",
  56935=>"001011011",
  56936=>"001000000",
  56937=>"010010000",
  56938=>"000011111",
  56939=>"010111111",
  56940=>"000111110",
  56941=>"000000000",
  56942=>"000000010",
  56943=>"100101101",
  56944=>"000000000",
  56945=>"000000000",
  56946=>"111111011",
  56947=>"001111111",
  56948=>"001011111",
  56949=>"110000000",
  56950=>"000000000",
  56951=>"010110010",
  56952=>"111111010",
  56953=>"000101000",
  56954=>"110111111",
  56955=>"001001000",
  56956=>"100101101",
  56957=>"011011100",
  56958=>"111111000",
  56959=>"001000000",
  56960=>"000000000",
  56961=>"001111110",
  56962=>"110110000",
  56963=>"000000000",
  56964=>"000100011",
  56965=>"000000000",
  56966=>"111111111",
  56967=>"111010111",
  56968=>"111111111",
  56969=>"100111111",
  56970=>"000001111",
  56971=>"000000000",
  56972=>"110111111",
  56973=>"111111000",
  56974=>"001000001",
  56975=>"110111001",
  56976=>"000000000",
  56977=>"011000001",
  56978=>"111111111",
  56979=>"111111101",
  56980=>"001000000",
  56981=>"000000001",
  56982=>"000010110",
  56983=>"000000000",
  56984=>"001000000",
  56985=>"111111111",
  56986=>"000111000",
  56987=>"111111100",
  56988=>"000100111",
  56989=>"111111000",
  56990=>"000000000",
  56991=>"000000000",
  56992=>"111111111",
  56993=>"100111111",
  56994=>"001001000",
  56995=>"000000000",
  56996=>"100001010",
  56997=>"000000000",
  56998=>"111000000",
  56999=>"001000001",
  57000=>"011111110",
  57001=>"000110011",
  57002=>"000110000",
  57003=>"111111111",
  57004=>"001110110",
  57005=>"000000000",
  57006=>"000000000",
  57007=>"000000000",
  57008=>"000010110",
  57009=>"000000010",
  57010=>"100110110",
  57011=>"111000000",
  57012=>"001000110",
  57013=>"110110100",
  57014=>"000000000",
  57015=>"111111111",
  57016=>"111111110",
  57017=>"000000000",
  57018=>"110100001",
  57019=>"000000001",
  57020=>"110111111",
  57021=>"111111111",
  57022=>"111111111",
  57023=>"100111111",
  57024=>"111000010",
  57025=>"111101101",
  57026=>"000000000",
  57027=>"000100110",
  57028=>"111111111",
  57029=>"000101111",
  57030=>"000000000",
  57031=>"000000011",
  57032=>"000010010",
  57033=>"000001011",
  57034=>"101101101",
  57035=>"000001001",
  57036=>"000000000",
  57037=>"101000000",
  57038=>"000000111",
  57039=>"000000000",
  57040=>"111101000",
  57041=>"111100100",
  57042=>"110100000",
  57043=>"111111111",
  57044=>"111111111",
  57045=>"111011011",
  57046=>"111111111",
  57047=>"100000000",
  57048=>"000000000",
  57049=>"001001100",
  57050=>"111111111",
  57051=>"000000011",
  57052=>"100110000",
  57053=>"100110000",
  57054=>"100100000",
  57055=>"100111111",
  57056=>"011111011",
  57057=>"111001011",
  57058=>"000000000",
  57059=>"000000000",
  57060=>"000000000",
  57061=>"111111111",
  57062=>"111001001",
  57063=>"111011001",
  57064=>"000000000",
  57065=>"000111111",
  57066=>"000011111",
  57067=>"100000000",
  57068=>"111111111",
  57069=>"111111111",
  57070=>"011111101",
  57071=>"111111011",
  57072=>"000000000",
  57073=>"000000000",
  57074=>"000010111",
  57075=>"001011011",
  57076=>"111101111",
  57077=>"110110110",
  57078=>"111111111",
  57079=>"000010010",
  57080=>"000000000",
  57081=>"110000000",
  57082=>"000000000",
  57083=>"111111011",
  57084=>"110110000",
  57085=>"011110110",
  57086=>"001001000",
  57087=>"100101111",
  57088=>"011011111",
  57089=>"100100111",
  57090=>"000000100",
  57091=>"111111111",
  57092=>"001001000",
  57093=>"001000000",
  57094=>"000000000",
  57095=>"000100100",
  57096=>"111111111",
  57097=>"111111101",
  57098=>"111011111",
  57099=>"111111111",
  57100=>"000000110",
  57101=>"000111111",
  57102=>"100100000",
  57103=>"000111111",
  57104=>"000000000",
  57105=>"000000000",
  57106=>"011000001",
  57107=>"101101100",
  57108=>"011000000",
  57109=>"000000111",
  57110=>"000010111",
  57111=>"000000101",
  57112=>"111111111",
  57113=>"011100100",
  57114=>"001101111",
  57115=>"000000000",
  57116=>"111111111",
  57117=>"011111111",
  57118=>"000000000",
  57119=>"111111111",
  57120=>"100100101",
  57121=>"000000000",
  57122=>"111111111",
  57123=>"000000000",
  57124=>"111111111",
  57125=>"100000111",
  57126=>"010111111",
  57127=>"000000011",
  57128=>"111101011",
  57129=>"100110000",
  57130=>"101111010",
  57131=>"011000101",
  57132=>"100000001",
  57133=>"110110111",
  57134=>"100000000",
  57135=>"000000000",
  57136=>"111111111",
  57137=>"011011001",
  57138=>"000001111",
  57139=>"000000000",
  57140=>"111111111",
  57141=>"111111011",
  57142=>"001001011",
  57143=>"001000000",
  57144=>"110100000",
  57145=>"111110000",
  57146=>"110111111",
  57147=>"000000110",
  57148=>"010001111",
  57149=>"001100100",
  57150=>"000000000",
  57151=>"010000000",
  57152=>"000100100",
  57153=>"001011111",
  57154=>"000011111",
  57155=>"000000000",
  57156=>"100111101",
  57157=>"111011111",
  57158=>"000000000",
  57159=>"111111111",
  57160=>"011111111",
  57161=>"011000000",
  57162=>"010111010",
  57163=>"000000000",
  57164=>"111111111",
  57165=>"000111101",
  57166=>"000000000",
  57167=>"000000100",
  57168=>"111111101",
  57169=>"000110100",
  57170=>"100100000",
  57171=>"000000000",
  57172=>"100000001",
  57173=>"111011011",
  57174=>"011100100",
  57175=>"111111111",
  57176=>"000000001",
  57177=>"000000000",
  57178=>"000000000",
  57179=>"111001010",
  57180=>"000000000",
  57181=>"000000111",
  57182=>"000000011",
  57183=>"111111111",
  57184=>"011110000",
  57185=>"000000000",
  57186=>"110110101",
  57187=>"000000000",
  57188=>"101111111",
  57189=>"000000010",
  57190=>"111000111",
  57191=>"001001000",
  57192=>"000001001",
  57193=>"000000000",
  57194=>"000000000",
  57195=>"111101111",
  57196=>"110110100",
  57197=>"110000011",
  57198=>"111000111",
  57199=>"111101100",
  57200=>"000000000",
  57201=>"111100101",
  57202=>"000000000",
  57203=>"111111101",
  57204=>"110110000",
  57205=>"100100110",
  57206=>"001111111",
  57207=>"000100000",
  57208=>"000000000",
  57209=>"010010111",
  57210=>"000000000",
  57211=>"111001000",
  57212=>"000000111",
  57213=>"111111111",
  57214=>"010000000",
  57215=>"000000000",
  57216=>"000000000",
  57217=>"101101110",
  57218=>"000001001",
  57219=>"000000000",
  57220=>"011011000",
  57221=>"100111001",
  57222=>"011001000",
  57223=>"000110001",
  57224=>"000000111",
  57225=>"000000000",
  57226=>"111110100",
  57227=>"000000010",
  57228=>"111111111",
  57229=>"000110010",
  57230=>"111000000",
  57231=>"000000000",
  57232=>"000000000",
  57233=>"000000000",
  57234=>"001000100",
  57235=>"010110111",
  57236=>"111111111",
  57237=>"011001001",
  57238=>"111111111",
  57239=>"100000100",
  57240=>"110110111",
  57241=>"100000000",
  57242=>"000100110",
  57243=>"001000000",
  57244=>"000001100",
  57245=>"111111000",
  57246=>"110110000",
  57247=>"000111111",
  57248=>"100100000",
  57249=>"100000000",
  57250=>"000000100",
  57251=>"001011111",
  57252=>"000100100",
  57253=>"000000000",
  57254=>"001000111",
  57255=>"101101111",
  57256=>"011001111",
  57257=>"001001000",
  57258=>"001111111",
  57259=>"100000000",
  57260=>"000000000",
  57261=>"101000000",
  57262=>"011111111",
  57263=>"000001000",
  57264=>"011101111",
  57265=>"111111111",
  57266=>"000000000",
  57267=>"111111111",
  57268=>"111111110",
  57269=>"111000000",
  57270=>"100100111",
  57271=>"111111110",
  57272=>"111110000",
  57273=>"111111111",
  57274=>"111111111",
  57275=>"000010000",
  57276=>"000111000",
  57277=>"111100110",
  57278=>"000100101",
  57279=>"111111111",
  57280=>"001010001",
  57281=>"001000000",
  57282=>"000000000",
  57283=>"000100100",
  57284=>"000000000",
  57285=>"001101111",
  57286=>"001111110",
  57287=>"000000100",
  57288=>"000000001",
  57289=>"000000000",
  57290=>"001111110",
  57291=>"010000110",
  57292=>"100000111",
  57293=>"100101111",
  57294=>"000000000",
  57295=>"011111111",
  57296=>"001111111",
  57297=>"010110100",
  57298=>"000000000",
  57299=>"011000111",
  57300=>"100000000",
  57301=>"001000000",
  57302=>"111011011",
  57303=>"001000011",
  57304=>"000011011",
  57305=>"000011111",
  57306=>"000000000",
  57307=>"111111111",
  57308=>"111111111",
  57309=>"100001001",
  57310=>"001011011",
  57311=>"101011011",
  57312=>"111111111",
  57313=>"010000011",
  57314=>"000001001",
  57315=>"000000000",
  57316=>"110111101",
  57317=>"000000000",
  57318=>"000000001",
  57319=>"000000000",
  57320=>"001000000",
  57321=>"000000000",
  57322=>"010110001",
  57323=>"111111111",
  57324=>"111111111",
  57325=>"111100000",
  57326=>"111111011",
  57327=>"110110110",
  57328=>"110110110",
  57329=>"111111111",
  57330=>"111000101",
  57331=>"000100110",
  57332=>"001000000",
  57333=>"011011000",
  57334=>"001011111",
  57335=>"001001101",
  57336=>"000000000",
  57337=>"100110110",
  57338=>"000000001",
  57339=>"111110110",
  57340=>"001001000",
  57341=>"111111111",
  57342=>"111111111",
  57343=>"000110110",
  57344=>"000000001",
  57345=>"100110110",
  57346=>"111111111",
  57347=>"111111111",
  57348=>"111111111",
  57349=>"110010010",
  57350=>"110000000",
  57351=>"000000000",
  57352=>"000000000",
  57353=>"100000001",
  57354=>"000011011",
  57355=>"000011111",
  57356=>"100110110",
  57357=>"110111111",
  57358=>"111000001",
  57359=>"111111111",
  57360=>"100000001",
  57361=>"000111001",
  57362=>"111011111",
  57363=>"110111011",
  57364=>"000000110",
  57365=>"010000000",
  57366=>"000000000",
  57367=>"111111011",
  57368=>"001011110",
  57369=>"111110111",
  57370=>"111111100",
  57371=>"111111010",
  57372=>"000000100",
  57373=>"111110110",
  57374=>"111111111",
  57375=>"100000001",
  57376=>"000000000",
  57377=>"110110011",
  57378=>"100000000",
  57379=>"010011001",
  57380=>"111011110",
  57381=>"111111111",
  57382=>"000000100",
  57383=>"000110111",
  57384=>"111000001",
  57385=>"011011111",
  57386=>"111111110",
  57387=>"011011011",
  57388=>"011111111",
  57389=>"111111000",
  57390=>"110110111",
  57391=>"000000000",
  57392=>"111111111",
  57393=>"000000100",
  57394=>"111101001",
  57395=>"000000000",
  57396=>"000000000",
  57397=>"011001001",
  57398=>"000011111",
  57399=>"100100101",
  57400=>"011011111",
  57401=>"001000011",
  57402=>"111111001",
  57403=>"000000000",
  57404=>"100100111",
  57405=>"011011001",
  57406=>"100100000",
  57407=>"001000000",
  57408=>"000100111",
  57409=>"000010000",
  57410=>"000110000",
  57411=>"111111111",
  57412=>"000000000",
  57413=>"000000011",
  57414=>"011000000",
  57415=>"111111101",
  57416=>"111001111",
  57417=>"000000000",
  57418=>"111111111",
  57419=>"111100110",
  57420=>"000000110",
  57421=>"110000000",
  57422=>"111101000",
  57423=>"000000101",
  57424=>"000000000",
  57425=>"011111011",
  57426=>"000000000",
  57427=>"110001011",
  57428=>"000000101",
  57429=>"111000000",
  57430=>"111110110",
  57431=>"000000000",
  57432=>"011001001",
  57433=>"111000000",
  57434=>"111110000",
  57435=>"100000000",
  57436=>"000000111",
  57437=>"000001111",
  57438=>"000000010",
  57439=>"000001111",
  57440=>"111111111",
  57441=>"001000000",
  57442=>"000001000",
  57443=>"000000000",
  57444=>"111111000",
  57445=>"000011000",
  57446=>"000000000",
  57447=>"111111111",
  57448=>"111111111",
  57449=>"111111011",
  57450=>"111000110",
  57451=>"000000000",
  57452=>"011011111",
  57453=>"000000100",
  57454=>"111111111",
  57455=>"000000000",
  57456=>"000000000",
  57457=>"000010111",
  57458=>"001001101",
  57459=>"000111101",
  57460=>"010000000",
  57461=>"010011111",
  57462=>"011011000",
  57463=>"010000000",
  57464=>"111111111",
  57465=>"111111100",
  57466=>"000000000",
  57467=>"111111011",
  57468=>"000100111",
  57469=>"111111111",
  57470=>"111111000",
  57471=>"000000000",
  57472=>"000000000",
  57473=>"000011000",
  57474=>"111111001",
  57475=>"100000100",
  57476=>"000000000",
  57477=>"000000000",
  57478=>"000010010",
  57479=>"011000000",
  57480=>"101000100",
  57481=>"000001001",
  57482=>"000000000",
  57483=>"111111111",
  57484=>"000000001",
  57485=>"111100110",
  57486=>"111111111",
  57487=>"000000110",
  57488=>"000000000",
  57489=>"001001111",
  57490=>"011111000",
  57491=>"111111000",
  57492=>"000001001",
  57493=>"000110110",
  57494=>"000000000",
  57495=>"111000000",
  57496=>"111111111",
  57497=>"000010110",
  57498=>"110100000",
  57499=>"111111111",
  57500=>"111100000",
  57501=>"000110111",
  57502=>"100100111",
  57503=>"111111110",
  57504=>"111001000",
  57505=>"000000000",
  57506=>"000000000",
  57507=>"101001000",
  57508=>"111111111",
  57509=>"111001111",
  57510=>"011000000",
  57511=>"100000100",
  57512=>"000000110",
  57513=>"000000000",
  57514=>"111111010",
  57515=>"111100110",
  57516=>"111001001",
  57517=>"111111101",
  57518=>"001011111",
  57519=>"001001000",
  57520=>"000000011",
  57521=>"011101101",
  57522=>"111111111",
  57523=>"000000000",
  57524=>"110111111",
  57525=>"000000000",
  57526=>"000000110",
  57527=>"111111101",
  57528=>"111111111",
  57529=>"111111011",
  57530=>"101111110",
  57531=>"101101001",
  57532=>"000000111",
  57533=>"111111111",
  57534=>"111111111",
  57535=>"001000000",
  57536=>"000000000",
  57537=>"011011011",
  57538=>"000000000",
  57539=>"110110010",
  57540=>"000000011",
  57541=>"001011111",
  57542=>"010010000",
  57543=>"011111110",
  57544=>"111111111",
  57545=>"000001001",
  57546=>"000000000",
  57547=>"000000000",
  57548=>"111100111",
  57549=>"111111111",
  57550=>"100111111",
  57551=>"000000000",
  57552=>"000000011",
  57553=>"111111100",
  57554=>"000100000",
  57555=>"111000000",
  57556=>"001000110",
  57557=>"111111110",
  57558=>"111010000",
  57559=>"111011111",
  57560=>"011111111",
  57561=>"011111000",
  57562=>"011010000",
  57563=>"111000000",
  57564=>"000100111",
  57565=>"100000000",
  57566=>"001011011",
  57567=>"111111011",
  57568=>"001000000",
  57569=>"000011011",
  57570=>"011011010",
  57571=>"111100000",
  57572=>"100100011",
  57573=>"100110110",
  57574=>"100100100",
  57575=>"110111111",
  57576=>"000000000",
  57577=>"000001001",
  57578=>"111011000",
  57579=>"111111111",
  57580=>"000000000",
  57581=>"111100000",
  57582=>"000010111",
  57583=>"000000000",
  57584=>"110111111",
  57585=>"110000001",
  57586=>"111111000",
  57587=>"111111011",
  57588=>"110111111",
  57589=>"000110111",
  57590=>"111111111",
  57591=>"000000000",
  57592=>"000110000",
  57593=>"111111111",
  57594=>"101000001",
  57595=>"111111111",
  57596=>"000000000",
  57597=>"001000111",
  57598=>"101000011",
  57599=>"000000000",
  57600=>"011000000",
  57601=>"111101111",
  57602=>"000000110",
  57603=>"110111100",
  57604=>"111111111",
  57605=>"111011111",
  57606=>"000000110",
  57607=>"000000110",
  57608=>"110111000",
  57609=>"011000000",
  57610=>"111000000",
  57611=>"111111111",
  57612=>"010010000",
  57613=>"001000011",
  57614=>"111111101",
  57615=>"111000000",
  57616=>"111110000",
  57617=>"111111011",
  57618=>"011001011",
  57619=>"001111011",
  57620=>"110101000",
  57621=>"000000001",
  57622=>"100110111",
  57623=>"111011001",
  57624=>"011001111",
  57625=>"000000100",
  57626=>"111111111",
  57627=>"000000011",
  57628=>"110110111",
  57629=>"000000000",
  57630=>"111111111",
  57631=>"001000000",
  57632=>"001001101",
  57633=>"000000000",
  57634=>"000110111",
  57635=>"100000111",
  57636=>"111011111",
  57637=>"011011000",
  57638=>"111111111",
  57639=>"000001010",
  57640=>"000111111",
  57641=>"000000000",
  57642=>"011001001",
  57643=>"000000001",
  57644=>"001110110",
  57645=>"001111111",
  57646=>"000000111",
  57647=>"100000100",
  57648=>"000000111",
  57649=>"101001000",
  57650=>"000000100",
  57651=>"011111111",
  57652=>"000000000",
  57653=>"111111101",
  57654=>"111100100",
  57655=>"000011111",
  57656=>"010110110",
  57657=>"111000000",
  57658=>"101100000",
  57659=>"000000000",
  57660=>"100110000",
  57661=>"000000000",
  57662=>"110111110",
  57663=>"101101001",
  57664=>"000000000",
  57665=>"001100110",
  57666=>"111110011",
  57667=>"111111111",
  57668=>"001000100",
  57669=>"111111111",
  57670=>"000000000",
  57671=>"110111111",
  57672=>"111111111",
  57673=>"000000000",
  57674=>"000000000",
  57675=>"000100100",
  57676=>"011101111",
  57677=>"111110111",
  57678=>"111111110",
  57679=>"110001111",
  57680=>"000111100",
  57681=>"100110011",
  57682=>"111001011",
  57683=>"101100100",
  57684=>"000001001",
  57685=>"011010011",
  57686=>"000000001",
  57687=>"001000011",
  57688=>"101000000",
  57689=>"111100110",
  57690=>"100001100",
  57691=>"110010111",
  57692=>"111111001",
  57693=>"000000000",
  57694=>"000111001",
  57695=>"111111111",
  57696=>"000000000",
  57697=>"000000101",
  57698=>"111111111",
  57699=>"111111111",
  57700=>"000000000",
  57701=>"111001101",
  57702=>"000110110",
  57703=>"000000000",
  57704=>"001001000",
  57705=>"110111110",
  57706=>"000000010",
  57707=>"100000011",
  57708=>"111111100",
  57709=>"111110110",
  57710=>"100111111",
  57711=>"000010010",
  57712=>"000000111",
  57713=>"110000000",
  57714=>"111101101",
  57715=>"001111111",
  57716=>"000010000",
  57717=>"111111001",
  57718=>"000000111",
  57719=>"000000000",
  57720=>"000000000",
  57721=>"000001011",
  57722=>"111111111",
  57723=>"001011001",
  57724=>"010000001",
  57725=>"001000001",
  57726=>"001000010",
  57727=>"111000000",
  57728=>"110111111",
  57729=>"001000000",
  57730=>"110110111",
  57731=>"111111111",
  57732=>"011111111",
  57733=>"111111111",
  57734=>"100000000",
  57735=>"100101101",
  57736=>"111111111",
  57737=>"010111010",
  57738=>"001000000",
  57739=>"111111010",
  57740=>"111100000",
  57741=>"111111111",
  57742=>"000001000",
  57743=>"000000000",
  57744=>"111111011",
  57745=>"110110111",
  57746=>"011001011",
  57747=>"111111110",
  57748=>"000000111",
  57749=>"000000000",
  57750=>"000000011",
  57751=>"110100000",
  57752=>"000001011",
  57753=>"100000000",
  57754=>"011000000",
  57755=>"001001001",
  57756=>"111111000",
  57757=>"111111111",
  57758=>"000111100",
  57759=>"111111111",
  57760=>"111111111",
  57761=>"111101111",
  57762=>"111111000",
  57763=>"111111111",
  57764=>"111010011",
  57765=>"000000000",
  57766=>"010111111",
  57767=>"111111100",
  57768=>"110000000",
  57769=>"000000000",
  57770=>"110110111",
  57771=>"001000000",
  57772=>"111111111",
  57773=>"111011011",
  57774=>"000000000",
  57775=>"001011011",
  57776=>"101000000",
  57777=>"111111100",
  57778=>"110110100",
  57779=>"001000000",
  57780=>"000000000",
  57781=>"111110110",
  57782=>"100110111",
  57783=>"000000100",
  57784=>"111000000",
  57785=>"100110111",
  57786=>"111110110",
  57787=>"111111101",
  57788=>"000000100",
  57789=>"000011000",
  57790=>"111000000",
  57791=>"100101101",
  57792=>"000000000",
  57793=>"000000000",
  57794=>"000000000",
  57795=>"000000000",
  57796=>"111000100",
  57797=>"011000111",
  57798=>"011000000",
  57799=>"111111000",
  57800=>"110010011",
  57801=>"111000000",
  57802=>"111000000",
  57803=>"000000011",
  57804=>"000110100",
  57805=>"110110111",
  57806=>"011000000",
  57807=>"010000110",
  57808=>"100000000",
  57809=>"000110111",
  57810=>"111111111",
  57811=>"111000110",
  57812=>"011111111",
  57813=>"111101111",
  57814=>"101000000",
  57815=>"000011011",
  57816=>"111100100",
  57817=>"001000000",
  57818=>"100000000",
  57819=>"000000000",
  57820=>"000110000",
  57821=>"000000110",
  57822=>"000000111",
  57823=>"000110110",
  57824=>"110001001",
  57825=>"111101111",
  57826=>"111111111",
  57827=>"111111111",
  57828=>"111111111",
  57829=>"111111111",
  57830=>"000000000",
  57831=>"011010001",
  57832=>"011001001",
  57833=>"000000100",
  57834=>"000000000",
  57835=>"001011011",
  57836=>"000111110",
  57837=>"000000001",
  57838=>"001011111",
  57839=>"111111111",
  57840=>"110111111",
  57841=>"000101111",
  57842=>"000001111",
  57843=>"100000000",
  57844=>"110000000",
  57845=>"111111111",
  57846=>"111111100",
  57847=>"011001111",
  57848=>"000100111",
  57849=>"001111111",
  57850=>"000110111",
  57851=>"111000000",
  57852=>"011011111",
  57853=>"101000000",
  57854=>"111011000",
  57855=>"000000000",
  57856=>"111111100",
  57857=>"110111111",
  57858=>"000000111",
  57859=>"100000000",
  57860=>"000000110",
  57861=>"010011111",
  57862=>"111111111",
  57863=>"111111111",
  57864=>"001000101",
  57865=>"111011010",
  57866=>"111010110",
  57867=>"000000000",
  57868=>"011010010",
  57869=>"111110111",
  57870=>"100111111",
  57871=>"101001001",
  57872=>"001000000",
  57873=>"111111100",
  57874=>"111111111",
  57875=>"010110000",
  57876=>"000110110",
  57877=>"111111000",
  57878=>"000000000",
  57879=>"000000000",
  57880=>"111111000",
  57881=>"011111111",
  57882=>"000000110",
  57883=>"110011000",
  57884=>"100110111",
  57885=>"011111011",
  57886=>"000000000",
  57887=>"111011000",
  57888=>"111111111",
  57889=>"111001000",
  57890=>"111111110",
  57891=>"011000000",
  57892=>"111111111",
  57893=>"111111011",
  57894=>"000001011",
  57895=>"000001001",
  57896=>"111111111",
  57897=>"010010000",
  57898=>"000000001",
  57899=>"111111111",
  57900=>"000001111",
  57901=>"111111111",
  57902=>"001001111",
  57903=>"111111111",
  57904=>"000000000",
  57905=>"000110010",
  57906=>"100000011",
  57907=>"111111000",
  57908=>"110000010",
  57909=>"111011111",
  57910=>"101000000",
  57911=>"111111100",
  57912=>"000000000",
  57913=>"000010000",
  57914=>"001111011",
  57915=>"100000000",
  57916=>"101000000",
  57917=>"100000000",
  57918=>"111111111",
  57919=>"111111111",
  57920=>"010111010",
  57921=>"000000110",
  57922=>"110100111",
  57923=>"111111111",
  57924=>"111001000",
  57925=>"111001001",
  57926=>"000000000",
  57927=>"000000011",
  57928=>"110001000",
  57929=>"111111111",
  57930=>"111111111",
  57931=>"000000000",
  57932=>"100000111",
  57933=>"000000000",
  57934=>"001110111",
  57935=>"111011001",
  57936=>"111111011",
  57937=>"111111111",
  57938=>"000000000",
  57939=>"000000011",
  57940=>"000000000",
  57941=>"000000100",
  57942=>"000000111",
  57943=>"111101111",
  57944=>"111111000",
  57945=>"111111111",
  57946=>"000000100",
  57947=>"011000110",
  57948=>"000111111",
  57949=>"100000000",
  57950=>"000101111",
  57951=>"111111011",
  57952=>"000000111",
  57953=>"010100110",
  57954=>"000000111",
  57955=>"000000000",
  57956=>"110110111",
  57957=>"000000000",
  57958=>"110111111",
  57959=>"000000000",
  57960=>"111111111",
  57961=>"111000000",
  57962=>"000111111",
  57963=>"000000000",
  57964=>"110111000",
  57965=>"000001011",
  57966=>"111101111",
  57967=>"111111111",
  57968=>"101000100",
  57969=>"000000010",
  57970=>"010010111",
  57971=>"010000000",
  57972=>"111111111",
  57973=>"111111111",
  57974=>"000000000",
  57975=>"110111001",
  57976=>"100100000",
  57977=>"010000000",
  57978=>"000011000",
  57979=>"111111111",
  57980=>"000000111",
  57981=>"001001111",
  57982=>"000000000",
  57983=>"111111001",
  57984=>"000000000",
  57985=>"001001000",
  57986=>"000000110",
  57987=>"111111000",
  57988=>"111111111",
  57989=>"011000111",
  57990=>"100100111",
  57991=>"000000000",
  57992=>"011010010",
  57993=>"000000000",
  57994=>"000000000",
  57995=>"111111000",
  57996=>"000000000",
  57997=>"111000100",
  57998=>"000000000",
  57999=>"111111110",
  58000=>"111000000",
  58001=>"010111000",
  58002=>"000010000",
  58003=>"111101111",
  58004=>"110000111",
  58005=>"000100110",
  58006=>"011111111",
  58007=>"011001001",
  58008=>"000000000",
  58009=>"111011001",
  58010=>"111010100",
  58011=>"000000111",
  58012=>"111111111",
  58013=>"111111111",
  58014=>"000000011",
  58015=>"111111111",
  58016=>"111111111",
  58017=>"000000000",
  58018=>"001000111",
  58019=>"011111111",
  58020=>"000000100",
  58021=>"111111111",
  58022=>"100111001",
  58023=>"100000111",
  58024=>"111111111",
  58025=>"100111111",
  58026=>"101000000",
  58027=>"111111000",
  58028=>"000111000",
  58029=>"011000111",
  58030=>"000000101",
  58031=>"000000000",
  58032=>"000001100",
  58033=>"111111111",
  58034=>"000111000",
  58035=>"111111001",
  58036=>"110100101",
  58037=>"000011000",
  58038=>"001011111",
  58039=>"000000000",
  58040=>"111110010",
  58041=>"010111111",
  58042=>"000000000",
  58043=>"000000000",
  58044=>"000000000",
  58045=>"011011000",
  58046=>"110101000",
  58047=>"000111111",
  58048=>"001001011",
  58049=>"000000000",
  58050=>"011111010",
  58051=>"000000111",
  58052=>"011111101",
  58053=>"111111111",
  58054=>"000100110",
  58055=>"000000000",
  58056=>"001011000",
  58057=>"111111111",
  58058=>"000000000",
  58059=>"111111000",
  58060=>"110000000",
  58061=>"111111111",
  58062=>"111111011",
  58063=>"101101000",
  58064=>"000001111",
  58065=>"011011011",
  58066=>"000000111",
  58067=>"001001011",
  58068=>"000000100",
  58069=>"100000011",
  58070=>"111000000",
  58071=>"110101000",
  58072=>"111110111",
  58073=>"111110100",
  58074=>"111111111",
  58075=>"000000111",
  58076=>"111111111",
  58077=>"100100110",
  58078=>"111100000",
  58079=>"111111111",
  58080=>"110110111",
  58081=>"000000000",
  58082=>"100111111",
  58083=>"111111111",
  58084=>"101101111",
  58085=>"100000000",
  58086=>"111011111",
  58087=>"111111110",
  58088=>"111111000",
  58089=>"111111110",
  58090=>"111111111",
  58091=>"110110111",
  58092=>"111100000",
  58093=>"100000111",
  58094=>"000000111",
  58095=>"111111100",
  58096=>"111010000",
  58097=>"000011111",
  58098=>"000111111",
  58099=>"010000100",
  58100=>"110110111",
  58101=>"111101000",
  58102=>"000000000",
  58103=>"111000000",
  58104=>"111111111",
  58105=>"000010010",
  58106=>"000000000",
  58107=>"000101110",
  58108=>"000000000",
  58109=>"000010000",
  58110=>"000000000",
  58111=>"111111111",
  58112=>"111111000",
  58113=>"000000000",
  58114=>"111111111",
  58115=>"111111111",
  58116=>"111111111",
  58117=>"110000000",
  58118=>"000111111",
  58119=>"000111111",
  58120=>"000000000",
  58121=>"100100000",
  58122=>"111111111",
  58123=>"100111111",
  58124=>"000000000",
  58125=>"111111111",
  58126=>"000000101",
  58127=>"000000000",
  58128=>"000000000",
  58129=>"000000110",
  58130=>"000000111",
  58131=>"000111111",
  58132=>"000100111",
  58133=>"111111111",
  58134=>"001101111",
  58135=>"111111111",
  58136=>"000000100",
  58137=>"000000100",
  58138=>"000000101",
  58139=>"001001001",
  58140=>"111111000",
  58141=>"110111010",
  58142=>"111111010",
  58143=>"000000100",
  58144=>"000000000",
  58145=>"111111010",
  58146=>"011111111",
  58147=>"000000000",
  58148=>"111111111",
  58149=>"111111110",
  58150=>"100000110",
  58151=>"010110000",
  58152=>"111111111",
  58153=>"111101001",
  58154=>"000000000",
  58155=>"111011111",
  58156=>"001000001",
  58157=>"000100100",
  58158=>"001000000",
  58159=>"000000100",
  58160=>"010001001",
  58161=>"111100000",
  58162=>"100100000",
  58163=>"000000100",
  58164=>"111000000",
  58165=>"100111111",
  58166=>"110011100",
  58167=>"000000000",
  58168=>"011010111",
  58169=>"111011111",
  58170=>"000000000",
  58171=>"001000000",
  58172=>"111111111",
  58173=>"000000111",
  58174=>"110111111",
  58175=>"100100000",
  58176=>"011011111",
  58177=>"000000110",
  58178=>"000110100",
  58179=>"100000111",
  58180=>"000000000",
  58181=>"111110010",
  58182=>"111000000",
  58183=>"000000111",
  58184=>"100000111",
  58185=>"110000000",
  58186=>"011000000",
  58187=>"000001100",
  58188=>"000100111",
  58189=>"111110000",
  58190=>"000000000",
  58191=>"000111111",
  58192=>"001111111",
  58193=>"110100110",
  58194=>"000111111",
  58195=>"110110110",
  58196=>"000000000",
  58197=>"110000011",
  58198=>"001001111",
  58199=>"000100101",
  58200=>"000011111",
  58201=>"111001000",
  58202=>"000000101",
  58203=>"000001001",
  58204=>"000000000",
  58205=>"110010111",
  58206=>"010111111",
  58207=>"000000000",
  58208=>"011011101",
  58209=>"000001001",
  58210=>"011011011",
  58211=>"111000111",
  58212=>"011111111",
  58213=>"000000000",
  58214=>"100000010",
  58215=>"001000000",
  58216=>"000100000",
  58217=>"000000010",
  58218=>"000000000",
  58219=>"100110110",
  58220=>"001000000",
  58221=>"011001000",
  58222=>"111111111",
  58223=>"000000000",
  58224=>"000000110",
  58225=>"100100110",
  58226=>"110111111",
  58227=>"000000100",
  58228=>"100100110",
  58229=>"110111110",
  58230=>"111011001",
  58231=>"111111000",
  58232=>"000000111",
  58233=>"111001000",
  58234=>"111111111",
  58235=>"111110111",
  58236=>"000000000",
  58237=>"111110000",
  58238=>"111110110",
  58239=>"111111111",
  58240=>"011011000",
  58241=>"111010000",
  58242=>"111110110",
  58243=>"000000100",
  58244=>"111111111",
  58245=>"111111111",
  58246=>"111110110",
  58247=>"111111111",
  58248=>"000000111",
  58249=>"111110000",
  58250=>"000000000",
  58251=>"010111111",
  58252=>"011000000",
  58253=>"000010000",
  58254=>"111111000",
  58255=>"000000110",
  58256=>"000000000",
  58257=>"001111111",
  58258=>"010000100",
  58259=>"111111100",
  58260=>"111011000",
  58261=>"000000001",
  58262=>"000000110",
  58263=>"011011111",
  58264=>"000000001",
  58265=>"111111000",
  58266=>"000101111",
  58267=>"010110111",
  58268=>"111111111",
  58269=>"000011111",
  58270=>"101100000",
  58271=>"100000110",
  58272=>"000000111",
  58273=>"011011011",
  58274=>"110111110",
  58275=>"000000000",
  58276=>"100110110",
  58277=>"000000111",
  58278=>"111100000",
  58279=>"111111101",
  58280=>"000000000",
  58281=>"010010110",
  58282=>"000000000",
  58283=>"000000000",
  58284=>"000000000",
  58285=>"111111111",
  58286=>"110010000",
  58287=>"000000000",
  58288=>"000000000",
  58289=>"111111001",
  58290=>"000111111",
  58291=>"111110000",
  58292=>"000000000",
  58293=>"000000000",
  58294=>"000000001",
  58295=>"011000000",
  58296=>"000001001",
  58297=>"000000010",
  58298=>"111111011",
  58299=>"001000101",
  58300=>"011001111",
  58301=>"111001011",
  58302=>"000000000",
  58303=>"000000000",
  58304=>"111111101",
  58305=>"100101111",
  58306=>"111111111",
  58307=>"110000000",
  58308=>"000000000",
  58309=>"100110111",
  58310=>"110111000",
  58311=>"000000000",
  58312=>"000000010",
  58313=>"111111000",
  58314=>"111010000",
  58315=>"111111111",
  58316=>"110111010",
  58317=>"111011010",
  58318=>"111111100",
  58319=>"000111111",
  58320=>"111111111",
  58321=>"000000111",
  58322=>"111110000",
  58323=>"111111111",
  58324=>"001001000",
  58325=>"110000000",
  58326=>"111000001",
  58327=>"110010000",
  58328=>"000000001",
  58329=>"111111100",
  58330=>"010011000",
  58331=>"000000000",
  58332=>"111000000",
  58333=>"011010000",
  58334=>"111110000",
  58335=>"000101111",
  58336=>"000000000",
  58337=>"111111111",
  58338=>"110101111",
  58339=>"000000100",
  58340=>"111000000",
  58341=>"101001000",
  58342=>"010000000",
  58343=>"000000101",
  58344=>"000000000",
  58345=>"111111000",
  58346=>"000000100",
  58347=>"000100111",
  58348=>"100000010",
  58349=>"110011111",
  58350=>"000000111",
  58351=>"110110000",
  58352=>"000000110",
  58353=>"000000111",
  58354=>"100001011",
  58355=>"011011010",
  58356=>"000000000",
  58357=>"000000011",
  58358=>"000000000",
  58359=>"111110000",
  58360=>"000000000",
  58361=>"000000110",
  58362=>"101100100",
  58363=>"000000000",
  58364=>"100101111",
  58365=>"111111001",
  58366=>"000001001",
  58367=>"000000110",
  58368=>"111111101",
  58369=>"000000001",
  58370=>"111101111",
  58371=>"000011000",
  58372=>"000000000",
  58373=>"101000001",
  58374=>"111111011",
  58375=>"111111111",
  58376=>"011111111",
  58377=>"101010010",
  58378=>"000011111",
  58379=>"111111110",
  58380=>"110110110",
  58381=>"111000100",
  58382=>"010011001",
  58383=>"111110100",
  58384=>"011001111",
  58385=>"011111111",
  58386=>"111111111",
  58387=>"001001111",
  58388=>"000000000",
  58389=>"111000111",
  58390=>"100110100",
  58391=>"000101111",
  58392=>"110000000",
  58393=>"011011010",
  58394=>"111000001",
  58395=>"001011011",
  58396=>"000000111",
  58397=>"111111111",
  58398=>"000010111",
  58399=>"000100110",
  58400=>"000001001",
  58401=>"111101111",
  58402=>"111000000",
  58403=>"101001001",
  58404=>"000000000",
  58405=>"000000000",
  58406=>"111000000",
  58407=>"000110111",
  58408=>"111111000",
  58409=>"101000000",
  58410=>"011001000",
  58411=>"101000001",
  58412=>"101000101",
  58413=>"000111100",
  58414=>"011010111",
  58415=>"010000000",
  58416=>"111000100",
  58417=>"111010000",
  58418=>"000000111",
  58419=>"000000000",
  58420=>"000110111",
  58421=>"000000000",
  58422=>"000000000",
  58423=>"000010011",
  58424=>"111111000",
  58425=>"000000001",
  58426=>"100000000",
  58427=>"001111111",
  58428=>"000000000",
  58429=>"111111011",
  58430=>"100110000",
  58431=>"000011111",
  58432=>"111100000",
  58433=>"111000001",
  58434=>"101000110",
  58435=>"110000101",
  58436=>"100000111",
  58437=>"000000000",
  58438=>"111000001",
  58439=>"111111111",
  58440=>"001111100",
  58441=>"000000000",
  58442=>"000000000",
  58443=>"101101101",
  58444=>"011111111",
  58445=>"001011111",
  58446=>"000111111",
  58447=>"111111000",
  58448=>"111111110",
  58449=>"101111011",
  58450=>"000000000",
  58451=>"010111110",
  58452=>"000000000",
  58453=>"000000000",
  58454=>"001101111",
  58455=>"000000000",
  58456=>"000010000",
  58457=>"000000000",
  58458=>"000000000",
  58459=>"011011001",
  58460=>"000000000",
  58461=>"000000111",
  58462=>"001000000",
  58463=>"100110100",
  58464=>"000000000",
  58465=>"000001111",
  58466=>"100000000",
  58467=>"011000000",
  58468=>"000000000",
  58469=>"001001001",
  58470=>"111111000",
  58471=>"001011111",
  58472=>"000000111",
  58473=>"110111011",
  58474=>"111001000",
  58475=>"011111111",
  58476=>"111111100",
  58477=>"111111001",
  58478=>"000000000",
  58479=>"000000000",
  58480=>"000111111",
  58481=>"100100001",
  58482=>"111111110",
  58483=>"001000001",
  58484=>"000000000",
  58485=>"011111110",
  58486=>"000000000",
  58487=>"000000000",
  58488=>"000001100",
  58489=>"111111111",
  58490=>"111111000",
  58491=>"000000000",
  58492=>"000111111",
  58493=>"011111110",
  58494=>"000010011",
  58495=>"000000100",
  58496=>"100111110",
  58497=>"110001001",
  58498=>"100000000",
  58499=>"110000000",
  58500=>"111111100",
  58501=>"001101111",
  58502=>"100100111",
  58503=>"110110111",
  58504=>"111101111",
  58505=>"000000001",
  58506=>"000000000",
  58507=>"111111000",
  58508=>"111110111",
  58509=>"010000000",
  58510=>"111111111",
  58511=>"111111111",
  58512=>"000111111",
  58513=>"100111110",
  58514=>"111011000",
  58515=>"011001001",
  58516=>"001111000",
  58517=>"100000011",
  58518=>"000000111",
  58519=>"111100101",
  58520=>"011111111",
  58521=>"111111111",
  58522=>"010000100",
  58523=>"000000111",
  58524=>"111000000",
  58525=>"000000101",
  58526=>"000001111",
  58527=>"111001111",
  58528=>"000000100",
  58529=>"000000000",
  58530=>"000000011",
  58531=>"111111111",
  58532=>"011000000",
  58533=>"111111010",
  58534=>"000111111",
  58535=>"000000000",
  58536=>"001000000",
  58537=>"000000001",
  58538=>"000000000",
  58539=>"111111010",
  58540=>"011011000",
  58541=>"001011010",
  58542=>"111111111",
  58543=>"001010000",
  58544=>"000000110",
  58545=>"111011001",
  58546=>"110111111",
  58547=>"000000100",
  58548=>"001001000",
  58549=>"000000000",
  58550=>"010111010",
  58551=>"111111111",
  58552=>"111110100",
  58553=>"111111111",
  58554=>"000000000",
  58555=>"111111111",
  58556=>"001001111",
  58557=>"110110110",
  58558=>"111111111",
  58559=>"000000110",
  58560=>"111111011",
  58561=>"111111110",
  58562=>"111111111",
  58563=>"000000101",
  58564=>"000000000",
  58565=>"100000000",
  58566=>"000000000",
  58567=>"000001000",
  58568=>"011111111",
  58569=>"001000000",
  58570=>"000010000",
  58571=>"000111111",
  58572=>"100100001",
  58573=>"111111111",
  58574=>"000010110",
  58575=>"000000001",
  58576=>"111101001",
  58577=>"011100000",
  58578=>"000000001",
  58579=>"111000000",
  58580=>"000011110",
  58581=>"100101111",
  58582=>"000100101",
  58583=>"011000000",
  58584=>"000000000",
  58585=>"011111001",
  58586=>"000000001",
  58587=>"000111111",
  58588=>"011111111",
  58589=>"000001111",
  58590=>"110110110",
  58591=>"000000000",
  58592=>"111011000",
  58593=>"011011000",
  58594=>"000000100",
  58595=>"011000100",
  58596=>"111011000",
  58597=>"111100000",
  58598=>"101111111",
  58599=>"000000101",
  58600=>"111011000",
  58601=>"001001111",
  58602=>"110110000",
  58603=>"100000000",
  58604=>"011111010",
  58605=>"000111110",
  58606=>"000000111",
  58607=>"001000111",
  58608=>"000000000",
  58609=>"110010110",
  58610=>"111111111",
  58611=>"111111010",
  58612=>"001001101",
  58613=>"111111111",
  58614=>"111000100",
  58615=>"100000000",
  58616=>"111000101",
  58617=>"111111111",
  58618=>"110111111",
  58619=>"111111111",
  58620=>"001000000",
  58621=>"000000110",
  58622=>"111111100",
  58623=>"111111111",
  58624=>"111111000",
  58625=>"000000111",
  58626=>"111111111",
  58627=>"111111111",
  58628=>"100000000",
  58629=>"001000000",
  58630=>"111000000",
  58631=>"000001111",
  58632=>"000000000",
  58633=>"000000001",
  58634=>"000000000",
  58635=>"011011000",
  58636=>"000000111",
  58637=>"111111111",
  58638=>"111111111",
  58639=>"000000010",
  58640=>"100111111",
  58641=>"000000000",
  58642=>"000000000",
  58643=>"000000000",
  58644=>"000000000",
  58645=>"000000111",
  58646=>"011000011",
  58647=>"111111111",
  58648=>"011011111",
  58649=>"011000001",
  58650=>"000000001",
  58651=>"000101111",
  58652=>"000111100",
  58653=>"011111111",
  58654=>"000000000",
  58655=>"111110111",
  58656=>"101100000",
  58657=>"000111111",
  58658=>"110011000",
  58659=>"111101001",
  58660=>"111001000",
  58661=>"111110010",
  58662=>"100111111",
  58663=>"001001001",
  58664=>"000000111",
  58665=>"010111111",
  58666=>"111111110",
  58667=>"111111000",
  58668=>"111110111",
  58669=>"000111111",
  58670=>"000000000",
  58671=>"001111100",
  58672=>"000000000",
  58673=>"111111111",
  58674=>"000000111",
  58675=>"111001000",
  58676=>"001001000",
  58677=>"000000001",
  58678=>"000000000",
  58679=>"111000000",
  58680=>"000000000",
  58681=>"111000100",
  58682=>"001111111",
  58683=>"000000001",
  58684=>"000000000",
  58685=>"111111111",
  58686=>"000000000",
  58687=>"111000111",
  58688=>"111101000",
  58689=>"000001000",
  58690=>"110000000",
  58691=>"000000000",
  58692=>"110000111",
  58693=>"000000001",
  58694=>"000000000",
  58695=>"111111111",
  58696=>"000000111",
  58697=>"000000000",
  58698=>"000000101",
  58699=>"101100000",
  58700=>"001001000",
  58701=>"000000011",
  58702=>"000000111",
  58703=>"000000111",
  58704=>"110000110",
  58705=>"001001111",
  58706=>"000101000",
  58707=>"001001011",
  58708=>"000000000",
  58709=>"111110011",
  58710=>"000110111",
  58711=>"000000111",
  58712=>"100000000",
  58713=>"100101111",
  58714=>"111111111",
  58715=>"000000100",
  58716=>"001000000",
  58717=>"000000000",
  58718=>"101001001",
  58719=>"000100111",
  58720=>"001000000",
  58721=>"001001111",
  58722=>"111110110",
  58723=>"000000000",
  58724=>"110110111",
  58725=>"000001001",
  58726=>"100100100",
  58727=>"001111111",
  58728=>"000110101",
  58729=>"111111111",
  58730=>"101101001",
  58731=>"101001000",
  58732=>"110000000",
  58733=>"111111111",
  58734=>"111000000",
  58735=>"000000000",
  58736=>"000000000",
  58737=>"000000110",
  58738=>"000000111",
  58739=>"111011011",
  58740=>"001001111",
  58741=>"001101101",
  58742=>"000000000",
  58743=>"110010110",
  58744=>"000000100",
  58745=>"111111110",
  58746=>"000000000",
  58747=>"101100001",
  58748=>"010111111",
  58749=>"111111010",
  58750=>"101101001",
  58751=>"111000000",
  58752=>"100101111",
  58753=>"001000111",
  58754=>"000000000",
  58755=>"000000000",
  58756=>"111101001",
  58757=>"111111001",
  58758=>"101001111",
  58759=>"111001000",
  58760=>"001001001",
  58761=>"001111111",
  58762=>"111101011",
  58763=>"111101001",
  58764=>"001001001",
  58765=>"000100000",
  58766=>"110110110",
  58767=>"000001001",
  58768=>"000000000",
  58769=>"000000000",
  58770=>"000000111",
  58771=>"100000000",
  58772=>"000000000",
  58773=>"000010000",
  58774=>"111111100",
  58775=>"010011111",
  58776=>"111101100",
  58777=>"001001001",
  58778=>"000000101",
  58779=>"111111110",
  58780=>"111111000",
  58781=>"100101000",
  58782=>"000111000",
  58783=>"111111001",
  58784=>"111101000",
  58785=>"110000111",
  58786=>"000000000",
  58787=>"000000000",
  58788=>"111111100",
  58789=>"111001111",
  58790=>"111001101",
  58791=>"100100000",
  58792=>"111000000",
  58793=>"111111011",
  58794=>"111111110",
  58795=>"000100110",
  58796=>"111111111",
  58797=>"000000111",
  58798=>"000001111",
  58799=>"001111111",
  58800=>"000000111",
  58801=>"011000000",
  58802=>"000001000",
  58803=>"111001001",
  58804=>"110111111",
  58805=>"111000000",
  58806=>"000111111",
  58807=>"111000000",
  58808=>"011001000",
  58809=>"111111011",
  58810=>"001000001",
  58811=>"011111111",
  58812=>"111000001",
  58813=>"111100100",
  58814=>"000111111",
  58815=>"111110100",
  58816=>"010010000",
  58817=>"111100000",
  58818=>"001000000",
  58819=>"000000111",
  58820=>"101100111",
  58821=>"000000111",
  58822=>"000000000",
  58823=>"111111111",
  58824=>"000000111",
  58825=>"101111111",
  58826=>"000000000",
  58827=>"000000110",
  58828=>"111111110",
  58829=>"000010110",
  58830=>"111111001",
  58831=>"111111101",
  58832=>"000111111",
  58833=>"000010110",
  58834=>"101000000",
  58835=>"111101111",
  58836=>"111110110",
  58837=>"111100100",
  58838=>"000000110",
  58839=>"111111110",
  58840=>"111010000",
  58841=>"001001000",
  58842=>"000111111",
  58843=>"011110111",
  58844=>"011111111",
  58845=>"010011000",
  58846=>"001001111",
  58847=>"000000111",
  58848=>"000000001",
  58849=>"001000111",
  58850=>"011000001",
  58851=>"000000000",
  58852=>"001011111",
  58853=>"101001100",
  58854=>"111111110",
  58855=>"000000000",
  58856=>"111111111",
  58857=>"111111111",
  58858=>"001000000",
  58859=>"000010111",
  58860=>"000110111",
  58861=>"110110110",
  58862=>"000010111",
  58863=>"000000000",
  58864=>"000111110",
  58865=>"000000000",
  58866=>"101000000",
  58867=>"000110000",
  58868=>"111111111",
  58869=>"111100100",
  58870=>"111111111",
  58871=>"111000000",
  58872=>"000000100",
  58873=>"011001001",
  58874=>"001000001",
  58875=>"111000100",
  58876=>"001001011",
  58877=>"111000000",
  58878=>"001001011",
  58879=>"000010011",
  58880=>"000011111",
  58881=>"010110111",
  58882=>"111001111",
  58883=>"010010111",
  58884=>"111111111",
  58885=>"111000000",
  58886=>"111111111",
  58887=>"000010010",
  58888=>"101111111",
  58889=>"111110000",
  58890=>"000000000",
  58891=>"111111010",
  58892=>"000110110",
  58893=>"000010011",
  58894=>"000000000",
  58895=>"000000000",
  58896=>"111111111",
  58897=>"111110000",
  58898=>"111111111",
  58899=>"001000111",
  58900=>"110111111",
  58901=>"111000111",
  58902=>"000000000",
  58903=>"111101110",
  58904=>"111111110",
  58905=>"000000000",
  58906=>"100101000",
  58907=>"110000000",
  58908=>"000000000",
  58909=>"001011111",
  58910=>"100100100",
  58911=>"111111111",
  58912=>"001111111",
  58913=>"100000000",
  58914=>"101111000",
  58915=>"000000000",
  58916=>"000000000",
  58917=>"000000000",
  58918=>"110111010",
  58919=>"111111000",
  58920=>"000000000",
  58921=>"000000000",
  58922=>"111101000",
  58923=>"101111111",
  58924=>"100100111",
  58925=>"000000000",
  58926=>"000000000",
  58927=>"001100000",
  58928=>"110111111",
  58929=>"111111010",
  58930=>"000000000",
  58931=>"111111110",
  58932=>"001111110",
  58933=>"001000010",
  58934=>"101111111",
  58935=>"000000000",
  58936=>"111111111",
  58937=>"000000100",
  58938=>"111111111",
  58939=>"000000000",
  58940=>"000000001",
  58941=>"101100111",
  58942=>"000011011",
  58943=>"000000000",
  58944=>"000000000",
  58945=>"000110000",
  58946=>"111111111",
  58947=>"111111000",
  58948=>"000100110",
  58949=>"000000000",
  58950=>"000000110",
  58951=>"011000000",
  58952=>"011011111",
  58953=>"011111111",
  58954=>"000000000",
  58955=>"000000100",
  58956=>"000001111",
  58957=>"111111111",
  58958=>"111111000",
  58959=>"000000000",
  58960=>"000000000",
  58961=>"000000000",
  58962=>"111111111",
  58963=>"111111000",
  58964=>"000000000",
  58965=>"111111111",
  58966=>"111000000",
  58967=>"000000000",
  58968=>"111001000",
  58969=>"100000100",
  58970=>"111111111",
  58971=>"111111111",
  58972=>"000011000",
  58973=>"000001001",
  58974=>"010000000",
  58975=>"111110111",
  58976=>"111111111",
  58977=>"111111111",
  58978=>"100000111",
  58979=>"111111111",
  58980=>"000000000",
  58981=>"111111111",
  58982=>"011011010",
  58983=>"111101101",
  58984=>"111111111",
  58985=>"001000000",
  58986=>"000000000",
  58987=>"000111111",
  58988=>"111000000",
  58989=>"000000000",
  58990=>"011011111",
  58991=>"100000000",
  58992=>"110000111",
  58993=>"111111111",
  58994=>"000000000",
  58995=>"000000000",
  58996=>"000000000",
  58997=>"000000000",
  58998=>"110110100",
  58999=>"111111000",
  59000=>"000001111",
  59001=>"000000111",
  59002=>"111111010",
  59003=>"000000000",
  59004=>"110110010",
  59005=>"000010000",
  59006=>"111111110",
  59007=>"000000000",
  59008=>"111001000",
  59009=>"000010010",
  59010=>"111110111",
  59011=>"111111001",
  59012=>"111111101",
  59013=>"001000111",
  59014=>"101111111",
  59015=>"111111000",
  59016=>"111111111",
  59017=>"000000010",
  59018=>"011111000",
  59019=>"110000000",
  59020=>"100000101",
  59021=>"000000000",
  59022=>"111111110",
  59023=>"111011000",
  59024=>"000000111",
  59025=>"000100100",
  59026=>"000000000",
  59027=>"111111111",
  59028=>"111111000",
  59029=>"001001011",
  59030=>"001000000",
  59031=>"000000000",
  59032=>"100000000",
  59033=>"001011111",
  59034=>"000000000",
  59035=>"111111111",
  59036=>"111111111",
  59037=>"111111111",
  59038=>"111111111",
  59039=>"000000000",
  59040=>"000000111",
  59041=>"011111111",
  59042=>"110000111",
  59043=>"111111111",
  59044=>"000000000",
  59045=>"001001101",
  59046=>"111111000",
  59047=>"000011111",
  59048=>"100011110",
  59049=>"111111111",
  59050=>"000000000",
  59051=>"000000100",
  59052=>"000000000",
  59053=>"100110100",
  59054=>"000000100",
  59055=>"111100001",
  59056=>"000001111",
  59057=>"111110010",
  59058=>"111111010",
  59059=>"000111111",
  59060=>"111111110",
  59061=>"111111111",
  59062=>"001000000",
  59063=>"001111111",
  59064=>"100100111",
  59065=>"000110111",
  59066=>"000000000",
  59067=>"111000000",
  59068=>"111111111",
  59069=>"000000000",
  59070=>"100111111",
  59071=>"110111111",
  59072=>"111011000",
  59073=>"000000000",
  59074=>"001000011",
  59075=>"100111001",
  59076=>"111111101",
  59077=>"000000000",
  59078=>"000000000",
  59079=>"000000000",
  59080=>"000000000",
  59081=>"000001000",
  59082=>"000000010",
  59083=>"111111111",
  59084=>"111111111",
  59085=>"001000000",
  59086=>"111110111",
  59087=>"110011000",
  59088=>"111100110",
  59089=>"000000000",
  59090=>"000000000",
  59091=>"000000100",
  59092=>"000001011",
  59093=>"011011111",
  59094=>"100101000",
  59095=>"010000000",
  59096=>"000000000",
  59097=>"001001101",
  59098=>"111011001",
  59099=>"000001001",
  59100=>"011111111",
  59101=>"011111111",
  59102=>"111111100",
  59103=>"101101111",
  59104=>"111111111",
  59105=>"111111000",
  59106=>"100000011",
  59107=>"000000111",
  59108=>"011000000",
  59109=>"111110111",
  59110=>"010011111",
  59111=>"111111111",
  59112=>"000000111",
  59113=>"000110111",
  59114=>"100111111",
  59115=>"000000000",
  59116=>"000000011",
  59117=>"111010001",
  59118=>"111111111",
  59119=>"111000000",
  59120=>"000110111",
  59121=>"000000101",
  59122=>"111111111",
  59123=>"001111111",
  59124=>"111111010",
  59125=>"011011111",
  59126=>"111111111",
  59127=>"000000000",
  59128=>"111111000",
  59129=>"111111111",
  59130=>"000000000",
  59131=>"000100000",
  59132=>"110010000",
  59133=>"111010111",
  59134=>"110010010",
  59135=>"000000000",
  59136=>"000000000",
  59137=>"010000000",
  59138=>"011111110",
  59139=>"000000100",
  59140=>"111111111",
  59141=>"011111111",
  59142=>"000000111",
  59143=>"111111011",
  59144=>"110011000",
  59145=>"000000000",
  59146=>"111111000",
  59147=>"000000000",
  59148=>"111101111",
  59149=>"000000011",
  59150=>"111111111",
  59151=>"111111000",
  59152=>"110111011",
  59153=>"000111111",
  59154=>"000000111",
  59155=>"111000100",
  59156=>"111111111",
  59157=>"111111111",
  59158=>"000111000",
  59159=>"111111111",
  59160=>"010000000",
  59161=>"000000000",
  59162=>"111111000",
  59163=>"111111111",
  59164=>"000000000",
  59165=>"111011000",
  59166=>"000111111",
  59167=>"111000000",
  59168=>"000000011",
  59169=>"111111111",
  59170=>"111000000",
  59171=>"111111111",
  59172=>"100000000",
  59173=>"000001010",
  59174=>"101110010",
  59175=>"000000000",
  59176=>"011001000",
  59177=>"000000000",
  59178=>"100000000",
  59179=>"000000000",
  59180=>"111110110",
  59181=>"110000000",
  59182=>"111111111",
  59183=>"111111111",
  59184=>"000000000",
  59185=>"111011010",
  59186=>"000100110",
  59187=>"111101110",
  59188=>"111111000",
  59189=>"000000100",
  59190=>"000001111",
  59191=>"000111000",
  59192=>"111111111",
  59193=>"111111100",
  59194=>"111001011",
  59195=>"000000000",
  59196=>"100000000",
  59197=>"000000111",
  59198=>"000001011",
  59199=>"000000000",
  59200=>"111101100",
  59201=>"111011010",
  59202=>"111111111",
  59203=>"000010111",
  59204=>"010110000",
  59205=>"000000000",
  59206=>"000111111",
  59207=>"111111111",
  59208=>"011001000",
  59209=>"111111111",
  59210=>"111111111",
  59211=>"111111011",
  59212=>"111001000",
  59213=>"000000000",
  59214=>"000000000",
  59215=>"111010100",
  59216=>"011001100",
  59217=>"101000101",
  59218=>"000000000",
  59219=>"111111111",
  59220=>"000000000",
  59221=>"011011001",
  59222=>"111110111",
  59223=>"010011011",
  59224=>"111111111",
  59225=>"000001011",
  59226=>"111111001",
  59227=>"000000000",
  59228=>"000110111",
  59229=>"000000000",
  59230=>"000100000",
  59231=>"111111110",
  59232=>"111111110",
  59233=>"000000000",
  59234=>"001000000",
  59235=>"111111111",
  59236=>"000011010",
  59237=>"111000111",
  59238=>"011001111",
  59239=>"111111000",
  59240=>"111111111",
  59241=>"000000000",
  59242=>"111111000",
  59243=>"100100111",
  59244=>"000000000",
  59245=>"110110100",
  59246=>"000000000",
  59247=>"111111000",
  59248=>"111001100",
  59249=>"111111111",
  59250=>"000010111",
  59251=>"011111111",
  59252=>"111111111",
  59253=>"111101111",
  59254=>"111110110",
  59255=>"011010000",
  59256=>"011001101",
  59257=>"111111111",
  59258=>"110110111",
  59259=>"000000000",
  59260=>"111011000",
  59261=>"111111111",
  59262=>"101011011",
  59263=>"001101101",
  59264=>"111111111",
  59265=>"100100000",
  59266=>"000000000",
  59267=>"001000000",
  59268=>"111111111",
  59269=>"000000100",
  59270=>"111111111",
  59271=>"111001111",
  59272=>"100000000",
  59273=>"110100011",
  59274=>"111111101",
  59275=>"000111111",
  59276=>"000000111",
  59277=>"101111111",
  59278=>"111110000",
  59279=>"110101000",
  59280=>"000000000",
  59281=>"111111111",
  59282=>"010000000",
  59283=>"000000000",
  59284=>"000000000",
  59285=>"010010000",
  59286=>"000110111",
  59287=>"001001010",
  59288=>"001101111",
  59289=>"110111111",
  59290=>"111111111",
  59291=>"111111100",
  59292=>"111111111",
  59293=>"111111111",
  59294=>"000000000",
  59295=>"111010010",
  59296=>"000000000",
  59297=>"111001011",
  59298=>"111111111",
  59299=>"000000000",
  59300=>"100010010",
  59301=>"000000101",
  59302=>"111111111",
  59303=>"111111111",
  59304=>"111111111",
  59305=>"000000000",
  59306=>"111011010",
  59307=>"000000011",
  59308=>"000000000",
  59309=>"011111110",
  59310=>"000000000",
  59311=>"010011111",
  59312=>"000000011",
  59313=>"001011000",
  59314=>"001111111",
  59315=>"111111111",
  59316=>"110000001",
  59317=>"000000000",
  59318=>"111111110",
  59319=>"011111000",
  59320=>"111001111",
  59321=>"001011011",
  59322=>"111001111",
  59323=>"000000000",
  59324=>"000000000",
  59325=>"000000001",
  59326=>"011110110",
  59327=>"110111110",
  59328=>"111111000",
  59329=>"111111111",
  59330=>"111111111",
  59331=>"000000011",
  59332=>"011010000",
  59333=>"000000110",
  59334=>"000011111",
  59335=>"000000100",
  59336=>"010110100",
  59337=>"000000000",
  59338=>"001001111",
  59339=>"000000011",
  59340=>"001000000",
  59341=>"111111111",
  59342=>"100000000",
  59343=>"111111111",
  59344=>"000000000",
  59345=>"001001001",
  59346=>"111111111",
  59347=>"111111011",
  59348=>"111111110",
  59349=>"110110111",
  59350=>"000010110",
  59351=>"000011001",
  59352=>"001000000",
  59353=>"000011000",
  59354=>"001001001",
  59355=>"110110011",
  59356=>"000000000",
  59357=>"111011001",
  59358=>"111111111",
  59359=>"000000001",
  59360=>"000000000",
  59361=>"000010000",
  59362=>"111111111",
  59363=>"111110111",
  59364=>"111111111",
  59365=>"000000000",
  59366=>"100100110",
  59367=>"000000000",
  59368=>"000000000",
  59369=>"111111111",
  59370=>"100000011",
  59371=>"001111111",
  59372=>"000111111",
  59373=>"010000000",
  59374=>"000000111",
  59375=>"000000000",
  59376=>"000000000",
  59377=>"111111111",
  59378=>"111111111",
  59379=>"110111011",
  59380=>"111111010",
  59381=>"000000100",
  59382=>"011011000",
  59383=>"100100111",
  59384=>"000000000",
  59385=>"111111011",
  59386=>"111111111",
  59387=>"111101111",
  59388=>"111111111",
  59389=>"100000111",
  59390=>"110110000",
  59391=>"011000000",
  59392=>"000000000",
  59393=>"111111111",
  59394=>"000000100",
  59395=>"110110111",
  59396=>"000111111",
  59397=>"111111000",
  59398=>"100000000",
  59399=>"111111111",
  59400=>"111111111",
  59401=>"000000000",
  59402=>"011111100",
  59403=>"001000000",
  59404=>"001110110",
  59405=>"101111111",
  59406=>"100100111",
  59407=>"000000010",
  59408=>"111000000",
  59409=>"110110110",
  59410=>"011000010",
  59411=>"110110010",
  59412=>"111111111",
  59413=>"111111011",
  59414=>"010110000",
  59415=>"111111111",
  59416=>"111111111",
  59417=>"000001001",
  59418=>"111111110",
  59419=>"100100000",
  59420=>"100000111",
  59421=>"001001001",
  59422=>"100100100",
  59423=>"110110110",
  59424=>"110110000",
  59425=>"000100000",
  59426=>"111011011",
  59427=>"101111111",
  59428=>"000000000",
  59429=>"111000000",
  59430=>"000001111",
  59431=>"000000110",
  59432=>"111111111",
  59433=>"011011000",
  59434=>"100100101",
  59435=>"010010000",
  59436=>"000000000",
  59437=>"111111111",
  59438=>"001001000",
  59439=>"011001000",
  59440=>"000000000",
  59441=>"000000000",
  59442=>"000100100",
  59443=>"111111111",
  59444=>"111010011",
  59445=>"001001011",
  59446=>"000000000",
  59447=>"101101111",
  59448=>"111011111",
  59449=>"110000000",
  59450=>"111111111",
  59451=>"111111111",
  59452=>"000000000",
  59453=>"000100010",
  59454=>"111111000",
  59455=>"000000000",
  59456=>"111000011",
  59457=>"110111101",
  59458=>"100000000",
  59459=>"111111011",
  59460=>"100110110",
  59461=>"000100000",
  59462=>"111111111",
  59463=>"000000000",
  59464=>"011011010",
  59465=>"111111111",
  59466=>"000000000",
  59467=>"001100000",
  59468=>"111111111",
  59469=>"110010000",
  59470=>"111111100",
  59471=>"101101000",
  59472=>"000000000",
  59473=>"000000000",
  59474=>"111111111",
  59475=>"011111111",
  59476=>"111111101",
  59477=>"100100100",
  59478=>"011011001",
  59479=>"110000000",
  59480=>"011111111",
  59481=>"001111001",
  59482=>"111111111",
  59483=>"111111111",
  59484=>"101000000",
  59485=>"000000000",
  59486=>"110111111",
  59487=>"011011000",
  59488=>"000000000",
  59489=>"001000000",
  59490=>"000000000",
  59491=>"000000000",
  59492=>"000010000",
  59493=>"111100100",
  59494=>"000000000",
  59495=>"000111001",
  59496=>"000000000",
  59497=>"111111111",
  59498=>"000001011",
  59499=>"000000000",
  59500=>"000001011",
  59501=>"000000000",
  59502=>"111101011",
  59503=>"111110010",
  59504=>"000000101",
  59505=>"000000001",
  59506=>"001000000",
  59507=>"110110000",
  59508=>"111111111",
  59509=>"000001011",
  59510=>"000000000",
  59511=>"000000001",
  59512=>"001000000",
  59513=>"101100000",
  59514=>"100100111",
  59515=>"111111100",
  59516=>"000000000",
  59517=>"111011111",
  59518=>"110111101",
  59519=>"111100000",
  59520=>"010111111",
  59521=>"000000010",
  59522=>"000000000",
  59523=>"000100111",
  59524=>"000000011",
  59525=>"000000000",
  59526=>"111111111",
  59527=>"000001000",
  59528=>"000110111",
  59529=>"000000000",
  59530=>"111111111",
  59531=>"000000000",
  59532=>"100111111",
  59533=>"111111100",
  59534=>"111111111",
  59535=>"111111100",
  59536=>"000000000",
  59537=>"101111011",
  59538=>"010111111",
  59539=>"000100100",
  59540=>"100110111",
  59541=>"010011000",
  59542=>"000011111",
  59543=>"111111000",
  59544=>"111111011",
  59545=>"111110000",
  59546=>"000000011",
  59547=>"000000001",
  59548=>"011001011",
  59549=>"000110000",
  59550=>"011111111",
  59551=>"011010110",
  59552=>"100000000",
  59553=>"000000000",
  59554=>"111111111",
  59555=>"000000000",
  59556=>"101100111",
  59557=>"111011100",
  59558=>"111000000",
  59559=>"111000001",
  59560=>"000001111",
  59561=>"000000000",
  59562=>"010000000",
  59563=>"000000000",
  59564=>"100110000",
  59565=>"000010111",
  59566=>"000000000",
  59567=>"000000000",
  59568=>"000000000",
  59569=>"100100000",
  59570=>"111111111",
  59571=>"110100101",
  59572=>"110110110",
  59573=>"000000000",
  59574=>"000000001",
  59575=>"000000001",
  59576=>"010111110",
  59577=>"000000000",
  59578=>"111110111",
  59579=>"111111111",
  59580=>"000000000",
  59581=>"111111000",
  59582=>"000000000",
  59583=>"000000000",
  59584=>"111011011",
  59585=>"000111000",
  59586=>"000000000",
  59587=>"111111100",
  59588=>"100100000",
  59589=>"000000000",
  59590=>"011000001",
  59591=>"111111011",
  59592=>"011111111",
  59593=>"111111111",
  59594=>"000110110",
  59595=>"010011111",
  59596=>"000011111",
  59597=>"100110111",
  59598=>"110111111",
  59599=>"110110100",
  59600=>"000100100",
  59601=>"000000010",
  59602=>"111111110",
  59603=>"000000000",
  59604=>"101101111",
  59605=>"111111111",
  59606=>"000011011",
  59607=>"101111111",
  59608=>"111111001",
  59609=>"101111001",
  59610=>"000000000",
  59611=>"111000111",
  59612=>"111111011",
  59613=>"111111111",
  59614=>"000010000",
  59615=>"111111110",
  59616=>"011001101",
  59617=>"011111111",
  59618=>"000000000",
  59619=>"111111111",
  59620=>"000001001",
  59621=>"110000000",
  59622=>"011111111",
  59623=>"111111111",
  59624=>"111111110",
  59625=>"001111111",
  59626=>"000000111",
  59627=>"111111111",
  59628=>"010001001",
  59629=>"011000001",
  59630=>"100111111",
  59631=>"111000000",
  59632=>"001011011",
  59633=>"100000000",
  59634=>"000000000",
  59635=>"001000011",
  59636=>"111111111",
  59637=>"111001001",
  59638=>"010000000",
  59639=>"011000000",
  59640=>"000000000",
  59641=>"111111111",
  59642=>"101101111",
  59643=>"111111111",
  59644=>"111111111",
  59645=>"100110110",
  59646=>"101100111",
  59647=>"011000000",
  59648=>"000000100",
  59649=>"000011011",
  59650=>"101110100",
  59651=>"111110111",
  59652=>"000100110",
  59653=>"000000011",
  59654=>"110000000",
  59655=>"011011000",
  59656=>"000000000",
  59657=>"100100111",
  59658=>"111111111",
  59659=>"000000000",
  59660=>"110110110",
  59661=>"001001001",
  59662=>"111111111",
  59663=>"000000011",
  59664=>"111111000",
  59665=>"000000010",
  59666=>"000000000",
  59667=>"000001111",
  59668=>"111111010",
  59669=>"111000000",
  59670=>"000010011",
  59671=>"111111111",
  59672=>"000000011",
  59673=>"111111111",
  59674=>"000000000",
  59675=>"000000000",
  59676=>"000000001",
  59677=>"100111000",
  59678=>"010010000",
  59679=>"111111000",
  59680=>"111101111",
  59681=>"000100110",
  59682=>"111011011",
  59683=>"000111111",
  59684=>"111110010",
  59685=>"001111011",
  59686=>"111111111",
  59687=>"111101000",
  59688=>"010010111",
  59689=>"101000000",
  59690=>"001000011",
  59691=>"011001000",
  59692=>"001001001",
  59693=>"111111111",
  59694=>"000000000",
  59695=>"110110111",
  59696=>"000000000",
  59697=>"100100101",
  59698=>"111101000",
  59699=>"000011011",
  59700=>"000000101",
  59701=>"111101000",
  59702=>"000000000",
  59703=>"101011000",
  59704=>"100000000",
  59705=>"111111111",
  59706=>"000010010",
  59707=>"011011001",
  59708=>"001001000",
  59709=>"111100001",
  59710=>"000110100",
  59711=>"110100100",
  59712=>"000000001",
  59713=>"000000000",
  59714=>"000111111",
  59715=>"000000000",
  59716=>"100111111",
  59717=>"001000000",
  59718=>"001001000",
  59719=>"111101111",
  59720=>"111111000",
  59721=>"000000000",
  59722=>"111111000",
  59723=>"000000011",
  59724=>"011111000",
  59725=>"110010000",
  59726=>"100100100",
  59727=>"000000110",
  59728=>"111111111",
  59729=>"110110110",
  59730=>"100111111",
  59731=>"000000110",
  59732=>"101100111",
  59733=>"011001011",
  59734=>"110111111",
  59735=>"100100110",
  59736=>"111111111",
  59737=>"111111111",
  59738=>"000111111",
  59739=>"100000110",
  59740=>"010000100",
  59741=>"011001111",
  59742=>"111011011",
  59743=>"111111110",
  59744=>"000000000",
  59745=>"000000011",
  59746=>"000000000",
  59747=>"111100000",
  59748=>"000000001",
  59749=>"000000100",
  59750=>"011000000",
  59751=>"111111111",
  59752=>"111100111",
  59753=>"000000000",
  59754=>"001001000",
  59755=>"111111111",
  59756=>"001001000",
  59757=>"111000000",
  59758=>"100111111",
  59759=>"000011111",
  59760=>"111111100",
  59761=>"111111001",
  59762=>"111000111",
  59763=>"111111111",
  59764=>"111111111",
  59765=>"001011000",
  59766=>"000010000",
  59767=>"111111110",
  59768=>"000001011",
  59769=>"000111111",
  59770=>"111111111",
  59771=>"111111111",
  59772=>"110100000",
  59773=>"000000010",
  59774=>"000100000",
  59775=>"000000000",
  59776=>"000000000",
  59777=>"000000000",
  59778=>"000000001",
  59779=>"000000000",
  59780=>"000000000",
  59781=>"001000000",
  59782=>"111100000",
  59783=>"111111000",
  59784=>"111101001",
  59785=>"110110001",
  59786=>"111111100",
  59787=>"000001001",
  59788=>"000000000",
  59789=>"000000000",
  59790=>"000100110",
  59791=>"001000000",
  59792=>"000000000",
  59793=>"111111111",
  59794=>"000000001",
  59795=>"111111111",
  59796=>"111110000",
  59797=>"000001000",
  59798=>"000000000",
  59799=>"001001001",
  59800=>"111111111",
  59801=>"100100100",
  59802=>"111111111",
  59803=>"001011111",
  59804=>"011001001",
  59805=>"111100100",
  59806=>"011000000",
  59807=>"000010011",
  59808=>"100110000",
  59809=>"011111000",
  59810=>"011000111",
  59811=>"000110111",
  59812=>"001000000",
  59813=>"010111111",
  59814=>"111111111",
  59815=>"011111111",
  59816=>"000010100",
  59817=>"111011111",
  59818=>"111010010",
  59819=>"111101111",
  59820=>"000000000",
  59821=>"111111011",
  59822=>"111110111",
  59823=>"111011000",
  59824=>"111000000",
  59825=>"110000100",
  59826=>"110110111",
  59827=>"000000000",
  59828=>"000001001",
  59829=>"111111000",
  59830=>"110110000",
  59831=>"000000000",
  59832=>"101111111",
  59833=>"111000100",
  59834=>"110100000",
  59835=>"000000000",
  59836=>"111111110",
  59837=>"111111100",
  59838=>"111111000",
  59839=>"001001001",
  59840=>"111111111",
  59841=>"000000101",
  59842=>"000000000",
  59843=>"000000000",
  59844=>"001111010",
  59845=>"000000000",
  59846=>"001111111",
  59847=>"000000001",
  59848=>"100101111",
  59849=>"111111010",
  59850=>"100000000",
  59851=>"001001111",
  59852=>"111111111",
  59853=>"000000000",
  59854=>"000000000",
  59855=>"000010000",
  59856=>"010000110",
  59857=>"000011011",
  59858=>"100100111",
  59859=>"000000000",
  59860=>"001000000",
  59861=>"110111110",
  59862=>"111111111",
  59863=>"000000001",
  59864=>"000000100",
  59865=>"111111011",
  59866=>"011111110",
  59867=>"100111111",
  59868=>"000011000",
  59869=>"000000000",
  59870=>"000110111",
  59871=>"010000000",
  59872=>"000000000",
  59873=>"111111111",
  59874=>"111101101",
  59875=>"000000000",
  59876=>"111000111",
  59877=>"110110110",
  59878=>"000000011",
  59879=>"000000000",
  59880=>"000100100",
  59881=>"000000000",
  59882=>"111011001",
  59883=>"111100000",
  59884=>"111111111",
  59885=>"111111111",
  59886=>"001101111",
  59887=>"111111110",
  59888=>"111111111",
  59889=>"111111001",
  59890=>"111111111",
  59891=>"000000000",
  59892=>"100101111",
  59893=>"000000000",
  59894=>"000000000",
  59895=>"100100100",
  59896=>"000000000",
  59897=>"000000000",
  59898=>"000001000",
  59899=>"000011111",
  59900=>"000001000",
  59901=>"111111010",
  59902=>"001000100",
  59903=>"111111111",
  59904=>"000000000",
  59905=>"011111011",
  59906=>"000000000",
  59907=>"000000110",
  59908=>"000000000",
  59909=>"111111011",
  59910=>"111101000",
  59911=>"011011111",
  59912=>"111001111",
  59913=>"000000101",
  59914=>"111111011",
  59915=>"000000000",
  59916=>"110110110",
  59917=>"111110110",
  59918=>"111011000",
  59919=>"000000000",
  59920=>"111100111",
  59921=>"100111111",
  59922=>"000000000",
  59923=>"100000101",
  59924=>"000000000",
  59925=>"111111100",
  59926=>"111111111",
  59927=>"100111111",
  59928=>"110111111",
  59929=>"001011011",
  59930=>"111100000",
  59931=>"000001000",
  59932=>"111111011",
  59933=>"000000000",
  59934=>"011111111",
  59935=>"000000000",
  59936=>"100000011",
  59937=>"111111110",
  59938=>"110011000",
  59939=>"110111111",
  59940=>"001111000",
  59941=>"110011110",
  59942=>"000010000",
  59943=>"000000110",
  59944=>"111111000",
  59945=>"000111111",
  59946=>"111111100",
  59947=>"111101011",
  59948=>"111111111",
  59949=>"111111000",
  59950=>"001000001",
  59951=>"111001001",
  59952=>"111111111",
  59953=>"000001111",
  59954=>"111111001",
  59955=>"011000010",
  59956=>"110000100",
  59957=>"011001001",
  59958=>"000000000",
  59959=>"000001001",
  59960=>"011111111",
  59961=>"011001001",
  59962=>"000000000",
  59963=>"000000101",
  59964=>"000000111",
  59965=>"111111011",
  59966=>"110100000",
  59967=>"000111011",
  59968=>"000000011",
  59969=>"000000000",
  59970=>"111111111",
  59971=>"000111111",
  59972=>"000100111",
  59973=>"111111111",
  59974=>"111110000",
  59975=>"111111111",
  59976=>"100000000",
  59977=>"000000000",
  59978=>"000001000",
  59979=>"111111111",
  59980=>"000111111",
  59981=>"110110111",
  59982=>"000110110",
  59983=>"011011010",
  59984=>"010010001",
  59985=>"100000000",
  59986=>"000110110",
  59987=>"110111111",
  59988=>"000000000",
  59989=>"001000000",
  59990=>"000011000",
  59991=>"000000000",
  59992=>"010100100",
  59993=>"000111111",
  59994=>"111111100",
  59995=>"000000000",
  59996=>"000000110",
  59997=>"000001011",
  59998=>"000000000",
  59999=>"111010010",
  60000=>"111000000",
  60001=>"000000101",
  60002=>"011010000",
  60003=>"111111111",
  60004=>"001111111",
  60005=>"011001111",
  60006=>"110011000",
  60007=>"110000000",
  60008=>"000000111",
  60009=>"111111000",
  60010=>"001111111",
  60011=>"110100100",
  60012=>"000011100",
  60013=>"001001000",
  60014=>"000111111",
  60015=>"000000111",
  60016=>"111000000",
  60017=>"000000001",
  60018=>"010010000",
  60019=>"011011111",
  60020=>"000011000",
  60021=>"111111000",
  60022=>"111111111",
  60023=>"001011111",
  60024=>"011001000",
  60025=>"011111000",
  60026=>"111101101",
  60027=>"000000000",
  60028=>"000111111",
  60029=>"111111000",
  60030=>"000001111",
  60031=>"111011010",
  60032=>"101000000",
  60033=>"010000000",
  60034=>"000000001",
  60035=>"111000000",
  60036=>"111000000",
  60037=>"000000000",
  60038=>"001111111",
  60039=>"000111111",
  60040=>"111111100",
  60041=>"000000000",
  60042=>"111111111",
  60043=>"000000010",
  60044=>"000011101",
  60045=>"000000000",
  60046=>"000111111",
  60047=>"000000111",
  60048=>"111111111",
  60049=>"000000000",
  60050=>"111111000",
  60051=>"111111111",
  60052=>"000110111",
  60053=>"110110000",
  60054=>"111111111",
  60055=>"101111111",
  60056=>"111001101",
  60057=>"000000000",
  60058=>"111000000",
  60059=>"010010110",
  60060=>"000000000",
  60061=>"000000111",
  60062=>"000000000",
  60063=>"000000101",
  60064=>"000000111",
  60065=>"000110111",
  60066=>"111111000",
  60067=>"011001000",
  60068=>"001010110",
  60069=>"111111011",
  60070=>"111011000",
  60071=>"001001111",
  60072=>"000000111",
  60073=>"111001001",
  60074=>"000000000",
  60075=>"111111111",
  60076=>"001010000",
  60077=>"000001001",
  60078=>"010110000",
  60079=>"000000000",
  60080=>"111111111",
  60081=>"000110110",
  60082=>"111011011",
  60083=>"000000111",
  60084=>"100100100",
  60085=>"111011000",
  60086=>"110111111",
  60087=>"111111111",
  60088=>"111110000",
  60089=>"001101111",
  60090=>"100000111",
  60091=>"111111111",
  60092=>"001000000",
  60093=>"011111111",
  60094=>"111000000",
  60095=>"000000111",
  60096=>"010000010",
  60097=>"111111110",
  60098=>"111111111",
  60099=>"111000000",
  60100=>"000000000",
  60101=>"000100100",
  60102=>"000110000",
  60103=>"000000000",
  60104=>"000111111",
  60105=>"000010000",
  60106=>"011111001",
  60107=>"100100111",
  60108=>"001000000",
  60109=>"000001111",
  60110=>"000000110",
  60111=>"000000010",
  60112=>"111111000",
  60113=>"000110100",
  60114=>"000000000",
  60115=>"111111111",
  60116=>"000111101",
  60117=>"010100111",
  60118=>"111111100",
  60119=>"000001001",
  60120=>"111111000",
  60121=>"011000000",
  60122=>"000000000",
  60123=>"111111111",
  60124=>"011011001",
  60125=>"111111111",
  60126=>"111111111",
  60127=>"000100000",
  60128=>"100100100",
  60129=>"111000000",
  60130=>"000000110",
  60131=>"000000000",
  60132=>"000100111",
  60133=>"000111000",
  60134=>"101001101",
  60135=>"010000000",
  60136=>"001000001",
  60137=>"111001111",
  60138=>"110110000",
  60139=>"101101111",
  60140=>"000100111",
  60141=>"000001000",
  60142=>"100000100",
  60143=>"000110011",
  60144=>"111111001",
  60145=>"101101100",
  60146=>"011111100",
  60147=>"000010110",
  60148=>"001100100",
  60149=>"111110000",
  60150=>"011011011",
  60151=>"111101000",
  60152=>"111101111",
  60153=>"000000000",
  60154=>"000110000",
  60155=>"000101111",
  60156=>"011111111",
  60157=>"000000000",
  60158=>"111111011",
  60159=>"000000000",
  60160=>"111111000",
  60161=>"111111110",
  60162=>"111111111",
  60163=>"000111111",
  60164=>"000101111",
  60165=>"000000000",
  60166=>"111100000",
  60167=>"010000101",
  60168=>"011111111",
  60169=>"000000111",
  60170=>"001001001",
  60171=>"011010000",
  60172=>"000000100",
  60173=>"000000001",
  60174=>"111111111",
  60175=>"000000000",
  60176=>"110100000",
  60177=>"110010000",
  60178=>"000111000",
  60179=>"000011111",
  60180=>"010000000",
  60181=>"000111111",
  60182=>"011011011",
  60183=>"011000000",
  60184=>"011111111",
  60185=>"111110111",
  60186=>"111111110",
  60187=>"000000010",
  60188=>"001001001",
  60189=>"000000000",
  60190=>"110000000",
  60191=>"111010000",
  60192=>"000001111",
  60193=>"010010100",
  60194=>"111111100",
  60195=>"011010000",
  60196=>"110111011",
  60197=>"111111111",
  60198=>"101111111",
  60199=>"000000000",
  60200=>"000111111",
  60201=>"010000000",
  60202=>"001011101",
  60203=>"111111101",
  60204=>"111110010",
  60205=>"100100111",
  60206=>"001111000",
  60207=>"000000000",
  60208=>"110111111",
  60209=>"000000000",
  60210=>"000000000",
  60211=>"001100101",
  60212=>"000000111",
  60213=>"000001000",
  60214=>"000100100",
  60215=>"111011111",
  60216=>"000000000",
  60217=>"000000000",
  60218=>"110110000",
  60219=>"000000100",
  60220=>"000111111",
  60221=>"000000000",
  60222=>"000000011",
  60223=>"110111000",
  60224=>"101111101",
  60225=>"111111111",
  60226=>"000000000",
  60227=>"111111000",
  60228=>"000000000",
  60229=>"000101111",
  60230=>"000000000",
  60231=>"111111001",
  60232=>"111011001",
  60233=>"000000000",
  60234=>"111111100",
  60235=>"000111001",
  60236=>"000000000",
  60237=>"011011011",
  60238=>"000000000",
  60239=>"001001001",
  60240=>"110100100",
  60241=>"000110111",
  60242=>"001111111",
  60243=>"111000000",
  60244=>"100000000",
  60245=>"011001101",
  60246=>"111000000",
  60247=>"000011011",
  60248=>"000000010",
  60249=>"111111111",
  60250=>"111111111",
  60251=>"001111111",
  60252=>"110110110",
  60253=>"010010011",
  60254=>"110100000",
  60255=>"110100000",
  60256=>"000000101",
  60257=>"111110000",
  60258=>"111111111",
  60259=>"000111111",
  60260=>"000000000",
  60261=>"000000000",
  60262=>"110000000",
  60263=>"111111000",
  60264=>"001001111",
  60265=>"000111111",
  60266=>"111111010",
  60267=>"000111011",
  60268=>"000110110",
  60269=>"111111111",
  60270=>"111111111",
  60271=>"000001111",
  60272=>"000001001",
  60273=>"000001000",
  60274=>"111000000",
  60275=>"110111111",
  60276=>"000111101",
  60277=>"111011000",
  60278=>"100110111",
  60279=>"000000000",
  60280=>"000000000",
  60281=>"000110111",
  60282=>"110111111",
  60283=>"000000011",
  60284=>"000111111",
  60285=>"000000000",
  60286=>"000110100",
  60287=>"101111000",
  60288=>"100000010",
  60289=>"110011010",
  60290=>"111011110",
  60291=>"000000000",
  60292=>"000000111",
  60293=>"101100111",
  60294=>"111110111",
  60295=>"110111111",
  60296=>"000000000",
  60297=>"100000001",
  60298=>"101000000",
  60299=>"111111111",
  60300=>"001000011",
  60301=>"001000111",
  60302=>"011011000",
  60303=>"110100101",
  60304=>"000000000",
  60305=>"000011000",
  60306=>"011011111",
  60307=>"011111111",
  60308=>"000000000",
  60309=>"010110111",
  60310=>"111111100",
  60311=>"000000000",
  60312=>"000000111",
  60313=>"111111111",
  60314=>"000000000",
  60315=>"000000000",
  60316=>"111000000",
  60317=>"000000000",
  60318=>"111111111",
  60319=>"101101000",
  60320=>"000001000",
  60321=>"110110011",
  60322=>"000001111",
  60323=>"000000110",
  60324=>"011111010",
  60325=>"001000000",
  60326=>"011001000",
  60327=>"111110000",
  60328=>"000000100",
  60329=>"111001000",
  60330=>"111111111",
  60331=>"101100000",
  60332=>"111111010",
  60333=>"000111111",
  60334=>"111001011",
  60335=>"110111011",
  60336=>"000100111",
  60337=>"111111111",
  60338=>"101110110",
  60339=>"000000000",
  60340=>"000000011",
  60341=>"111111000",
  60342=>"100000011",
  60343=>"111111000",
  60344=>"000000111",
  60345=>"110111111",
  60346=>"000011001",
  60347=>"111111001",
  60348=>"000000110",
  60349=>"010100110",
  60350=>"000100100",
  60351=>"101001100",
  60352=>"011010010",
  60353=>"111111010",
  60354=>"010111111",
  60355=>"000001001",
  60356=>"000000000",
  60357=>"001001001",
  60358=>"111111101",
  60359=>"101101101",
  60360=>"101000000",
  60361=>"001011111",
  60362=>"000110111",
  60363=>"000000000",
  60364=>"000000000",
  60365=>"011011000",
  60366=>"000000000",
  60367=>"111111100",
  60368=>"011111111",
  60369=>"101111100",
  60370=>"000001000",
  60371=>"101101001",
  60372=>"000000000",
  60373=>"000000000",
  60374=>"000000000",
  60375=>"111011001",
  60376=>"000010000",
  60377=>"000000000",
  60378=>"000000000",
  60379=>"000000000",
  60380=>"000000010",
  60381=>"011000111",
  60382=>"000011111",
  60383=>"100000010",
  60384=>"111111111",
  60385=>"000111111",
  60386=>"000000000",
  60387=>"000000000",
  60388=>"111111111",
  60389=>"100100000",
  60390=>"000000000",
  60391=>"100110111",
  60392=>"111111011",
  60393=>"111111111",
  60394=>"111110101",
  60395=>"000011111",
  60396=>"111010000",
  60397=>"000000100",
  60398=>"110110010",
  60399=>"111110110",
  60400=>"110111111",
  60401=>"111110100",
  60402=>"000001000",
  60403=>"010000100",
  60404=>"000110111",
  60405=>"000000000",
  60406=>"111111111",
  60407=>"111011111",
  60408=>"001001111",
  60409=>"100111000",
  60410=>"111111000",
  60411=>"111111000",
  60412=>"001011001",
  60413=>"010000011",
  60414=>"000000000",
  60415=>"000001101",
  60416=>"000000000",
  60417=>"111111111",
  60418=>"010000111",
  60419=>"111011011",
  60420=>"000000101",
  60421=>"011110100",
  60422=>"011111111",
  60423=>"000000000",
  60424=>"111111111",
  60425=>"000000001",
  60426=>"111111000",
  60427=>"111101000",
  60428=>"011001011",
  60429=>"111111111",
  60430=>"001011111",
  60431=>"111111111",
  60432=>"000000100",
  60433=>"101111111",
  60434=>"000001111",
  60435=>"010111111",
  60436=>"000000111",
  60437=>"111111111",
  60438=>"100111110",
  60439=>"111110100",
  60440=>"000000000",
  60441=>"000100101",
  60442=>"111111111",
  60443=>"101111111",
  60444=>"111111111",
  60445=>"111111111",
  60446=>"000000101",
  60447=>"000000000",
  60448=>"110111111",
  60449=>"111111111",
  60450=>"001011111",
  60451=>"000000000",
  60452=>"000000000",
  60453=>"100100111",
  60454=>"000110000",
  60455=>"111111111",
  60456=>"001001111",
  60457=>"111111111",
  60458=>"111111100",
  60459=>"111111111",
  60460=>"000000111",
  60461=>"000000000",
  60462=>"111110111",
  60463=>"000011000",
  60464=>"110100110",
  60465=>"000000101",
  60466=>"000001001",
  60467=>"000000000",
  60468=>"111111110",
  60469=>"010000111",
  60470=>"001000000",
  60471=>"000000000",
  60472=>"111111111",
  60473=>"000000100",
  60474=>"111111111",
  60475=>"111111000",
  60476=>"111101100",
  60477=>"001001000",
  60478=>"000000001",
  60479=>"000000000",
  60480=>"001001111",
  60481=>"110111100",
  60482=>"011111001",
  60483=>"000000000",
  60484=>"011001001",
  60485=>"011011111",
  60486=>"011000000",
  60487=>"000000000",
  60488=>"110111111",
  60489=>"111111111",
  60490=>"111110000",
  60491=>"111111111",
  60492=>"111111110",
  60493=>"100111111",
  60494=>"000000000",
  60495=>"001101001",
  60496=>"100000111",
  60497=>"000111110",
  60498=>"000000000",
  60499=>"001001101",
  60500=>"000000000",
  60501=>"101001111",
  60502=>"111111111",
  60503=>"100111111",
  60504=>"111111111",
  60505=>"000000000",
  60506=>"111000010",
  60507=>"000000101",
  60508=>"111011011",
  60509=>"010111111",
  60510=>"000000000",
  60511=>"011010000",
  60512=>"000000000",
  60513=>"000010110",
  60514=>"111111111",
  60515=>"000100000",
  60516=>"110111111",
  60517=>"101101000",
  60518=>"000111111",
  60519=>"111111111",
  60520=>"111111110",
  60521=>"010000000",
  60522=>"110000000",
  60523=>"111111111",
  60524=>"000000000",
  60525=>"100101111",
  60526=>"100111111",
  60527=>"000000101",
  60528=>"000100111",
  60529=>"000010111",
  60530=>"000010011",
  60531=>"000000111",
  60532=>"010000000",
  60533=>"000111100",
  60534=>"111001001",
  60535=>"000000000",
  60536=>"000110111",
  60537=>"111100100",
  60538=>"000000000",
  60539=>"000000111",
  60540=>"000110110",
  60541=>"001000000",
  60542=>"000000000",
  60543=>"000000000",
  60544=>"001000100",
  60545=>"101011000",
  60546=>"000000000",
  60547=>"000011011",
  60548=>"000011001",
  60549=>"000000111",
  60550=>"000000000",
  60551=>"000111111",
  60552=>"111111111",
  60553=>"111001000",
  60554=>"111001011",
  60555=>"000000000",
  60556=>"111011000",
  60557=>"111111111",
  60558=>"111111000",
  60559=>"000001001",
  60560=>"111111111",
  60561=>"000000000",
  60562=>"000000000",
  60563=>"001001011",
  60564=>"000100100",
  60565=>"000000001",
  60566=>"111111111",
  60567=>"111110111",
  60568=>"100011001",
  60569=>"111000000",
  60570=>"111111111",
  60571=>"011001111",
  60572=>"111001000",
  60573=>"011010101",
  60574=>"000000000",
  60575=>"000001000",
  60576=>"111000100",
  60577=>"000000000",
  60578=>"111111111",
  60579=>"011111011",
  60580=>"111111111",
  60581=>"000111111",
  60582=>"100000000",
  60583=>"000000000",
  60584=>"110000000",
  60585=>"000000000",
  60586=>"111101111",
  60587=>"000000010",
  60588=>"111111111",
  60589=>"000000000",
  60590=>"000000111",
  60591=>"100111111",
  60592=>"111111000",
  60593=>"000000000",
  60594=>"011111000",
  60595=>"101000000",
  60596=>"111111000",
  60597=>"000000010",
  60598=>"011101111",
  60599=>"111111111",
  60600=>"111100110",
  60601=>"111111111",
  60602=>"001001011",
  60603=>"111001001",
  60604=>"000000000",
  60605=>"111111111",
  60606=>"110110110",
  60607=>"110111011",
  60608=>"100000100",
  60609=>"111111111",
  60610=>"000000000",
  60611=>"111111111",
  60612=>"111111111",
  60613=>"000000000",
  60614=>"110110111",
  60615=>"111111111",
  60616=>"000000000",
  60617=>"000000111",
  60618=>"000000000",
  60619=>"000000001",
  60620=>"000011011",
  60621=>"111111111",
  60622=>"100000001",
  60623=>"000000000",
  60624=>"001000000",
  60625=>"111111111",
  60626=>"001001111",
  60627=>"111111111",
  60628=>"101111111",
  60629=>"110000101",
  60630=>"001001000",
  60631=>"111111111",
  60632=>"000110000",
  60633=>"000000000",
  60634=>"111111111",
  60635=>"111111111",
  60636=>"111111111",
  60637=>"100000000",
  60638=>"000000001",
  60639=>"000000000",
  60640=>"000000000",
  60641=>"000011010",
  60642=>"000000000",
  60643=>"111111111",
  60644=>"000000000",
  60645=>"111101100",
  60646=>"111111110",
  60647=>"000000000",
  60648=>"011111111",
  60649=>"000000000",
  60650=>"111111111",
  60651=>"110100111",
  60652=>"000000000",
  60653=>"000000100",
  60654=>"000001000",
  60655=>"111111000",
  60656=>"110110110",
  60657=>"010000000",
  60658=>"111001001",
  60659=>"001000000",
  60660=>"000111011",
  60661=>"111000000",
  60662=>"000000000",
  60663=>"111011010",
  60664=>"111111111",
  60665=>"111111111",
  60666=>"000000000",
  60667=>"000000000",
  60668=>"001001111",
  60669=>"000001001",
  60670=>"000000000",
  60671=>"111111111",
  60672=>"001000001",
  60673=>"001111101",
  60674=>"000000000",
  60675=>"000000111",
  60676=>"111100000",
  60677=>"100100011",
  60678=>"100100111",
  60679=>"000000111",
  60680=>"111111111",
  60681=>"111111011",
  60682=>"011011001",
  60683=>"000000000",
  60684=>"110111010",
  60685=>"111101111",
  60686=>"000000101",
  60687=>"011111110",
  60688=>"000000000",
  60689=>"111000001",
  60690=>"111111111",
  60691=>"001111110",
  60692=>"111111110",
  60693=>"001001001",
  60694=>"011111001",
  60695=>"000100100",
  60696=>"000100100",
  60697=>"111111111",
  60698=>"111111111",
  60699=>"111000000",
  60700=>"111011011",
  60701=>"111011111",
  60702=>"111000000",
  60703=>"000000101",
  60704=>"000000000",
  60705=>"111111111",
  60706=>"111011000",
  60707=>"111111111",
  60708=>"000001001",
  60709=>"111111011",
  60710=>"110110111",
  60711=>"001111111",
  60712=>"010010111",
  60713=>"000000000",
  60714=>"001000000",
  60715=>"000000000",
  60716=>"000000000",
  60717=>"000111000",
  60718=>"111001000",
  60719=>"000000000",
  60720=>"000000000",
  60721=>"100111100",
  60722=>"111000000",
  60723=>"000000000",
  60724=>"000000000",
  60725=>"000000000",
  60726=>"110100100",
  60727=>"111101001",
  60728=>"000000000",
  60729=>"110111111",
  60730=>"000000000",
  60731=>"111111111",
  60732=>"011011101",
  60733=>"111111111",
  60734=>"001111111",
  60735=>"100101000",
  60736=>"001111111",
  60737=>"000000001",
  60738=>"000000001",
  60739=>"100100000",
  60740=>"111100000",
  60741=>"000000110",
  60742=>"000000000",
  60743=>"100110111",
  60744=>"000000000",
  60745=>"000000000",
  60746=>"000000000",
  60747=>"000000100",
  60748=>"000000000",
  60749=>"111111111",
  60750=>"111001000",
  60751=>"110110111",
  60752=>"100101011",
  60753=>"011000000",
  60754=>"000000000",
  60755=>"111111111",
  60756=>"110111111",
  60757=>"011011011",
  60758=>"000001000",
  60759=>"000000111",
  60760=>"000000001",
  60761=>"000000000",
  60762=>"000101101",
  60763=>"111111111",
  60764=>"111111111",
  60765=>"111111111",
  60766=>"110100000",
  60767=>"011011000",
  60768=>"000000000",
  60769=>"000000000",
  60770=>"001011110",
  60771=>"010111111",
  60772=>"011011111",
  60773=>"000001001",
  60774=>"110100100",
  60775=>"000000000",
  60776=>"001001000",
  60777=>"000111111",
  60778=>"011110000",
  60779=>"011011111",
  60780=>"100100110",
  60781=>"001000000",
  60782=>"111000000",
  60783=>"000000000",
  60784=>"111011011",
  60785=>"001000111",
  60786=>"000000011",
  60787=>"111011111",
  60788=>"000010000",
  60789=>"000000000",
  60790=>"010010110",
  60791=>"000101111",
  60792=>"000000000",
  60793=>"111111111",
  60794=>"100000000",
  60795=>"111111011",
  60796=>"000000000",
  60797=>"111111111",
  60798=>"000101111",
  60799=>"111111111",
  60800=>"011011011",
  60801=>"111000110",
  60802=>"100100101",
  60803=>"111111111",
  60804=>"110000000",
  60805=>"000011111",
  60806=>"111110100",
  60807=>"000000000",
  60808=>"111111111",
  60809=>"011011010",
  60810=>"000000000",
  60811=>"111111111",
  60812=>"001001111",
  60813=>"111011111",
  60814=>"001001000",
  60815=>"000000000",
  60816=>"000000000",
  60817=>"001000001",
  60818=>"111111111",
  60819=>"111000000",
  60820=>"011001000",
  60821=>"000000000",
  60822=>"111111111",
  60823=>"011000000",
  60824=>"110000000",
  60825=>"111010010",
  60826=>"000000110",
  60827=>"111111111",
  60828=>"111110000",
  60829=>"111101100",
  60830=>"000011111",
  60831=>"111111111",
  60832=>"000000000",
  60833=>"111011011",
  60834=>"011110111",
  60835=>"111111111",
  60836=>"001101111",
  60837=>"000000000",
  60838=>"000000000",
  60839=>"100000100",
  60840=>"011000000",
  60841=>"111111111",
  60842=>"111111111",
  60843=>"000110111",
  60844=>"010010010",
  60845=>"001000111",
  60846=>"111100000",
  60847=>"000000000",
  60848=>"111111111",
  60849=>"000000000",
  60850=>"000011111",
  60851=>"000000000",
  60852=>"111000000",
  60853=>"110111111",
  60854=>"000000000",
  60855=>"111111110",
  60856=>"000110111",
  60857=>"111111111",
  60858=>"011111111",
  60859=>"000000000",
  60860=>"000000000",
  60861=>"111111100",
  60862=>"000000000",
  60863=>"000000001",
  60864=>"000000111",
  60865=>"000000000",
  60866=>"000000000",
  60867=>"000000000",
  60868=>"111110111",
  60869=>"110111111",
  60870=>"111000000",
  60871=>"000000000",
  60872=>"000000001",
  60873=>"000000000",
  60874=>"000000000",
  60875=>"000000111",
  60876=>"000000000",
  60877=>"000000000",
  60878=>"111111111",
  60879=>"111000000",
  60880=>"001100100",
  60881=>"000100111",
  60882=>"000000000",
  60883=>"000000000",
  60884=>"001011111",
  60885=>"111101000",
  60886=>"111111010",
  60887=>"110111111",
  60888=>"111111111",
  60889=>"000100000",
  60890=>"111111111",
  60891=>"001000000",
  60892=>"111101101",
  60893=>"110110111",
  60894=>"000010010",
  60895=>"000111110",
  60896=>"000100110",
  60897=>"000000001",
  60898=>"111001001",
  60899=>"000000000",
  60900=>"111111111",
  60901=>"111101111",
  60902=>"000101111",
  60903=>"110000000",
  60904=>"001111111",
  60905=>"111101110",
  60906=>"100110000",
  60907=>"001111111",
  60908=>"010000011",
  60909=>"000000000",
  60910=>"110110111",
  60911=>"000000111",
  60912=>"000000000",
  60913=>"000100000",
  60914=>"100110000",
  60915=>"000000000",
  60916=>"111111111",
  60917=>"001000000",
  60918=>"111111111",
  60919=>"111100100",
  60920=>"000000000",
  60921=>"100000000",
  60922=>"110110111",
  60923=>"111011010",
  60924=>"111111101",
  60925=>"100111111",
  60926=>"111000000",
  60927=>"000000000",
  60928=>"110111000",
  60929=>"000100110",
  60930=>"000100011",
  60931=>"000001000",
  60932=>"000000000",
  60933=>"000111010",
  60934=>"000000000",
  60935=>"111111111",
  60936=>"100000000",
  60937=>"111111001",
  60938=>"000100110",
  60939=>"000000000",
  60940=>"001011000",
  60941=>"011011001",
  60942=>"000000111",
  60943=>"100000101",
  60944=>"111111111",
  60945=>"110111011",
  60946=>"000000111",
  60947=>"100000111",
  60948=>"111000000",
  60949=>"100100100",
  60950=>"000001111",
  60951=>"000000000",
  60952=>"000000011",
  60953=>"000101111",
  60954=>"100000000",
  60955=>"000100111",
  60956=>"111111111",
  60957=>"000000000",
  60958=>"100111111",
  60959=>"111111000",
  60960=>"111000000",
  60961=>"000011111",
  60962=>"001011000",
  60963=>"001001001",
  60964=>"110000111",
  60965=>"111111011",
  60966=>"000000000",
  60967=>"110010111",
  60968=>"110111000",
  60969=>"000010010",
  60970=>"000000000",
  60971=>"000000001",
  60972=>"100110111",
  60973=>"000000000",
  60974=>"001000000",
  60975=>"011010000",
  60976=>"111001001",
  60977=>"011011111",
  60978=>"111111001",
  60979=>"001001000",
  60980=>"000000000",
  60981=>"011111111",
  60982=>"001000000",
  60983=>"001011000",
  60984=>"111000111",
  60985=>"110001000",
  60986=>"000001000",
  60987=>"000000000",
  60988=>"111100000",
  60989=>"000000000",
  60990=>"101011001",
  60991=>"000000000",
  60992=>"000000000",
  60993=>"111111000",
  60994=>"111000000",
  60995=>"111110000",
  60996=>"001001011",
  60997=>"011011011",
  60998=>"110111000",
  60999=>"011111111",
  61000=>"000000011",
  61001=>"010111111",
  61002=>"000000100",
  61003=>"111111111",
  61004=>"001100100",
  61005=>"111011011",
  61006=>"101111011",
  61007=>"011000111",
  61008=>"000000000",
  61009=>"111111011",
  61010=>"111000111",
  61011=>"110111111",
  61012=>"111111000",
  61013=>"000000111",
  61014=>"001001011",
  61015=>"111000111",
  61016=>"000000000",
  61017=>"001101101",
  61018=>"111010000",
  61019=>"111111000",
  61020=>"111111111",
  61021=>"111111111",
  61022=>"000000011",
  61023=>"111111100",
  61024=>"000000000",
  61025=>"101100111",
  61026=>"111111000",
  61027=>"000000111",
  61028=>"000000101",
  61029=>"111000000",
  61030=>"111101100",
  61031=>"011111000",
  61032=>"111111000",
  61033=>"010000001",
  61034=>"110000111",
  61035=>"000111000",
  61036=>"110110111",
  61037=>"111111001",
  61038=>"111111111",
  61039=>"000000111",
  61040=>"001000000",
  61041=>"000000001",
  61042=>"111111111",
  61043=>"011111111",
  61044=>"111111000",
  61045=>"111111111",
  61046=>"000000011",
  61047=>"001101111",
  61048=>"111001111",
  61049=>"000000111",
  61050=>"111111011",
  61051=>"000000000",
  61052=>"000111101",
  61053=>"110111111",
  61054=>"000111000",
  61055=>"000001000",
  61056=>"100000010",
  61057=>"000000000",
  61058=>"110110111",
  61059=>"000000111",
  61060=>"111111111",
  61061=>"111000111",
  61062=>"110110110",
  61063=>"000001001",
  61064=>"111000000",
  61065=>"000000000",
  61066=>"000000111",
  61067=>"100000111",
  61068=>"111111000",
  61069=>"111111111",
  61070=>"111110111",
  61071=>"111111010",
  61072=>"111111111",
  61073=>"001111000",
  61074=>"111100000",
  61075=>"111111001",
  61076=>"000000000",
  61077=>"000000000",
  61078=>"000010011",
  61079=>"000111111",
  61080=>"000000001",
  61081=>"111111111",
  61082=>"000000000",
  61083=>"000111000",
  61084=>"000000000",
  61085=>"100001000",
  61086=>"101111000",
  61087=>"000000000",
  61088=>"110000000",
  61089=>"111110000",
  61090=>"111111000",
  61091=>"111111111",
  61092=>"100111111",
  61093=>"100000000",
  61094=>"000000011",
  61095=>"111111111",
  61096=>"111111111",
  61097=>"100000111",
  61098=>"000000111",
  61099=>"110111111",
  61100=>"001000100",
  61101=>"110010000",
  61102=>"111111101",
  61103=>"111111000",
  61104=>"111111000",
  61105=>"001001011",
  61106=>"111111010",
  61107=>"111000000",
  61108=>"110111111",
  61109=>"110000000",
  61110=>"011001001",
  61111=>"000000111",
  61112=>"111111100",
  61113=>"000000111",
  61114=>"000000001",
  61115=>"111111111",
  61116=>"111111111",
  61117=>"000100111",
  61118=>"000111111",
  61119=>"011011011",
  61120=>"100000000",
  61121=>"111111100",
  61122=>"100100111",
  61123=>"110111000",
  61124=>"111100000",
  61125=>"000111111",
  61126=>"110111111",
  61127=>"000000000",
  61128=>"000000100",
  61129=>"000100111",
  61130=>"000000000",
  61131=>"000000000",
  61132=>"000100100",
  61133=>"000010111",
  61134=>"111111110",
  61135=>"111001111",
  61136=>"011011010",
  61137=>"000000000",
  61138=>"111000000",
  61139=>"111110111",
  61140=>"000000000",
  61141=>"001000000",
  61142=>"000000011",
  61143=>"000111111",
  61144=>"000011000",
  61145=>"111111111",
  61146=>"001111111",
  61147=>"100100100",
  61148=>"111111111",
  61149=>"111011111",
  61150=>"111111011",
  61151=>"101000111",
  61152=>"111111000",
  61153=>"010010000",
  61154=>"011001000",
  61155=>"111000001",
  61156=>"000000101",
  61157=>"111110000",
  61158=>"000000111",
  61159=>"001111111",
  61160=>"110110011",
  61161=>"000001111",
  61162=>"111111001",
  61163=>"101110101",
  61164=>"111011000",
  61165=>"000000000",
  61166=>"001000111",
  61167=>"100110000",
  61168=>"111111111",
  61169=>"000000100",
  61170=>"111111111",
  61171=>"000000110",
  61172=>"000000000",
  61173=>"111111001",
  61174=>"011011001",
  61175=>"111111000",
  61176=>"111000111",
  61177=>"111011111",
  61178=>"100000111",
  61179=>"110000000",
  61180=>"001011011",
  61181=>"000000001",
  61182=>"111100001",
  61183=>"111111111",
  61184=>"111011000",
  61185=>"001000000",
  61186=>"000001001",
  61187=>"000000111",
  61188=>"101100111",
  61189=>"011001000",
  61190=>"000111111",
  61191=>"111111111",
  61192=>"000000000",
  61193=>"001000000",
  61194=>"000000000",
  61195=>"011011000",
  61196=>"000000110",
  61197=>"111011110",
  61198=>"000110000",
  61199=>"100000111",
  61200=>"001000000",
  61201=>"000000001",
  61202=>"011000110",
  61203=>"111000011",
  61204=>"011000000",
  61205=>"001000000",
  61206=>"111111110",
  61207=>"000000001",
  61208=>"000111111",
  61209=>"100100111",
  61210=>"110001100",
  61211=>"111000000",
  61212=>"011011111",
  61213=>"000000000",
  61214=>"000000111",
  61215=>"000000111",
  61216=>"000010010",
  61217=>"000101011",
  61218=>"000000000",
  61219=>"111111111",
  61220=>"000000000",
  61221=>"000100100",
  61222=>"000000000",
  61223=>"001001000",
  61224=>"110000001",
  61225=>"111111111",
  61226=>"110111111",
  61227=>"011000010",
  61228=>"000000000",
  61229=>"101100000",
  61230=>"000001000",
  61231=>"000101110",
  61232=>"010000001",
  61233=>"111111111",
  61234=>"111110100",
  61235=>"000000100",
  61236=>"000000000",
  61237=>"011011001",
  61238=>"111011011",
  61239=>"111000000",
  61240=>"000000000",
  61241=>"000000000",
  61242=>"111111111",
  61243=>"111000000",
  61244=>"110000110",
  61245=>"111111111",
  61246=>"000000111",
  61247=>"100111111",
  61248=>"111000000",
  61249=>"110011111",
  61250=>"001000000",
  61251=>"000001011",
  61252=>"000000000",
  61253=>"000000011",
  61254=>"110110111",
  61255=>"000000000",
  61256=>"111000110",
  61257=>"000000000",
  61258=>"000000000",
  61259=>"001100000",
  61260=>"110100000",
  61261=>"111111000",
  61262=>"000000000",
  61263=>"000111111",
  61264=>"111111000",
  61265=>"000000111",
  61266=>"111110111",
  61267=>"000010000",
  61268=>"000000111",
  61269=>"000000110",
  61270=>"111000000",
  61271=>"111011011",
  61272=>"100100111",
  61273=>"110011010",
  61274=>"000010110",
  61275=>"000000111",
  61276=>"111100100",
  61277=>"100000000",
  61278=>"101000000",
  61279=>"111100000",
  61280=>"111001000",
  61281=>"000000000",
  61282=>"001001101",
  61283=>"000000000",
  61284=>"000000010",
  61285=>"000000000",
  61286=>"000000000",
  61287=>"000000000",
  61288=>"101000000",
  61289=>"000001111",
  61290=>"011011111",
  61291=>"111111000",
  61292=>"100100110",
  61293=>"111111111",
  61294=>"100110111",
  61295=>"001000001",
  61296=>"111001000",
  61297=>"000000000",
  61298=>"000000001",
  61299=>"000110011",
  61300=>"111000000",
  61301=>"111101000",
  61302=>"111101000",
  61303=>"000000000",
  61304=>"000000111",
  61305=>"011011001",
  61306=>"100101101",
  61307=>"000000000",
  61308=>"010111111",
  61309=>"000000111",
  61310=>"111100000",
  61311=>"000101111",
  61312=>"110111111",
  61313=>"100111111",
  61314=>"110010010",
  61315=>"111000010",
  61316=>"000000000",
  61317=>"010010000",
  61318=>"111111111",
  61319=>"000000111",
  61320=>"111101111",
  61321=>"001000000",
  61322=>"000000000",
  61323=>"111111000",
  61324=>"111111000",
  61325=>"000100001",
  61326=>"000001001",
  61327=>"000101111",
  61328=>"001101000",
  61329=>"111111111",
  61330=>"111111110",
  61331=>"000000111",
  61332=>"111000000",
  61333=>"000000000",
  61334=>"110110111",
  61335=>"000000100",
  61336=>"000000000",
  61337=>"111111001",
  61338=>"000000111",
  61339=>"111111111",
  61340=>"000000100",
  61341=>"111011001",
  61342=>"111000000",
  61343=>"010000000",
  61344=>"111000000",
  61345=>"001011111",
  61346=>"000010101",
  61347=>"010010011",
  61348=>"000000001",
  61349=>"111111000",
  61350=>"000111110",
  61351=>"010010001",
  61352=>"000110000",
  61353=>"000111011",
  61354=>"111111110",
  61355=>"000000000",
  61356=>"000000000",
  61357=>"110000000",
  61358=>"100001001",
  61359=>"111000001",
  61360=>"111111111",
  61361=>"010110000",
  61362=>"111011000",
  61363=>"000110110",
  61364=>"000110000",
  61365=>"100110000",
  61366=>"111111111",
  61367=>"000010000",
  61368=>"010000010",
  61369=>"111111111",
  61370=>"000000000",
  61371=>"111100000",
  61372=>"110111111",
  61373=>"111111111",
  61374=>"011011001",
  61375=>"101111001",
  61376=>"011111111",
  61377=>"000111111",
  61378=>"111011011",
  61379=>"000011001",
  61380=>"100000111",
  61381=>"001001001",
  61382=>"010000001",
  61383=>"000011000",
  61384=>"111111000",
  61385=>"000000111",
  61386=>"000000000",
  61387=>"001000000",
  61388=>"000001101",
  61389=>"000000000",
  61390=>"111111000",
  61391=>"111111111",
  61392=>"001111100",
  61393=>"111111100",
  61394=>"111111001",
  61395=>"000000000",
  61396=>"000000111",
  61397=>"000000000",
  61398=>"000000010",
  61399=>"011110110",
  61400=>"000000111",
  61401=>"101000000",
  61402=>"000000000",
  61403=>"111001000",
  61404=>"000000000",
  61405=>"110000100",
  61406=>"000000000",
  61407=>"101001001",
  61408=>"100110111",
  61409=>"111000000",
  61410=>"111000111",
  61411=>"001001001",
  61412=>"110111000",
  61413=>"000000111",
  61414=>"011010100",
  61415=>"110111110",
  61416=>"100100000",
  61417=>"110111001",
  61418=>"010000100",
  61419=>"100111000",
  61420=>"000001111",
  61421=>"000000011",
  61422=>"111000111",
  61423=>"110111111",
  61424=>"000000001",
  61425=>"111100000",
  61426=>"011111100",
  61427=>"001001101",
  61428=>"000000000",
  61429=>"000100000",
  61430=>"000001001",
  61431=>"010010000",
  61432=>"000000000",
  61433=>"010111000",
  61434=>"111111000",
  61435=>"000000000",
  61436=>"000000001",
  61437=>"100000011",
  61438=>"000001000",
  61439=>"000000111",
  61440=>"011010100",
  61441=>"000000000",
  61442=>"111111111",
  61443=>"000000000",
  61444=>"001111111",
  61445=>"110010000",
  61446=>"000000000",
  61447=>"111111111",
  61448=>"111110000",
  61449=>"111100100",
  61450=>"111000000",
  61451=>"100101111",
  61452=>"100100110",
  61453=>"111101000",
  61454=>"101111111",
  61455=>"000000000",
  61456=>"000011111",
  61457=>"000000000",
  61458=>"000000000",
  61459=>"111111111",
  61460=>"000100111",
  61461=>"111111111",
  61462=>"110100111",
  61463=>"110100110",
  61464=>"001111111",
  61465=>"001001100",
  61466=>"110101111",
  61467=>"111111001",
  61468=>"111111000",
  61469=>"111000000",
  61470=>"000111111",
  61471=>"000000011",
  61472=>"111111001",
  61473=>"111111111",
  61474=>"100000000",
  61475=>"111000000",
  61476=>"100100100",
  61477=>"111111100",
  61478=>"111101111",
  61479=>"110100000",
  61480=>"001011011",
  61481=>"011000000",
  61482=>"111001001",
  61483=>"000000010",
  61484=>"000000111",
  61485=>"000000000",
  61486=>"000000000",
  61487=>"111001000",
  61488=>"001000000",
  61489=>"101100100",
  61490=>"110111111",
  61491=>"000000010",
  61492=>"001101111",
  61493=>"110110110",
  61494=>"111000000",
  61495=>"111000110",
  61496=>"111111011",
  61497=>"000000001",
  61498=>"111000000",
  61499=>"100001111",
  61500=>"111111011",
  61501=>"111111001",
  61502=>"000111111",
  61503=>"111000000",
  61504=>"111111111",
  61505=>"111111000",
  61506=>"111111100",
  61507=>"101000000",
  61508=>"111101101",
  61509=>"001011010",
  61510=>"111110000",
  61511=>"111111111",
  61512=>"111111001",
  61513=>"111111111",
  61514=>"000111111",
  61515=>"000000000",
  61516=>"111111000",
  61517=>"111111010",
  61518=>"000000000",
  61519=>"000000000",
  61520=>"100000000",
  61521=>"111001000",
  61522=>"001000011",
  61523=>"111100000",
  61524=>"111100111",
  61525=>"000000000",
  61526=>"111000000",
  61527=>"000111111",
  61528=>"000000000",
  61529=>"111000000",
  61530=>"111000000",
  61531=>"000010000",
  61532=>"000110111",
  61533=>"000111111",
  61534=>"100100111",
  61535=>"111111111",
  61536=>"000000000",
  61537=>"000000010",
  61538=>"000000111",
  61539=>"000000111",
  61540=>"000000011",
  61541=>"011000000",
  61542=>"111111111",
  61543=>"000000000",
  61544=>"110101111",
  61545=>"001111111",
  61546=>"111000000",
  61547=>"110000000",
  61548=>"000100111",
  61549=>"000011111",
  61550=>"111111111",
  61551=>"110111111",
  61552=>"000000000",
  61553=>"001000111",
  61554=>"110111001",
  61555=>"000010111",
  61556=>"010000000",
  61557=>"000000000",
  61558=>"000000000",
  61559=>"000000101",
  61560=>"110110100",
  61561=>"100000000",
  61562=>"000001111",
  61563=>"000000000",
  61564=>"000000110",
  61565=>"101000100",
  61566=>"000000011",
  61567=>"000000001",
  61568=>"000111111",
  61569=>"111100000",
  61570=>"111000000",
  61571=>"100100000",
  61572=>"111000000",
  61573=>"001000000",
  61574=>"111000110",
  61575=>"000000010",
  61576=>"001101000",
  61577=>"111111111",
  61578=>"000100111",
  61579=>"000000111",
  61580=>"001011001",
  61581=>"111000000",
  61582=>"111111111",
  61583=>"000111111",
  61584=>"111000000",
  61585=>"010110010",
  61586=>"111111111",
  61587=>"011000000",
  61588=>"111111111",
  61589=>"000000111",
  61590=>"111111000",
  61591=>"111000000",
  61592=>"101101000",
  61593=>"111111111",
  61594=>"111000000",
  61595=>"000101111",
  61596=>"111000000",
  61597=>"000000001",
  61598=>"000000000",
  61599=>"111111111",
  61600=>"110000000",
  61601=>"000001111",
  61602=>"000111000",
  61603=>"111111111",
  61604=>"000001001",
  61605=>"100110100",
  61606=>"001000000",
  61607=>"000000011",
  61608=>"000010110",
  61609=>"000000000",
  61610=>"000000100",
  61611=>"111111111",
  61612=>"000111111",
  61613=>"000110111",
  61614=>"100000000",
  61615=>"001101111",
  61616=>"000000000",
  61617=>"011011011",
  61618=>"111111111",
  61619=>"111111000",
  61620=>"001000111",
  61621=>"010111111",
  61622=>"000011111",
  61623=>"010111111",
  61624=>"100000001",
  61625=>"000000000",
  61626=>"000000000",
  61627=>"111000000",
  61628=>"000000100",
  61629=>"110000000",
  61630=>"100000111",
  61631=>"110111011",
  61632=>"101111111",
  61633=>"001000000",
  61634=>"000000000",
  61635=>"000100000",
  61636=>"111001011",
  61637=>"000000000",
  61638=>"000000000",
  61639=>"111111111",
  61640=>"000111111",
  61641=>"000111111",
  61642=>"000111110",
  61643=>"111111000",
  61644=>"000100111",
  61645=>"100000000",
  61646=>"111111001",
  61647=>"000010111",
  61648=>"101000000",
  61649=>"001101111",
  61650=>"000111111",
  61651=>"000001111",
  61652=>"111100000",
  61653=>"111111111",
  61654=>"000111111",
  61655=>"011111111",
  61656=>"000110111",
  61657=>"101111111",
  61658=>"111111000",
  61659=>"101111111",
  61660=>"000000000",
  61661=>"111111111",
  61662=>"000000010",
  61663=>"111000000",
  61664=>"111001000",
  61665=>"010011010",
  61666=>"000111111",
  61667=>"100100000",
  61668=>"111000000",
  61669=>"110111100",
  61670=>"000111111",
  61671=>"111111111",
  61672=>"111111111",
  61673=>"000000001",
  61674=>"000000101",
  61675=>"100101100",
  61676=>"000111111",
  61677=>"000000001",
  61678=>"010111101",
  61679=>"111111000",
  61680=>"100000000",
  61681=>"000111111",
  61682=>"000000111",
  61683=>"000011000",
  61684=>"111111000",
  61685=>"110111111",
  61686=>"110010010",
  61687=>"000000000",
  61688=>"000000000",
  61689=>"000000000",
  61690=>"111111000",
  61691=>"000000110",
  61692=>"000100100",
  61693=>"000010111",
  61694=>"000000000",
  61695=>"110000000",
  61696=>"001000000",
  61697=>"001111111",
  61698=>"000001000",
  61699=>"000111000",
  61700=>"000000000",
  61701=>"111111111",
  61702=>"000000000",
  61703=>"111111111",
  61704=>"000000000",
  61705=>"000001111",
  61706=>"000000000",
  61707=>"011111111",
  61708=>"011000111",
  61709=>"100000010",
  61710=>"000011111",
  61711=>"000000000",
  61712=>"000000000",
  61713=>"000000100",
  61714=>"111000000",
  61715=>"100001000",
  61716=>"111111111",
  61717=>"111000110",
  61718=>"001100100",
  61719=>"110111110",
  61720=>"000000000",
  61721=>"111111111",
  61722=>"111000000",
  61723=>"000000000",
  61724=>"000111000",
  61725=>"111101000",
  61726=>"000000000",
  61727=>"000000000",
  61728=>"001111111",
  61729=>"111000000",
  61730=>"111000000",
  61731=>"111110000",
  61732=>"101100000",
  61733=>"000111100",
  61734=>"111111111",
  61735=>"011111111",
  61736=>"000111111",
  61737=>"111001000",
  61738=>"000110110",
  61739=>"000000111",
  61740=>"000011111",
  61741=>"001011010",
  61742=>"000000111",
  61743=>"000000111",
  61744=>"000000110",
  61745=>"110101011",
  61746=>"000100111",
  61747=>"011011001",
  61748=>"111100000",
  61749=>"111111111",
  61750=>"111010000",
  61751=>"000000000",
  61752=>"110110000",
  61753=>"000000000",
  61754=>"000110111",
  61755=>"101111111",
  61756=>"100000000",
  61757=>"111111000",
  61758=>"100100000",
  61759=>"000000110",
  61760=>"000000111",
  61761=>"000101000",
  61762=>"000000000",
  61763=>"111000000",
  61764=>"001000001",
  61765=>"000000001",
  61766=>"000001001",
  61767=>"100100110",
  61768=>"000000000",
  61769=>"000000000",
  61770=>"000111100",
  61771=>"001011111",
  61772=>"000111111",
  61773=>"100100010",
  61774=>"111111000",
  61775=>"000000100",
  61776=>"000011111",
  61777=>"111111111",
  61778=>"000000000",
  61779=>"000000010",
  61780=>"100000000",
  61781=>"001001011",
  61782=>"111000000",
  61783=>"111000000",
  61784=>"000000101",
  61785=>"000001000",
  61786=>"001111011",
  61787=>"000000000",
  61788=>"001000000",
  61789=>"111111111",
  61790=>"111000000",
  61791=>"000010110",
  61792=>"111111110",
  61793=>"111101000",
  61794=>"000010110",
  61795=>"111000000",
  61796=>"110100000",
  61797=>"000001111",
  61798=>"000101111",
  61799=>"000000000",
  61800=>"000110111",
  61801=>"100100000",
  61802=>"000000000",
  61803=>"101000000",
  61804=>"000000000",
  61805=>"000000000",
  61806=>"111111111",
  61807=>"000111111",
  61808=>"000000110",
  61809=>"111001000",
  61810=>"000000000",
  61811=>"000111111",
  61812=>"111111111",
  61813=>"001000011",
  61814=>"000000000",
  61815=>"000100001",
  61816=>"000000111",
  61817=>"111111111",
  61818=>"111111111",
  61819=>"110110111",
  61820=>"000000000",
  61821=>"111011000",
  61822=>"111111111",
  61823=>"000000000",
  61824=>"000111111",
  61825=>"111111111",
  61826=>"100111111",
  61827=>"111111110",
  61828=>"000111111",
  61829=>"011101011",
  61830=>"000010000",
  61831=>"100100000",
  61832=>"111000000",
  61833=>"000000000",
  61834=>"111011000",
  61835=>"000111111",
  61836=>"111111111",
  61837=>"000000000",
  61838=>"101100111",
  61839=>"000000111",
  61840=>"000110000",
  61841=>"101011111",
  61842=>"111111011",
  61843=>"000000000",
  61844=>"000101111",
  61845=>"000010010",
  61846=>"101100111",
  61847=>"001000000",
  61848=>"011000100",
  61849=>"111111110",
  61850=>"111111111",
  61851=>"000000111",
  61852=>"000001111",
  61853=>"011000000",
  61854=>"000000000",
  61855=>"111110110",
  61856=>"000111000",
  61857=>"011001011",
  61858=>"000101111",
  61859=>"000111111",
  61860=>"101111111",
  61861=>"100111100",
  61862=>"111101000",
  61863=>"111111001",
  61864=>"101000111",
  61865=>"000000000",
  61866=>"111111111",
  61867=>"111000010",
  61868=>"000000110",
  61869=>"111000000",
  61870=>"000110000",
  61871=>"000000000",
  61872=>"111000000",
  61873=>"111111000",
  61874=>"111111110",
  61875=>"000000000",
  61876=>"000000001",
  61877=>"111111111",
  61878=>"000100111",
  61879=>"000111101",
  61880=>"111111000",
  61881=>"111111111",
  61882=>"111111110",
  61883=>"100000011",
  61884=>"111111001",
  61885=>"111111111",
  61886=>"101000000",
  61887=>"100100100",
  61888=>"001000000",
  61889=>"110000000",
  61890=>"000000111",
  61891=>"111000000",
  61892=>"000001001",
  61893=>"000000000",
  61894=>"111010000",
  61895=>"000110110",
  61896=>"000000000",
  61897=>"111110110",
  61898=>"101001000",
  61899=>"111100000",
  61900=>"011111111",
  61901=>"000000111",
  61902=>"100111100",
  61903=>"111111001",
  61904=>"001000001",
  61905=>"100000001",
  61906=>"100111111",
  61907=>"111111111",
  61908=>"001111111",
  61909=>"100000000",
  61910=>"000010111",
  61911=>"000001101",
  61912=>"101000000",
  61913=>"100100000",
  61914=>"001000011",
  61915=>"000000101",
  61916=>"000000001",
  61917=>"011111111",
  61918=>"000000100",
  61919=>"001011001",
  61920=>"101000110",
  61921=>"111111111",
  61922=>"001000000",
  61923=>"111111111",
  61924=>"111111111",
  61925=>"000000110",
  61926=>"000010111",
  61927=>"000000001",
  61928=>"101111110",
  61929=>"000111111",
  61930=>"111011000",
  61931=>"100111111",
  61932=>"111111111",
  61933=>"001001001",
  61934=>"111111111",
  61935=>"000000000",
  61936=>"111100000",
  61937=>"000111000",
  61938=>"000000000",
  61939=>"101101111",
  61940=>"000001010",
  61941=>"011001111",
  61942=>"111111011",
  61943=>"111000000",
  61944=>"000000000",
  61945=>"001001000",
  61946=>"100100000",
  61947=>"000000111",
  61948=>"110111111",
  61949=>"111001000",
  61950=>"001000000",
  61951=>"000000011",
  61952=>"000001101",
  61953=>"000000000",
  61954=>"111101111",
  61955=>"111111111",
  61956=>"000001110",
  61957=>"111111111",
  61958=>"000100000",
  61959=>"111111111",
  61960=>"000010011",
  61961=>"001101111",
  61962=>"100111111",
  61963=>"000111111",
  61964=>"000000000",
  61965=>"000000100",
  61966=>"000000000",
  61967=>"000000000",
  61968=>"110110111",
  61969=>"000001000",
  61970=>"110111111",
  61971=>"000000000",
  61972=>"001000000",
  61973=>"000000000",
  61974=>"000100000",
  61975=>"111111111",
  61976=>"000000000",
  61977=>"000000100",
  61978=>"000000000",
  61979=>"010001010",
  61980=>"111111111",
  61981=>"100000000",
  61982=>"000000000",
  61983=>"000000000",
  61984=>"000000000",
  61985=>"111111111",
  61986=>"010000000",
  61987=>"000000000",
  61988=>"000000111",
  61989=>"111110000",
  61990=>"110111110",
  61991=>"011000000",
  61992=>"011111001",
  61993=>"000000000",
  61994=>"111111111",
  61995=>"001111000",
  61996=>"111111011",
  61997=>"000001000",
  61998=>"101101100",
  61999=>"000110110",
  62000=>"000000000",
  62001=>"000111000",
  62002=>"110110111",
  62003=>"000000000",
  62004=>"110111111",
  62005=>"101101000",
  62006=>"010110100",
  62007=>"111111111",
  62008=>"001011111",
  62009=>"011010000",
  62010=>"100101101",
  62011=>"000000000",
  62012=>"000101101",
  62013=>"000000000",
  62014=>"000110111",
  62015=>"111111001",
  62016=>"000000000",
  62017=>"010110010",
  62018=>"011000000",
  62019=>"001010000",
  62020=>"000001001",
  62021=>"110111111",
  62022=>"000000000",
  62023=>"111111000",
  62024=>"011001001",
  62025=>"111101101",
  62026=>"111111111",
  62027=>"111110000",
  62028=>"101001000",
  62029=>"101111111",
  62030=>"000000100",
  62031=>"111111111",
  62032=>"111111110",
  62033=>"000000110",
  62034=>"000000000",
  62035=>"011111111",
  62036=>"000000000",
  62037=>"000000000",
  62038=>"111111111",
  62039=>"111111100",
  62040=>"011111110",
  62041=>"000000000",
  62042=>"100100001",
  62043=>"000000000",
  62044=>"011011000",
  62045=>"110111111",
  62046=>"000111111",
  62047=>"000000000",
  62048=>"000000001",
  62049=>"000000000",
  62050=>"001010100",
  62051=>"000000000",
  62052=>"111111111",
  62053=>"000000000",
  62054=>"111100000",
  62055=>"000000000",
  62056=>"000000000",
  62057=>"111111111",
  62058=>"000000111",
  62059=>"010000011",
  62060=>"001011011",
  62061=>"111111111",
  62062=>"111111111",
  62063=>"011111111",
  62064=>"111100100",
  62065=>"001001001",
  62066=>"111111111",
  62067=>"111111010",
  62068=>"000000000",
  62069=>"001001000",
  62070=>"011000111",
  62071=>"111111111",
  62072=>"000000100",
  62073=>"100000000",
  62074=>"111111111",
  62075=>"000000000",
  62076=>"111111111",
  62077=>"000100100",
  62078=>"101000000",
  62079=>"000000000",
  62080=>"000111111",
  62081=>"011011000",
  62082=>"000000000",
  62083=>"000000011",
  62084=>"000000000",
  62085=>"000000000",
  62086=>"010010111",
  62087=>"000011111",
  62088=>"111000000",
  62089=>"000011111",
  62090=>"111011000",
  62091=>"111000000",
  62092=>"000000000",
  62093=>"111111111",
  62094=>"111110111",
  62095=>"000100110",
  62096=>"111111111",
  62097=>"000000000",
  62098=>"111101111",
  62099=>"000000100",
  62100=>"111111111",
  62101=>"000000000",
  62102=>"111000000",
  62103=>"111111101",
  62104=>"111111111",
  62105=>"111101111",
  62106=>"000111111",
  62107=>"000000000",
  62108=>"111111000",
  62109=>"000101111",
  62110=>"100000111",
  62111=>"000000000",
  62112=>"000000000",
  62113=>"111111111",
  62114=>"001001111",
  62115=>"111111111",
  62116=>"111001000",
  62117=>"000000111",
  62118=>"010100111",
  62119=>"001111011",
  62120=>"001000111",
  62121=>"111111111",
  62122=>"000001111",
  62123=>"111000000",
  62124=>"111011000",
  62125=>"001000110",
  62126=>"111001000",
  62127=>"000000100",
  62128=>"000000000",
  62129=>"000000000",
  62130=>"110100100",
  62131=>"111101000",
  62132=>"000000000",
  62133=>"111100101",
  62134=>"111111111",
  62135=>"111111111",
  62136=>"111111110",
  62137=>"000000000",
  62138=>"000000000",
  62139=>"000000100",
  62140=>"111111111",
  62141=>"011111000",
  62142=>"111111111",
  62143=>"010000001",
  62144=>"000000000",
  62145=>"000000111",
  62146=>"000000100",
  62147=>"000000000",
  62148=>"000011111",
  62149=>"111111111",
  62150=>"000000111",
  62151=>"000110111",
  62152=>"000111100",
  62153=>"111111111",
  62154=>"101100000",
  62155=>"111111001",
  62156=>"100110111",
  62157=>"000000000",
  62158=>"111111101",
  62159=>"000000000",
  62160=>"001000000",
  62161=>"000000100",
  62162=>"111111111",
  62163=>"111111111",
  62164=>"111111000",
  62165=>"111111111",
  62166=>"100111111",
  62167=>"000001111",
  62168=>"111111111",
  62169=>"011011111",
  62170=>"011000000",
  62171=>"000000001",
  62172=>"101101111",
  62173=>"001000000",
  62174=>"001001010",
  62175=>"000000000",
  62176=>"000000000",
  62177=>"000000000",
  62178=>"011000000",
  62179=>"101001001",
  62180=>"000000000",
  62181=>"000000000",
  62182=>"011011000",
  62183=>"000000000",
  62184=>"000000000",
  62185=>"111111111",
  62186=>"000000000",
  62187=>"000000000",
  62188=>"110100000",
  62189=>"111111111",
  62190=>"001010111",
  62191=>"000000100",
  62192=>"010110111",
  62193=>"011000000",
  62194=>"000111111",
  62195=>"111001001",
  62196=>"111111111",
  62197=>"000000000",
  62198=>"111101111",
  62199=>"000000111",
  62200=>"111111111",
  62201=>"000000000",
  62202=>"000000000",
  62203=>"111111100",
  62204=>"000011001",
  62205=>"111001101",
  62206=>"000000000",
  62207=>"111111111",
  62208=>"010000000",
  62209=>"001011011",
  62210=>"000010111",
  62211=>"111000000",
  62212=>"000001001",
  62213=>"110000110",
  62214=>"110110000",
  62215=>"101100000",
  62216=>"111111111",
  62217=>"000000000",
  62218=>"000000100",
  62219=>"000001111",
  62220=>"111000101",
  62221=>"100000000",
  62222=>"000000011",
  62223=>"111110110",
  62224=>"011001001",
  62225=>"001111111",
  62226=>"110000000",
  62227=>"000000100",
  62228=>"000110111",
  62229=>"000000000",
  62230=>"000000100",
  62231=>"111111110",
  62232=>"000000000",
  62233=>"100111111",
  62234=>"000000000",
  62235=>"010011111",
  62236=>"100111011",
  62237=>"100000000",
  62238=>"000011011",
  62239=>"111111001",
  62240=>"110110111",
  62241=>"001000000",
  62242=>"000000000",
  62243=>"101000000",
  62244=>"111111001",
  62245=>"000000000",
  62246=>"000000000",
  62247=>"101111111",
  62248=>"000000000",
  62249=>"000110110",
  62250=>"001000111",
  62251=>"000000000",
  62252=>"000000000",
  62253=>"111111111",
  62254=>"000000000",
  62255=>"000000000",
  62256=>"100100100",
  62257=>"111111111",
  62258=>"111010110",
  62259=>"000000000",
  62260=>"011111111",
  62261=>"000000100",
  62262=>"001011111",
  62263=>"000000000",
  62264=>"100100101",
  62265=>"111111111",
  62266=>"000000111",
  62267=>"000010010",
  62268=>"111111111",
  62269=>"100100100",
  62270=>"111111111",
  62271=>"111010000",
  62272=>"111000000",
  62273=>"000001001",
  62274=>"111111110",
  62275=>"111111001",
  62276=>"001001001",
  62277=>"011011000",
  62278=>"100111111",
  62279=>"000100000",
  62280=>"000000000",
  62281=>"000011000",
  62282=>"000000000",
  62283=>"001001000",
  62284=>"001001101",
  62285=>"010000000",
  62286=>"011111111",
  62287=>"011111111",
  62288=>"000000000",
  62289=>"111000000",
  62290=>"111000000",
  62291=>"001001111",
  62292=>"000000000",
  62293=>"011011011",
  62294=>"000000110",
  62295=>"110100111",
  62296=>"111111111",
  62297=>"000000000",
  62298=>"111010000",
  62299=>"100000000",
  62300=>"000111111",
  62301=>"111111111",
  62302=>"000000100",
  62303=>"101001001",
  62304=>"111111111",
  62305=>"111111001",
  62306=>"011000000",
  62307=>"111111111",
  62308=>"000111111",
  62309=>"111000100",
  62310=>"111111111",
  62311=>"000000000",
  62312=>"000000000",
  62313=>"011010110",
  62314=>"100001111",
  62315=>"111111101",
  62316=>"001001001",
  62317=>"111111111",
  62318=>"000000000",
  62319=>"111111000",
  62320=>"000111111",
  62321=>"100111100",
  62322=>"100000000",
  62323=>"000000000",
  62324=>"100110000",
  62325=>"111110000",
  62326=>"100100110",
  62327=>"000001001",
  62328=>"111111111",
  62329=>"011111110",
  62330=>"000000000",
  62331=>"000000000",
  62332=>"111111100",
  62333=>"000000000",
  62334=>"111111111",
  62335=>"000110000",
  62336=>"001000101",
  62337=>"000000000",
  62338=>"111111111",
  62339=>"011001000",
  62340=>"111111111",
  62341=>"000000000",
  62342=>"000000000",
  62343=>"101111111",
  62344=>"000001000",
  62345=>"101111100",
  62346=>"110110110",
  62347=>"000010111",
  62348=>"111111111",
  62349=>"111111000",
  62350=>"010000000",
  62351=>"000000000",
  62352=>"000000000",
  62353=>"111111111",
  62354=>"111111001",
  62355=>"111111111",
  62356=>"111111001",
  62357=>"000000011",
  62358=>"000001111",
  62359=>"111001000",
  62360=>"000111111",
  62361=>"001000000",
  62362=>"000000000",
  62363=>"001001111",
  62364=>"111101111",
  62365=>"000000000",
  62366=>"100000000",
  62367=>"111111100",
  62368=>"000000000",
  62369=>"111111111",
  62370=>"111110000",
  62371=>"011011001",
  62372=>"111111100",
  62373=>"000000001",
  62374=>"000000000",
  62375=>"111111111",
  62376=>"001000000",
  62377=>"001000000",
  62378=>"000011011",
  62379=>"000000000",
  62380=>"000000000",
  62381=>"000000000",
  62382=>"010010000",
  62383=>"000000100",
  62384=>"111110000",
  62385=>"001111111",
  62386=>"001110111",
  62387=>"000000000",
  62388=>"001111111",
  62389=>"111111001",
  62390=>"011110111",
  62391=>"110000101",
  62392=>"001000000",
  62393=>"001000100",
  62394=>"000001000",
  62395=>"111111111",
  62396=>"000000000",
  62397=>"000000000",
  62398=>"000000000",
  62399=>"110111000",
  62400=>"111000000",
  62401=>"111111111",
  62402=>"000000000",
  62403=>"111111111",
  62404=>"111001001",
  62405=>"111111111",
  62406=>"111110001",
  62407=>"110010000",
  62408=>"000000000",
  62409=>"011011001",
  62410=>"000100000",
  62411=>"000000001",
  62412=>"111000000",
  62413=>"111011101",
  62414=>"011000000",
  62415=>"000000000",
  62416=>"000000101",
  62417=>"111111101",
  62418=>"000001001",
  62419=>"111011111",
  62420=>"111110100",
  62421=>"101111111",
  62422=>"000000000",
  62423=>"000000000",
  62424=>"110000000",
  62425=>"111111111",
  62426=>"000000111",
  62427=>"110111111",
  62428=>"100001001",
  62429=>"111111111",
  62430=>"111111011",
  62431=>"000000000",
  62432=>"011111100",
  62433=>"000011101",
  62434=>"000000110",
  62435=>"000101100",
  62436=>"111111001",
  62437=>"111111100",
  62438=>"000000000",
  62439=>"111111111",
  62440=>"001001000",
  62441=>"110111111",
  62442=>"001000100",
  62443=>"101000000",
  62444=>"000111001",
  62445=>"100000000",
  62446=>"000111111",
  62447=>"000111111",
  62448=>"111101001",
  62449=>"110110110",
  62450=>"111101000",
  62451=>"000000000",
  62452=>"011001000",
  62453=>"111111111",
  62454=>"000000111",
  62455=>"100111111",
  62456=>"000000000",
  62457=>"100101001",
  62458=>"000011000",
  62459=>"000000000",
  62460=>"100000000",
  62461=>"000100000",
  62462=>"011000000",
  62463=>"000000000",
  62464=>"001101101",
  62465=>"111111111",
  62466=>"001101111",
  62467=>"111110100",
  62468=>"001111111",
  62469=>"010010001",
  62470=>"000000000",
  62471=>"100000000",
  62472=>"000000000",
  62473=>"001011011",
  62474=>"111111111",
  62475=>"000000010",
  62476=>"110110110",
  62477=>"011110111",
  62478=>"010010000",
  62479=>"010011111",
  62480=>"001000000",
  62481=>"000000000",
  62482=>"111101111",
  62483=>"000000001",
  62484=>"000000000",
  62485=>"110000011",
  62486=>"000000011",
  62487=>"000001110",
  62488=>"000000000",
  62489=>"111101101",
  62490=>"000010000",
  62491=>"000001001",
  62492=>"110111111",
  62493=>"000110000",
  62494=>"111111111",
  62495=>"110111100",
  62496=>"110010000",
  62497=>"111011000",
  62498=>"101111001",
  62499=>"000011011",
  62500=>"000000000",
  62501=>"001000000",
  62502=>"011010100",
  62503=>"111111111",
  62504=>"000011011",
  62505=>"111111111",
  62506=>"000000100",
  62507=>"111111111",
  62508=>"111111000",
  62509=>"000000111",
  62510=>"010010000",
  62511=>"011000000",
  62512=>"111011001",
  62513=>"000000000",
  62514=>"100111101",
  62515=>"000111000",
  62516=>"010110100",
  62517=>"111111100",
  62518=>"000000001",
  62519=>"001001000",
  62520=>"111111111",
  62521=>"110000001",
  62522=>"100111110",
  62523=>"001000101",
  62524=>"001000000",
  62525=>"100000000",
  62526=>"011010000",
  62527=>"111111111",
  62528=>"111111111",
  62529=>"000000001",
  62530=>"000000000",
  62531=>"100100111",
  62532=>"111111011",
  62533=>"000000000",
  62534=>"110000000",
  62535=>"111111111",
  62536=>"000110000",
  62537=>"101101111",
  62538=>"000000000",
  62539=>"001000001",
  62540=>"000000000",
  62541=>"011011001",
  62542=>"110000000",
  62543=>"000000000",
  62544=>"000000001",
  62545=>"111011011",
  62546=>"000100110",
  62547=>"100000001",
  62548=>"110111111",
  62549=>"110100000",
  62550=>"011110111",
  62551=>"000000000",
  62552=>"000000000",
  62553=>"000000000",
  62554=>"011011111",
  62555=>"011111110",
  62556=>"000000000",
  62557=>"000000000",
  62558=>"111111111",
  62559=>"010000111",
  62560=>"000000000",
  62561=>"100101000",
  62562=>"111111111",
  62563=>"011111111",
  62564=>"101101000",
  62565=>"111111111",
  62566=>"111111100",
  62567=>"000000000",
  62568=>"001000000",
  62569=>"111111011",
  62570=>"011111111",
  62571=>"000011111",
  62572=>"000001001",
  62573=>"000000000",
  62574=>"000001000",
  62575=>"000011001",
  62576=>"000001000",
  62577=>"000000001",
  62578=>"111111111",
  62579=>"000000111",
  62580=>"100001111",
  62581=>"001011000",
  62582=>"111111001",
  62583=>"000000000",
  62584=>"000100111",
  62585=>"000010000",
  62586=>"101000000",
  62587=>"000000001",
  62588=>"110000000",
  62589=>"000000000",
  62590=>"110010000",
  62591=>"000000000",
  62592=>"000111111",
  62593=>"111111000",
  62594=>"000011111",
  62595=>"000000000",
  62596=>"110110111",
  62597=>"111001001",
  62598=>"111111110",
  62599=>"010111010",
  62600=>"000110111",
  62601=>"111111111",
  62602=>"111111111",
  62603=>"111110111",
  62604=>"111110100",
  62605=>"110110000",
  62606=>"100111111",
  62607=>"000110000",
  62608=>"111100000",
  62609=>"000010110",
  62610=>"001000000",
  62611=>"011100111",
  62612=>"110110101",
  62613=>"111111110",
  62614=>"001001101",
  62615=>"001001001",
  62616=>"001011111",
  62617=>"111111101",
  62618=>"101000000",
  62619=>"001101000",
  62620=>"011000011",
  62621=>"000000111",
  62622=>"111111111",
  62623=>"001010011",
  62624=>"000001111",
  62625=>"110111111",
  62626=>"000010000",
  62627=>"000000000",
  62628=>"111111101",
  62629=>"110010010",
  62630=>"111001000",
  62631=>"001001011",
  62632=>"111111111",
  62633=>"000000001",
  62634=>"000000000",
  62635=>"111001011",
  62636=>"111011011",
  62637=>"111101101",
  62638=>"000000000",
  62639=>"110011011",
  62640=>"000001111",
  62641=>"110111011",
  62642=>"111111110",
  62643=>"000000000",
  62644=>"001101111",
  62645=>"000000000",
  62646=>"011111110",
  62647=>"000000010",
  62648=>"000000000",
  62649=>"101001101",
  62650=>"100001000",
  62651=>"111111111",
  62652=>"111010010",
  62653=>"111110100",
  62654=>"000000000",
  62655=>"111111101",
  62656=>"111111111",
  62657=>"110111111",
  62658=>"011010000",
  62659=>"000000111",
  62660=>"100000000",
  62661=>"000000111",
  62662=>"111011001",
  62663=>"111111111",
  62664=>"001111111",
  62665=>"011000111",
  62666=>"110110000",
  62667=>"111011011",
  62668=>"111111000",
  62669=>"111111110",
  62670=>"111111001",
  62671=>"000000110",
  62672=>"111100000",
  62673=>"000001010",
  62674=>"111111111",
  62675=>"000011011",
  62676=>"110111101",
  62677=>"001111110",
  62678=>"000000111",
  62679=>"110000000",
  62680=>"100000000",
  62681=>"111111111",
  62682=>"100100100",
  62683=>"000110110",
  62684=>"000000111",
  62685=>"100011001",
  62686=>"111111111",
  62687=>"110110110",
  62688=>"111111000",
  62689=>"011000001",
  62690=>"101001100",
  62691=>"000000111",
  62692=>"000001000",
  62693=>"101000000",
  62694=>"111111111",
  62695=>"010011000",
  62696=>"011000000",
  62697=>"100111111",
  62698=>"011000000",
  62699=>"110110000",
  62700=>"110111111",
  62701=>"111111111",
  62702=>"110111111",
  62703=>"111111000",
  62704=>"111010000",
  62705=>"000001111",
  62706=>"001011011",
  62707=>"011110000",
  62708=>"000000110",
  62709=>"011111111",
  62710=>"001001101",
  62711=>"111111111",
  62712=>"001000000",
  62713=>"111101000",
  62714=>"000101111",
  62715=>"011010110",
  62716=>"010010100",
  62717=>"111110100",
  62718=>"000000000",
  62719=>"000101011",
  62720=>"001001100",
  62721=>"111101100",
  62722=>"000000111",
  62723=>"111111011",
  62724=>"011001000",
  62725=>"001001000",
  62726=>"111111111",
  62727=>"000111001",
  62728=>"000110111",
  62729=>"111111111",
  62730=>"010010000",
  62731=>"110111111",
  62732=>"000000100",
  62733=>"111010001",
  62734=>"111111110",
  62735=>"111111111",
  62736=>"100000000",
  62737=>"001111111",
  62738=>"100000000",
  62739=>"000110000",
  62740=>"000000001",
  62741=>"101001011",
  62742=>"001001110",
  62743=>"000000000",
  62744=>"000000011",
  62745=>"000000000",
  62746=>"000000000",
  62747=>"000001000",
  62748=>"111111111",
  62749=>"011100000",
  62750=>"111111111",
  62751=>"110110110",
  62752=>"000111111",
  62753=>"101100000",
  62754=>"010001101",
  62755=>"111110000",
  62756=>"110110010",
  62757=>"000111111",
  62758=>"000110110",
  62759=>"000011011",
  62760=>"000000000",
  62761=>"100111111",
  62762=>"111110000",
  62763=>"000000000",
  62764=>"000011011",
  62765=>"011111111",
  62766=>"000000000",
  62767=>"000000000",
  62768=>"100100000",
  62769=>"000000000",
  62770=>"000000111",
  62771=>"010000000",
  62772=>"111111111",
  62773=>"100100110",
  62774=>"111111011",
  62775=>"000000000",
  62776=>"011000000",
  62777=>"000000000",
  62778=>"000000000",
  62779=>"111111011",
  62780=>"111011111",
  62781=>"000001000",
  62782=>"110110110",
  62783=>"100110100",
  62784=>"000001111",
  62785=>"110100111",
  62786=>"011111111",
  62787=>"001000000",
  62788=>"111010100",
  62789=>"000000100",
  62790=>"000000000",
  62791=>"111111111",
  62792=>"111110001",
  62793=>"000000000",
  62794=>"111110000",
  62795=>"000000100",
  62796=>"011000000",
  62797=>"111100111",
  62798=>"000110110",
  62799=>"000101101",
  62800=>"000100101",
  62801=>"111111101",
  62802=>"000000000",
  62803=>"000000000",
  62804=>"000000000",
  62805=>"001111111",
  62806=>"111000001",
  62807=>"100111111",
  62808=>"110111111",
  62809=>"000100111",
  62810=>"010100111",
  62811=>"000000000",
  62812=>"101101111",
  62813=>"000000010",
  62814=>"000100000",
  62815=>"111001000",
  62816=>"001001000",
  62817=>"000000000",
  62818=>"010100100",
  62819=>"101101000",
  62820=>"100000000",
  62821=>"000011111",
  62822=>"111001011",
  62823=>"000000000",
  62824=>"101000101",
  62825=>"000000001",
  62826=>"111100000",
  62827=>"011010000",
  62828=>"000100001",
  62829=>"111111010",
  62830=>"000000101",
  62831=>"111101110",
  62832=>"000000000",
  62833=>"111111111",
  62834=>"000000000",
  62835=>"010010000",
  62836=>"000001001",
  62837=>"000000000",
  62838=>"111111011",
  62839=>"000000001",
  62840=>"000000000",
  62841=>"111111111",
  62842=>"000000000",
  62843=>"000000000",
  62844=>"011011010",
  62845=>"011001000",
  62846=>"000100000",
  62847=>"001101111",
  62848=>"000000000",
  62849=>"110111001",
  62850=>"000110100",
  62851=>"111111111",
  62852=>"000111100",
  62853=>"000000000",
  62854=>"000000000",
  62855=>"111110100",
  62856=>"100000000",
  62857=>"110111011",
  62858=>"001000000",
  62859=>"001001001",
  62860=>"000111111",
  62861=>"100110111",
  62862=>"000000000",
  62863=>"000000000",
  62864=>"000000000",
  62865=>"010110110",
  62866=>"011011001",
  62867=>"110110111",
  62868=>"111111000",
  62869=>"000000000",
  62870=>"000010010",
  62871=>"111111100",
  62872=>"000000000",
  62873=>"000110001",
  62874=>"111111111",
  62875=>"111111111",
  62876=>"000000111",
  62877=>"110010000",
  62878=>"111111010",
  62879=>"000000000",
  62880=>"000000000",
  62881=>"010001000",
  62882=>"001000000",
  62883=>"000000000",
  62884=>"000110000",
  62885=>"000110111",
  62886=>"000000000",
  62887=>"101111111",
  62888=>"000000000",
  62889=>"110110001",
  62890=>"111001000",
  62891=>"110000000",
  62892=>"000000000",
  62893=>"110110111",
  62894=>"011011111",
  62895=>"111111111",
  62896=>"111001001",
  62897=>"101111111",
  62898=>"000000110",
  62899=>"001011110",
  62900=>"100010000",
  62901=>"110110000",
  62902=>"111111111",
  62903=>"000000000",
  62904=>"111111111",
  62905=>"111111111",
  62906=>"010000100",
  62907=>"000001001",
  62908=>"010010000",
  62909=>"111111111",
  62910=>"111011000",
  62911=>"100010100",
  62912=>"110111111",
  62913=>"111111111",
  62914=>"000000000",
  62915=>"011111111",
  62916=>"000000001",
  62917=>"111111111",
  62918=>"100000001",
  62919=>"001000110",
  62920=>"011001001",
  62921=>"111111110",
  62922=>"001111011",
  62923=>"000000000",
  62924=>"111000000",
  62925=>"000000000",
  62926=>"111110011",
  62927=>"100111101",
  62928=>"000000000",
  62929=>"011011001",
  62930=>"111111111",
  62931=>"001000000",
  62932=>"000000000",
  62933=>"000011111",
  62934=>"111111111",
  62935=>"111011001",
  62936=>"000000000",
  62937=>"001011111",
  62938=>"111111111",
  62939=>"000000000",
  62940=>"000111111",
  62941=>"000000000",
  62942=>"000100110",
  62943=>"110110101",
  62944=>"001001011",
  62945=>"111111111",
  62946=>"000100110",
  62947=>"101111001",
  62948=>"000010100",
  62949=>"101111111",
  62950=>"000011110",
  62951=>"001000011",
  62952=>"111110111",
  62953=>"111011011",
  62954=>"000110111",
  62955=>"111111111",
  62956=>"011000100",
  62957=>"111111111",
  62958=>"110000110",
  62959=>"000000000",
  62960=>"111011001",
  62961=>"111111001",
  62962=>"000000000",
  62963=>"011111111",
  62964=>"000010010",
  62965=>"000001011",
  62966=>"101111111",
  62967=>"101101001",
  62968=>"111111111",
  62969=>"100000100",
  62970=>"001000000",
  62971=>"000000000",
  62972=>"110111111",
  62973=>"100111111",
  62974=>"110110110",
  62975=>"011111111",
  62976=>"111111110",
  62977=>"010111111",
  62978=>"111111111",
  62979=>"010100111",
  62980=>"011111111",
  62981=>"010110100",
  62982=>"011011001",
  62983=>"111111000",
  62984=>"000111111",
  62985=>"000000110",
  62986=>"000000000",
  62987=>"111001000",
  62988=>"000100100",
  62989=>"111000111",
  62990=>"000110000",
  62991=>"000000000",
  62992=>"100100000",
  62993=>"000110110",
  62994=>"000000111",
  62995=>"000000000",
  62996=>"000110111",
  62997=>"111110111",
  62998=>"110111111",
  62999=>"111111001",
  63000=>"101111110",
  63001=>"100111100",
  63002=>"111100000",
  63003=>"110100010",
  63004=>"000000000",
  63005=>"111111110",
  63006=>"011001000",
  63007=>"000000000",
  63008=>"000110111",
  63009=>"111111111",
  63010=>"100110111",
  63011=>"101000000",
  63012=>"010010011",
  63013=>"111000000",
  63014=>"111000000",
  63015=>"111010111",
  63016=>"000000000",
  63017=>"111111100",
  63018=>"110100100",
  63019=>"111111001",
  63020=>"001111111",
  63021=>"000101111",
  63022=>"111100100",
  63023=>"000000100",
  63024=>"000000000",
  63025=>"111010010",
  63026=>"000000101",
  63027=>"000000001",
  63028=>"111001000",
  63029=>"101100100",
  63030=>"000100000",
  63031=>"110111000",
  63032=>"000111111",
  63033=>"100000100",
  63034=>"011011011",
  63035=>"000110111",
  63036=>"111000000",
  63037=>"001000000",
  63038=>"111111111",
  63039=>"010000111",
  63040=>"111111101",
  63041=>"010000110",
  63042=>"111111000",
  63043=>"011111000",
  63044=>"000000110",
  63045=>"110111111",
  63046=>"111111000",
  63047=>"000000100",
  63048=>"111111111",
  63049=>"000001111",
  63050=>"111111111",
  63051=>"000110110",
  63052=>"000000000",
  63053=>"000000000",
  63054=>"110100100",
  63055=>"000000000",
  63056=>"011111001",
  63057=>"110100111",
  63058=>"111111010",
  63059=>"000001001",
  63060=>"111000000",
  63061=>"000000111",
  63062=>"000000000",
  63063=>"100011011",
  63064=>"001001000",
  63065=>"000000000",
  63066=>"000011000",
  63067=>"111000000",
  63068=>"000000000",
  63069=>"000000000",
  63070=>"011111111",
  63071=>"001000111",
  63072=>"000000000",
  63073=>"000000000",
  63074=>"000000111",
  63075=>"111111111",
  63076=>"000011111",
  63077=>"000000000",
  63078=>"011000000",
  63079=>"111111111",
  63080=>"000000110",
  63081=>"000000010",
  63082=>"111010100",
  63083=>"001011000",
  63084=>"111110000",
  63085=>"011000000",
  63086=>"111110110",
  63087=>"111111111",
  63088=>"111111110",
  63089=>"000010000",
  63090=>"111111011",
  63091=>"111111111",
  63092=>"111001000",
  63093=>"000110111",
  63094=>"000110111",
  63095=>"111000111",
  63096=>"110000100",
  63097=>"111010000",
  63098=>"111001000",
  63099=>"111111111",
  63100=>"101000000",
  63101=>"111111010",
  63102=>"111000011",
  63103=>"000000000",
  63104=>"000000111",
  63105=>"001000000",
  63106=>"011000010",
  63107=>"100100000",
  63108=>"111111010",
  63109=>"111101111",
  63110=>"001111111",
  63111=>"101101000",
  63112=>"111111111",
  63113=>"000111111",
  63114=>"000000111",
  63115=>"000000000",
  63116=>"111111000",
  63117=>"111111111",
  63118=>"110000000",
  63119=>"111000000",
  63120=>"001100111",
  63121=>"111111000",
  63122=>"000000110",
  63123=>"100000000",
  63124=>"111111111",
  63125=>"111111111",
  63126=>"110111111",
  63127=>"100100000",
  63128=>"111001001",
  63129=>"000000111",
  63130=>"110110111",
  63131=>"011000000",
  63132=>"111111111",
  63133=>"001000100",
  63134=>"111111111",
  63135=>"000000000",
  63136=>"011000010",
  63137=>"000110110",
  63138=>"100110000",
  63139=>"000000111",
  63140=>"000000000",
  63141=>"000000000",
  63142=>"111111000",
  63143=>"110111001",
  63144=>"111011111",
  63145=>"000000000",
  63146=>"000000111",
  63147=>"001111111",
  63148=>"111111111",
  63149=>"100001111",
  63150=>"000000110",
  63151=>"000110000",
  63152=>"111011001",
  63153=>"011011111",
  63154=>"010111010",
  63155=>"000000010",
  63156=>"111000100",
  63157=>"010110111",
  63158=>"000000011",
  63159=>"100001001",
  63160=>"000000011",
  63161=>"111111111",
  63162=>"111011011",
  63163=>"111000000",
  63164=>"000000110",
  63165=>"000000111",
  63166=>"000111111",
  63167=>"011000000",
  63168=>"000001000",
  63169=>"111011000",
  63170=>"111111111",
  63171=>"111111000",
  63172=>"000010010",
  63173=>"000011011",
  63174=>"000011001",
  63175=>"111111000",
  63176=>"111000000",
  63177=>"000110111",
  63178=>"111111001",
  63179=>"000000011",
  63180=>"110111111",
  63181=>"000100000",
  63182=>"000111111",
  63183=>"111000000",
  63184=>"000000001",
  63185=>"110010000",
  63186=>"111111111",
  63187=>"000000011",
  63188=>"110111111",
  63189=>"000000110",
  63190=>"000000000",
  63191=>"100001000",
  63192=>"111110000",
  63193=>"000010010",
  63194=>"011000111",
  63195=>"111111111",
  63196=>"000111111",
  63197=>"000000110",
  63198=>"000111000",
  63199=>"011111111",
  63200=>"000000000",
  63201=>"011111000",
  63202=>"111111000",
  63203=>"011111111",
  63204=>"011111111",
  63205=>"100000000",
  63206=>"000000000",
  63207=>"111100000",
  63208=>"000000000",
  63209=>"000011111",
  63210=>"000111111",
  63211=>"000000000",
  63212=>"000000011",
  63213=>"111111111",
  63214=>"111111111",
  63215=>"000000111",
  63216=>"101111101",
  63217=>"001011111",
  63218=>"100000001",
  63219=>"000000000",
  63220=>"000011111",
  63221=>"100000000",
  63222=>"111111111",
  63223=>"110110000",
  63224=>"000000000",
  63225=>"011000000",
  63226=>"000000000",
  63227=>"000011111",
  63228=>"111100110",
  63229=>"000000001",
  63230=>"011000000",
  63231=>"111100000",
  63232=>"010000111",
  63233=>"110110110",
  63234=>"111111000",
  63235=>"000110000",
  63236=>"111010000",
  63237=>"000000101",
  63238=>"100100111",
  63239=>"000111111",
  63240=>"111000000",
  63241=>"001011011",
  63242=>"110110000",
  63243=>"110111111",
  63244=>"110110000",
  63245=>"100000111",
  63246=>"111111000",
  63247=>"000000111",
  63248=>"000000111",
  63249=>"000000000",
  63250=>"000000110",
  63251=>"000001111",
  63252=>"111000001",
  63253=>"011111100",
  63254=>"110110000",
  63255=>"111111111",
  63256=>"001001000",
  63257=>"111111111",
  63258=>"001000000",
  63259=>"111111111",
  63260=>"000110111",
  63261=>"000011011",
  63262=>"111111101",
  63263=>"000000111",
  63264=>"100111111",
  63265=>"111111110",
  63266=>"011111111",
  63267=>"011000000",
  63268=>"111111100",
  63269=>"111000000",
  63270=>"111001001",
  63271=>"000000110",
  63272=>"111111111",
  63273=>"000000010",
  63274=>"000000111",
  63275=>"000111111",
  63276=>"001000000",
  63277=>"100001111",
  63278=>"010000111",
  63279=>"000000000",
  63280=>"111111000",
  63281=>"111111000",
  63282=>"000000011",
  63283=>"111011000",
  63284=>"000111111",
  63285=>"111000001",
  63286=>"111111000",
  63287=>"110110111",
  63288=>"110100000",
  63289=>"111111101",
  63290=>"010010010",
  63291=>"000000111",
  63292=>"000000110",
  63293=>"000000000",
  63294=>"100101111",
  63295=>"000000000",
  63296=>"111100000",
  63297=>"000000000",
  63298=>"111101001",
  63299=>"000000111",
  63300=>"000000000",
  63301=>"000000001",
  63302=>"000001001",
  63303=>"111111000",
  63304=>"111000000",
  63305=>"110111111",
  63306=>"111000000",
  63307=>"111111100",
  63308=>"000000000",
  63309=>"010000000",
  63310=>"110000000",
  63311=>"011011000",
  63312=>"001001111",
  63313=>"000000010",
  63314=>"111010000",
  63315=>"000000000",
  63316=>"000000000",
  63317=>"011011001",
  63318=>"000000000",
  63319=>"111111000",
  63320=>"111011000",
  63321=>"000000000",
  63322=>"110111010",
  63323=>"011000000",
  63324=>"110000000",
  63325=>"000000000",
  63326=>"000000000",
  63327=>"000010100",
  63328=>"010110110",
  63329=>"000000000",
  63330=>"100110111",
  63331=>"111000000",
  63332=>"000100111",
  63333=>"000000000",
  63334=>"111110000",
  63335=>"111111000",
  63336=>"110100000",
  63337=>"011001000",
  63338=>"001001100",
  63339=>"000110110",
  63340=>"001111111",
  63341=>"000001111",
  63342=>"000000111",
  63343=>"011000000",
  63344=>"111110000",
  63345=>"001111111",
  63346=>"110111111",
  63347=>"001001011",
  63348=>"111111111",
  63349=>"111100000",
  63350=>"111110100",
  63351=>"011000000",
  63352=>"001000000",
  63353=>"111111111",
  63354=>"111011000",
  63355=>"111100000",
  63356=>"111001011",
  63357=>"111000000",
  63358=>"000000011",
  63359=>"000111011",
  63360=>"111111000",
  63361=>"000000000",
  63362=>"111111011",
  63363=>"000000000",
  63364=>"000000000",
  63365=>"000001001",
  63366=>"000000100",
  63367=>"000111111",
  63368=>"010011000",
  63369=>"011011011",
  63370=>"011111011",
  63371=>"010111011",
  63372=>"000100111",
  63373=>"110110010",
  63374=>"000011001",
  63375=>"111000101",
  63376=>"111111000",
  63377=>"100110111",
  63378=>"111011000",
  63379=>"000000011",
  63380=>"110110100",
  63381=>"000001011",
  63382=>"000000000",
  63383=>"111100110",
  63384=>"000000110",
  63385=>"111001000",
  63386=>"110110111",
  63387=>"111001001",
  63388=>"000000111",
  63389=>"011111111",
  63390=>"000000000",
  63391=>"000000000",
  63392=>"111011001",
  63393=>"101100100",
  63394=>"000111011",
  63395=>"000011100",
  63396=>"111100111",
  63397=>"001111111",
  63398=>"111000000",
  63399=>"001000011",
  63400=>"100000000",
  63401=>"111101000",
  63402=>"000111111",
  63403=>"000110000",
  63404=>"000010000",
  63405=>"011000001",
  63406=>"011000000",
  63407=>"111111111",
  63408=>"000000111",
  63409=>"000000010",
  63410=>"011000000",
  63411=>"111001000",
  63412=>"111111000",
  63413=>"111111111",
  63414=>"111111000",
  63415=>"000000000",
  63416=>"111000000",
  63417=>"000111111",
  63418=>"111111111",
  63419=>"110111000",
  63420=>"111100001",
  63421=>"011011110",
  63422=>"000000000",
  63423=>"110000011",
  63424=>"000000111",
  63425=>"000000000",
  63426=>"111111000",
  63427=>"000000111",
  63428=>"111000111",
  63429=>"001001111",
  63430=>"000101010",
  63431=>"000000100",
  63432=>"110000001",
  63433=>"011000000",
  63434=>"000000000",
  63435=>"000000111",
  63436=>"000000000",
  63437=>"000000000",
  63438=>"100000000",
  63439=>"111111100",
  63440=>"111001001",
  63441=>"111111000",
  63442=>"111111000",
  63443=>"111110001",
  63444=>"001000000",
  63445=>"000111111",
  63446=>"011111000",
  63447=>"000011011",
  63448=>"111111111",
  63449=>"000000100",
  63450=>"000000000",
  63451=>"011000000",
  63452=>"111011111",
  63453=>"000001000",
  63454=>"100100000",
  63455=>"011000011",
  63456=>"011110000",
  63457=>"111111000",
  63458=>"000000011",
  63459=>"100111110",
  63460=>"111000000",
  63461=>"000110111",
  63462=>"000000000",
  63463=>"000000111",
  63464=>"111111111",
  63465=>"110000000",
  63466=>"111100100",
  63467=>"000000000",
  63468=>"111101111",
  63469=>"000000110",
  63470=>"000110101",
  63471=>"111000000",
  63472=>"000000111",
  63473=>"110100010",
  63474=>"101100111",
  63475=>"011011000",
  63476=>"111011111",
  63477=>"111111000",
  63478=>"111111000",
  63479=>"000001000",
  63480=>"001000000",
  63481=>"011001000",
  63482=>"110111111",
  63483=>"111111111",
  63484=>"100111111",
  63485=>"111100100",
  63486=>"111110010",
  63487=>"111000000",
  63488=>"001111100",
  63489=>"000000000",
  63490=>"101000110",
  63491=>"000000100",
  63492=>"001000111",
  63493=>"001111111",
  63494=>"000000000",
  63495=>"111100000",
  63496=>"111111001",
  63497=>"111111000",
  63498=>"000000000",
  63499=>"111111111",
  63500=>"000000000",
  63501=>"111100010",
  63502=>"111111000",
  63503=>"001111111",
  63504=>"010110111",
  63505=>"111111111",
  63506=>"111111111",
  63507=>"110110110",
  63508=>"000000000",
  63509=>"111000000",
  63510=>"000000010",
  63511=>"000000001",
  63512=>"110111111",
  63513=>"111111111",
  63514=>"000111111",
  63515=>"000011011",
  63516=>"011111000",
  63517=>"000000111",
  63518=>"111111111",
  63519=>"100000010",
  63520=>"000000000",
  63521=>"110110000",
  63522=>"111111111",
  63523=>"000000000",
  63524=>"111111111",
  63525=>"011000000",
  63526=>"011111011",
  63527=>"100001000",
  63528=>"111111001",
  63529=>"111111111",
  63530=>"111111111",
  63531=>"001001111",
  63532=>"111111111",
  63533=>"011111111",
  63534=>"000000101",
  63535=>"000100110",
  63536=>"000110000",
  63537=>"111111111",
  63538=>"111011011",
  63539=>"111111111",
  63540=>"000000111",
  63541=>"111011111",
  63542=>"101000111",
  63543=>"101001001",
  63544=>"111000000",
  63545=>"101110110",
  63546=>"000000000",
  63547=>"000000010",
  63548=>"000000101",
  63549=>"000001001",
  63550=>"110010000",
  63551=>"001000000",
  63552=>"111011000",
  63553=>"000010010",
  63554=>"111101000",
  63555=>"111111111",
  63556=>"111111111",
  63557=>"001001111",
  63558=>"111111000",
  63559=>"000111111",
  63560=>"000000010",
  63561=>"100100111",
  63562=>"111110000",
  63563=>"111000000",
  63564=>"111111000",
  63565=>"101000001",
  63566=>"011111000",
  63567=>"000001111",
  63568=>"000000000",
  63569=>"001111011",
  63570=>"010000000",
  63571=>"110010110",
  63572=>"001001111",
  63573=>"110000110",
  63574=>"101101000",
  63575=>"000000000",
  63576=>"000101110",
  63577=>"111111111",
  63578=>"000000000",
  63579=>"100100000",
  63580=>"000000000",
  63581=>"111111000",
  63582=>"111111111",
  63583=>"000110100",
  63584=>"111111000",
  63585=>"111100100",
  63586=>"011111111",
  63587=>"000000000",
  63588=>"010000001",
  63589=>"000000100",
  63590=>"000000000",
  63591=>"111111111",
  63592=>"100000110",
  63593=>"111110000",
  63594=>"000000010",
  63595=>"000111111",
  63596=>"101001000",
  63597=>"100100000",
  63598=>"111111000",
  63599=>"111001001",
  63600=>"000011011",
  63601=>"011011110",
  63602=>"001111110",
  63603=>"000100111",
  63604=>"001001011",
  63605=>"111111111",
  63606=>"000000000",
  63607=>"011001111",
  63608=>"000000000",
  63609=>"000000000",
  63610=>"111101000",
  63611=>"000000000",
  63612=>"111111111",
  63613=>"111000000",
  63614=>"000000000",
  63615=>"111100000",
  63616=>"110110110",
  63617=>"101100111",
  63618=>"000000000",
  63619=>"000100110",
  63620=>"111111100",
  63621=>"111111110",
  63622=>"000011111",
  63623=>"000111111",
  63624=>"000010110",
  63625=>"001001000",
  63626=>"000000000",
  63627=>"000000000",
  63628=>"111111111",
  63629=>"001000011",
  63630=>"111000000",
  63631=>"001000000",
  63632=>"111110000",
  63633=>"000000000",
  63634=>"111110000",
  63635=>"000000000",
  63636=>"001000110",
  63637=>"001100110",
  63638=>"110101001",
  63639=>"110110111",
  63640=>"100111100",
  63641=>"111100000",
  63642=>"000111111",
  63643=>"000000000",
  63644=>"111100111",
  63645=>"011111111",
  63646=>"111100001",
  63647=>"000111111",
  63648=>"111111001",
  63649=>"110000000",
  63650=>"000000000",
  63651=>"100000100",
  63652=>"111001111",
  63653=>"101000111",
  63654=>"111111111",
  63655=>"001101111",
  63656=>"100101000",
  63657=>"111111111",
  63658=>"111111111",
  63659=>"111001000",
  63660=>"000000000",
  63661=>"111111110",
  63662=>"001100111",
  63663=>"000010111",
  63664=>"111111111",
  63665=>"111000100",
  63666=>"001001001",
  63667=>"000000101",
  63668=>"010010000",
  63669=>"110000000",
  63670=>"001000000",
  63671=>"011000000",
  63672=>"000011111",
  63673=>"000000000",
  63674=>"111101101",
  63675=>"000111011",
  63676=>"000000000",
  63677=>"111011000",
  63678=>"000100111",
  63679=>"101101100",
  63680=>"111111010",
  63681=>"111110000",
  63682=>"001001001",
  63683=>"111111111",
  63684=>"111111000",
  63685=>"011000000",
  63686=>"000000000",
  63687=>"111110111",
  63688=>"000110111",
  63689=>"111111110",
  63690=>"011110100",
  63691=>"111111110",
  63692=>"100100000",
  63693=>"111101111",
  63694=>"000100000",
  63695=>"111001000",
  63696=>"000011111",
  63697=>"111111011",
  63698=>"111111111",
  63699=>"111000000",
  63700=>"101001111",
  63701=>"000000111",
  63702=>"111000000",
  63703=>"000110010",
  63704=>"100000000",
  63705=>"111111001",
  63706=>"000000000",
  63707=>"111111110",
  63708=>"100000011",
  63709=>"000000100",
  63710=>"001000000",
  63711=>"111111111",
  63712=>"000000000",
  63713=>"011111111",
  63714=>"111111111",
  63715=>"100000000",
  63716=>"001000100",
  63717=>"001000000",
  63718=>"111000000",
  63719=>"011111101",
  63720=>"111111111",
  63721=>"111111100",
  63722=>"111111111",
  63723=>"111110010",
  63724=>"000110111",
  63725=>"000010110",
  63726=>"111111111",
  63727=>"111011000",
  63728=>"011011000",
  63729=>"000000000",
  63730=>"000000001",
  63731=>"000110111",
  63732=>"111111111",
  63733=>"000010010",
  63734=>"111111011",
  63735=>"111111111",
  63736=>"111110000",
  63737=>"001001011",
  63738=>"111111111",
  63739=>"111111111",
  63740=>"100110000",
  63741=>"000000110",
  63742=>"101000000",
  63743=>"001101100",
  63744=>"001001000",
  63745=>"000010000",
  63746=>"111111111",
  63747=>"111110000",
  63748=>"000000000",
  63749=>"001000000",
  63750=>"000000111",
  63751=>"010000001",
  63752=>"101111110",
  63753=>"000000000",
  63754=>"000000010",
  63755=>"001111111",
  63756=>"100000000",
  63757=>"000000000",
  63758=>"100100000",
  63759=>"000111001",
  63760=>"110110100",
  63761=>"000000001",
  63762=>"000000000",
  63763=>"011111111",
  63764=>"110110110",
  63765=>"000000000",
  63766=>"000100110",
  63767=>"000001011",
  63768=>"001111111",
  63769=>"111111111",
  63770=>"000000000",
  63771=>"111111111",
  63772=>"111001000",
  63773=>"111111011",
  63774=>"111111111",
  63775=>"111010000",
  63776=>"110111111",
  63777=>"101101000",
  63778=>"101101111",
  63779=>"000111110",
  63780=>"000000000",
  63781=>"000000001",
  63782=>"000000011",
  63783=>"000000111",
  63784=>"010010010",
  63785=>"001001001",
  63786=>"001000000",
  63787=>"000011111",
  63788=>"000000000",
  63789=>"000000000",
  63790=>"000100000",
  63791=>"111110110",
  63792=>"111001001",
  63793=>"001001111",
  63794=>"000000111",
  63795=>"011000000",
  63796=>"110111111",
  63797=>"111111011",
  63798=>"111000000",
  63799=>"011000000",
  63800=>"000000000",
  63801=>"111110110",
  63802=>"111111001",
  63803=>"110000000",
  63804=>"000000000",
  63805=>"000000000",
  63806=>"111111111",
  63807=>"000000000",
  63808=>"000000000",
  63809=>"111111111",
  63810=>"000000011",
  63811=>"000000000",
  63812=>"000111011",
  63813=>"000000000",
  63814=>"110000000",
  63815=>"110110110",
  63816=>"000000000",
  63817=>"000000000",
  63818=>"110000000",
  63819=>"011010000",
  63820=>"000110110",
  63821=>"100000000",
  63822=>"101111111",
  63823=>"000000111",
  63824=>"001000100",
  63825=>"000000001",
  63826=>"100100000",
  63827=>"111111111",
  63828=>"001101101",
  63829=>"111111111",
  63830=>"111100000",
  63831=>"000110111",
  63832=>"001001011",
  63833=>"000000000",
  63834=>"111111000",
  63835=>"101001000",
  63836=>"001111000",
  63837=>"111111111",
  63838=>"111000000",
  63839=>"110110011",
  63840=>"111100001",
  63841=>"001000100",
  63842=>"111000001",
  63843=>"010000000",
  63844=>"001011111",
  63845=>"001011011",
  63846=>"000000110",
  63847=>"000000000",
  63848=>"001000000",
  63849=>"010111111",
  63850=>"111111101",
  63851=>"011111111",
  63852=>"001111001",
  63853=>"110000000",
  63854=>"111000000",
  63855=>"000000000",
  63856=>"110110010",
  63857=>"111000000",
  63858=>"000011000",
  63859=>"110110110",
  63860=>"111111001",
  63861=>"001011110",
  63862=>"001111001",
  63863=>"100100111",
  63864=>"111111111",
  63865=>"111111000",
  63866=>"000001111",
  63867=>"111000111",
  63868=>"110110111",
  63869=>"000000000",
  63870=>"001000000",
  63871=>"000000111",
  63872=>"011011011",
  63873=>"111111110",
  63874=>"110110111",
  63875=>"000000000",
  63876=>"100000000",
  63877=>"010011010",
  63878=>"000000000",
  63879=>"000010000",
  63880=>"000000000",
  63881=>"011010110",
  63882=>"111111100",
  63883=>"111111111",
  63884=>"000111111",
  63885=>"000100111",
  63886=>"000000000",
  63887=>"000000010",
  63888=>"000000000",
  63889=>"001000000",
  63890=>"010110111",
  63891=>"001001101",
  63892=>"111111111",
  63893=>"000000000",
  63894=>"111111111",
  63895=>"111111111",
  63896=>"011111111",
  63897=>"111111110",
  63898=>"011111000",
  63899=>"101101111",
  63900=>"111100000",
  63901=>"111101000",
  63902=>"001011111",
  63903=>"100111111",
  63904=>"111101011",
  63905=>"011111000",
  63906=>"001001000",
  63907=>"110110000",
  63908=>"000110100",
  63909=>"000000000",
  63910=>"111111000",
  63911=>"000100000",
  63912=>"011111010",
  63913=>"011000001",
  63914=>"110111111",
  63915=>"111111111",
  63916=>"000000111",
  63917=>"100110000",
  63918=>"111110100",
  63919=>"101000111",
  63920=>"000000000",
  63921=>"111000110",
  63922=>"111110111",
  63923=>"001000000",
  63924=>"111111000",
  63925=>"000000001",
  63926=>"011111111",
  63927=>"010010100",
  63928=>"000100000",
  63929=>"001111111",
  63930=>"000000001",
  63931=>"100100100",
  63932=>"000000000",
  63933=>"111111011",
  63934=>"000000000",
  63935=>"000000010",
  63936=>"111111100",
  63937=>"000000000",
  63938=>"111111111",
  63939=>"000000000",
  63940=>"110110111",
  63941=>"111110100",
  63942=>"101111111",
  63943=>"111111111",
  63944=>"000000101",
  63945=>"000000000",
  63946=>"000010000",
  63947=>"110110000",
  63948=>"000000000",
  63949=>"111111111",
  63950=>"000000000",
  63951=>"000000000",
  63952=>"000000000",
  63953=>"110100110",
  63954=>"000000000",
  63955=>"111010000",
  63956=>"111111111",
  63957=>"111111111",
  63958=>"000000000",
  63959=>"100010111",
  63960=>"000001000",
  63961=>"111001001",
  63962=>"000010000",
  63963=>"111111111",
  63964=>"111111011",
  63965=>"111110111",
  63966=>"000000000",
  63967=>"110100110",
  63968=>"000000011",
  63969=>"111000000",
  63970=>"001111010",
  63971=>"000000011",
  63972=>"000000010",
  63973=>"000111111",
  63974=>"011011001",
  63975=>"000000000",
  63976=>"011111000",
  63977=>"111000010",
  63978=>"011010000",
  63979=>"111111111",
  63980=>"111111001",
  63981=>"101101111",
  63982=>"000000000",
  63983=>"111110100",
  63984=>"111111111",
  63985=>"111000000",
  63986=>"011011111",
  63987=>"000000000",
  63988=>"111111010",
  63989=>"001001000",
  63990=>"111111111",
  63991=>"111000000",
  63992=>"010011111",
  63993=>"001000110",
  63994=>"011010111",
  63995=>"111110000",
  63996=>"111111000",
  63997=>"111111110",
  63998=>"000000000",
  63999=>"000000000",
  64000=>"111111111",
  64001=>"000000111",
  64002=>"000000101",
  64003=>"100000000",
  64004=>"010010111",
  64005=>"000000001",
  64006=>"000000000",
  64007=>"100101001",
  64008=>"110011011",
  64009=>"000001111",
  64010=>"110000000",
  64011=>"111110111",
  64012=>"000000000",
  64013=>"111111111",
  64014=>"100100000",
  64015=>"111111111",
  64016=>"000000000",
  64017=>"000000000",
  64018=>"100000000",
  64019=>"000000000",
  64020=>"111111111",
  64021=>"000001011",
  64022=>"011111111",
  64023=>"110111111",
  64024=>"111111111",
  64025=>"000011011",
  64026=>"111111111",
  64027=>"001000000",
  64028=>"001011111",
  64029=>"111111111",
  64030=>"000000000",
  64031=>"011100110",
  64032=>"100000000",
  64033=>"000100100",
  64034=>"001000000",
  64035=>"111111111",
  64036=>"001000000",
  64037=>"100100100",
  64038=>"111101111",
  64039=>"110100111",
  64040=>"000100111",
  64041=>"000000000",
  64042=>"000000000",
  64043=>"000000000",
  64044=>"111111111",
  64045=>"111111001",
  64046=>"000000000",
  64047=>"001000011",
  64048=>"111111111",
  64049=>"111011011",
  64050=>"001011011",
  64051=>"000000000",
  64052=>"001001001",
  64053=>"000000000",
  64054=>"111110111",
  64055=>"100100111",
  64056=>"000000001",
  64057=>"000000110",
  64058=>"000000000",
  64059=>"000000000",
  64060=>"100100111",
  64061=>"111010000",
  64062=>"101000111",
  64063=>"111111000",
  64064=>"011111010",
  64065=>"101100100",
  64066=>"111110110",
  64067=>"011111011",
  64068=>"000000100",
  64069=>"111111011",
  64070=>"110000000",
  64071=>"111111111",
  64072=>"000000000",
  64073=>"111111111",
  64074=>"000000000",
  64075=>"011111100",
  64076=>"111011000",
  64077=>"100110000",
  64078=>"000000001",
  64079=>"000011111",
  64080=>"111011111",
  64081=>"001001000",
  64082=>"111111111",
  64083=>"000000000",
  64084=>"000000000",
  64085=>"111111100",
  64086=>"111001011",
  64087=>"101111111",
  64088=>"111111111",
  64089=>"101000000",
  64090=>"111111001",
  64091=>"000000000",
  64092=>"111011011",
  64093=>"000000000",
  64094=>"110110111",
  64095=>"111111111",
  64096=>"000000000",
  64097=>"110111000",
  64098=>"000000000",
  64099=>"000000111",
  64100=>"000000111",
  64101=>"111111011",
  64102=>"011111111",
  64103=>"011000000",
  64104=>"110000000",
  64105=>"111000000",
  64106=>"000101001",
  64107=>"111110000",
  64108=>"001011110",
  64109=>"000000010",
  64110=>"111111111",
  64111=>"111111111",
  64112=>"111111111",
  64113=>"001111000",
  64114=>"001001001",
  64115=>"110111111",
  64116=>"000000000",
  64117=>"000000000",
  64118=>"111111011",
  64119=>"001000000",
  64120=>"100000100",
  64121=>"010110000",
  64122=>"011000000",
  64123=>"000000000",
  64124=>"110110110",
  64125=>"001000000",
  64126=>"000000000",
  64127=>"000000000",
  64128=>"000101111",
  64129=>"010000010",
  64130=>"101011111",
  64131=>"000011000",
  64132=>"011011110",
  64133=>"111111100",
  64134=>"111110111",
  64135=>"111011011",
  64136=>"000000000",
  64137=>"111111111",
  64138=>"111001111",
  64139=>"011111111",
  64140=>"000000111",
  64141=>"111000000",
  64142=>"011111111",
  64143=>"011111111",
  64144=>"000000000",
  64145=>"000000000",
  64146=>"001011011",
  64147=>"111111111",
  64148=>"100011111",
  64149=>"001100110",
  64150=>"101101000",
  64151=>"111111111",
  64152=>"111111000",
  64153=>"000000000",
  64154=>"001000000",
  64155=>"111111011",
  64156=>"111111000",
  64157=>"010110110",
  64158=>"111111111",
  64159=>"111111111",
  64160=>"001000000",
  64161=>"000000000",
  64162=>"000000000",
  64163=>"000000110",
  64164=>"110000000",
  64165=>"001101111",
  64166=>"000000000",
  64167=>"100000000",
  64168=>"011111101",
  64169=>"000011111",
  64170=>"111111111",
  64171=>"001000000",
  64172=>"111111111",
  64173=>"111111111",
  64174=>"100100101",
  64175=>"000000111",
  64176=>"000111111",
  64177=>"000000010",
  64178=>"100000000",
  64179=>"111000000",
  64180=>"000000000",
  64181=>"001000111",
  64182=>"000000100",
  64183=>"111111001",
  64184=>"011101111",
  64185=>"000000000",
  64186=>"111100000",
  64187=>"100100100",
  64188=>"010000000",
  64189=>"000000000",
  64190=>"000000000",
  64191=>"000011010",
  64192=>"001000101",
  64193=>"010000000",
  64194=>"111111111",
  64195=>"111111111",
  64196=>"111101001",
  64197=>"111111111",
  64198=>"111111111",
  64199=>"011011111",
  64200=>"000010000",
  64201=>"000000100",
  64202=>"110100000",
  64203=>"000000000",
  64204=>"000000001",
  64205=>"000000000",
  64206=>"000001000",
  64207=>"111111010",
  64208=>"001000010",
  64209=>"001001111",
  64210=>"000101111",
  64211=>"000100100",
  64212=>"001000011",
  64213=>"000101000",
  64214=>"111111111",
  64215=>"101101111",
  64216=>"001000011",
  64217=>"111001000",
  64218=>"111000111",
  64219=>"001011011",
  64220=>"001100001",
  64221=>"000000000",
  64222=>"110111111",
  64223=>"100100101",
  64224=>"100000000",
  64225=>"000000000",
  64226=>"100111111",
  64227=>"111011011",
  64228=>"010010000",
  64229=>"000000111",
  64230=>"111110110",
  64231=>"110111110",
  64232=>"000001011",
  64233=>"000100000",
  64234=>"001001000",
  64235=>"000000000",
  64236=>"110000100",
  64237=>"111111111",
  64238=>"000111111",
  64239=>"111101111",
  64240=>"110111100",
  64241=>"110110100",
  64242=>"111111111",
  64243=>"110101101",
  64244=>"111111000",
  64245=>"111111011",
  64246=>"000000000",
  64247=>"111111111",
  64248=>"111111111",
  64249=>"111111111",
  64250=>"111011011",
  64251=>"001001001",
  64252=>"000001001",
  64253=>"000000001",
  64254=>"000000000",
  64255=>"111011111",
  64256=>"100000000",
  64257=>"111000000",
  64258=>"000100110",
  64259=>"111111100",
  64260=>"010000000",
  64261=>"000000000",
  64262=>"000000000",
  64263=>"001001011",
  64264=>"011111100",
  64265=>"000000000",
  64266=>"111110110",
  64267=>"111111111",
  64268=>"101101001",
  64269=>"111111011",
  64270=>"000000100",
  64271=>"001011011",
  64272=>"111111101",
  64273=>"100010000",
  64274=>"000000000",
  64275=>"111011001",
  64276=>"111100000",
  64277=>"111111110",
  64278=>"000000000",
  64279=>"001010110",
  64280=>"000000000",
  64281=>"000000100",
  64282=>"111000000",
  64283=>"001001111",
  64284=>"110111111",
  64285=>"111110000",
  64286=>"000100111",
  64287=>"000000111",
  64288=>"111000011",
  64289=>"111111111",
  64290=>"000000000",
  64291=>"100000000",
  64292=>"000000000",
  64293=>"000000000",
  64294=>"001011111",
  64295=>"001100000",
  64296=>"000000001",
  64297=>"111111111",
  64298=>"000000101",
  64299=>"111111111",
  64300=>"111111110",
  64301=>"000001000",
  64302=>"111000111",
  64303=>"111111000",
  64304=>"000000000",
  64305=>"010110000",
  64306=>"110111001",
  64307=>"000000000",
  64308=>"011011111",
  64309=>"000000000",
  64310=>"111001111",
  64311=>"111111111",
  64312=>"000000001",
  64313=>"111111111",
  64314=>"000000000",
  64315=>"100000111",
  64316=>"000000110",
  64317=>"000011111",
  64318=>"111011011",
  64319=>"111101111",
  64320=>"111111000",
  64321=>"111111000",
  64322=>"101101111",
  64323=>"111111111",
  64324=>"000000000",
  64325=>"000000010",
  64326=>"000000000",
  64327=>"001001011",
  64328=>"000000000",
  64329=>"111000111",
  64330=>"000110111",
  64331=>"000000100",
  64332=>"111100111",
  64333=>"000100000",
  64334=>"001011010",
  64335=>"001000000",
  64336=>"000000110",
  64337=>"000010011",
  64338=>"000000000",
  64339=>"000000000",
  64340=>"000000000",
  64341=>"011011011",
  64342=>"111111111",
  64343=>"011111111",
  64344=>"000100000",
  64345=>"111000000",
  64346=>"001111000",
  64347=>"000000001",
  64348=>"111111000",
  64349=>"111111111",
  64350=>"001101111",
  64351=>"001001000",
  64352=>"000000000",
  64353=>"001010010",
  64354=>"001000001",
  64355=>"111111111",
  64356=>"000000111",
  64357=>"110111111",
  64358=>"111111111",
  64359=>"100100101",
  64360=>"100100000",
  64361=>"000000000",
  64362=>"100111111",
  64363=>"111110100",
  64364=>"000000011",
  64365=>"111111111",
  64366=>"111111111",
  64367=>"000000111",
  64368=>"001111111",
  64369=>"011011111",
  64370=>"111100000",
  64371=>"000000000",
  64372=>"111100011",
  64373=>"000000000",
  64374=>"000111111",
  64375=>"000000000",
  64376=>"000000110",
  64377=>"000111000",
  64378=>"101101111",
  64379=>"111111111",
  64380=>"111111011",
  64381=>"111111111",
  64382=>"000101111",
  64383=>"110100100",
  64384=>"100000000",
  64385=>"011001001",
  64386=>"111111000",
  64387=>"111111111",
  64388=>"011110000",
  64389=>"111000000",
  64390=>"000000000",
  64391=>"000000000",
  64392=>"001001111",
  64393=>"100100110",
  64394=>"000000010",
  64395=>"000000000",
  64396=>"111111111",
  64397=>"000000000",
  64398=>"111111111",
  64399=>"000000000",
  64400=>"000000000",
  64401=>"111011010",
  64402=>"000001111",
  64403=>"000000000",
  64404=>"111111111",
  64405=>"000000000",
  64406=>"110000110",
  64407=>"111000011",
  64408=>"001001111",
  64409=>"011011000",
  64410=>"010010011",
  64411=>"000000000",
  64412=>"111111111",
  64413=>"011111111",
  64414=>"100111111",
  64415=>"000000000",
  64416=>"011011011",
  64417=>"111111111",
  64418=>"100101001",
  64419=>"111111111",
  64420=>"111111111",
  64421=>"111111111",
  64422=>"000000101",
  64423=>"011111111",
  64424=>"100000001",
  64425=>"101111111",
  64426=>"000000000",
  64427=>"101101111",
  64428=>"111101000",
  64429=>"111111111",
  64430=>"111000000",
  64431=>"000000000",
  64432=>"000000111",
  64433=>"000000000",
  64434=>"111111111",
  64435=>"111000000",
  64436=>"011011010",
  64437=>"101000000",
  64438=>"000100111",
  64439=>"111001000",
  64440=>"000000000",
  64441=>"000000000",
  64442=>"001000000",
  64443=>"000100000",
  64444=>"001001001",
  64445=>"111111111",
  64446=>"111001011",
  64447=>"000000000",
  64448=>"000010000",
  64449=>"111111111",
  64450=>"000000000",
  64451=>"111111111",
  64452=>"111001011",
  64453=>"010011011",
  64454=>"111111111",
  64455=>"111111111",
  64456=>"100000000",
  64457=>"111011010",
  64458=>"000000000",
  64459=>"111111111",
  64460=>"111111000",
  64461=>"111111111",
  64462=>"111000000",
  64463=>"000000000",
  64464=>"000001111",
  64465=>"111111111",
  64466=>"110000000",
  64467=>"000000000",
  64468=>"100000110",
  64469=>"111000000",
  64470=>"011111111",
  64471=>"100100000",
  64472=>"000111110",
  64473=>"111111111",
  64474=>"000000110",
  64475=>"000000011",
  64476=>"000100000",
  64477=>"111001101",
  64478=>"111111011",
  64479=>"000001001",
  64480=>"100000000",
  64481=>"111111111",
  64482=>"011011011",
  64483=>"101111111",
  64484=>"111111001",
  64485=>"111111001",
  64486=>"001001111",
  64487=>"111111111",
  64488=>"000000000",
  64489=>"100001001",
  64490=>"000000000",
  64491=>"111111011",
  64492=>"011000111",
  64493=>"011011011",
  64494=>"111111111",
  64495=>"000000101",
  64496=>"110111111",
  64497=>"000000000",
  64498=>"000000110",
  64499=>"001001111",
  64500=>"000000000",
  64501=>"110100000",
  64502=>"110111111",
  64503=>"100110110",
  64504=>"111111110",
  64505=>"000010011",
  64506=>"111111000",
  64507=>"000000000",
  64508=>"111011111",
  64509=>"000000100",
  64510=>"101001010",
  64511=>"000110111",
  64512=>"100110110",
  64513=>"000000000",
  64514=>"111101100",
  64515=>"001000001",
  64516=>"010111110",
  64517=>"101001000",
  64518=>"111111000",
  64519=>"001001001",
  64520=>"101001111",
  64521=>"110110000",
  64522=>"101000001",
  64523=>"100000000",
  64524=>"110110110",
  64525=>"011001100",
  64526=>"000000000",
  64527=>"111111110",
  64528=>"101100111",
  64529=>"010111011",
  64530=>"000000000",
  64531=>"000000000",
  64532=>"000000100",
  64533=>"111111110",
  64534=>"101111111",
  64535=>"100100110",
  64536=>"001000000",
  64537=>"001000001",
  64538=>"000000000",
  64539=>"111111101",
  64540=>"001000111",
  64541=>"110001000",
  64542=>"000000001",
  64543=>"001111110",
  64544=>"111111111",
  64545=>"000000111",
  64546=>"000011000",
  64547=>"101100111",
  64548=>"000110110",
  64549=>"111110000",
  64550=>"001001111",
  64551=>"000000110",
  64552=>"000011111",
  64553=>"000000000",
  64554=>"000000001",
  64555=>"111111111",
  64556=>"111111011",
  64557=>"111111000",
  64558=>"100000001",
  64559=>"000000000",
  64560=>"001000111",
  64561=>"010111010",
  64562=>"000000000",
  64563=>"000000111",
  64564=>"100000000",
  64565=>"110010010",
  64566=>"000000000",
  64567=>"110111001",
  64568=>"000011111",
  64569=>"111111111",
  64570=>"000111111",
  64571=>"000000000",
  64572=>"100000001",
  64573=>"010111010",
  64574=>"000100100",
  64575=>"000000101",
  64576=>"011011011",
  64577=>"100101111",
  64578=>"000000001",
  64579=>"001111111",
  64580=>"000000000",
  64581=>"000000100",
  64582=>"000000011",
  64583=>"000000000",
  64584=>"111111101",
  64585=>"001001101",
  64586=>"000000001",
  64587=>"000000000",
  64588=>"010111111",
  64589=>"100100000",
  64590=>"100000000",
  64591=>"101101101",
  64592=>"111111111",
  64593=>"111111111",
  64594=>"000000101",
  64595=>"110110010",
  64596=>"111000000",
  64597=>"000000000",
  64598=>"010000011",
  64599=>"000000100",
  64600=>"000001001",
  64601=>"101100101",
  64602=>"010010011",
  64603=>"110110111",
  64604=>"011011011",
  64605=>"000000111",
  64606=>"000000111",
  64607=>"000011011",
  64608=>"100000000",
  64609=>"111011001",
  64610=>"010111110",
  64611=>"010000000",
  64612=>"110110000",
  64613=>"011000000",
  64614=>"111110000",
  64615=>"111000000",
  64616=>"100000110",
  64617=>"001000000",
  64618=>"011010111",
  64619=>"000000000",
  64620=>"000000001",
  64621=>"000001010",
  64622=>"000000000",
  64623=>"000011001",
  64624=>"111111111",
  64625=>"000000001",
  64626=>"011011110",
  64627=>"000111111",
  64628=>"000000000",
  64629=>"010110110",
  64630=>"111111101",
  64631=>"001111111",
  64632=>"000000011",
  64633=>"010110111",
  64634=>"111000000",
  64635=>"000000000",
  64636=>"101111101",
  64637=>"011001100",
  64638=>"000000000",
  64639=>"001011111",
  64640=>"100000101",
  64641=>"000000001",
  64642=>"000100000",
  64643=>"111111010",
  64644=>"011110010",
  64645=>"101000000",
  64646=>"000000111",
  64647=>"010000000",
  64648=>"111010111",
  64649=>"111100000",
  64650=>"111111111",
  64651=>"111111111",
  64652=>"000000000",
  64653=>"101000000",
  64654=>"110100101",
  64655=>"111111111",
  64656=>"000000001",
  64657=>"111000000",
  64658=>"000010111",
  64659=>"110000000",
  64660=>"000000110",
  64661=>"111011011",
  64662=>"000000000",
  64663=>"101000111",
  64664=>"101000000",
  64665=>"001000000",
  64666=>"110111111",
  64667=>"010000000",
  64668=>"111111100",
  64669=>"111111001",
  64670=>"000000000",
  64671=>"111110110",
  64672=>"011111111",
  64673=>"101100001",
  64674=>"011011001",
  64675=>"111111111",
  64676=>"000110011",
  64677=>"100111001",
  64678=>"101001101",
  64679=>"100111101",
  64680=>"000000101",
  64681=>"011000000",
  64682=>"000000000",
  64683=>"111100000",
  64684=>"000011111",
  64685=>"111100111",
  64686=>"000000000",
  64687=>"010100000",
  64688=>"110111001",
  64689=>"111111111",
  64690=>"111111111",
  64691=>"111111101",
  64692=>"110110000",
  64693=>"111111000",
  64694=>"000011111",
  64695=>"000000000",
  64696=>"100110111",
  64697=>"110111111",
  64698=>"001000000",
  64699=>"110110111",
  64700=>"000000000",
  64701=>"111110010",
  64702=>"101100000",
  64703=>"011111110",
  64704=>"100101111",
  64705=>"000000000",
  64706=>"000000000",
  64707=>"001000000",
  64708=>"100000101",
  64709=>"001001011",
  64710=>"000000111",
  64711=>"111111110",
  64712=>"010010111",
  64713=>"111111111",
  64714=>"111011011",
  64715=>"000101111",
  64716=>"111111100",
  64717=>"000001001",
  64718=>"000100110",
  64719=>"011011011",
  64720=>"011000000",
  64721=>"000000000",
  64722=>"011001001",
  64723=>"000000000",
  64724=>"111001000",
  64725=>"011111110",
  64726=>"000000000",
  64727=>"000000101",
  64728=>"000000000",
  64729=>"000000111",
  64730=>"111111101",
  64731=>"000000000",
  64732=>"111010001",
  64733=>"011000000",
  64734=>"111111111",
  64735=>"001011001",
  64736=>"111111111",
  64737=>"000000000",
  64738=>"001111111",
  64739=>"110111000",
  64740=>"000111000",
  64741=>"111111111",
  64742=>"000000000",
  64743=>"111110101",
  64744=>"111001000",
  64745=>"010111111",
  64746=>"001000001",
  64747=>"001111111",
  64748=>"100000000",
  64749=>"000101111",
  64750=>"100101111",
  64751=>"111111101",
  64752=>"100100100",
  64753=>"111111111",
  64754=>"000000010",
  64755=>"000010111",
  64756=>"111111111",
  64757=>"110110111",
  64758=>"000000000",
  64759=>"111111111",
  64760=>"111111111",
  64761=>"101111111",
  64762=>"000000000",
  64763=>"101000000",
  64764=>"011011011",
  64765=>"011010110",
  64766=>"111111111",
  64767=>"111111000",
  64768=>"111111011",
  64769=>"000000000",
  64770=>"000000000",
  64771=>"111111110",
  64772=>"000000000",
  64773=>"100110110",
  64774=>"111111111",
  64775=>"111011011",
  64776=>"001111111",
  64777=>"111100100",
  64778=>"111001101",
  64779=>"111111000",
  64780=>"101000111",
  64781=>"101100111",
  64782=>"110111111",
  64783=>"000000010",
  64784=>"111101100",
  64785=>"000000001",
  64786=>"100000111",
  64787=>"000000001",
  64788=>"000000110",
  64789=>"010111111",
  64790=>"001111001",
  64791=>"000000100",
  64792=>"111111110",
  64793=>"111111111",
  64794=>"100100000",
  64795=>"010010010",
  64796=>"000000111",
  64797=>"111111111",
  64798=>"000000000",
  64799=>"111111111",
  64800=>"000000000",
  64801=>"000011111",
  64802=>"111111111",
  64803=>"111111111",
  64804=>"110111011",
  64805=>"111111111",
  64806=>"011111111",
  64807=>"100111111",
  64808=>"111011011",
  64809=>"001000101",
  64810=>"010111010",
  64811=>"110000000",
  64812=>"110000000",
  64813=>"100111111",
  64814=>"001101101",
  64815=>"111110000",
  64816=>"110111110",
  64817=>"011111111",
  64818=>"000000000",
  64819=>"011000000",
  64820=>"000000000",
  64821=>"010011111",
  64822=>"100111111",
  64823=>"000000101",
  64824=>"110111110",
  64825=>"101000000",
  64826=>"101000000",
  64827=>"011000000",
  64828=>"000000000",
  64829=>"111111000",
  64830=>"000001000",
  64831=>"000000000",
  64832=>"011101000",
  64833=>"000000111",
  64834=>"111111010",
  64835=>"001101111",
  64836=>"000001111",
  64837=>"000000000",
  64838=>"000010010",
  64839=>"001001000",
  64840=>"000000000",
  64841=>"000000000",
  64842=>"010111111",
  64843=>"000000100",
  64844=>"001000000",
  64845=>"000000000",
  64846=>"000000101",
  64847=>"011011000",
  64848=>"011011110",
  64849=>"000100000",
  64850=>"000110110",
  64851=>"000011111",
  64852=>"001111111",
  64853=>"011011001",
  64854=>"010011000",
  64855=>"000101101",
  64856=>"111111100",
  64857=>"001000100",
  64858=>"111110010",
  64859=>"111001000",
  64860=>"111100000",
  64861=>"011111010",
  64862=>"000101111",
  64863=>"100000000",
  64864=>"111000000",
  64865=>"000000000",
  64866=>"000000000",
  64867=>"111111000",
  64868=>"000110110",
  64869=>"000000000",
  64870=>"001001101",
  64871=>"000000000",
  64872=>"001000111",
  64873=>"011000101",
  64874=>"110011010",
  64875=>"000111111",
  64876=>"110110110",
  64877=>"000000011",
  64878=>"001111111",
  64879=>"100000000",
  64880=>"000000001",
  64881=>"111111111",
  64882=>"111111010",
  64883=>"011011000",
  64884=>"000000001",
  64885=>"000000000",
  64886=>"000000101",
  64887=>"001111000",
  64888=>"100111001",
  64889=>"000000111",
  64890=>"111111111",
  64891=>"011011110",
  64892=>"000000001",
  64893=>"111111111",
  64894=>"000000111",
  64895=>"000100011",
  64896=>"110110110",
  64897=>"011011111",
  64898=>"100001011",
  64899=>"100100001",
  64900=>"011111111",
  64901=>"111101111",
  64902=>"111111111",
  64903=>"000000101",
  64904=>"101001000",
  64905=>"001000000",
  64906=>"000000000",
  64907=>"100110100",
  64908=>"111111001",
  64909=>"111111111",
  64910=>"111111010",
  64911=>"111111110",
  64912=>"000000000",
  64913=>"000000001",
  64914=>"110000011",
  64915=>"110000000",
  64916=>"111010011",
  64917=>"000111011",
  64918=>"000000001",
  64919=>"110000000",
  64920=>"001000000",
  64921=>"111000000",
  64922=>"000000000",
  64923=>"111111010",
  64924=>"000000000",
  64925=>"010011111",
  64926=>"111001001",
  64927=>"000000111",
  64928=>"000000000",
  64929=>"000101111",
  64930=>"111000000",
  64931=>"001101111",
  64932=>"111111110",
  64933=>"000111111",
  64934=>"000000101",
  64935=>"111111111",
  64936=>"111111111",
  64937=>"000000001",
  64938=>"111111111",
  64939=>"001000000",
  64940=>"000000000",
  64941=>"000000000",
  64942=>"111111000",
  64943=>"000000100",
  64944=>"010110111",
  64945=>"111011000",
  64946=>"000000110",
  64947=>"000000000",
  64948=>"001001101",
  64949=>"111111111",
  64950=>"000100101",
  64951=>"111111111",
  64952=>"000000000",
  64953=>"001000000",
  64954=>"000000000",
  64955=>"011111111",
  64956=>"000000010",
  64957=>"111111111",
  64958=>"111100000",
  64959=>"100000100",
  64960=>"000000101",
  64961=>"001111111",
  64962=>"000000000",
  64963=>"110110000",
  64964=>"111111011",
  64965=>"000110111",
  64966=>"010010010",
  64967=>"000000000",
  64968=>"111000000",
  64969=>"010111011",
  64970=>"101000101",
  64971=>"010000000",
  64972=>"000000000",
  64973=>"000110111",
  64974=>"110000010",
  64975=>"101000000",
  64976=>"111111000",
  64977=>"011011011",
  64978=>"000011011",
  64979=>"000000011",
  64980=>"111111001",
  64981=>"110111111",
  64982=>"010111100",
  64983=>"011011001",
  64984=>"101111111",
  64985=>"101101101",
  64986=>"001111111",
  64987=>"111011011",
  64988=>"111111100",
  64989=>"010001000",
  64990=>"000000001",
  64991=>"100100111",
  64992=>"010111000",
  64993=>"011001000",
  64994=>"101000000",
  64995=>"111111100",
  64996=>"111000000",
  64997=>"111111001",
  64998=>"000101111",
  64999=>"101111001",
  65000=>"000001000",
  65001=>"111011011",
  65002=>"111100101",
  65003=>"000100111",
  65004=>"111001000",
  65005=>"011011110",
  65006=>"111111111",
  65007=>"111000000",
  65008=>"000000000",
  65009=>"000011000",
  65010=>"011001000",
  65011=>"000000001",
  65012=>"000000001",
  65013=>"001000000",
  65014=>"011111111",
  65015=>"000000000",
  65016=>"011011110",
  65017=>"001000000",
  65018=>"010111010",
  65019=>"000000000",
  65020=>"000000000",
  65021=>"110111110",
  65022=>"111110000",
  65023=>"001001111",
  65024=>"001001001",
  65025=>"100111000",
  65026=>"000000000",
  65027=>"000000000",
  65028=>"000100000",
  65029=>"111011011",
  65030=>"000000111",
  65031=>"111111100",
  65032=>"010001000",
  65033=>"000100111",
  65034=>"111111110",
  65035=>"000100100",
  65036=>"001000100",
  65037=>"110110110",
  65038=>"000011111",
  65039=>"111000111",
  65040=>"111000000",
  65041=>"100100100",
  65042=>"001100000",
  65043=>"100000000",
  65044=>"011000000",
  65045=>"010010111",
  65046=>"011011111",
  65047=>"000001011",
  65048=>"000100111",
  65049=>"000100100",
  65050=>"010000011",
  65051=>"000000101",
  65052=>"000000010",
  65053=>"000111111",
  65054=>"001111111",
  65055=>"000000000",
  65056=>"010010001",
  65057=>"110110000",
  65058=>"111001000",
  65059=>"111010000",
  65060=>"000000000",
  65061=>"000000000",
  65062=>"011010011",
  65063=>"000000000",
  65064=>"111100111",
  65065=>"111111101",
  65066=>"010000000",
  65067=>"011001001",
  65068=>"011111110",
  65069=>"001000000",
  65070=>"000000000",
  65071=>"000000000",
  65072=>"000000000",
  65073=>"100111111",
  65074=>"001001001",
  65075=>"000000000",
  65076=>"110110110",
  65077=>"111111011",
  65078=>"101000000",
  65079=>"101011011",
  65080=>"001001111",
  65081=>"011111111",
  65082=>"000011110",
  65083=>"011111100",
  65084=>"000000000",
  65085=>"111101111",
  65086=>"111111111",
  65087=>"001001111",
  65088=>"000000000",
  65089=>"110000000",
  65090=>"110000000",
  65091=>"111111111",
  65092=>"111111111",
  65093=>"100000000",
  65094=>"100100000",
  65095=>"000000000",
  65096=>"111111011",
  65097=>"001000000",
  65098=>"111001000",
  65099=>"000000001",
  65100=>"111111111",
  65101=>"001011011",
  65102=>"010110100",
  65103=>"000000000",
  65104=>"111111000",
  65105=>"110110000",
  65106=>"010110111",
  65107=>"001001111",
  65108=>"000000000",
  65109=>"100001011",
  65110=>"101110100",
  65111=>"000000000",
  65112=>"100100000",
  65113=>"000000000",
  65114=>"111101001",
  65115=>"011000000",
  65116=>"011111111",
  65117=>"001001000",
  65118=>"011111111",
  65119=>"101100100",
  65120=>"000000110",
  65121=>"111100001",
  65122=>"110110111",
  65123=>"000010110",
  65124=>"100110100",
  65125=>"111100100",
  65126=>"100110000",
  65127=>"100000000",
  65128=>"001011000",
  65129=>"001001000",
  65130=>"111111110",
  65131=>"011011001",
  65132=>"001001000",
  65133=>"111001010",
  65134=>"011000000",
  65135=>"111001000",
  65136=>"000100110",
  65137=>"000011111",
  65138=>"011011111",
  65139=>"011111110",
  65140=>"111111001",
  65141=>"001111111",
  65142=>"111111111",
  65143=>"111111111",
  65144=>"011010100",
  65145=>"011111101",
  65146=>"001111110",
  65147=>"000000000",
  65148=>"000000000",
  65149=>"111100000",
  65150=>"110110111",
  65151=>"011011011",
  65152=>"100100100",
  65153=>"000000000",
  65154=>"111111000",
  65155=>"100110010",
  65156=>"111100111",
  65157=>"000000000",
  65158=>"100100000",
  65159=>"000000000",
  65160=>"000101000",
  65161=>"000000000",
  65162=>"000100100",
  65163=>"100111111",
  65164=>"111110000",
  65165=>"111111111",
  65166=>"100000011",
  65167=>"000000000",
  65168=>"111110000",
  65169=>"000100100",
  65170=>"011000000",
  65171=>"110000001",
  65172=>"010010000",
  65173=>"000010001",
  65174=>"111111010",
  65175=>"001000000",
  65176=>"111111111",
  65177=>"110100100",
  65178=>"111101111",
  65179=>"111111111",
  65180=>"011011011",
  65181=>"111011011",
  65182=>"001001001",
  65183=>"100000000",
  65184=>"011011111",
  65185=>"101110110",
  65186=>"001011111",
  65187=>"111100110",
  65188=>"011011001",
  65189=>"100101101",
  65190=>"111110000",
  65191=>"001000000",
  65192=>"011111111",
  65193=>"111111111",
  65194=>"000000000",
  65195=>"000000000",
  65196=>"111111110",
  65197=>"011011100",
  65198=>"111111101",
  65199=>"000000000",
  65200=>"111111111",
  65201=>"000110100",
  65202=>"111111011",
  65203=>"111111111",
  65204=>"111001001",
  65205=>"111011111",
  65206=>"000001111",
  65207=>"000000100",
  65208=>"000000000",
  65209=>"000000000",
  65210=>"011011001",
  65211=>"011011011",
  65212=>"001001001",
  65213=>"000000100",
  65214=>"000000001",
  65215=>"001001000",
  65216=>"000000000",
  65217=>"000110110",
  65218=>"111101111",
  65219=>"000111111",
  65220=>"111100000",
  65221=>"010000000",
  65222=>"010011100",
  65223=>"000100100",
  65224=>"110000000",
  65225=>"000111001",
  65226=>"001100001",
  65227=>"000100111",
  65228=>"001100000",
  65229=>"110011111",
  65230=>"011000000",
  65231=>"000000001",
  65232=>"110110010",
  65233=>"001111001",
  65234=>"100100000",
  65235=>"000000000",
  65236=>"111111000",
  65237=>"001001001",
  65238=>"011011000",
  65239=>"111111111",
  65240=>"001000100",
  65241=>"111100100",
  65242=>"000000000",
  65243=>"001000000",
  65244=>"001000001",
  65245=>"011011011",
  65246=>"111111000",
  65247=>"001000001",
  65248=>"000000000",
  65249=>"110010111",
  65250=>"000000000",
  65251=>"111100111",
  65252=>"011111111",
  65253=>"110110110",
  65254=>"001111111",
  65255=>"011111111",
  65256=>"100111111",
  65257=>"000000100",
  65258=>"101100101",
  65259=>"111000000",
  65260=>"000011001",
  65261=>"011110110",
  65262=>"111100100",
  65263=>"000000111",
  65264=>"100000000",
  65265=>"000000000",
  65266=>"010010110",
  65267=>"001001000",
  65268=>"111111001",
  65269=>"111011001",
  65270=>"100111111",
  65271=>"001011001",
  65272=>"000000000",
  65273=>"000000000",
  65274=>"100100001",
  65275=>"111010110",
  65276=>"010001001",
  65277=>"001001001",
  65278=>"011011011",
  65279=>"000000010",
  65280=>"001000000",
  65281=>"011000000",
  65282=>"001001001",
  65283=>"001111011",
  65284=>"001001111",
  65285=>"110010111",
  65286=>"000010000",
  65287=>"100000011",
  65288=>"111100100",
  65289=>"000000001",
  65290=>"101111111",
  65291=>"100110111",
  65292=>"001001101",
  65293=>"000001001",
  65294=>"111111111",
  65295=>"011011000",
  65296=>"011011001",
  65297=>"000111111",
  65298=>"000000111",
  65299=>"111010000",
  65300=>"111111111",
  65301=>"011010110",
  65302=>"100111110",
  65303=>"000010111",
  65304=>"000000101",
  65305=>"001010000",
  65306=>"000000001",
  65307=>"100110111",
  65308=>"000000000",
  65309=>"001111111",
  65310=>"111111001",
  65311=>"100100110",
  65312=>"011011000",
  65313=>"110110000",
  65314=>"000000000",
  65315=>"111001111",
  65316=>"110111011",
  65317=>"110110111",
  65318=>"111110001",
  65319=>"010101111",
  65320=>"100100000",
  65321=>"001001000",
  65322=>"001001001",
  65323=>"010010011",
  65324=>"000110111",
  65325=>"110100000",
  65326=>"110110000",
  65327=>"000000111",
  65328=>"000000001",
  65329=>"001000100",
  65330=>"000000000",
  65331=>"110110011",
  65332=>"110000000",
  65333=>"011000000",
  65334=>"011011001",
  65335=>"010010000",
  65336=>"000000000",
  65337=>"111001101",
  65338=>"010110111",
  65339=>"100111111",
  65340=>"111001001",
  65341=>"001000100",
  65342=>"001011000",
  65343=>"111101111",
  65344=>"000010111",
  65345=>"011011111",
  65346=>"100111111",
  65347=>"110110010",
  65348=>"000000110",
  65349=>"111100100",
  65350=>"000000000",
  65351=>"000101111",
  65352=>"111111111",
  65353=>"000000000",
  65354=>"001111000",
  65355=>"111111001",
  65356=>"011111011",
  65357=>"111001011",
  65358=>"111111111",
  65359=>"100101111",
  65360=>"101101101",
  65361=>"011000001",
  65362=>"100000000",
  65363=>"111011011",
  65364=>"100100100",
  65365=>"011011011",
  65366=>"000111011",
  65367=>"000000000",
  65368=>"111111111",
  65369=>"100000000",
  65370=>"000000000",
  65371=>"110100000",
  65372=>"110010111",
  65373=>"110110110",
  65374=>"010000000",
  65375=>"110111111",
  65376=>"111111111",
  65377=>"101001111",
  65378=>"100000101",
  65379=>"111101111",
  65380=>"111110100",
  65381=>"011111111",
  65382=>"000000000",
  65383=>"000111111",
  65384=>"001010000",
  65385=>"000010010",
  65386=>"000000000",
  65387=>"000000000",
  65388=>"111111100",
  65389=>"011010111",
  65390=>"010000000",
  65391=>"000000000",
  65392=>"111101001",
  65393=>"111110000",
  65394=>"111111111",
  65395=>"111111011",
  65396=>"001101101",
  65397=>"111111011",
  65398=>"001001111",
  65399=>"101001111",
  65400=>"001000000",
  65401=>"011111111",
  65402=>"000000000",
  65403=>"011011000",
  65404=>"011111110",
  65405=>"001011011",
  65406=>"000000000",
  65407=>"111110000",
  65408=>"000111111",
  65409=>"111110001",
  65410=>"001001000",
  65411=>"110100110",
  65412=>"011000000",
  65413=>"110110010",
  65414=>"111011011",
  65415=>"000001001",
  65416=>"000000000",
  65417=>"011111111",
  65418=>"001100100",
  65419=>"000000000",
  65420=>"101101111",
  65421=>"100000001",
  65422=>"111111111",
  65423=>"000000110",
  65424=>"100000000",
  65425=>"001000000",
  65426=>"000100100",
  65427=>"111011111",
  65428=>"000000011",
  65429=>"110010011",
  65430=>"110010000",
  65431=>"001001001",
  65432=>"110100100",
  65433=>"111111011",
  65434=>"000000000",
  65435=>"000000000",
  65436=>"000100111",
  65437=>"100100111",
  65438=>"011011011",
  65439=>"111111111",
  65440=>"111011011",
  65441=>"000000000",
  65442=>"000001001",
  65443=>"111001011",
  65444=>"000001001",
  65445=>"011000000",
  65446=>"000100001",
  65447=>"111110100",
  65448=>"100100110",
  65449=>"110111111",
  65450=>"101100101",
  65451=>"111000001",
  65452=>"000000000",
  65453=>"110100000",
  65454=>"001001010",
  65455=>"001100100",
  65456=>"011111010",
  65457=>"011011111",
  65458=>"000100111",
  65459=>"000001111",
  65460=>"000000000",
  65461=>"111111111",
  65462=>"111111001",
  65463=>"111111001",
  65464=>"001011001",
  65465=>"111111111",
  65466=>"011011001",
  65467=>"100100100",
  65468=>"110101000",
  65469=>"111100000",
  65470=>"011000000",
  65471=>"000010111",
  65472=>"111111110",
  65473=>"110111111",
  65474=>"000000000",
  65475=>"000000001",
  65476=>"111110011",
  65477=>"101101111",
  65478=>"111111011",
  65479=>"111111110",
  65480=>"001101101",
  65481=>"000000110",
  65482=>"010000010",
  65483=>"001001001",
  65484=>"110000000",
  65485=>"011101111",
  65486=>"100111011",
  65487=>"000011111",
  65488=>"000110111",
  65489=>"101111001",
  65490=>"111111111",
  65491=>"100000001",
  65492=>"111011111",
  65493=>"111111110",
  65494=>"001000000",
  65495=>"110100001",
  65496=>"000000000",
  65497=>"111110100",
  65498=>"110010000",
  65499=>"111111110",
  65500=>"000000100",
  65501=>"111111011",
  65502=>"000111101",
  65503=>"000000011",
  65504=>"110110110",
  65505=>"100110110",
  65506=>"111011111",
  65507=>"000000000",
  65508=>"111111110",
  65509=>"110000000",
  65510=>"110100000",
  65511=>"001000000",
  65512=>"000100111",
  65513=>"011011111",
  65514=>"000001111",
  65515=>"100111011",
  65516=>"100100000",
  65517=>"100100000",
  65518=>"111111111",
  65519=>"001000000",
  65520=>"100101111",
  65521=>"111100111",
  65522=>"100110100",
  65523=>"011000000",
  65524=>"001000000",
  65525=>"000011000",
  65526=>"001101111",
  65527=>"110111111",
  65528=>"010000000",
  65529=>"111101101",
  65530=>"111100100",
  65531=>"011010000",
  65532=>"000000000",
  65533=>"111011011",
  65534=>"000000110",
  65535=>"000000000");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;