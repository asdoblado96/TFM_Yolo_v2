LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L7_5_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(7) - 1 DOWNTO 0));
END L7_5_WROM;

ARCHITECTURE RTL OF L7_5_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"001001111",
  1=>"000000000",
  2=>"000000101",
  3=>"000000101",
  4=>"111001111",
  5=>"000000000",
  6=>"110111110",
  7=>"101100101",
  8=>"101111111",
  9=>"111011010",
  10=>"111111000",
  11=>"000000100",
  12=>"000000100",
  13=>"101001001",
  14=>"111100100",
  15=>"111111111",
  16=>"100000111",
  17=>"111111111",
  18=>"000010000",
  19=>"111111111",
  20=>"000001000",
  21=>"111110111",
  22=>"111111011",
  23=>"110000100",
  24=>"111101111",
  25=>"001001000",
  26=>"011111111",
  27=>"000000000",
  28=>"111001100",
  29=>"111111111",
  30=>"010110000",
  31=>"110010111",
  32=>"000001001",
  33=>"000001101",
  34=>"100010010",
  35=>"000000111",
  36=>"000111110",
  37=>"111001000",
  38=>"010010000",
  39=>"111111111",
  40=>"111001111",
  41=>"111001001",
  42=>"000000000",
  43=>"111111111",
  44=>"111111011",
  45=>"000010000",
  46=>"111111111",
  47=>"000000000",
  48=>"001000111",
  49=>"000010000",
  50=>"011011000",
  51=>"111000101",
  52=>"000000000",
  53=>"000000001",
  54=>"010000100",
  55=>"101001001",
  56=>"000000001",
  57=>"010000000",
  58=>"111111111",
  59=>"100000000",
  60=>"101111111",
  61=>"111011111",
  62=>"011111110",
  63=>"000000010",
  64=>"001001001",
  65=>"101100111",
  66=>"011111111",
  67=>"111111111",
  68=>"111011111",
  69=>"011111000",
  70=>"011000000",
  71=>"000000111",
  72=>"110100110",
  73=>"111111111",
  74=>"101000111",
  75=>"000000000",
  76=>"000000000",
  77=>"000000000",
  78=>"111000000",
  79=>"011111010",
  80=>"100111100",
  81=>"101101101",
  82=>"000001000",
  83=>"111111111",
  84=>"111000000",
  85=>"000000000",
  86=>"011011011",
  87=>"101000001",
  88=>"000000000",
  89=>"111111111",
  90=>"111111111",
  91=>"001001111",
  92=>"000011010",
  93=>"100110000",
  94=>"110111111",
  95=>"110000111",
  96=>"111111111",
  97=>"011000001",
  98=>"010010000",
  99=>"000000000",
  100=>"001000000",
  101=>"001000001",
  102=>"111110000",
  103=>"000000000",
  104=>"001000000",
  105=>"000000000",
  106=>"000101000",
  107=>"010000000",
  108=>"111001111",
  109=>"000000000",
  110=>"000000000",
  111=>"011001001",
  112=>"000000000",
  113=>"110010000",
  114=>"010111010",
  115=>"010000000",
  116=>"111111111",
  117=>"110000001",
  118=>"010010000",
  119=>"000000000",
  120=>"111111000",
  121=>"101111110",
  122=>"111111000",
  123=>"000110000",
  124=>"111111111",
  125=>"000000000",
  126=>"110000000",
  127=>"111111111",
  128=>"000000000",
  129=>"000000000",
  130=>"000000000",
  131=>"111000111",
  132=>"000000000",
  133=>"100000111",
  134=>"111111111",
  135=>"011111010",
  136=>"111111111",
  137=>"111101111",
  138=>"000111010",
  139=>"010000000",
  140=>"111110111",
  141=>"000000000",
  142=>"111011111",
  143=>"000000010",
  144=>"111111111",
  145=>"000010010",
  146=>"111111111",
  147=>"011000000",
  148=>"110000000",
  149=>"111100110",
  150=>"001001011",
  151=>"111111111",
  152=>"000111111",
  153=>"000001000",
  154=>"101000000",
  155=>"001111111",
  156=>"111100110",
  157=>"011010000",
  158=>"100000111",
  159=>"101000001",
  160=>"111110000",
  161=>"111000001",
  162=>"000000000",
  163=>"111111101",
  164=>"100100000",
  165=>"000100100",
  166=>"000000000",
  167=>"110100110",
  168=>"000000110",
  169=>"000010010",
  170=>"010111010",
  171=>"111111011",
  172=>"111101001",
  173=>"011001111",
  174=>"000000010",
  175=>"011000000",
  176=>"110010111",
  177=>"110000000",
  178=>"111111110",
  179=>"000000000",
  180=>"111101000",
  181=>"000111011",
  182=>"111001000",
  183=>"000000011",
  184=>"001000001",
  185=>"111111111",
  186=>"111111111",
  187=>"001001111",
  188=>"000111000",
  189=>"001000000",
  190=>"000000000",
  191=>"011000101",
  192=>"000000000",
  193=>"111101111",
  194=>"011111111",
  195=>"111111000",
  196=>"111111010",
  197=>"000010000",
  198=>"000000000",
  199=>"100111111",
  200=>"000000000",
  201=>"000000111",
  202=>"111000000",
  203=>"010000000",
  204=>"100000000",
  205=>"000000000",
  206=>"111111111",
  207=>"110111000",
  208=>"111011000",
  209=>"000000000",
  210=>"111000011",
  211=>"000001000",
  212=>"101111111",
  213=>"100110111",
  214=>"000000000",
  215=>"110100000",
  216=>"000000101",
  217=>"110111111",
  218=>"000000000",
  219=>"000010000",
  220=>"111111111",
  221=>"000000011",
  222=>"010000000",
  223=>"111001000",
  224=>"010111111",
  225=>"001000100",
  226=>"000110110",
  227=>"001011000",
  228=>"000000000",
  229=>"100100100",
  230=>"111111011",
  231=>"111011001",
  232=>"001001001",
  233=>"000000000",
  234=>"110000100",
  235=>"000000011",
  236=>"000000000",
  237=>"111111111",
  238=>"000000100",
  239=>"111111111",
  240=>"110010010",
  241=>"111011111",
  242=>"000000000",
  243=>"011011000",
  244=>"000100111",
  245=>"111001011",
  246=>"000000010",
  247=>"101001101",
  248=>"010000000",
  249=>"111111010",
  250=>"000000000",
  251=>"001101111",
  252=>"000001000",
  253=>"001001011",
  254=>"000110000",
  255=>"110110111",
  256=>"010111000",
  257=>"000001001",
  258=>"010111000",
  259=>"111010000",
  260=>"011111101",
  261=>"001001000",
  262=>"111100000",
  263=>"111111111",
  264=>"000000000",
  265=>"010111010",
  266=>"111111111",
  267=>"110111111",
  268=>"001000001",
  269=>"111111000",
  270=>"101000000",
  271=>"001101111",
  272=>"000000000",
  273=>"101000111",
  274=>"111101111",
  275=>"111111111",
  276=>"000000000",
  277=>"000000000",
  278=>"000001011",
  279=>"111000001",
  280=>"011011111",
  281=>"111111111",
  282=>"110000000",
  283=>"000000000",
  284=>"011001001",
  285=>"011011000",
  286=>"011011000",
  287=>"000011000",
  288=>"111101111",
  289=>"100110000",
  290=>"101111111",
  291=>"111000011",
  292=>"111100100",
  293=>"000000000",
  294=>"100001001",
  295=>"111111100",
  296=>"000000000",
  297=>"101000100",
  298=>"111111000",
  299=>"110111000",
  300=>"000010110",
  301=>"111011011",
  302=>"000000000",
  303=>"000111110",
  304=>"001000011",
  305=>"000000000",
  306=>"000000000",
  307=>"000000100",
  308=>"100000100",
  309=>"111111111",
  310=>"111111111",
  311=>"010111111",
  312=>"001000000",
  313=>"000000101",
  314=>"111111111",
  315=>"000000001",
  316=>"010011000",
  317=>"001001111",
  318=>"001101101",
  319=>"111011011",
  320=>"001000000",
  321=>"000000111",
  322=>"000000000",
  323=>"110000000",
  324=>"000101111",
  325=>"000101000",
  326=>"000110000",
  327=>"111010000",
  328=>"000000000",
  329=>"000000000",
  330=>"111101111",
  331=>"000000000",
  332=>"000000001",
  333=>"000000001",
  334=>"101001001",
  335=>"010000111",
  336=>"111011011",
  337=>"100100110",
  338=>"001000011",
  339=>"111000100",
  340=>"000000000",
  341=>"111000111",
  342=>"000000000",
  343=>"111111111",
  344=>"111111010",
  345=>"110111110",
  346=>"101111111",
  347=>"111111111",
  348=>"000000000",
  349=>"101000000",
  350=>"110001011",
  351=>"111111111",
  352=>"000000000",
  353=>"111111110",
  354=>"000000111",
  355=>"110111010",
  356=>"000000000",
  357=>"000000000",
  358=>"000000011",
  359=>"110100000",
  360=>"011000000",
  361=>"000000111",
  362=>"000000000",
  363=>"111111111",
  364=>"111011111",
  365=>"011000001",
  366=>"000111110",
  367=>"111111111",
  368=>"100000111",
  369=>"000000000",
  370=>"111111111",
  371=>"000000100",
  372=>"110110000",
  373=>"010010000",
  374=>"000000000",
  375=>"000000000",
  376=>"000111111",
  377=>"111111111",
  378=>"111111111",
  379=>"000000000",
  380=>"000000111",
  381=>"111001111",
  382=>"111000000",
  383=>"011111000",
  384=>"000000100",
  385=>"000000001",
  386=>"110111001",
  387=>"111111110",
  388=>"000110000",
  389=>"110111110",
  390=>"000000000",
  391=>"000110001",
  392=>"011111111",
  393=>"000000000",
  394=>"100000000",
  395=>"000000001",
  396=>"111111111",
  397=>"000000000",
  398=>"000000011",
  399=>"000000000",
  400=>"000000000",
  401=>"111111111",
  402=>"000001001",
  403=>"000010000",
  404=>"000000000",
  405=>"000000001",
  406=>"000000000",
  407=>"100000000",
  408=>"101100100",
  409=>"111010000",
  410=>"000000000",
  411=>"001000100",
  412=>"001111111",
  413=>"000000000",
  414=>"001011011",
  415=>"000000000",
  416=>"110000000",
  417=>"011000000",
  418=>"111111111",
  419=>"000111110",
  420=>"111101111",
  421=>"100100101",
  422=>"111111111",
  423=>"001000000",
  424=>"111111001",
  425=>"111111110",
  426=>"000000111",
  427=>"000000000",
  428=>"000010010",
  429=>"111000000",
  430=>"001100111",
  431=>"000101111",
  432=>"000000111",
  433=>"000000100",
  434=>"000000000",
  435=>"110001001",
  436=>"111101101",
  437=>"000000000",
  438=>"111000001",
  439=>"010000000",
  440=>"000000001",
  441=>"000000000",
  442=>"110100111",
  443=>"100001011",
  444=>"000000000",
  445=>"000000000",
  446=>"000110111",
  447=>"000111011",
  448=>"000101101",
  449=>"111111111",
  450=>"000000001",
  451=>"111111000",
  452=>"000000000",
  453=>"010011000",
  454=>"000010000",
  455=>"000011000",
  456=>"000011000",
  457=>"001001000",
  458=>"111110110",
  459=>"111001001",
  460=>"101101111",
  461=>"000000000",
  462=>"000000000",
  463=>"001001101",
  464=>"111111101",
  465=>"000000000",
  466=>"100110100",
  467=>"011111000",
  468=>"000000111",
  469=>"011010000",
  470=>"000000000",
  471=>"010000000",
  472=>"000000000",
  473=>"111000001",
  474=>"011000000",
  475=>"111000000",
  476=>"000000000",
  477=>"011000000",
  478=>"000000011",
  479=>"111010010",
  480=>"000000000",
  481=>"000010001",
  482=>"111111111",
  483=>"100000111",
  484=>"111000000",
  485=>"111101001",
  486=>"000000000",
  487=>"011111111",
  488=>"111001111",
  489=>"000000000",
  490=>"010000000",
  491=>"111000111",
  492=>"011000111",
  493=>"010000011",
  494=>"000000001",
  495=>"111101111",
  496=>"011111011",
  497=>"000000000",
  498=>"111101111",
  499=>"101101100",
  500=>"000000000",
  501=>"000000000",
  502=>"111000000",
  503=>"100000000",
  504=>"111111111",
  505=>"001111110",
  506=>"000010000",
  507=>"000011000",
  508=>"001001111",
  509=>"000000110",
  510=>"000000000",
  511=>"111111111",
  512=>"001001000",
  513=>"100000000",
  514=>"101000100",
  515=>"001000001",
  516=>"001001000",
  517=>"111111011",
  518=>"000000000",
  519=>"000000000",
  520=>"000000000",
  521=>"000111111",
  522=>"000000000",
  523=>"001000000",
  524=>"111000000",
  525=>"000000000",
  526=>"000000000",
  527=>"000000000",
  528=>"100100011",
  529=>"000001000",
  530=>"111011011",
  531=>"000000000",
  532=>"111111111",
  533=>"111111111",
  534=>"000010000",
  535=>"111111110",
  536=>"000011111",
  537=>"000000000",
  538=>"111111111",
  539=>"111111111",
  540=>"100110111",
  541=>"111100100",
  542=>"000000000",
  543=>"110110111",
  544=>"111001000",
  545=>"000101111",
  546=>"110100100",
  547=>"101000000",
  548=>"111111111",
  549=>"001001001",
  550=>"110111111",
  551=>"111111111",
  552=>"000000000",
  553=>"110000100",
  554=>"000000000",
  555=>"000000000",
  556=>"000000000",
  557=>"000000000",
  558=>"111111011",
  559=>"111110110",
  560=>"000100111",
  561=>"000000110",
  562=>"100100110",
  563=>"000001001",
  564=>"111111111",
  565=>"000000000",
  566=>"000000110",
  567=>"001111111",
  568=>"111111111",
  569=>"011000110",
  570=>"000000111",
  571=>"011111111",
  572=>"111000101",
  573=>"001011111",
  574=>"111111001",
  575=>"000000000",
  576=>"000000000",
  577=>"000010000",
  578=>"101000000",
  579=>"110110111",
  580=>"100100100",
  581=>"000000000",
  582=>"111010110",
  583=>"000000000",
  584=>"011011111",
  585=>"111111111",
  586=>"000000011",
  587=>"001011011",
  588=>"111111111",
  589=>"011011111",
  590=>"010011010",
  591=>"000010001",
  592=>"011000000",
  593=>"000000000",
  594=>"000000001",
  595=>"010000000",
  596=>"111111111",
  597=>"000000010",
  598=>"111111111",
  599=>"111100111",
  600=>"111111111",
  601=>"111101111",
  602=>"000100111",
  603=>"111111011",
  604=>"000000000",
  605=>"111111111",
  606=>"000000000",
  607=>"100100000",
  608=>"001111001",
  609=>"000000000",
  610=>"000101111",
  611=>"010100000",
  612=>"111000000",
  613=>"000000000",
  614=>"001000111",
  615=>"000000000",
  616=>"111001000",
  617=>"000000000",
  618=>"011011111",
  619=>"000111000",
  620=>"001111111",
  621=>"001111111",
  622=>"111100110",
  623=>"111110000",
  624=>"011000000",
  625=>"000010110",
  626=>"111111000",
  627=>"111110110",
  628=>"000000011",
  629=>"000000000",
  630=>"111111111",
  631=>"000001000",
  632=>"111110110",
  633=>"001000000",
  634=>"000000000",
  635=>"000000000",
  636=>"110110110",
  637=>"000000100",
  638=>"100000100",
  639=>"111111000",
  640=>"000000000",
  641=>"010010110",
  642=>"111111111",
  643=>"000000100",
  644=>"111111111",
  645=>"110000010",
  646=>"001011111",
  647=>"000000000",
  648=>"011000101",
  649=>"000000000",
  650=>"111111111",
  651=>"000000110",
  652=>"000011001",
  653=>"000000000",
  654=>"111011000",
  655=>"000000000",
  656=>"000000111",
  657=>"001001001",
  658=>"000000000",
  659=>"111111111",
  660=>"000000000",
  661=>"111100000",
  662=>"000011000",
  663=>"000000111",
  664=>"110101111",
  665=>"100111111",
  666=>"000000000",
  667=>"000111111",
  668=>"000000100",
  669=>"000010011",
  670=>"111100100",
  671=>"000000000",
  672=>"010110110",
  673=>"111111000",
  674=>"000110111",
  675=>"100110111",
  676=>"000000100",
  677=>"000000000",
  678=>"111111111",
  679=>"011011010",
  680=>"010111011",
  681=>"000000000",
  682=>"000000100",
  683=>"111111111",
  684=>"111111111",
  685=>"000000011",
  686=>"001111111",
  687=>"000000000",
  688=>"011011000",
  689=>"000010111",
  690=>"000011111",
  691=>"000000000",
  692=>"111000111",
  693=>"100110011",
  694=>"100111111",
  695=>"000101111",
  696=>"111000000",
  697=>"000000000",
  698=>"100100000",
  699=>"100000000",
  700=>"101111101",
  701=>"111100111",
  702=>"110111111",
  703=>"011000010",
  704=>"101100101",
  705=>"000000000",
  706=>"011111111",
  707=>"111111111",
  708=>"000111000",
  709=>"111111111",
  710=>"000111111",
  711=>"101111111",
  712=>"000000111",
  713=>"111000000",
  714=>"111000000",
  715=>"000011111",
  716=>"111111111",
  717=>"011111111",
  718=>"110111111",
  719=>"000000000",
  720=>"011001000",
  721=>"000000000",
  722=>"111000000",
  723=>"111000000",
  724=>"100000110",
  725=>"110010010",
  726=>"111111111",
  727=>"100000000",
  728=>"011000000",
  729=>"001111100",
  730=>"111110111",
  731=>"111111000",
  732=>"000000000",
  733=>"111111111",
  734=>"000001000",
  735=>"011111111",
  736=>"000000000",
  737=>"111110110",
  738=>"000011111",
  739=>"011111111",
  740=>"111111111",
  741=>"111111111",
  742=>"000000010",
  743=>"100111001",
  744=>"000000001",
  745=>"001111111",
  746=>"011011000",
  747=>"011010111",
  748=>"011001000",
  749=>"000111111",
  750=>"000111111",
  751=>"111111000",
  752=>"001001011",
  753=>"111111111",
  754=>"111110111",
  755=>"000010000",
  756=>"000000000",
  757=>"000000000",
  758=>"111111101",
  759=>"111111111",
  760=>"000000000",
  761=>"000000000",
  762=>"000000000",
  763=>"111011000",
  764=>"100000000",
  765=>"100000001",
  766=>"111010000",
  767=>"001001000",
  768=>"111111111",
  769=>"111111111",
  770=>"011111111",
  771=>"000000000",
  772=>"111000000",
  773=>"111111111",
  774=>"110111111",
  775=>"000010000",
  776=>"111111111",
  777=>"111111000",
  778=>"111111111",
  779=>"000000100",
  780=>"111100100",
  781=>"100000000",
  782=>"100111011",
  783=>"000001000",
  784=>"000000000",
  785=>"111111100",
  786=>"101001001",
  787=>"111111111",
  788=>"111111111",
  789=>"011110001",
  790=>"111111011",
  791=>"111111111",
  792=>"100110110",
  793=>"111111111",
  794=>"111000000",
  795=>"111111111",
  796=>"000000111",
  797=>"111111111",
  798=>"111111111",
  799=>"000000000",
  800=>"001000000",
  801=>"100000000",
  802=>"011000000",
  803=>"000000000",
  804=>"100100111",
  805=>"011000101",
  806=>"000000111",
  807=>"100100100",
  808=>"111111111",
  809=>"011010000",
  810=>"111111111",
  811=>"000111111",
  812=>"111111101",
  813=>"111111111",
  814=>"000000000",
  815=>"111111111",
  816=>"000000000",
  817=>"000000000",
  818=>"000000100",
  819=>"000000000",
  820=>"000000000",
  821=>"111000100",
  822=>"000000000",
  823=>"111111111",
  824=>"000000000",
  825=>"111000011",
  826=>"000000001",
  827=>"000000000",
  828=>"000100100",
  829=>"000000110",
  830=>"000000000",
  831=>"000000000",
  832=>"000100000",
  833=>"111111000",
  834=>"111111111",
  835=>"111111111",
  836=>"011001000",
  837=>"111111111",
  838=>"111100100",
  839=>"000000000",
  840=>"000000000",
  841=>"110110000",
  842=>"000000000",
  843=>"111111111",
  844=>"100000000",
  845=>"000100000",
  846=>"000000000",
  847=>"111111111",
  848=>"001000010",
  849=>"111110111",
  850=>"001000000",
  851=>"000000000",
  852=>"110110111",
  853=>"111111011",
  854=>"100000000",
  855=>"111111111",
  856=>"111111111",
  857=>"111111000",
  858=>"111111000",
  859=>"000101101",
  860=>"000000000",
  861=>"000001111",
  862=>"000000000",
  863=>"011111111",
  864=>"000000000",
  865=>"000000000",
  866=>"000000000",
  867=>"111111111",
  868=>"101111110",
  869=>"000010011",
  870=>"111111110",
  871=>"111011000",
  872=>"111111110",
  873=>"111000000",
  874=>"111111100",
  875=>"010010111",
  876=>"110110000",
  877=>"010110110",
  878=>"000000000",
  879=>"000000000",
  880=>"111000000",
  881=>"000000000",
  882=>"110111111",
  883=>"011011010",
  884=>"010000000",
  885=>"010000000",
  886=>"111011111",
  887=>"111111110",
  888=>"111111111",
  889=>"000111111",
  890=>"111111111",
  891=>"000000000",
  892=>"000000000",
  893=>"111111111",
  894=>"110000000",
  895=>"110111111",
  896=>"111111111",
  897=>"000000000",
  898=>"001011001",
  899=>"001101111",
  900=>"111011111",
  901=>"000000011",
  902=>"011111111",
  903=>"001001001",
  904=>"111111111",
  905=>"010110110",
  906=>"111111111",
  907=>"111111111",
  908=>"111111111",
  909=>"000111111",
  910=>"000000001",
  911=>"000000000",
  912=>"000000000",
  913=>"110110110",
  914=>"000001001",
  915=>"000011111",
  916=>"001000000",
  917=>"000000000",
  918=>"000000111",
  919=>"111010010",
  920=>"000001111",
  921=>"110111111",
  922=>"000100000",
  923=>"000000100",
  924=>"111111111",
  925=>"111111000",
  926=>"000000000",
  927=>"000000001",
  928=>"000110111",
  929=>"001001011",
  930=>"111111111",
  931=>"111110111",
  932=>"000000101",
  933=>"000000000",
  934=>"111111111",
  935=>"000111011",
  936=>"111111111",
  937=>"111011101",
  938=>"110000111",
  939=>"000000000",
  940=>"111111111",
  941=>"000000001",
  942=>"111011101",
  943=>"111111111",
  944=>"111111111",
  945=>"100100000",
  946=>"011001111",
  947=>"011000011",
  948=>"000000101",
  949=>"111100000",
  950=>"000000100",
  951=>"010101000",
  952=>"000010111",
  953=>"111011111",
  954=>"010000111",
  955=>"111111111",
  956=>"000000000",
  957=>"111111111",
  958=>"000000000",
  959=>"100100000",
  960=>"000000000",
  961=>"110110110",
  962=>"000000000",
  963=>"001000000",
  964=>"111111110",
  965=>"000000000",
  966=>"000000000",
  967=>"000000000",
  968=>"111110000",
  969=>"000000000",
  970=>"100100000",
  971=>"111111111",
  972=>"110011000",
  973=>"010010111",
  974=>"111000000",
  975=>"111111110",
  976=>"111110110",
  977=>"111111111",
  978=>"111111010",
  979=>"111111111",
  980=>"000000000",
  981=>"000000100",
  982=>"011101001",
  983=>"001000100",
  984=>"110100100",
  985=>"011011111",
  986=>"110110000",
  987=>"111111111",
  988=>"100100110",
  989=>"111111011",
  990=>"100110000",
  991=>"110100100",
  992=>"110111110",
  993=>"111111111",
  994=>"000111011",
  995=>"000000000",
  996=>"100100111",
  997=>"110100101",
  998=>"111000000",
  999=>"000000000",
  1000=>"111111010",
  1001=>"111111111",
  1002=>"000000000",
  1003=>"000001001",
  1004=>"101111101",
  1005=>"000000000",
  1006=>"001101111",
  1007=>"000100110",
  1008=>"100000000",
  1009=>"001000100",
  1010=>"000000100",
  1011=>"000010000",
  1012=>"100000000",
  1013=>"111111111",
  1014=>"011111000",
  1015=>"110110011",
  1016=>"000000000",
  1017=>"011111111",
  1018=>"101101100",
  1019=>"000000001",
  1020=>"111000000",
  1021=>"101001110",
  1022=>"111011111",
  1023=>"000100111",
  1024=>"111111111",
  1025=>"110111111",
  1026=>"000111111",
  1027=>"100100000",
  1028=>"000111111",
  1029=>"111011001",
  1030=>"111011111",
  1031=>"111110000",
  1032=>"011111111",
  1033=>"000010111",
  1034=>"110111111",
  1035=>"000000001",
  1036=>"101001000",
  1037=>"111000000",
  1038=>"001000000",
  1039=>"101110110",
  1040=>"011111111",
  1041=>"111111111",
  1042=>"110011010",
  1043=>"111111111",
  1044=>"000001111",
  1045=>"100100000",
  1046=>"000011000",
  1047=>"000000000",
  1048=>"000000101",
  1049=>"100010000",
  1050=>"000000111",
  1051=>"000000100",
  1052=>"000000000",
  1053=>"101001111",
  1054=>"111011000",
  1055=>"000110000",
  1056=>"000000000",
  1057=>"000001011",
  1058=>"111011000",
  1059=>"111111001",
  1060=>"100111111",
  1061=>"111000000",
  1062=>"000000000",
  1063=>"000100101",
  1064=>"111111011",
  1065=>"000100111",
  1066=>"000100000",
  1067=>"000000111",
  1068=>"011001000",
  1069=>"000000000",
  1070=>"011011000",
  1071=>"110110111",
  1072=>"011111001",
  1073=>"111111000",
  1074=>"000011111",
  1075=>"000000000",
  1076=>"000000000",
  1077=>"100100000",
  1078=>"110100000",
  1079=>"000000000",
  1080=>"000000011",
  1081=>"110000110",
  1082=>"000000001",
  1083=>"101101111",
  1084=>"011111111",
  1085=>"000000000",
  1086=>"000000000",
  1087=>"111111111",
  1088=>"101000000",
  1089=>"110110110",
  1090=>"111111111",
  1091=>"111100000",
  1092=>"111011001",
  1093=>"110111100",
  1094=>"111111111",
  1095=>"111110000",
  1096=>"011001001",
  1097=>"000000000",
  1098=>"000110111",
  1099=>"000000111",
  1100=>"111111000",
  1101=>"000110000",
  1102=>"101110111",
  1103=>"011000000",
  1104=>"000000000",
  1105=>"111111011",
  1106=>"110100111",
  1107=>"111000000",
  1108=>"000001000",
  1109=>"100100000",
  1110=>"011011100",
  1111=>"000000000",
  1112=>"000000000",
  1113=>"111111111",
  1114=>"010000000",
  1115=>"001101111",
  1116=>"101111111",
  1117=>"000110000",
  1118=>"011111111",
  1119=>"111111111",
  1120=>"111111111",
  1121=>"111111111",
  1122=>"001001001",
  1123=>"111111011",
  1124=>"111001001",
  1125=>"111111111",
  1126=>"001001111",
  1127=>"000000000",
  1128=>"111010001",
  1129=>"111011110",
  1130=>"111111100",
  1131=>"000111111",
  1132=>"111111111",
  1133=>"000111111",
  1134=>"000011111",
  1135=>"000010000",
  1136=>"001001111",
  1137=>"011000000",
  1138=>"000000001",
  1139=>"111111111",
  1140=>"111001011",
  1141=>"111111111",
  1142=>"111111011",
  1143=>"111000000",
  1144=>"000000000",
  1145=>"000000000",
  1146=>"000010010",
  1147=>"000000000",
  1148=>"001000000",
  1149=>"111111111",
  1150=>"000110110",
  1151=>"000000000",
  1152=>"110000000",
  1153=>"001000000",
  1154=>"111111111",
  1155=>"000100101",
  1156=>"000000000",
  1157=>"111100000",
  1158=>"010110111",
  1159=>"111111001",
  1160=>"001001011",
  1161=>"100111111",
  1162=>"111001000",
  1163=>"100111111",
  1164=>"000000000",
  1165=>"111111111",
  1166=>"111111001",
  1167=>"111111111",
  1168=>"111111011",
  1169=>"111011001",
  1170=>"111000000",
  1171=>"000101111",
  1172=>"001000010",
  1173=>"000111111",
  1174=>"000000111",
  1175=>"000111111",
  1176=>"000000000",
  1177=>"000110111",
  1178=>"000000000",
  1179=>"111111111",
  1180=>"000001010",
  1181=>"000001101",
  1182=>"111011111",
  1183=>"111111110",
  1184=>"000000000",
  1185=>"111111111",
  1186=>"111111111",
  1187=>"000110111",
  1188=>"000000111",
  1189=>"000000011",
  1190=>"000011111",
  1191=>"000000000",
  1192=>"001000110",
  1193=>"000000000",
  1194=>"110010010",
  1195=>"001111111",
  1196=>"011010010",
  1197=>"011011011",
  1198=>"000000000",
  1199=>"111101000",
  1200=>"100000100",
  1201=>"000001001",
  1202=>"000001001",
  1203=>"000111110",
  1204=>"100100100",
  1205=>"011011111",
  1206=>"111111111",
  1207=>"000000000",
  1208=>"000000000",
  1209=>"000000000",
  1210=>"100000000",
  1211=>"000000000",
  1212=>"000000000",
  1213=>"111111111",
  1214=>"111111010",
  1215=>"000001001",
  1216=>"111111111",
  1217=>"001111011",
  1218=>"111111111",
  1219=>"011111111",
  1220=>"100000001",
  1221=>"011011000",
  1222=>"001000000",
  1223=>"111111111",
  1224=>"000000000",
  1225=>"001000000",
  1226=>"011001001",
  1227=>"000000000",
  1228=>"111110110",
  1229=>"000001000",
  1230=>"111000000",
  1231=>"110000111",
  1232=>"001111111",
  1233=>"000000000",
  1234=>"001001111",
  1235=>"000000000",
  1236=>"111111100",
  1237=>"000000000",
  1238=>"000010010",
  1239=>"111111111",
  1240=>"111111111",
  1241=>"100100100",
  1242=>"111001111",
  1243=>"110000000",
  1244=>"111111101",
  1245=>"000000000",
  1246=>"000001000",
  1247=>"000000000",
  1248=>"000000000",
  1249=>"010111011",
  1250=>"110111111",
  1251=>"111111111",
  1252=>"101111111",
  1253=>"000000010",
  1254=>"111111001",
  1255=>"111111001",
  1256=>"000001011",
  1257=>"000000100",
  1258=>"111111110",
  1259=>"000100000",
  1260=>"110000000",
  1261=>"101111111",
  1262=>"111111111",
  1263=>"000000000",
  1264=>"100100110",
  1265=>"111111111",
  1266=>"000000000",
  1267=>"110000000",
  1268=>"000000011",
  1269=>"111111111",
  1270=>"000000000",
  1271=>"000000000",
  1272=>"011000001",
  1273=>"000000000",
  1274=>"001001000",
  1275=>"110000000",
  1276=>"000010000",
  1277=>"110110010",
  1278=>"000000110",
  1279=>"000000000",
  1280=>"000000000",
  1281=>"001011011",
  1282=>"110111111",
  1283=>"111111111",
  1284=>"000000100",
  1285=>"100110111",
  1286=>"010000000",
  1287=>"000000111",
  1288=>"111111111",
  1289=>"000111111",
  1290=>"010111111",
  1291=>"001111111",
  1292=>"000000000",
  1293=>"111111011",
  1294=>"111110100",
  1295=>"111000000",
  1296=>"100111111",
  1297=>"111101101",
  1298=>"100110100",
  1299=>"000001000",
  1300=>"011001000",
  1301=>"101000000",
  1302=>"001011111",
  1303=>"000000001",
  1304=>"001111111",
  1305=>"111111111",
  1306=>"100100000",
  1307=>"000000000",
  1308=>"000100111",
  1309=>"000000010",
  1310=>"000000000",
  1311=>"111111000",
  1312=>"101001001",
  1313=>"000000000",
  1314=>"111111000",
  1315=>"110100000",
  1316=>"111111111",
  1317=>"111111000",
  1318=>"000000011",
  1319=>"111011011",
  1320=>"111111111",
  1321=>"000000000",
  1322=>"011000000",
  1323=>"000000000",
  1324=>"000000000",
  1325=>"011011010",
  1326=>"111111110",
  1327=>"000000000",
  1328=>"000000000",
  1329=>"100011011",
  1330=>"111101100",
  1331=>"000010011",
  1332=>"000000110",
  1333=>"111111111",
  1334=>"000011011",
  1335=>"000000000",
  1336=>"000000000",
  1337=>"000000000",
  1338=>"100111111",
  1339=>"011000000",
  1340=>"001011111",
  1341=>"011010100",
  1342=>"111111111",
  1343=>"000000000",
  1344=>"000000000",
  1345=>"001000111",
  1346=>"111111000",
  1347=>"000000000",
  1348=>"111111111",
  1349=>"000000000",
  1350=>"111111100",
  1351=>"111111111",
  1352=>"111000000",
  1353=>"000000001",
  1354=>"011010110",
  1355=>"000001000",
  1356=>"001001000",
  1357=>"000111000",
  1358=>"011000000",
  1359=>"000000100",
  1360=>"000000011",
  1361=>"111000000",
  1362=>"110111000",
  1363=>"001000110",
  1364=>"000000100",
  1365=>"010110111",
  1366=>"011011011",
  1367=>"111111111",
  1368=>"000111000",
  1369=>"010010000",
  1370=>"111100100",
  1371=>"000110000",
  1372=>"111101001",
  1373=>"111111011",
  1374=>"110011000",
  1375=>"110010000",
  1376=>"111110000",
  1377=>"000001000",
  1378=>"111111011",
  1379=>"111111111",
  1380=>"001011011",
  1381=>"000000110",
  1382=>"010000000",
  1383=>"000000000",
  1384=>"000000000",
  1385=>"000000010",
  1386=>"000000111",
  1387=>"000000101",
  1388=>"000001111",
  1389=>"001011100",
  1390=>"110111111",
  1391=>"011011001",
  1392=>"110110111",
  1393=>"011000010",
  1394=>"000110100",
  1395=>"000011011",
  1396=>"110100000",
  1397=>"110110111",
  1398=>"111101000",
  1399=>"000000000",
  1400=>"111100111",
  1401=>"111110111",
  1402=>"000000000",
  1403=>"000000000",
  1404=>"100011011",
  1405=>"010111110",
  1406=>"100110110",
  1407=>"111111111",
  1408=>"001101000",
  1409=>"000111010",
  1410=>"111001001",
  1411=>"000000011",
  1412=>"001110111",
  1413=>"000000000",
  1414=>"101111110",
  1415=>"000110100",
  1416=>"100100111",
  1417=>"000000000",
  1418=>"111111111",
  1419=>"111111111",
  1420=>"000011000",
  1421=>"111001000",
  1422=>"000011001",
  1423=>"000010111",
  1424=>"000000111",
  1425=>"111111110",
  1426=>"111111010",
  1427=>"111100100",
  1428=>"000101011",
  1429=>"000111000",
  1430=>"011000111",
  1431=>"111110111",
  1432=>"001011001",
  1433=>"011010000",
  1434=>"111110111",
  1435=>"100100110",
  1436=>"000000101",
  1437=>"111111111",
  1438=>"000000000",
  1439=>"100100111",
  1440=>"000000000",
  1441=>"000100100",
  1442=>"111111111",
  1443=>"000000000",
  1444=>"111111110",
  1445=>"110111000",
  1446=>"000000000",
  1447=>"000000100",
  1448=>"011000000",
  1449=>"000001000",
  1450=>"011111111",
  1451=>"111111111",
  1452=>"111101100",
  1453=>"111111111",
  1454=>"101011000",
  1455=>"100100100",
  1456=>"111111000",
  1457=>"100100111",
  1458=>"111111111",
  1459=>"000000000",
  1460=>"111111111",
  1461=>"000000000",
  1462=>"110111000",
  1463=>"100110000",
  1464=>"111100000",
  1465=>"111111111",
  1466=>"111100000",
  1467=>"000010010",
  1468=>"000000001",
  1469=>"111000000",
  1470=>"000000000",
  1471=>"011011000",
  1472=>"000010111",
  1473=>"000000000",
  1474=>"011011000",
  1475=>"000001001",
  1476=>"010000000",
  1477=>"111000000",
  1478=>"000000000",
  1479=>"000000000",
  1480=>"000000000",
  1481=>"110110000",
  1482=>"110010111",
  1483=>"110000000",
  1484=>"010000000",
  1485=>"000001001",
  1486=>"111000110",
  1487=>"111100100",
  1488=>"000111111",
  1489=>"000000000",
  1490=>"000011111",
  1491=>"111111111",
  1492=>"000000100",
  1493=>"111111100",
  1494=>"000111111",
  1495=>"000000000",
  1496=>"111111000",
  1497=>"100000000",
  1498=>"011001111",
  1499=>"100100000",
  1500=>"000000001",
  1501=>"000000000",
  1502=>"100100001",
  1503=>"000000000",
  1504=>"000111111",
  1505=>"000010000",
  1506=>"000111111",
  1507=>"000000000",
  1508=>"001011010",
  1509=>"000000000",
  1510=>"111111011",
  1511=>"111000000",
  1512=>"001000111",
  1513=>"100111110",
  1514=>"001111111",
  1515=>"111111111",
  1516=>"111111111",
  1517=>"111111111",
  1518=>"000000111",
  1519=>"111010000",
  1520=>"000000000",
  1521=>"111111111",
  1522=>"001000000",
  1523=>"111000000",
  1524=>"010111111",
  1525=>"111111000",
  1526=>"000000000",
  1527=>"000000000",
  1528=>"000000000",
  1529=>"111111100",
  1530=>"111111111",
  1531=>"001111111",
  1532=>"000000000",
  1533=>"111111001",
  1534=>"111111111",
  1535=>"001000000",
  1536=>"000000000",
  1537=>"111111110",
  1538=>"000000000",
  1539=>"111111111",
  1540=>"111111111",
  1541=>"011001000",
  1542=>"111100000",
  1543=>"100000000",
  1544=>"110110000",
  1545=>"111101111",
  1546=>"000000000",
  1547=>"000001100",
  1548=>"100000000",
  1549=>"111111101",
  1550=>"111111110",
  1551=>"111101000",
  1552=>"000000000",
  1553=>"111001000",
  1554=>"001111111",
  1555=>"111111111",
  1556=>"000111111",
  1557=>"101111111",
  1558=>"000010111",
  1559=>"001000000",
  1560=>"111111111",
  1561=>"100100001",
  1562=>"100000110",
  1563=>"011011011",
  1564=>"110110010",
  1565=>"010000000",
  1566=>"000010011",
  1567=>"001001001",
  1568=>"000000000",
  1569=>"110111111",
  1570=>"100000000",
  1571=>"111011000",
  1572=>"100101001",
  1573=>"000110111",
  1574=>"000000000",
  1575=>"000111011",
  1576=>"111111111",
  1577=>"000011011",
  1578=>"000100001",
  1579=>"111111111",
  1580=>"101111111",
  1581=>"000000000",
  1582=>"111111111",
  1583=>"111111111",
  1584=>"000111100",
  1585=>"111111111",
  1586=>"000111111",
  1587=>"110110110",
  1588=>"000001001",
  1589=>"111000000",
  1590=>"111001001",
  1591=>"111001101",
  1592=>"000000001",
  1593=>"101101111",
  1594=>"000000000",
  1595=>"100000100",
  1596=>"000000000",
  1597=>"011111111",
  1598=>"011111010",
  1599=>"111111111",
  1600=>"100100000",
  1601=>"111110110",
  1602=>"100001111",
  1603=>"000000111",
  1604=>"111111110",
  1605=>"001011101",
  1606=>"110110000",
  1607=>"000100000",
  1608=>"000000000",
  1609=>"111110110",
  1610=>"000000000",
  1611=>"111111111",
  1612=>"001000100",
  1613=>"111111111",
  1614=>"100111111",
  1615=>"001001001",
  1616=>"000000100",
  1617=>"000110000",
  1618=>"001001000",
  1619=>"001001001",
  1620=>"001000101",
  1621=>"111111000",
  1622=>"010000010",
  1623=>"111111111",
  1624=>"001001100",
  1625=>"000000000",
  1626=>"000000000",
  1627=>"110110000",
  1628=>"111111111",
  1629=>"000000000",
  1630=>"000010011",
  1631=>"010111111",
  1632=>"000010110",
  1633=>"001010000",
  1634=>"100111011",
  1635=>"110111010",
  1636=>"011011000",
  1637=>"011101101",
  1638=>"111000000",
  1639=>"111101101",
  1640=>"000010111",
  1641=>"111000001",
  1642=>"111100110",
  1643=>"111010000",
  1644=>"111001001",
  1645=>"100010111",
  1646=>"111111111",
  1647=>"111101000",
  1648=>"000000100",
  1649=>"001111111",
  1650=>"111100100",
  1651=>"111111011",
  1652=>"101101101",
  1653=>"110111111",
  1654=>"110110000",
  1655=>"111100000",
  1656=>"011011000",
  1657=>"111001111",
  1658=>"111010000",
  1659=>"000111111",
  1660=>"111011010",
  1661=>"111001000",
  1662=>"000001001",
  1663=>"111101101",
  1664=>"111111111",
  1665=>"000000000",
  1666=>"000000000",
  1667=>"000000100",
  1668=>"111111111",
  1669=>"011000000",
  1670=>"000000000",
  1671=>"000000000",
  1672=>"111111010",
  1673=>"000011111",
  1674=>"111111000",
  1675=>"011000001",
  1676=>"000010111",
  1677=>"001000111",
  1678=>"011011110",
  1679=>"101100000",
  1680=>"000000000",
  1681=>"101111111",
  1682=>"111111111",
  1683=>"111101101",
  1684=>"111111011",
  1685=>"001111111",
  1686=>"111000101",
  1687=>"000000000",
  1688=>"010010011",
  1689=>"000110111",
  1690=>"111111111",
  1691=>"000000000",
  1692=>"110110110",
  1693=>"000000100",
  1694=>"000000000",
  1695=>"111111111",
  1696=>"110111110",
  1697=>"111100000",
  1698=>"111111110",
  1699=>"011011000",
  1700=>"111111100",
  1701=>"111111111",
  1702=>"000000001",
  1703=>"000000000",
  1704=>"110110000",
  1705=>"001001100",
  1706=>"000111111",
  1707=>"000000000",
  1708=>"111111011",
  1709=>"100100000",
  1710=>"000000000",
  1711=>"000100100",
  1712=>"000111111",
  1713=>"101101101",
  1714=>"000000000",
  1715=>"000000000",
  1716=>"111111011",
  1717=>"000000110",
  1718=>"111111111",
  1719=>"111111000",
  1720=>"000000000",
  1721=>"000000101",
  1722=>"100101111",
  1723=>"110111111",
  1724=>"000110111",
  1725=>"111111110",
  1726=>"000000100",
  1727=>"111111111",
  1728=>"101101000",
  1729=>"111111001",
  1730=>"101100100",
  1731=>"001101111",
  1732=>"101001000",
  1733=>"101101111",
  1734=>"110000110",
  1735=>"000011111",
  1736=>"000000000",
  1737=>"111011000",
  1738=>"111111001",
  1739=>"000000000",
  1740=>"000001011",
  1741=>"111111000",
  1742=>"111000000",
  1743=>"111100000",
  1744=>"111111110",
  1745=>"111111010",
  1746=>"001000000",
  1747=>"001000000",
  1748=>"111111101",
  1749=>"100110111",
  1750=>"000000000",
  1751=>"000000000",
  1752=>"111111000",
  1753=>"000000000",
  1754=>"110111111",
  1755=>"001111101",
  1756=>"000000000",
  1757=>"000000000",
  1758=>"000100101",
  1759=>"000100100",
  1760=>"001000000",
  1761=>"000010111",
  1762=>"000000111",
  1763=>"111111100",
  1764=>"111000000",
  1765=>"000011011",
  1766=>"110111000",
  1767=>"000000000",
  1768=>"001000001",
  1769=>"011111111",
  1770=>"111111111",
  1771=>"111111011",
  1772=>"111111111",
  1773=>"000000000",
  1774=>"000111001",
  1775=>"011011000",
  1776=>"111000101",
  1777=>"010111111",
  1778=>"000000000",
  1779=>"000011011",
  1780=>"111001001",
  1781=>"110111011",
  1782=>"110111111",
  1783=>"000000000",
  1784=>"001000110",
  1785=>"000000000",
  1786=>"000010011",
  1787=>"000000000",
  1788=>"001011011",
  1789=>"100000000",
  1790=>"001001001",
  1791=>"000000101",
  1792=>"000000000",
  1793=>"110010000",
  1794=>"000000000",
  1795=>"111110000",
  1796=>"111111111",
  1797=>"111101101",
  1798=>"111111100",
  1799=>"111111111",
  1800=>"000001000",
  1801=>"111111101",
  1802=>"001001000",
  1803=>"110110111",
  1804=>"111011000",
  1805=>"000000100",
  1806=>"111111111",
  1807=>"011011001",
  1808=>"001111101",
  1809=>"000000000",
  1810=>"100110111",
  1811=>"111000000",
  1812=>"001111000",
  1813=>"000000000",
  1814=>"011011011",
  1815=>"000100111",
  1816=>"001001101",
  1817=>"111111111",
  1818=>"000000101",
  1819=>"110000000",
  1820=>"110110000",
  1821=>"000000000",
  1822=>"001000000",
  1823=>"011011001",
  1824=>"100000000",
  1825=>"011011000",
  1826=>"100110111",
  1827=>"000000000",
  1828=>"000011100",
  1829=>"111111111",
  1830=>"000000000",
  1831=>"000000000",
  1832=>"100100000",
  1833=>"011111111",
  1834=>"111111111",
  1835=>"111111110",
  1836=>"001100000",
  1837=>"000000000",
  1838=>"000000000",
  1839=>"101000000",
  1840=>"110110101",
  1841=>"000000000",
  1842=>"011111001",
  1843=>"111111000",
  1844=>"000000000",
  1845=>"000000000",
  1846=>"000111011",
  1847=>"010111011",
  1848=>"111111000",
  1849=>"111111110",
  1850=>"111111100",
  1851=>"011000000",
  1852=>"000000001",
  1853=>"101110100",
  1854=>"001001101",
  1855=>"000001000",
  1856=>"111111111",
  1857=>"111111111",
  1858=>"000000000",
  1859=>"000100000",
  1860=>"001111111",
  1861=>"000000011",
  1862=>"111111111",
  1863=>"000000000",
  1864=>"000000001",
  1865=>"011111010",
  1866=>"000000000",
  1867=>"111111101",
  1868=>"100100000",
  1869=>"111111001",
  1870=>"111111111",
  1871=>"111001001",
  1872=>"001011011",
  1873=>"111001111",
  1874=>"000000000",
  1875=>"100100111",
  1876=>"000000000",
  1877=>"011011111",
  1878=>"000000000",
  1879=>"100000000",
  1880=>"000000000",
  1881=>"000000000",
  1882=>"111111111",
  1883=>"010000000",
  1884=>"111110110",
  1885=>"000000000",
  1886=>"110110000",
  1887=>"001010111",
  1888=>"001000100",
  1889=>"000000000",
  1890=>"101110010",
  1891=>"000000000",
  1892=>"110000110",
  1893=>"000101111",
  1894=>"111000000",
  1895=>"111111000",
  1896=>"011011001",
  1897=>"111111110",
  1898=>"001000111",
  1899=>"111111110",
  1900=>"111101001",
  1901=>"000110000",
  1902=>"100000000",
  1903=>"101111001",
  1904=>"000000000",
  1905=>"110100111",
  1906=>"111111111",
  1907=>"111111110",
  1908=>"110110100",
  1909=>"001001011",
  1910=>"000000000",
  1911=>"000000000",
  1912=>"110000000",
  1913=>"110000000",
  1914=>"000000011",
  1915=>"001001001",
  1916=>"111111111",
  1917=>"000000000",
  1918=>"000010111",
  1919=>"101100001",
  1920=>"110100000",
  1921=>"000000100",
  1922=>"111111111",
  1923=>"010000100",
  1924=>"000011011",
  1925=>"000000000",
  1926=>"111100000",
  1927=>"000000000",
  1928=>"000000000",
  1929=>"111111000",
  1930=>"000000000",
  1931=>"000000000",
  1932=>"111111111",
  1933=>"101111001",
  1934=>"111111111",
  1935=>"000000110",
  1936=>"000000111",
  1937=>"111111111",
  1938=>"101000000",
  1939=>"111111001",
  1940=>"000101111",
  1941=>"110110110",
  1942=>"111001000",
  1943=>"000110100",
  1944=>"000000111",
  1945=>"000000100",
  1946=>"111111110",
  1947=>"111111100",
  1948=>"011011001",
  1949=>"011111000",
  1950=>"101000101",
  1951=>"000000111",
  1952=>"011000000",
  1953=>"111000000",
  1954=>"000000000",
  1955=>"010010111",
  1956=>"011111110",
  1957=>"000000000",
  1958=>"000000000",
  1959=>"000001001",
  1960=>"000000000",
  1961=>"010111111",
  1962=>"111111111",
  1963=>"000000001",
  1964=>"000000000",
  1965=>"011111111",
  1966=>"010111000",
  1967=>"111011011",
  1968=>"111000100",
  1969=>"100001000",
  1970=>"100101000",
  1971=>"101111111",
  1972=>"001111111",
  1973=>"001011111",
  1974=>"100000000",
  1975=>"111111111",
  1976=>"111110000",
  1977=>"100100000",
  1978=>"001000101",
  1979=>"011111111",
  1980=>"010000010",
  1981=>"001000000",
  1982=>"100100100",
  1983=>"110110100",
  1984=>"001000000",
  1985=>"000000000",
  1986=>"000000000",
  1987=>"111111000",
  1988=>"011110000",
  1989=>"100110111",
  1990=>"111111111",
  1991=>"010000000",
  1992=>"000000000",
  1993=>"111111111",
  1994=>"000000000",
  1995=>"000011011",
  1996=>"110110011",
  1997=>"111111111",
  1998=>"000111111",
  1999=>"110110000",
  2000=>"111100111",
  2001=>"100111001",
  2002=>"000100101",
  2003=>"000111111",
  2004=>"111110111",
  2005=>"111111000",
  2006=>"000000011",
  2007=>"001101100",
  2008=>"000000001",
  2009=>"000011101",
  2010=>"111001111",
  2011=>"000011111",
  2012=>"001001001",
  2013=>"000000000",
  2014=>"111000000",
  2015=>"110111100",
  2016=>"011001000",
  2017=>"000111111",
  2018=>"000000001",
  2019=>"101101111",
  2020=>"111111111",
  2021=>"111110110",
  2022=>"000000000",
  2023=>"111111111",
  2024=>"111111111",
  2025=>"111111111",
  2026=>"000000000",
  2027=>"000000000",
  2028=>"000000000",
  2029=>"000001000",
  2030=>"000111111",
  2031=>"111001011",
  2032=>"111101111",
  2033=>"111111111",
  2034=>"001001011",
  2035=>"111010111",
  2036=>"101111111",
  2037=>"100110000",
  2038=>"011011001",
  2039=>"011011000",
  2040=>"000000000",
  2041=>"001111111",
  2042=>"010111010",
  2043=>"111111111",
  2044=>"111111100",
  2045=>"000001001",
  2046=>"000000100",
  2047=>"000000000",
  2048=>"111000000",
  2049=>"111000000",
  2050=>"111111111",
  2051=>"111111111",
  2052=>"000000000",
  2053=>"000100011",
  2054=>"111111000",
  2055=>"000000111",
  2056=>"111001111",
  2057=>"100000000",
  2058=>"000001111",
  2059=>"001111111",
  2060=>"110110010",
  2061=>"111111000",
  2062=>"111111000",
  2063=>"111000000",
  2064=>"001000000",
  2065=>"001001000",
  2066=>"111000000",
  2067=>"000000000",
  2068=>"111111000",
  2069=>"000000101",
  2070=>"111111111",
  2071=>"111111111",
  2072=>"011111111",
  2073=>"101001001",
  2074=>"111101111",
  2075=>"000000001",
  2076=>"000000111",
  2077=>"111000000",
  2078=>"001100000",
  2079=>"010110110",
  2080=>"100111111",
  2081=>"111111111",
  2082=>"111111000",
  2083=>"110000000",
  2084=>"111111111",
  2085=>"101100111",
  2086=>"111111101",
  2087=>"111111001",
  2088=>"000000100",
  2089=>"000000000",
  2090=>"000000010",
  2091=>"000000010",
  2092=>"000000000",
  2093=>"100000000",
  2094=>"111011011",
  2095=>"100100111",
  2096=>"000000000",
  2097=>"011111011",
  2098=>"011110111",
  2099=>"000110111",
  2100=>"000111111",
  2101=>"111111111",
  2102=>"000000000",
  2103=>"000010111",
  2104=>"000000111",
  2105=>"001000000",
  2106=>"000001011",
  2107=>"000000000",
  2108=>"000000000",
  2109=>"111111100",
  2110=>"000000000",
  2111=>"111111000",
  2112=>"000010000",
  2113=>"111100110",
  2114=>"000001111",
  2115=>"111011111",
  2116=>"000011011",
  2117=>"111111111",
  2118=>"111100111",
  2119=>"111111000",
  2120=>"100111111",
  2121=>"111100111",
  2122=>"000111111",
  2123=>"111011010",
  2124=>"011110111",
  2125=>"000000011",
  2126=>"000000000",
  2127=>"111111010",
  2128=>"000000001",
  2129=>"111100000",
  2130=>"000000111",
  2131=>"000000111",
  2132=>"000000000",
  2133=>"000001011",
  2134=>"000000011",
  2135=>"100000000",
  2136=>"000000111",
  2137=>"111000000",
  2138=>"000111111",
  2139=>"111000010",
  2140=>"000000000",
  2141=>"000111111",
  2142=>"011110110",
  2143=>"111111111",
  2144=>"110100000",
  2145=>"110100000",
  2146=>"001111100",
  2147=>"111111111",
  2148=>"000001111",
  2149=>"110101101",
  2150=>"111000000",
  2151=>"000000110",
  2152=>"100000000",
  2153=>"111111111",
  2154=>"100000010",
  2155=>"011000110",
  2156=>"011010000",
  2157=>"111111000",
  2158=>"111011111",
  2159=>"001000000",
  2160=>"000100000",
  2161=>"111111000",
  2162=>"000100110",
  2163=>"100110100",
  2164=>"111100110",
  2165=>"111111111",
  2166=>"100000000",
  2167=>"111111111",
  2168=>"100101100",
  2169=>"111111111",
  2170=>"110111110",
  2171=>"111000000",
  2172=>"001011111",
  2173=>"111111111",
  2174=>"000000000",
  2175=>"000000110",
  2176=>"000000111",
  2177=>"000000000",
  2178=>"000100111",
  2179=>"000000111",
  2180=>"111111111",
  2181=>"111111100",
  2182=>"001000000",
  2183=>"111111011",
  2184=>"000000111",
  2185=>"000000100",
  2186=>"111111111",
  2187=>"000000000",
  2188=>"000000000",
  2189=>"111111000",
  2190=>"111111000",
  2191=>"111011000",
  2192=>"000000111",
  2193=>"111101110",
  2194=>"000000000",
  2195=>"111111111",
  2196=>"100000101",
  2197=>"000000001",
  2198=>"000000000",
  2199=>"111000100",
  2200=>"111000100",
  2201=>"001000000",
  2202=>"111111111",
  2203=>"000000111",
  2204=>"000000000",
  2205=>"000000001",
  2206=>"000000101",
  2207=>"111110000",
  2208=>"000000000",
  2209=>"001000000",
  2210=>"000000001",
  2211=>"111010000",
  2212=>"100000001",
  2213=>"001000000",
  2214=>"110111111",
  2215=>"110110110",
  2216=>"000110101",
  2217=>"011000000",
  2218=>"000000000",
  2219=>"011111111",
  2220=>"011011111",
  2221=>"111100000",
  2222=>"111111000",
  2223=>"001001000",
  2224=>"111110111",
  2225=>"011001000",
  2226=>"010111111",
  2227=>"000000000",
  2228=>"000000101",
  2229=>"111111101",
  2230=>"011000000",
  2231=>"000111000",
  2232=>"110000000",
  2233=>"110000000",
  2234=>"011000000",
  2235=>"111000111",
  2236=>"000000000",
  2237=>"000110110",
  2238=>"000110111",
  2239=>"000000111",
  2240=>"000000000",
  2241=>"000000000",
  2242=>"111111111",
  2243=>"000000000",
  2244=>"000000000",
  2245=>"111111110",
  2246=>"110111111",
  2247=>"000101111",
  2248=>"111011010",
  2249=>"001000000",
  2250=>"000000000",
  2251=>"111000000",
  2252=>"001000110",
  2253=>"101000000",
  2254=>"111111111",
  2255=>"000000100",
  2256=>"001000001",
  2257=>"001001001",
  2258=>"100100101",
  2259=>"111111110",
  2260=>"000000000",
  2261=>"011110110",
  2262=>"000000000",
  2263=>"100101101",
  2264=>"000000001",
  2265=>"111100000",
  2266=>"000000000",
  2267=>"100111111",
  2268=>"000000111",
  2269=>"010110111",
  2270=>"000000000",
  2271=>"000000000",
  2272=>"111111111",
  2273=>"100000000",
  2274=>"000000111",
  2275=>"110000000",
  2276=>"111111010",
  2277=>"111000000",
  2278=>"100110111",
  2279=>"000000000",
  2280=>"111111000",
  2281=>"111111111",
  2282=>"110100001",
  2283=>"111111000",
  2284=>"000000000",
  2285=>"000000000",
  2286=>"000000000",
  2287=>"000000111",
  2288=>"111111101",
  2289=>"111111111",
  2290=>"111000000",
  2291=>"000110101",
  2292=>"011000000",
  2293=>"000000000",
  2294=>"000001111",
  2295=>"000000000",
  2296=>"110111111",
  2297=>"011001111",
  2298=>"111000000",
  2299=>"111111000",
  2300=>"001001011",
  2301=>"010011111",
  2302=>"111010000",
  2303=>"001000000",
  2304=>"111111100",
  2305=>"011011001",
  2306=>"000000010",
  2307=>"111010000",
  2308=>"000000000",
  2309=>"000000000",
  2310=>"111111111",
  2311=>"100000111",
  2312=>"000100111",
  2313=>"000000000",
  2314=>"000000001",
  2315=>"111001000",
  2316=>"111000000",
  2317=>"000010110",
  2318=>"000111111",
  2319=>"111111000",
  2320=>"100000110",
  2321=>"101001111",
  2322=>"111000111",
  2323=>"000000000",
  2324=>"111110000",
  2325=>"001001011",
  2326=>"011001011",
  2327=>"111110000",
  2328=>"111111111",
  2329=>"000111110",
  2330=>"111010000",
  2331=>"111000000",
  2332=>"000010011",
  2333=>"000000001",
  2334=>"000000000",
  2335=>"000111111",
  2336=>"110110111",
  2337=>"000000000",
  2338=>"000000000",
  2339=>"000000111",
  2340=>"111111111",
  2341=>"001111111",
  2342=>"100110000",
  2343=>"100100100",
  2344=>"011001001",
  2345=>"111111000",
  2346=>"000000000",
  2347=>"111111100",
  2348=>"001001111",
  2349=>"001101111",
  2350=>"111000111",
  2351=>"000000001",
  2352=>"000000000",
  2353=>"000000000",
  2354=>"111111111",
  2355=>"000000100",
  2356=>"111111100",
  2357=>"111111000",
  2358=>"000000000",
  2359=>"011001000",
  2360=>"111111111",
  2361=>"100100100",
  2362=>"111111000",
  2363=>"000000110",
  2364=>"001000000",
  2365=>"111001011",
  2366=>"000010000",
  2367=>"110111111",
  2368=>"000000000",
  2369=>"011111111",
  2370=>"000000000",
  2371=>"111000000",
  2372=>"111110000",
  2373=>"111000000",
  2374=>"000001000",
  2375=>"111111001",
  2376=>"111111111",
  2377=>"011001111",
  2378=>"011000000",
  2379=>"000100000",
  2380=>"000000111",
  2381=>"111111111",
  2382=>"101101111",
  2383=>"100000000",
  2384=>"111111001",
  2385=>"000100111",
  2386=>"110100011",
  2387=>"010010000",
  2388=>"000000000",
  2389=>"000000011",
  2390=>"000000000",
  2391=>"000000000",
  2392=>"000000000",
  2393=>"111110001",
  2394=>"111011001",
  2395=>"111111111",
  2396=>"000100101",
  2397=>"011111001",
  2398=>"111000000",
  2399=>"111111111",
  2400=>"110000000",
  2401=>"011111111",
  2402=>"110010000",
  2403=>"001000000",
  2404=>"001000000",
  2405=>"000000000",
  2406=>"000000110",
  2407=>"000001001",
  2408=>"011000000",
  2409=>"111111111",
  2410=>"000000100",
  2411=>"111111111",
  2412=>"000000000",
  2413=>"110010100",
  2414=>"000010000",
  2415=>"001011011",
  2416=>"000000011",
  2417=>"000000110",
  2418=>"000000101",
  2419=>"111111101",
  2420=>"000000000",
  2421=>"001001000",
  2422=>"000000111",
  2423=>"011000000",
  2424=>"111001111",
  2425=>"111001011",
  2426=>"000000000",
  2427=>"110111000",
  2428=>"111111111",
  2429=>"001001111",
  2430=>"100100100",
  2431=>"000000000",
  2432=>"110111111",
  2433=>"001110000",
  2434=>"011111111",
  2435=>"111000000",
  2436=>"100101000",
  2437=>"111111110",
  2438=>"111000000",
  2439=>"100100000",
  2440=>"100000000",
  2441=>"000000000",
  2442=>"111000000",
  2443=>"111111110",
  2444=>"111111001",
  2445=>"011101011",
  2446=>"000010000",
  2447=>"010011000",
  2448=>"000000011",
  2449=>"111111010",
  2450=>"111111111",
  2451=>"100000000",
  2452=>"000000000",
  2453=>"000000000",
  2454=>"111111110",
  2455=>"000000010",
  2456=>"000011111",
  2457=>"001000001",
  2458=>"111000100",
  2459=>"111010000",
  2460=>"000000101",
  2461=>"111111010",
  2462=>"101101000",
  2463=>"000111111",
  2464=>"000000000",
  2465=>"111011010",
  2466=>"111010000",
  2467=>"001000111",
  2468=>"111111000",
  2469=>"000000000",
  2470=>"000000011",
  2471=>"000000000",
  2472=>"111100100",
  2473=>"000001111",
  2474=>"111111111",
  2475=>"101111111",
  2476=>"111101000",
  2477=>"111000000",
  2478=>"000010111",
  2479=>"000000111",
  2480=>"000100110",
  2481=>"000111111",
  2482=>"011000110",
  2483=>"000010111",
  2484=>"110111111",
  2485=>"111111010",
  2486=>"111010000",
  2487=>"011000000",
  2488=>"000000000",
  2489=>"111111100",
  2490=>"011111011",
  2491=>"001011101",
  2492=>"111111101",
  2493=>"011010000",
  2494=>"000100100",
  2495=>"111110000",
  2496=>"100100000",
  2497=>"001000111",
  2498=>"111111000",
  2499=>"111000000",
  2500=>"000000000",
  2501=>"000000111",
  2502=>"000100111",
  2503=>"101101100",
  2504=>"001111111",
  2505=>"111111100",
  2506=>"001000000",
  2507=>"111001000",
  2508=>"111001001",
  2509=>"000000111",
  2510=>"000100000",
  2511=>"110110000",
  2512=>"000100100",
  2513=>"001111111",
  2514=>"100000101",
  2515=>"000111110",
  2516=>"010100000",
  2517=>"000000000",
  2518=>"000000000",
  2519=>"001111110",
  2520=>"111111001",
  2521=>"000000000",
  2522=>"111111111",
  2523=>"111111111",
  2524=>"111111000",
  2525=>"000000101",
  2526=>"111111111",
  2527=>"110000001",
  2528=>"100100111",
  2529=>"000011010",
  2530=>"110111111",
  2531=>"000000000",
  2532=>"000111011",
  2533=>"111111111",
  2534=>"111111111",
  2535=>"100111011",
  2536=>"000111111",
  2537=>"000111111",
  2538=>"111101100",
  2539=>"001111111",
  2540=>"111000101",
  2541=>"000000000",
  2542=>"100100000",
  2543=>"111111111",
  2544=>"000000011",
  2545=>"000000011",
  2546=>"000000111",
  2547=>"000111111",
  2548=>"111000000",
  2549=>"001000000",
  2550=>"000110000",
  2551=>"111111100",
  2552=>"010111111",
  2553=>"100000100",
  2554=>"001011000",
  2555=>"100100111",
  2556=>"101000000",
  2557=>"000000000",
  2558=>"000001111",
  2559=>"011001111",
  2560=>"001011000",
  2561=>"111111000",
  2562=>"000000000",
  2563=>"101000000",
  2564=>"000011010",
  2565=>"001001000",
  2566=>"000000010",
  2567=>"101101000",
  2568=>"111101001",
  2569=>"111111000",
  2570=>"000111111",
  2571=>"111001011",
  2572=>"000000000",
  2573=>"111011000",
  2574=>"101000000",
  2575=>"010010000",
  2576=>"001000111",
  2577=>"111111111",
  2578=>"000000000",
  2579=>"000000111",
  2580=>"111111000",
  2581=>"111111100",
  2582=>"111000000",
  2583=>"110111101",
  2584=>"111111110",
  2585=>"000011111",
  2586=>"111111100",
  2587=>"111110000",
  2588=>"000111111",
  2589=>"001000000",
  2590=>"000000110",
  2591=>"010011011",
  2592=>"100100000",
  2593=>"000000111",
  2594=>"100100000",
  2595=>"001111011",
  2596=>"111001111",
  2597=>"000111111",
  2598=>"111111001",
  2599=>"000001000",
  2600=>"111001000",
  2601=>"111111000",
  2602=>"111011000",
  2603=>"001111000",
  2604=>"000000000",
  2605=>"111111111",
  2606=>"111100110",
  2607=>"110111111",
  2608=>"100111111",
  2609=>"000000111",
  2610=>"110000011",
  2611=>"011111010",
  2612=>"110000011",
  2613=>"000000001",
  2614=>"111111111",
  2615=>"111010000",
  2616=>"111111111",
  2617=>"000000000",
  2618=>"000000000",
  2619=>"000110000",
  2620=>"000000111",
  2621=>"001111110",
  2622=>"111110110",
  2623=>"001111011",
  2624=>"000000000",
  2625=>"111111000",
  2626=>"000100111",
  2627=>"000011101",
  2628=>"100100110",
  2629=>"111111111",
  2630=>"111111000",
  2631=>"111111111",
  2632=>"000100111",
  2633=>"000000000",
  2634=>"001111111",
  2635=>"000000110",
  2636=>"111111111",
  2637=>"000000110",
  2638=>"111011000",
  2639=>"111111111",
  2640=>"111111011",
  2641=>"000101000",
  2642=>"111111010",
  2643=>"111010001",
  2644=>"000000000",
  2645=>"111000110",
  2646=>"011111111",
  2647=>"111111000",
  2648=>"000000100",
  2649=>"000000010",
  2650=>"101101001",
  2651=>"111111111",
  2652=>"111111000",
  2653=>"111111100",
  2654=>"111111000",
  2655=>"110111111",
  2656=>"111000000",
  2657=>"111010000",
  2658=>"000000000",
  2659=>"010000111",
  2660=>"001111100",
  2661=>"000000101",
  2662=>"000000000",
  2663=>"000000111",
  2664=>"000000000",
  2665=>"001100111",
  2666=>"000100000",
  2667=>"100100000",
  2668=>"111011000",
  2669=>"111000000",
  2670=>"111111111",
  2671=>"111100111",
  2672=>"000000010",
  2673=>"000000110",
  2674=>"111001001",
  2675=>"100000111",
  2676=>"111111111",
  2677=>"011111111",
  2678=>"100100111",
  2679=>"111111110",
  2680=>"000000000",
  2681=>"111010000",
  2682=>"110111111",
  2683=>"000000000",
  2684=>"011011011",
  2685=>"000000000",
  2686=>"100111111",
  2687=>"111110000",
  2688=>"000000000",
  2689=>"010000000",
  2690=>"000000111",
  2691=>"111010010",
  2692=>"011011010",
  2693=>"011010111",
  2694=>"111111001",
  2695=>"000111011",
  2696=>"000000000",
  2697=>"000000000",
  2698=>"100110000",
  2699=>"000100010",
  2700=>"000000111",
  2701=>"111110100",
  2702=>"110110000",
  2703=>"001001100",
  2704=>"110100111",
  2705=>"111111111",
  2706=>"000000011",
  2707=>"111011111",
  2708=>"000000000",
  2709=>"111111101",
  2710=>"111000000",
  2711=>"000000000",
  2712=>"010110000",
  2713=>"111100110",
  2714=>"111000000",
  2715=>"111110000",
  2716=>"111111000",
  2717=>"011111000",
  2718=>"010000110",
  2719=>"000101101",
  2720=>"100111111",
  2721=>"000000000",
  2722=>"000101111",
  2723=>"111111111",
  2724=>"000000000",
  2725=>"000100000",
  2726=>"110011111",
  2727=>"001000100",
  2728=>"000011000",
  2729=>"000000000",
  2730=>"111001001",
  2731=>"000100111",
  2732=>"000100101",
  2733=>"000001001",
  2734=>"111111111",
  2735=>"100111000",
  2736=>"000110000",
  2737=>"000010110",
  2738=>"111111110",
  2739=>"000000000",
  2740=>"110010000",
  2741=>"000000000",
  2742=>"111111111",
  2743=>"111000000",
  2744=>"111111110",
  2745=>"000000110",
  2746=>"111000000",
  2747=>"011100000",
  2748=>"010111111",
  2749=>"000001111",
  2750=>"111110000",
  2751=>"111111111",
  2752=>"010011010",
  2753=>"111111111",
  2754=>"001000000",
  2755=>"111000010",
  2756=>"000000000",
  2757=>"111111111",
  2758=>"101000000",
  2759=>"101111111",
  2760=>"000111110",
  2761=>"111111111",
  2762=>"000000000",
  2763=>"111111111",
  2764=>"011011000",
  2765=>"010011111",
  2766=>"111111010",
  2767=>"000000000",
  2768=>"000000000",
  2769=>"111111010",
  2770=>"111111000",
  2771=>"000000000",
  2772=>"111111111",
  2773=>"110111111",
  2774=>"000000000",
  2775=>"010010000",
  2776=>"111111011",
  2777=>"001011001",
  2778=>"000000111",
  2779=>"000000000",
  2780=>"111101000",
  2781=>"000000111",
  2782=>"000001001",
  2783=>"111111000",
  2784=>"011000000",
  2785=>"111111111",
  2786=>"000111111",
  2787=>"011011011",
  2788=>"000000101",
  2789=>"100010000",
  2790=>"110111111",
  2791=>"100111111",
  2792=>"000001111",
  2793=>"000110110",
  2794=>"111110101",
  2795=>"000110111",
  2796=>"110000000",
  2797=>"000000110",
  2798=>"111111111",
  2799=>"000111111",
  2800=>"000000000",
  2801=>"000111111",
  2802=>"000000000",
  2803=>"001001000",
  2804=>"101101101",
  2805=>"000011011",
  2806=>"110111110",
  2807=>"111111111",
  2808=>"000000100",
  2809=>"000000001",
  2810=>"000000000",
  2811=>"111100000",
  2812=>"111101111",
  2813=>"000000100",
  2814=>"000000000",
  2815=>"111000000",
  2816=>"000000000",
  2817=>"110100100",
  2818=>"111110000",
  2819=>"101000000",
  2820=>"000000000",
  2821=>"111111010",
  2822=>"001110110",
  2823=>"100110100",
  2824=>"111111111",
  2825=>"111111111",
  2826=>"111111000",
  2827=>"111100000",
  2828=>"111001111",
  2829=>"000001100",
  2830=>"000100110",
  2831=>"011111000",
  2832=>"000111110",
  2833=>"110100000",
  2834=>"000000000",
  2835=>"111001011",
  2836=>"000000000",
  2837=>"000000111",
  2838=>"111011001",
  2839=>"110000000",
  2840=>"110111011",
  2841=>"000100111",
  2842=>"000000000",
  2843=>"111111000",
  2844=>"111011110",
  2845=>"111000111",
  2846=>"000000000",
  2847=>"000000000",
  2848=>"111001001",
  2849=>"000000000",
  2850=>"011111111",
  2851=>"111111010",
  2852=>"001000000",
  2853=>"000011000",
  2854=>"110111001",
  2855=>"011001000",
  2856=>"000000000",
  2857=>"000000000",
  2858=>"100101001",
  2859=>"000000000",
  2860=>"101111111",
  2861=>"000000000",
  2862=>"000000000",
  2863=>"100111111",
  2864=>"000001000",
  2865=>"000000110",
  2866=>"010000000",
  2867=>"100100111",
  2868=>"110000000",
  2869=>"010011011",
  2870=>"000000001",
  2871=>"001000000",
  2872=>"000000001",
  2873=>"100100111",
  2874=>"100111111",
  2875=>"000000001",
  2876=>"111110110",
  2877=>"001111111",
  2878=>"111101111",
  2879=>"111110000",
  2880=>"000000101",
  2881=>"001000111",
  2882=>"111111111",
  2883=>"000100001",
  2884=>"000010000",
  2885=>"001001001",
  2886=>"010111111",
  2887=>"111111000",
  2888=>"111111111",
  2889=>"111111000",
  2890=>"110111010",
  2891=>"010000111",
  2892=>"111111000",
  2893=>"001000100",
  2894=>"000111111",
  2895=>"001111111",
  2896=>"110001111",
  2897=>"000111111",
  2898=>"111111111",
  2899=>"010010111",
  2900=>"000000011",
  2901=>"000000000",
  2902=>"110000001",
  2903=>"000000000",
  2904=>"111011000",
  2905=>"111000000",
  2906=>"111111111",
  2907=>"000111011",
  2908=>"010110111",
  2909=>"111100000",
  2910=>"010010000",
  2911=>"100000111",
  2912=>"111111111",
  2913=>"111111111",
  2914=>"000101100",
  2915=>"000000111",
  2916=>"011111110",
  2917=>"000000000",
  2918=>"111010001",
  2919=>"111111000",
  2920=>"000000001",
  2921=>"011000100",
  2922=>"111111000",
  2923=>"000101100",
  2924=>"110011011",
  2925=>"001011111",
  2926=>"000000000",
  2927=>"000001000",
  2928=>"001011000",
  2929=>"111000111",
  2930=>"111111000",
  2931=>"111111111",
  2932=>"110000111",
  2933=>"011000000",
  2934=>"000000011",
  2935=>"111100001",
  2936=>"111000000",
  2937=>"111111111",
  2938=>"000000000",
  2939=>"110101101",
  2940=>"001111101",
  2941=>"000001111",
  2942=>"110111000",
  2943=>"000000000",
  2944=>"110000000",
  2945=>"111111111",
  2946=>"101001001",
  2947=>"000000100",
  2948=>"000000000",
  2949=>"000000000",
  2950=>"000000000",
  2951=>"100111111",
  2952=>"000010000",
  2953=>"000000001",
  2954=>"110100001",
  2955=>"111111101",
  2956=>"111111111",
  2957=>"001111111",
  2958=>"000010000",
  2959=>"011000000",
  2960=>"000000000",
  2961=>"111111000",
  2962=>"000011011",
  2963=>"011011011",
  2964=>"101111000",
  2965=>"000000000",
  2966=>"000000000",
  2967=>"111001000",
  2968=>"100000000",
  2969=>"000111111",
  2970=>"000100110",
  2971=>"100100000",
  2972=>"111110000",
  2973=>"000000000",
  2974=>"111111111",
  2975=>"000000000",
  2976=>"111111101",
  2977=>"111110100",
  2978=>"000111110",
  2979=>"001100000",
  2980=>"011100000",
  2981=>"000000000",
  2982=>"000000000",
  2983=>"000000000",
  2984=>"000000000",
  2985=>"000000001",
  2986=>"000000001",
  2987=>"000110111",
  2988=>"000011001",
  2989=>"000110100",
  2990=>"111001111",
  2991=>"111111111",
  2992=>"000000011",
  2993=>"000000000",
  2994=>"100110000",
  2995=>"000011111",
  2996=>"000000000",
  2997=>"000000000",
  2998=>"000000011",
  2999=>"000001111",
  3000=>"000001111",
  3001=>"111111111",
  3002=>"110111111",
  3003=>"000001000",
  3004=>"000000000",
  3005=>"111111111",
  3006=>"000000000",
  3007=>"111111101",
  3008=>"111111000",
  3009=>"000101000",
  3010=>"110000000",
  3011=>"111011000",
  3012=>"000000000",
  3013=>"110000001",
  3014=>"000111000",
  3015=>"101000000",
  3016=>"000000000",
  3017=>"000000110",
  3018=>"010000000",
  3019=>"000000111",
  3020=>"000010000",
  3021=>"000111000",
  3022=>"000000000",
  3023=>"000111000",
  3024=>"010011000",
  3025=>"000100101",
  3026=>"000000000",
  3027=>"111000111",
  3028=>"000000100",
  3029=>"000001000",
  3030=>"000000001",
  3031=>"000000000",
  3032=>"000000111",
  3033=>"000111110",
  3034=>"111000001",
  3035=>"000000111",
  3036=>"000000000",
  3037=>"000000000",
  3038=>"111111000",
  3039=>"011000000",
  3040=>"010110111",
  3041=>"111111000",
  3042=>"000000011",
  3043=>"111111011",
  3044=>"000000111",
  3045=>"000100100",
  3046=>"001010000",
  3047=>"000000011",
  3048=>"111111111",
  3049=>"111111111",
  3050=>"000000101",
  3051=>"101101111",
  3052=>"111111101",
  3053=>"000000000",
  3054=>"111111010",
  3055=>"011111111",
  3056=>"110111111",
  3057=>"111111111",
  3058=>"000001011",
  3059=>"110111110",
  3060=>"000111110",
  3061=>"000000000",
  3062=>"000111111",
  3063=>"000100110",
  3064=>"111111010",
  3065=>"000000000",
  3066=>"001111011",
  3067=>"111111001",
  3068=>"000000000",
  3069=>"111111101",
  3070=>"000000000",
  3071=>"100001001",
  3072=>"100100111",
  3073=>"000000000",
  3074=>"000100000",
  3075=>"000000100",
  3076=>"100000000",
  3077=>"000000100",
  3078=>"000000000",
  3079=>"111000000",
  3080=>"111011000",
  3081=>"111111111",
  3082=>"001000000",
  3083=>"000001101",
  3084=>"000100110",
  3085=>"000000000",
  3086=>"100100101",
  3087=>"111111110",
  3088=>"000000000",
  3089=>"000110100",
  3090=>"111000000",
  3091=>"000000000",
  3092=>"001001001",
  3093=>"111101111",
  3094=>"000111001",
  3095=>"011101111",
  3096=>"111111111",
  3097=>"111110110",
  3098=>"101000111",
  3099=>"111011001",
  3100=>"000000000",
  3101=>"111111100",
  3102=>"011111111",
  3103=>"111111000",
  3104=>"001000000",
  3105=>"111111000",
  3106=>"100001011",
  3107=>"000000000",
  3108=>"001000000",
  3109=>"111111111",
  3110=>"111100000",
  3111=>"111000011",
  3112=>"111111111",
  3113=>"100100111",
  3114=>"000000011",
  3115=>"000000000",
  3116=>"110011011",
  3117=>"000000000",
  3118=>"000111111",
  3119=>"011011111",
  3120=>"011100100",
  3121=>"000000000",
  3122=>"000000000",
  3123=>"111100100",
  3124=>"000000100",
  3125=>"000011111",
  3126=>"001000000",
  3127=>"101011111",
  3128=>"111101000",
  3129=>"000000111",
  3130=>"011011011",
  3131=>"111110010",
  3132=>"000101111",
  3133=>"111111111",
  3134=>"000000001",
  3135=>"111011010",
  3136=>"111111111",
  3137=>"111111111",
  3138=>"001000011",
  3139=>"000000011",
  3140=>"111111111",
  3141=>"111111111",
  3142=>"111000000",
  3143=>"000000101",
  3144=>"111111101",
  3145=>"111111111",
  3146=>"000000000",
  3147=>"111111111",
  3148=>"001111111",
  3149=>"100111000",
  3150=>"100000000",
  3151=>"111111001",
  3152=>"000000000",
  3153=>"011011111",
  3154=>"111111111",
  3155=>"000000101",
  3156=>"100100111",
  3157=>"111000000",
  3158=>"000000000",
  3159=>"111110111",
  3160=>"100000000",
  3161=>"001000000",
  3162=>"111111000",
  3163=>"111101101",
  3164=>"000000000",
  3165=>"111000100",
  3166=>"100100000",
  3167=>"111111000",
  3168=>"111000000",
  3169=>"000000000",
  3170=>"000100111",
  3171=>"111111111",
  3172=>"111011111",
  3173=>"000100110",
  3174=>"111111111",
  3175=>"000000011",
  3176=>"111111000",
  3177=>"111101111",
  3178=>"001001001",
  3179=>"100000000",
  3180=>"000000000",
  3181=>"000000000",
  3182=>"111111111",
  3183=>"111111111",
  3184=>"101111111",
  3185=>"001111000",
  3186=>"100100111",
  3187=>"111000111",
  3188=>"000000000",
  3189=>"110000001",
  3190=>"101111111",
  3191=>"000000111",
  3192=>"110110110",
  3193=>"110000001",
  3194=>"000000000",
  3195=>"111000111",
  3196=>"010110110",
  3197=>"100100101",
  3198=>"000000000",
  3199=>"111111111",
  3200=>"000000000",
  3201=>"000000111",
  3202=>"010000000",
  3203=>"110000000",
  3204=>"000000000",
  3205=>"000111111",
  3206=>"000000100",
  3207=>"000111000",
  3208=>"000000000",
  3209=>"111000110",
  3210=>"110111111",
  3211=>"010000000",
  3212=>"000000001",
  3213=>"000000000",
  3214=>"000000010",
  3215=>"110110111",
  3216=>"000000011",
  3217=>"100100000",
  3218=>"001111110",
  3219=>"111111000",
  3220=>"100110111",
  3221=>"111111000",
  3222=>"000000000",
  3223=>"000000000",
  3224=>"000000000",
  3225=>"111111111",
  3226=>"101000000",
  3227=>"000011111",
  3228=>"011010111",
  3229=>"000000000",
  3230=>"011111110",
  3231=>"101100000",
  3232=>"010111111",
  3233=>"001111111",
  3234=>"010010010",
  3235=>"111111000",
  3236=>"000000000",
  3237=>"000010000",
  3238=>"000000000",
  3239=>"101001111",
  3240=>"100111111",
  3241=>"000000001",
  3242=>"111111111",
  3243=>"111111111",
  3244=>"000000011",
  3245=>"011111111",
  3246=>"111111111",
  3247=>"111111011",
  3248=>"111111010",
  3249=>"111110000",
  3250=>"111111111",
  3251=>"000000000",
  3252=>"001111111",
  3253=>"000000001",
  3254=>"000000111",
  3255=>"111101001",
  3256=>"111111100",
  3257=>"000010111",
  3258=>"000011010",
  3259=>"000001001",
  3260=>"001000000",
  3261=>"001000000",
  3262=>"111110000",
  3263=>"000000000",
  3264=>"000100000",
  3265=>"000000111",
  3266=>"111001001",
  3267=>"110111000",
  3268=>"010000000",
  3269=>"111001001",
  3270=>"111111110",
  3271=>"110000000",
  3272=>"000000000",
  3273=>"000000000",
  3274=>"100110110",
  3275=>"111011000",
  3276=>"001011000",
  3277=>"011011011",
  3278=>"111100000",
  3279=>"000000000",
  3280=>"100110000",
  3281=>"111110000",
  3282=>"111000000",
  3283=>"000000000",
  3284=>"000011111",
  3285=>"000000000",
  3286=>"000100111",
  3287=>"010000001",
  3288=>"111111111",
  3289=>"111101001",
  3290=>"100000111",
  3291=>"011111111",
  3292=>"100000000",
  3293=>"000000000",
  3294=>"000001111",
  3295=>"000000001",
  3296=>"000000111",
  3297=>"000000000",
  3298=>"110110110",
  3299=>"111111111",
  3300=>"111111111",
  3301=>"111110100",
  3302=>"110000100",
  3303=>"111101100",
  3304=>"100111000",
  3305=>"011011110",
  3306=>"111111111",
  3307=>"000000010",
  3308=>"011011000",
  3309=>"111000000",
  3310=>"000010111",
  3311=>"110000000",
  3312=>"110011011",
  3313=>"111111111",
  3314=>"111111111",
  3315=>"000001001",
  3316=>"011111011",
  3317=>"111101001",
  3318=>"111111111",
  3319=>"111111111",
  3320=>"000000001",
  3321=>"110110110",
  3322=>"000000000",
  3323=>"111000000",
  3324=>"111111111",
  3325=>"001001000",
  3326=>"000100111",
  3327=>"001101111",
  3328=>"000000000",
  3329=>"100100100",
  3330=>"000000000",
  3331=>"000000000",
  3332=>"000000000",
  3333=>"000110011",
  3334=>"000000000",
  3335=>"000000000",
  3336=>"100110101",
  3337=>"000000000",
  3338=>"000000000",
  3339=>"000000000",
  3340=>"101000001",
  3341=>"000000000",
  3342=>"110111000",
  3343=>"111111111",
  3344=>"100000000",
  3345=>"001011011",
  3346=>"111000000",
  3347=>"000111111",
  3348=>"000000000",
  3349=>"000000000",
  3350=>"111110100",
  3351=>"110110000",
  3352=>"111111111",
  3353=>"011111111",
  3354=>"111111110",
  3355=>"111111111",
  3356=>"000000100",
  3357=>"000000000",
  3358=>"010010000",
  3359=>"111000000",
  3360=>"000100111",
  3361=>"000000000",
  3362=>"001101111",
  3363=>"100100000",
  3364=>"111010000",
  3365=>"000100001",
  3366=>"001001001",
  3367=>"000000000",
  3368=>"111111111",
  3369=>"100110111",
  3370=>"001000000",
  3371=>"000000000",
  3372=>"101111110",
  3373=>"101011111",
  3374=>"101111111",
  3375=>"111111110",
  3376=>"110111111",
  3377=>"111111110",
  3378=>"111111010",
  3379=>"111111011",
  3380=>"001000001",
  3381=>"111111111",
  3382=>"000110100",
  3383=>"001111111",
  3384=>"011011111",
  3385=>"000000000",
  3386=>"000000000",
  3387=>"000111111",
  3388=>"000000011",
  3389=>"000001111",
  3390=>"100110000",
  3391=>"100101100",
  3392=>"000011111",
  3393=>"111111110",
  3394=>"111011011",
  3395=>"000000000",
  3396=>"000000000",
  3397=>"111111111",
  3398=>"010111110",
  3399=>"001101111",
  3400=>"000000000",
  3401=>"000000000",
  3402=>"111101001",
  3403=>"111011101",
  3404=>"000011001",
  3405=>"011111111",
  3406=>"000001001",
  3407=>"111010011",
  3408=>"111011111",
  3409=>"011111011",
  3410=>"111110100",
  3411=>"000000010",
  3412=>"000000100",
  3413=>"011011000",
  3414=>"000000000",
  3415=>"101001111",
  3416=>"111110010",
  3417=>"110100000",
  3418=>"000000000",
  3419=>"000001111",
  3420=>"011001101",
  3421=>"111111111",
  3422=>"111111111",
  3423=>"001000000",
  3424=>"000001111",
  3425=>"101001000",
  3426=>"101111011",
  3427=>"000000000",
  3428=>"011011001",
  3429=>"000000000",
  3430=>"000000000",
  3431=>"111111111",
  3432=>"111111111",
  3433=>"000000000",
  3434=>"000000000",
  3435=>"111100110",
  3436=>"111010000",
  3437=>"000011000",
  3438=>"111111000",
  3439=>"011111100",
  3440=>"011000110",
  3441=>"000111111",
  3442=>"000000000",
  3443=>"111110000",
  3444=>"011001001",
  3445=>"100110000",
  3446=>"010110000",
  3447=>"111111000",
  3448=>"011001001",
  3449=>"000000001",
  3450=>"000110111",
  3451=>"000100000",
  3452=>"000000000",
  3453=>"110110110",
  3454=>"000000000",
  3455=>"000001000",
  3456=>"000100111",
  3457=>"000011111",
  3458=>"111110000",
  3459=>"111011001",
  3460=>"111111111",
  3461=>"010010010",
  3462=>"001000011",
  3463=>"111001001",
  3464=>"011111111",
  3465=>"000000111",
  3466=>"110000100",
  3467=>"111111010",
  3468=>"000000111",
  3469=>"100100100",
  3470=>"111111111",
  3471=>"000000010",
  3472=>"000000000",
  3473=>"000000011",
  3474=>"001001111",
  3475=>"000000000",
  3476=>"000000000",
  3477=>"000000000",
  3478=>"000110111",
  3479=>"011011111",
  3480=>"111111011",
  3481=>"111001000",
  3482=>"111111000",
  3483=>"001000000",
  3484=>"111011110",
  3485=>"000001000",
  3486=>"100111111",
  3487=>"111011000",
  3488=>"100000000",
  3489=>"111100100",
  3490=>"000110110",
  3491=>"000011111",
  3492=>"100101000",
  3493=>"000000001",
  3494=>"111111111",
  3495=>"100110111",
  3496=>"111011001",
  3497=>"000000000",
  3498=>"000000000",
  3499=>"000000000",
  3500=>"000000000",
  3501=>"000000110",
  3502=>"001011111",
  3503=>"111111111",
  3504=>"111111111",
  3505=>"000000000",
  3506=>"000110001",
  3507=>"000011111",
  3508=>"000000000",
  3509=>"111011011",
  3510=>"001111111",
  3511=>"000001011",
  3512=>"000000111",
  3513=>"000110000",
  3514=>"000010111",
  3515=>"000000000",
  3516=>"111111111",
  3517=>"111100000",
  3518=>"000000101",
  3519=>"000100100",
  3520=>"000000011",
  3521=>"011011001",
  3522=>"000000001",
  3523=>"000000000",
  3524=>"100111011",
  3525=>"001111111",
  3526=>"000011110",
  3527=>"000000101",
  3528=>"000110000",
  3529=>"000111000",
  3530=>"000000000",
  3531=>"101111111",
  3532=>"001101111",
  3533=>"000010111",
  3534=>"111111111",
  3535=>"110110111",
  3536=>"011000011",
  3537=>"011011000",
  3538=>"110111110",
  3539=>"111000000",
  3540=>"000011111",
  3541=>"100000010",
  3542=>"111100000",
  3543=>"000010111",
  3544=>"000011000",
  3545=>"111011010",
  3546=>"100100000",
  3547=>"110000000",
  3548=>"000000000",
  3549=>"000000000",
  3550=>"100110100",
  3551=>"000000111",
  3552=>"000000000",
  3553=>"111111001",
  3554=>"111000000",
  3555=>"111111111",
  3556=>"000111111",
  3557=>"111000110",
  3558=>"000000001",
  3559=>"111000000",
  3560=>"011001001",
  3561=>"000000100",
  3562=>"000000111",
  3563=>"110111111",
  3564=>"001001001",
  3565=>"110100100",
  3566=>"011111111",
  3567=>"001111000",
  3568=>"111110000",
  3569=>"111111010",
  3570=>"111111111",
  3571=>"000000000",
  3572=>"000000000",
  3573=>"111011011",
  3574=>"111111111",
  3575=>"001001000",
  3576=>"111111100",
  3577=>"111000000",
  3578=>"100000001",
  3579=>"111001111",
  3580=>"000010000",
  3581=>"111101111",
  3582=>"111111111",
  3583=>"111111111",
  3584=>"010110110",
  3585=>"000000000",
  3586=>"111111000",
  3587=>"111111111",
  3588=>"010000111",
  3589=>"111111111",
  3590=>"000000000",
  3591=>"010111000",
  3592=>"000000000",
  3593=>"110100000",
  3594=>"000001000",
  3595=>"110111111",
  3596=>"000000000",
  3597=>"000001011",
  3598=>"110110000",
  3599=>"000000000",
  3600=>"000001111",
  3601=>"111111110",
  3602=>"000000000",
  3603=>"000000110",
  3604=>"000000000",
  3605=>"111111000",
  3606=>"111111111",
  3607=>"000000000",
  3608=>"011000100",
  3609=>"001001001",
  3610=>"000000000",
  3611=>"111111111",
  3612=>"111111111",
  3613=>"000000000",
  3614=>"111111111",
  3615=>"000000011",
  3616=>"001011110",
  3617=>"111111100",
  3618=>"001011111",
  3619=>"111000000",
  3620=>"111111111",
  3621=>"000110100",
  3622=>"111111111",
  3623=>"111101111",
  3624=>"110110111",
  3625=>"000000000",
  3626=>"111111111",
  3627=>"010000000",
  3628=>"000011111",
  3629=>"111110000",
  3630=>"000000101",
  3631=>"100000001",
  3632=>"011111111",
  3633=>"000000000",
  3634=>"110110100",
  3635=>"111000000",
  3636=>"000100110",
  3637=>"010010000",
  3638=>"001001111",
  3639=>"110011011",
  3640=>"111111111",
  3641=>"011011111",
  3642=>"111111111",
  3643=>"000000000",
  3644=>"000000000",
  3645=>"111001000",
  3646=>"000000000",
  3647=>"001111000",
  3648=>"001011001",
  3649=>"100111101",
  3650=>"001111111",
  3651=>"000011111",
  3652=>"010111000",
  3653=>"000000000",
  3654=>"111000000",
  3655=>"111111111",
  3656=>"011111000",
  3657=>"111111110",
  3658=>"000001101",
  3659=>"110010000",
  3660=>"001001111",
  3661=>"011001000",
  3662=>"000000000",
  3663=>"111111111",
  3664=>"111001000",
  3665=>"111011111",
  3666=>"000111111",
  3667=>"110110110",
  3668=>"000000000",
  3669=>"110111111",
  3670=>"001000000",
  3671=>"000000000",
  3672=>"110000000",
  3673=>"000111001",
  3674=>"011101001",
  3675=>"001011111",
  3676=>"111010000",
  3677=>"000001000",
  3678=>"001001001",
  3679=>"100010111",
  3680=>"001000000",
  3681=>"011010110",
  3682=>"111000000",
  3683=>"000000001",
  3684=>"011111001",
  3685=>"111111111",
  3686=>"000000000",
  3687=>"000000000",
  3688=>"100110110",
  3689=>"000100110",
  3690=>"110111000",
  3691=>"111000000",
  3692=>"000000000",
  3693=>"000000000",
  3694=>"000000101",
  3695=>"110111110",
  3696=>"000000100",
  3697=>"111111111",
  3698=>"111111111",
  3699=>"000000000",
  3700=>"111000000",
  3701=>"111111111",
  3702=>"011011110",
  3703=>"000111000",
  3704=>"000000000",
  3705=>"000000111",
  3706=>"000000000",
  3707=>"111001011",
  3708=>"011111111",
  3709=>"000000000",
  3710=>"110110111",
  3711=>"001000111",
  3712=>"111111111",
  3713=>"011000000",
  3714=>"111111000",
  3715=>"011001000",
  3716=>"111011001",
  3717=>"000000000",
  3718=>"000000000",
  3719=>"111111011",
  3720=>"111010000",
  3721=>"111111111",
  3722=>"111000000",
  3723=>"011000000",
  3724=>"110111000",
  3725=>"000010111",
  3726=>"111111111",
  3727=>"000000000",
  3728=>"000000000",
  3729=>"000110111",
  3730=>"111111000",
  3731=>"110000000",
  3732=>"000000000",
  3733=>"000000000",
  3734=>"111111111",
  3735=>"000000000",
  3736=>"000000000",
  3737=>"000000111",
  3738=>"000000000",
  3739=>"111111000",
  3740=>"110000010",
  3741=>"111111111",
  3742=>"111000000",
  3743=>"111111111",
  3744=>"110110111",
  3745=>"001000000",
  3746=>"111111111",
  3747=>"000111111",
  3748=>"000011000",
  3749=>"101000000",
  3750=>"000010111",
  3751=>"000000111",
  3752=>"001001100",
  3753=>"111111111",
  3754=>"000000000",
  3755=>"001001111",
  3756=>"101000000",
  3757=>"000110101",
  3758=>"110111111",
  3759=>"000000000",
  3760=>"000000000",
  3761=>"111111111",
  3762=>"110111111",
  3763=>"100111111",
  3764=>"111111111",
  3765=>"001111111",
  3766=>"011111111",
  3767=>"110000000",
  3768=>"000100111",
  3769=>"111111111",
  3770=>"000000000",
  3771=>"001001001",
  3772=>"000000000",
  3773=>"111111111",
  3774=>"000000000",
  3775=>"000000000",
  3776=>"001000000",
  3777=>"111111111",
  3778=>"110100100",
  3779=>"000010000",
  3780=>"111111111",
  3781=>"111111111",
  3782=>"000000010",
  3783=>"010011011",
  3784=>"000111111",
  3785=>"111000001",
  3786=>"000000000",
  3787=>"000100000",
  3788=>"011111100",
  3789=>"111100111",
  3790=>"111000000",
  3791=>"000000000",
  3792=>"111111111",
  3793=>"100000000",
  3794=>"000000000",
  3795=>"110000000",
  3796=>"000000100",
  3797=>"011000000",
  3798=>"101000000",
  3799=>"110000100",
  3800=>"111111111",
  3801=>"111111111",
  3802=>"000000010",
  3803=>"000111011",
  3804=>"111011011",
  3805=>"111101111",
  3806=>"111111111",
  3807=>"110000000",
  3808=>"010111010",
  3809=>"111111000",
  3810=>"011011000",
  3811=>"000000000",
  3812=>"100000000",
  3813=>"100100110",
  3814=>"010111111",
  3815=>"110111111",
  3816=>"111111111",
  3817=>"000100111",
  3818=>"001001111",
  3819=>"000010000",
  3820=>"000000000",
  3821=>"111111111",
  3822=>"111101000",
  3823=>"000000000",
  3824=>"111010110",
  3825=>"111100101",
  3826=>"000000000",
  3827=>"000000101",
  3828=>"100101111",
  3829=>"111011111",
  3830=>"110001111",
  3831=>"000001000",
  3832=>"110000001",
  3833=>"000000000",
  3834=>"111111111",
  3835=>"001101000",
  3836=>"010110110",
  3837=>"011111000",
  3838=>"000010000",
  3839=>"111111000",
  3840=>"111111110",
  3841=>"001000001",
  3842=>"000000000",
  3843=>"111000000",
  3844=>"000000000",
  3845=>"000000000",
  3846=>"111111111",
  3847=>"101100000",
  3848=>"000000110",
  3849=>"111111111",
  3850=>"111111111",
  3851=>"000000000",
  3852=>"111000000",
  3853=>"000000000",
  3854=>"010010011",
  3855=>"111001001",
  3856=>"000000000",
  3857=>"111111111",
  3858=>"001000000",
  3859=>"111101000",
  3860=>"000011011",
  3861=>"000000000",
  3862=>"000000011",
  3863=>"000000000",
  3864=>"111111111",
  3865=>"000110111",
  3866=>"010010000",
  3867=>"111100000",
  3868=>"001001001",
  3869=>"111111111",
  3870=>"111111110",
  3871=>"011001100",
  3872=>"100100000",
  3873=>"111110011",
  3874=>"000100110",
  3875=>"011010110",
  3876=>"110110100",
  3877=>"000100100",
  3878=>"000001111",
  3879=>"111111111",
  3880=>"000111111",
  3881=>"000000111",
  3882=>"001001101",
  3883=>"000110000",
  3884=>"100100100",
  3885=>"001000000",
  3886=>"111111010",
  3887=>"000000000",
  3888=>"011111111",
  3889=>"110111111",
  3890=>"000111111",
  3891=>"000000000",
  3892=>"111111011",
  3893=>"000001000",
  3894=>"000000111",
  3895=>"111111111",
  3896=>"000000000",
  3897=>"111111111",
  3898=>"000000110",
  3899=>"110000111",
  3900=>"111111110",
  3901=>"000000000",
  3902=>"111001111",
  3903=>"011111011",
  3904=>"111101111",
  3905=>"111011111",
  3906=>"001111111",
  3907=>"000000000",
  3908=>"000011011",
  3909=>"000000111",
  3910=>"000000111",
  3911=>"000000000",
  3912=>"111111111",
  3913=>"000111111",
  3914=>"111111110",
  3915=>"111011011",
  3916=>"111001111",
  3917=>"000000000",
  3918=>"111000001",
  3919=>"111111111",
  3920=>"010110111",
  3921=>"000000000",
  3922=>"111011110",
  3923=>"000000000",
  3924=>"000000001",
  3925=>"000000100",
  3926=>"111011010",
  3927=>"100100100",
  3928=>"000111111",
  3929=>"001000000",
  3930=>"010000000",
  3931=>"000000000",
  3932=>"110111111",
  3933=>"000111110",
  3934=>"111111111",
  3935=>"111001100",
  3936=>"101000000",
  3937=>"000000111",
  3938=>"001111111",
  3939=>"000000001",
  3940=>"000000010",
  3941=>"000000000",
  3942=>"111110111",
  3943=>"000000000",
  3944=>"110110110",
  3945=>"111111010",
  3946=>"011000111",
  3947=>"111101101",
  3948=>"011000010",
  3949=>"011111000",
  3950=>"000000000",
  3951=>"111111001",
  3952=>"111111111",
  3953=>"100000000",
  3954=>"111100000",
  3955=>"000000100",
  3956=>"110001101",
  3957=>"111111111",
  3958=>"111101111",
  3959=>"001111000",
  3960=>"111111111",
  3961=>"000111111",
  3962=>"110000000",
  3963=>"111111111",
  3964=>"111111001",
  3965=>"100000000",
  3966=>"000000000",
  3967=>"000000111",
  3968=>"110110110",
  3969=>"000000000",
  3970=>"000000000",
  3971=>"100100000",
  3972=>"010111000",
  3973=>"100100100",
  3974=>"101101111",
  3975=>"001111111",
  3976=>"000000000",
  3977=>"000000000",
  3978=>"111000000",
  3979=>"000111101",
  3980=>"010110110",
  3981=>"000010111",
  3982=>"000000011",
  3983=>"000000011",
  3984=>"000000000",
  3985=>"000000000",
  3986=>"000001000",
  3987=>"111111111",
  3988=>"101101000",
  3989=>"000000000",
  3990=>"111001001",
  3991=>"011000001",
  3992=>"111110100",
  3993=>"011001000",
  3994=>"000000000",
  3995=>"110111111",
  3996=>"000000111",
  3997=>"000110111",
  3998=>"001000110",
  3999=>"110110110",
  4000=>"000000000",
  4001=>"110110101",
  4002=>"000000000",
  4003=>"001000000",
  4004=>"001100101",
  4005=>"111111111",
  4006=>"101101000",
  4007=>"010010111",
  4008=>"000000000",
  4009=>"000000000",
  4010=>"001101100",
  4011=>"000000000",
  4012=>"001000001",
  4013=>"001000000",
  4014=>"111111111",
  4015=>"111111101",
  4016=>"101101000",
  4017=>"000000000",
  4018=>"111001000",
  4019=>"000000000",
  4020=>"000111001",
  4021=>"111111101",
  4022=>"111111001",
  4023=>"000000111",
  4024=>"000000100",
  4025=>"110110110",
  4026=>"000111110",
  4027=>"111111001",
  4028=>"101000000",
  4029=>"111111111",
  4030=>"000000000",
  4031=>"000011011",
  4032=>"000000001",
  4033=>"111111000",
  4034=>"111111111",
  4035=>"111101000",
  4036=>"001000000",
  4037=>"011111111",
  4038=>"000000011",
  4039=>"000000000",
  4040=>"000101111",
  4041=>"010111110",
  4042=>"001000001",
  4043=>"000000111",
  4044=>"011111111",
  4045=>"000111111",
  4046=>"100011000",
  4047=>"111111111",
  4048=>"111111111",
  4049=>"111111111",
  4050=>"000000000",
  4051=>"011111111",
  4052=>"000000010",
  4053=>"000000000",
  4054=>"111111001",
  4055=>"011011001",
  4056=>"000000001",
  4057=>"001000000",
  4058=>"000100111",
  4059=>"111111011",
  4060=>"111111011",
  4061=>"011101111",
  4062=>"111111111",
  4063=>"000000000",
  4064=>"011011010",
  4065=>"011011000",
  4066=>"000000001",
  4067=>"111100000",
  4068=>"111111111",
  4069=>"111111111",
  4070=>"111111111",
  4071=>"111111111",
  4072=>"111111111",
  4073=>"111111111",
  4074=>"101001110",
  4075=>"111101000",
  4076=>"101111111",
  4077=>"010000100",
  4078=>"111001000",
  4079=>"001001001",
  4080=>"000000000",
  4081=>"000111111",
  4082=>"100110010",
  4083=>"111111011",
  4084=>"000000000",
  4085=>"110111111",
  4086=>"000000100",
  4087=>"001111101",
  4088=>"111111111",
  4089=>"001011111",
  4090=>"111111100",
  4091=>"000000001",
  4092=>"111101000",
  4093=>"001000000",
  4094=>"011011011",
  4095=>"000000100",
  4096=>"000000010",
  4097=>"001001000",
  4098=>"000000101",
  4099=>"111001000",
  4100=>"001001001",
  4101=>"101000101",
  4102=>"000111111",
  4103=>"100101100",
  4104=>"111111111",
  4105=>"000010000",
  4106=>"100110100",
  4107=>"111000000",
  4108=>"000001001",
  4109=>"000000100",
  4110=>"000011101",
  4111=>"110011000",
  4112=>"000000000",
  4113=>"000001101",
  4114=>"000111111",
  4115=>"000000111",
  4116=>"000000000",
  4117=>"000001000",
  4118=>"000000000",
  4119=>"111011011",
  4120=>"110111001",
  4121=>"111110100",
  4122=>"000000111",
  4123=>"011110000",
  4124=>"111111111",
  4125=>"111001001",
  4126=>"110100000",
  4127=>"001011111",
  4128=>"000000000",
  4129=>"000000000",
  4130=>"100000111",
  4131=>"010000000",
  4132=>"111111111",
  4133=>"000000000",
  4134=>"000000111",
  4135=>"110111111",
  4136=>"001011011",
  4137=>"101101000",
  4138=>"011001111",
  4139=>"100000000",
  4140=>"110110110",
  4141=>"000000000",
  4142=>"010111010",
  4143=>"000100000",
  4144=>"101000001",
  4145=>"000000011",
  4146=>"000001000",
  4147=>"111000000",
  4148=>"110100100",
  4149=>"000000110",
  4150=>"000001111",
  4151=>"000000000",
  4152=>"000001011",
  4153=>"111111100",
  4154=>"101111111",
  4155=>"010111111",
  4156=>"101001000",
  4157=>"000111111",
  4158=>"011111111",
  4159=>"000000100",
  4160=>"001001000",
  4161=>"000000000",
  4162=>"110111100",
  4163=>"100101100",
  4164=>"000000110",
  4165=>"111111100",
  4166=>"111111111",
  4167=>"000000110",
  4168=>"100100111",
  4169=>"001000011",
  4170=>"111111111",
  4171=>"000011011",
  4172=>"000000111",
  4173=>"011111111",
  4174=>"011011111",
  4175=>"000000000",
  4176=>"111111001",
  4177=>"000000000",
  4178=>"000100100",
  4179=>"000001000",
  4180=>"011111011",
  4181=>"000000000",
  4182=>"110111111",
  4183=>"000000000",
  4184=>"111111101",
  4185=>"101000110",
  4186=>"111101111",
  4187=>"000000000",
  4188=>"111111111",
  4189=>"100100001",
  4190=>"111111111",
  4191=>"001001100",
  4192=>"100100110",
  4193=>"010100111",
  4194=>"111100100",
  4195=>"110110111",
  4196=>"000110000",
  4197=>"000000111",
  4198=>"011000000",
  4199=>"111111111",
  4200=>"110100100",
  4201=>"000000100",
  4202=>"100101110",
  4203=>"111111000",
  4204=>"110001111",
  4205=>"000000111",
  4206=>"111101000",
  4207=>"001011001",
  4208=>"110100100",
  4209=>"100000000",
  4210=>"000100111",
  4211=>"011111101",
  4212=>"111111000",
  4213=>"000111111",
  4214=>"011001111",
  4215=>"111111000",
  4216=>"111111111",
  4217=>"000000100",
  4218=>"000111111",
  4219=>"011001001",
  4220=>"110111000",
  4221=>"000000000",
  4222=>"111111110",
  4223=>"111111111",
  4224=>"001111011",
  4225=>"010110111",
  4226=>"110111111",
  4227=>"111011111",
  4228=>"000000101",
  4229=>"111111110",
  4230=>"111111111",
  4231=>"111000000",
  4232=>"000000000",
  4233=>"000000000",
  4234=>"000111100",
  4235=>"100000000",
  4236=>"100000000",
  4237=>"010111000",
  4238=>"110110110",
  4239=>"001000001",
  4240=>"110100110",
  4241=>"111000110",
  4242=>"111011000",
  4243=>"111111101",
  4244=>"111111101",
  4245=>"011111011",
  4246=>"111111111",
  4247=>"111111100",
  4248=>"000001111",
  4249=>"111010111",
  4250=>"011011011",
  4251=>"101111001",
  4252=>"000000000",
  4253=>"011011001",
  4254=>"111111101",
  4255=>"100000100",
  4256=>"000000000",
  4257=>"100100100",
  4258=>"100101101",
  4259=>"111111111",
  4260=>"000011011",
  4261=>"000000111",
  4262=>"110110111",
  4263=>"111100001",
  4264=>"111000000",
  4265=>"011111111",
  4266=>"111111111",
  4267=>"111011001",
  4268=>"100011111",
  4269=>"110100100",
  4270=>"011011000",
  4271=>"000000000",
  4272=>"110111110",
  4273=>"000100101",
  4274=>"010110010",
  4275=>"010111111",
  4276=>"000000111",
  4277=>"000010011",
  4278=>"100100100",
  4279=>"000000110",
  4280=>"000000100",
  4281=>"110100000",
  4282=>"000000111",
  4283=>"000000101",
  4284=>"001001001",
  4285=>"000000011",
  4286=>"111111111",
  4287=>"111111111",
  4288=>"111111111",
  4289=>"111111111",
  4290=>"111111111",
  4291=>"000000111",
  4292=>"110000000",
  4293=>"111111100",
  4294=>"000000100",
  4295=>"000000000",
  4296=>"000000101",
  4297=>"000111111",
  4298=>"001001101",
  4299=>"111111111",
  4300=>"100111111",
  4301=>"100111111",
  4302=>"010111111",
  4303=>"000000111",
  4304=>"011111111",
  4305=>"000100100",
  4306=>"110111111",
  4307=>"101101111",
  4308=>"001001001",
  4309=>"000000001",
  4310=>"111111111",
  4311=>"010100100",
  4312=>"101111101",
  4313=>"001000000",
  4314=>"000000000",
  4315=>"111111111",
  4316=>"000110000",
  4317=>"000000110",
  4318=>"101000110",
  4319=>"000010000",
  4320=>"000000000",
  4321=>"110110010",
  4322=>"111011001",
  4323=>"111000001",
  4324=>"000000100",
  4325=>"111111101",
  4326=>"000001011",
  4327=>"101111111",
  4328=>"000000110",
  4329=>"111000000",
  4330=>"111111011",
  4331=>"111111111",
  4332=>"000000000",
  4333=>"000000000",
  4334=>"010000000",
  4335=>"111111111",
  4336=>"100000000",
  4337=>"000000100",
  4338=>"111111001",
  4339=>"100110011",
  4340=>"001011111",
  4341=>"110111011",
  4342=>"101110111",
  4343=>"000100111",
  4344=>"100000111",
  4345=>"000001000",
  4346=>"100000111",
  4347=>"000111011",
  4348=>"000000100",
  4349=>"000000000",
  4350=>"000000001",
  4351=>"000100111",
  4352=>"111011000",
  4353=>"110110110",
  4354=>"110111111",
  4355=>"001000000",
  4356=>"000110100",
  4357=>"000000000",
  4358=>"111000000",
  4359=>"101010010",
  4360=>"000000111",
  4361=>"000000110",
  4362=>"000000001",
  4363=>"000100111",
  4364=>"110100111",
  4365=>"110110010",
  4366=>"011000000",
  4367=>"000000000",
  4368=>"001111111",
  4369=>"000111111",
  4370=>"111111111",
  4371=>"000100110",
  4372=>"111111000",
  4373=>"011001000",
  4374=>"001000000",
  4375=>"000000101",
  4376=>"000000000",
  4377=>"000000000",
  4378=>"111110100",
  4379=>"000000000",
  4380=>"001000000",
  4381=>"111111111",
  4382=>"000101111",
  4383=>"011000111",
  4384=>"001001011",
  4385=>"111111110",
  4386=>"111011011",
  4387=>"000000000",
  4388=>"000000000",
  4389=>"111111111",
  4390=>"110110110",
  4391=>"100000110",
  4392=>"111111111",
  4393=>"000000000",
  4394=>"011000000",
  4395=>"111111111",
  4396=>"110111010",
  4397=>"110111110",
  4398=>"000011000",
  4399=>"000000000",
  4400=>"111111100",
  4401=>"000000001",
  4402=>"100100000",
  4403=>"000011011",
  4404=>"110001010",
  4405=>"111111001",
  4406=>"011100100",
  4407=>"000000001",
  4408=>"100000000",
  4409=>"001000000",
  4410=>"111011011",
  4411=>"000001011",
  4412=>"111110100",
  4413=>"001101101",
  4414=>"000000100",
  4415=>"111111110",
  4416=>"110100100",
  4417=>"000110000",
  4418=>"111111001",
  4419=>"100110111",
  4420=>"000000101",
  4421=>"111010111",
  4422=>"111011000",
  4423=>"000000111",
  4424=>"100100111",
  4425=>"011111111",
  4426=>"111110100",
  4427=>"000000000",
  4428=>"000011001",
  4429=>"000001001",
  4430=>"111111111",
  4431=>"100001000",
  4432=>"111111001",
  4433=>"111011110",
  4434=>"000000111",
  4435=>"001011000",
  4436=>"111100101",
  4437=>"001111011",
  4438=>"110110111",
  4439=>"000000000",
  4440=>"110110000",
  4441=>"000100111",
  4442=>"000111111",
  4443=>"110111000",
  4444=>"111111111",
  4445=>"000000111",
  4446=>"110111100",
  4447=>"111011011",
  4448=>"000110010",
  4449=>"110000111",
  4450=>"100000100",
  4451=>"100000111",
  4452=>"001111111",
  4453=>"111111111",
  4454=>"111000001",
  4455=>"000011001",
  4456=>"100100000",
  4457=>"111000000",
  4458=>"000000111",
  4459=>"111100001",
  4460=>"100001001",
  4461=>"000110111",
  4462=>"000000000",
  4463=>"100000100",
  4464=>"100110101",
  4465=>"000001000",
  4466=>"111111000",
  4467=>"010000000",
  4468=>"000000011",
  4469=>"111111111",
  4470=>"111111111",
  4471=>"111111101",
  4472=>"111111111",
  4473=>"011000000",
  4474=>"111111111",
  4475=>"100000000",
  4476=>"111111111",
  4477=>"000100111",
  4478=>"011011000",
  4479=>"000000000",
  4480=>"000000000",
  4481=>"100100101",
  4482=>"000000011",
  4483=>"111001011",
  4484=>"000001011",
  4485=>"000000100",
  4486=>"001000000",
  4487=>"000000101",
  4488=>"000100100",
  4489=>"111111111",
  4490=>"111101001",
  4491=>"111111000",
  4492=>"111011111",
  4493=>"110110011",
  4494=>"111111000",
  4495=>"000000000",
  4496=>"000000000",
  4497=>"110000000",
  4498=>"000000000",
  4499=>"000011000",
  4500=>"000000000",
  4501=>"010010000",
  4502=>"111110111",
  4503=>"110111000",
  4504=>"000110111",
  4505=>"101100101",
  4506=>"000000010",
  4507=>"010000000",
  4508=>"001001000",
  4509=>"111111100",
  4510=>"100000000",
  4511=>"000000000",
  4512=>"000000100",
  4513=>"001100100",
  4514=>"000000011",
  4515=>"111111111",
  4516=>"100110101",
  4517=>"111110110",
  4518=>"000000000",
  4519=>"111111111",
  4520=>"111111111",
  4521=>"110000100",
  4522=>"111001111",
  4523=>"110000000",
  4524=>"111001000",
  4525=>"100100110",
  4526=>"110100100",
  4527=>"111111110",
  4528=>"101111110",
  4529=>"011001011",
  4530=>"000111111",
  4531=>"111111111",
  4532=>"100100100",
  4533=>"000000000",
  4534=>"000000101",
  4535=>"001111000",
  4536=>"011011000",
  4537=>"011011011",
  4538=>"000101111",
  4539=>"100100000",
  4540=>"101111111",
  4541=>"110000000",
  4542=>"000100100",
  4543=>"110100100",
  4544=>"000001111",
  4545=>"000100000",
  4546=>"111100100",
  4547=>"000100100",
  4548=>"100110111",
  4549=>"111011001",
  4550=>"111110110",
  4551=>"000000100",
  4552=>"101000111",
  4553=>"110111111",
  4554=>"111100101",
  4555=>"111111111",
  4556=>"111111000",
  4557=>"001111000",
  4558=>"100111100",
  4559=>"111111011",
  4560=>"000110000",
  4561=>"100100000",
  4562=>"111001111",
  4563=>"110011000",
  4564=>"001001001",
  4565=>"111100100",
  4566=>"111111000",
  4567=>"111111111",
  4568=>"110000000",
  4569=>"010011011",
  4570=>"111111011",
  4571=>"001000111",
  4572=>"001001111",
  4573=>"001000000",
  4574=>"111111001",
  4575=>"000100010",
  4576=>"111111110",
  4577=>"000000000",
  4578=>"000000111",
  4579=>"111001001",
  4580=>"000000101",
  4581=>"111111111",
  4582=>"111111111",
  4583=>"111011001",
  4584=>"111111100",
  4585=>"111001100",
  4586=>"000000000",
  4587=>"100111000",
  4588=>"111111000",
  4589=>"111011100",
  4590=>"000000000",
  4591=>"000000000",
  4592=>"110111010",
  4593=>"110111111",
  4594=>"000100101",
  4595=>"000000000",
  4596=>"000000000",
  4597=>"111111111",
  4598=>"110000000",
  4599=>"111111100",
  4600=>"111111000",
  4601=>"100000000",
  4602=>"111111111",
  4603=>"111111111",
  4604=>"000000000",
  4605=>"000000001",
  4606=>"100100111",
  4607=>"100000111",
  4608=>"111111111",
  4609=>"000000000",
  4610=>"000000000",
  4611=>"000111111",
  4612=>"100000000",
  4613=>"101101000",
  4614=>"011111001",
  4615=>"000000001",
  4616=>"000000000",
  4617=>"101001001",
  4618=>"111111111",
  4619=>"100111011",
  4620=>"100110100",
  4621=>"110100100",
  4622=>"000000101",
  4623=>"100000000",
  4624=>"000000000",
  4625=>"000111111",
  4626=>"110111111",
  4627=>"000000000",
  4628=>"000000000",
  4629=>"111000000",
  4630=>"101101111",
  4631=>"001010011",
  4632=>"100000000",
  4633=>"010000010",
  4634=>"111101000",
  4635=>"001110110",
  4636=>"000110110",
  4637=>"100000000",
  4638=>"001011111",
  4639=>"000000000",
  4640=>"111110111",
  4641=>"111111111",
  4642=>"111111101",
  4643=>"111111111",
  4644=>"111111000",
  4645=>"111010000",
  4646=>"000000000",
  4647=>"000000011",
  4648=>"111100100",
  4649=>"111111111",
  4650=>"000111111",
  4651=>"001000000",
  4652=>"000000000",
  4653=>"111111100",
  4654=>"000000000",
  4655=>"011111111",
  4656=>"110110011",
  4657=>"000000000",
  4658=>"000111111",
  4659=>"111111111",
  4660=>"000000000",
  4661=>"110110110",
  4662=>"000000000",
  4663=>"111111011",
  4664=>"111011001",
  4665=>"000000000",
  4666=>"100000000",
  4667=>"000000111",
  4668=>"000000000",
  4669=>"111111111",
  4670=>"001010000",
  4671=>"101000000",
  4672=>"001111100",
  4673=>"111011111",
  4674=>"000000011",
  4675=>"011010000",
  4676=>"000000000",
  4677=>"000000000",
  4678=>"111111110",
  4679=>"111111111",
  4680=>"111111111",
  4681=>"001000000",
  4682=>"111111111",
  4683=>"011111110",
  4684=>"011001100",
  4685=>"100100000",
  4686=>"000000000",
  4687=>"111110110",
  4688=>"111111100",
  4689=>"000000000",
  4690=>"000110000",
  4691=>"111100111",
  4692=>"000000000",
  4693=>"000000000",
  4694=>"111110111",
  4695=>"001000000",
  4696=>"111111011",
  4697=>"000000000",
  4698=>"001111111",
  4699=>"001000000",
  4700=>"110110111",
  4701=>"111000000",
  4702=>"111000000",
  4703=>"000011001",
  4704=>"000000000",
  4705=>"110100000",
  4706=>"000000000",
  4707=>"111001100",
  4708=>"000101110",
  4709=>"010110111",
  4710=>"111111111",
  4711=>"000000111",
  4712=>"111101111",
  4713=>"000000000",
  4714=>"011111110",
  4715=>"110000000",
  4716=>"000100110",
  4717=>"000010000",
  4718=>"000000000",
  4719=>"111111100",
  4720=>"000000000",
  4721=>"010110111",
  4722=>"011010110",
  4723=>"111111011",
  4724=>"000000001",
  4725=>"000000000",
  4726=>"000111111",
  4727=>"000000000",
  4728=>"000000000",
  4729=>"000000000",
  4730=>"000110111",
  4731=>"111111100",
  4732=>"001001011",
  4733=>"001111111",
  4734=>"000000000",
  4735=>"100000001",
  4736=>"111000000",
  4737=>"111110000",
  4738=>"111111110",
  4739=>"111110111",
  4740=>"100000000",
  4741=>"000000000",
  4742=>"100001001",
  4743=>"110111111",
  4744=>"111100000",
  4745=>"000000000",
  4746=>"111111111",
  4747=>"111111111",
  4748=>"000000100",
  4749=>"111111111",
  4750=>"001111111",
  4751=>"110110000",
  4752=>"111111111",
  4753=>"111010000",
  4754=>"110111101",
  4755=>"001001000",
  4756=>"000000110",
  4757=>"000000000",
  4758=>"111111110",
  4759=>"011000000",
  4760=>"000000110",
  4761=>"111111111",
  4762=>"000000000",
  4763=>"111110110",
  4764=>"011000000",
  4765=>"000100110",
  4766=>"011000000",
  4767=>"000000011",
  4768=>"000000011",
  4769=>"111001010",
  4770=>"011111111",
  4771=>"111111111",
  4772=>"000000100",
  4773=>"010010000",
  4774=>"000000111",
  4775=>"100100111",
  4776=>"000100111",
  4777=>"000000100",
  4778=>"111000000",
  4779=>"111111111",
  4780=>"111100100",
  4781=>"000000101",
  4782=>"001111111",
  4783=>"000000000",
  4784=>"000000111",
  4785=>"000000000",
  4786=>"110111111",
  4787=>"000000000",
  4788=>"001111111",
  4789=>"011111111",
  4790=>"110111111",
  4791=>"001001001",
  4792=>"111111110",
  4793=>"000000000",
  4794=>"001011001",
  4795=>"011110111",
  4796=>"111111100",
  4797=>"111111111",
  4798=>"000111111",
  4799=>"000011010",
  4800=>"010111111",
  4801=>"000000000",
  4802=>"001001011",
  4803=>"000001111",
  4804=>"111111111",
  4805=>"000000000",
  4806=>"111000101",
  4807=>"100110000",
  4808=>"000000000",
  4809=>"001011011",
  4810=>"111000000",
  4811=>"000000000",
  4812=>"000000000",
  4813=>"111101000",
  4814=>"000111111",
  4815=>"101000000",
  4816=>"111100100",
  4817=>"100000000",
  4818=>"000000111",
  4819=>"100100110",
  4820=>"011101101",
  4821=>"111110110",
  4822=>"001001001",
  4823=>"011011111",
  4824=>"100110110",
  4825=>"011111111",
  4826=>"111100000",
  4827=>"000100000",
  4828=>"100000000",
  4829=>"000000110",
  4830=>"111111111",
  4831=>"111101000",
  4832=>"111111111",
  4833=>"001011000",
  4834=>"011000000",
  4835=>"000110111",
  4836=>"111111111",
  4837=>"000000000",
  4838=>"111111111",
  4839=>"000000000",
  4840=>"111111001",
  4841=>"110101111",
  4842=>"001000000",
  4843=>"110000000",
  4844=>"111111110",
  4845=>"111111111",
  4846=>"111110000",
  4847=>"000000110",
  4848=>"110010000",
  4849=>"000000000",
  4850=>"000000000",
  4851=>"011010000",
  4852=>"010111110",
  4853=>"000000000",
  4854=>"110000000",
  4855=>"101001111",
  4856=>"001000100",
  4857=>"111011011",
  4858=>"111111111",
  4859=>"001001001",
  4860=>"011011010",
  4861=>"011001000",
  4862=>"011110110",
  4863=>"000100111",
  4864=>"001001000",
  4865=>"100100101",
  4866=>"111111111",
  4867=>"111001000",
  4868=>"000000000",
  4869=>"000110000",
  4870=>"111111000",
  4871=>"011001000",
  4872=>"000010111",
  4873=>"011111111",
  4874=>"111111111",
  4875=>"000000010",
  4876=>"110110111",
  4877=>"000100110",
  4878=>"000000111",
  4879=>"111111111",
  4880=>"000000111",
  4881=>"101011111",
  4882=>"000000000",
  4883=>"000000000",
  4884=>"011010000",
  4885=>"000011111",
  4886=>"000100001",
  4887=>"011111111",
  4888=>"111111111",
  4889=>"000000000",
  4890=>"111000000",
  4891=>"000110000",
  4892=>"000011111",
  4893=>"000000111",
  4894=>"001000000",
  4895=>"011111111",
  4896=>"111111111",
  4897=>"111111011",
  4898=>"111111111",
  4899=>"111000100",
  4900=>"100100100",
  4901=>"000000000",
  4902=>"110000011",
  4903=>"100000000",
  4904=>"111111111",
  4905=>"000000000",
  4906=>"101111111",
  4907=>"111101001",
  4908=>"000111011",
  4909=>"011101100",
  4910=>"000111100",
  4911=>"110100111",
  4912=>"111011010",
  4913=>"111111100",
  4914=>"111011111",
  4915=>"100111101",
  4916=>"000000110",
  4917=>"111110110",
  4918=>"000000111",
  4919=>"000000000",
  4920=>"111001000",
  4921=>"100000000",
  4922=>"111111111",
  4923=>"001000111",
  4924=>"111111110",
  4925=>"010111110",
  4926=>"001111111",
  4927=>"000000001",
  4928=>"111111111",
  4929=>"000000000",
  4930=>"110110111",
  4931=>"000111111",
  4932=>"000000010",
  4933=>"111110101",
  4934=>"111001001",
  4935=>"000000000",
  4936=>"000000000",
  4937=>"000000000",
  4938=>"111111110",
  4939=>"000001001",
  4940=>"100111100",
  4941=>"111110000",
  4942=>"000011111",
  4943=>"110111111",
  4944=>"000001000",
  4945=>"111111111",
  4946=>"000000100",
  4947=>"000000000",
  4948=>"000110001",
  4949=>"110111111",
  4950=>"010000000",
  4951=>"000001000",
  4952=>"000000111",
  4953=>"110100111",
  4954=>"111111111",
  4955=>"000000000",
  4956=>"111111111",
  4957=>"010000000",
  4958=>"001000000",
  4959=>"001001111",
  4960=>"100111111",
  4961=>"111001001",
  4962=>"000111011",
  4963=>"000111111",
  4964=>"111111111",
  4965=>"000000001",
  4966=>"000000111",
  4967=>"001011111",
  4968=>"001111011",
  4969=>"111111001",
  4970=>"000000000",
  4971=>"000001011",
  4972=>"110110110",
  4973=>"000010111",
  4974=>"000000000",
  4975=>"000100100",
  4976=>"110000000",
  4977=>"111000000",
  4978=>"101111111",
  4979=>"111110110",
  4980=>"000000110",
  4981=>"000001010",
  4982=>"110000000",
  4983=>"111110000",
  4984=>"000000001",
  4985=>"111000000",
  4986=>"000000000",
  4987=>"000000000",
  4988=>"100101111",
  4989=>"000110110",
  4990=>"000000011",
  4991=>"000000000",
  4992=>"001001001",
  4993=>"000111111",
  4994=>"000000000",
  4995=>"000000000",
  4996=>"110110011",
  4997=>"000000000",
  4998=>"111111111",
  4999=>"001001000",
  5000=>"111111101",
  5001=>"111111111",
  5002=>"111111100",
  5003=>"000000000",
  5004=>"011000000",
  5005=>"110110100",
  5006=>"110100000",
  5007=>"000000000",
  5008=>"000001111",
  5009=>"111111111",
  5010=>"101000000",
  5011=>"100111111",
  5012=>"000000000",
  5013=>"001000001",
  5014=>"001111000",
  5015=>"011111001",
  5016=>"000001011",
  5017=>"111001000",
  5018=>"101001001",
  5019=>"111011000",
  5020=>"100110100",
  5021=>"000101100",
  5022=>"000011011",
  5023=>"100000101",
  5024=>"100000000",
  5025=>"011110111",
  5026=>"011111111",
  5027=>"111111111",
  5028=>"100110000",
  5029=>"011000000",
  5030=>"000111111",
  5031=>"111111111",
  5032=>"000000000",
  5033=>"111110110",
  5034=>"010110000",
  5035=>"111000000",
  5036=>"000000000",
  5037=>"001000001",
  5038=>"111000110",
  5039=>"000000000",
  5040=>"111111111",
  5041=>"000000100",
  5042=>"100000000",
  5043=>"011100100",
  5044=>"000010110",
  5045=>"000000000",
  5046=>"000000000",
  5047=>"000011011",
  5048=>"101111000",
  5049=>"000100110",
  5050=>"111100100",
  5051=>"000001001",
  5052=>"000000111",
  5053=>"000111011",
  5054=>"111100000",
  5055=>"001111111",
  5056=>"111111111",
  5057=>"000000000",
  5058=>"111000111",
  5059=>"001000000",
  5060=>"000000001",
  5061=>"111011111",
  5062=>"001110000",
  5063=>"000000100",
  5064=>"001011111",
  5065=>"000001111",
  5066=>"011011010",
  5067=>"111110000",
  5068=>"000000000",
  5069=>"001000111",
  5070=>"101111110",
  5071=>"111000000",
  5072=>"001001001",
  5073=>"000011001",
  5074=>"000110111",
  5075=>"000000000",
  5076=>"111111100",
  5077=>"111111111",
  5078=>"011111011",
  5079=>"111111111",
  5080=>"011010000",
  5081=>"111110110",
  5082=>"001011111",
  5083=>"000000010",
  5084=>"001000000",
  5085=>"011010010",
  5086=>"000000100",
  5087=>"101110110",
  5088=>"001111111",
  5089=>"000000000",
  5090=>"001000011",
  5091=>"000000111",
  5092=>"101100000",
  5093=>"111111000",
  5094=>"101000000",
  5095=>"111110100",
  5096=>"101001001",
  5097=>"011000000",
  5098=>"101000001",
  5099=>"001000000",
  5100=>"001001111",
  5101=>"010000000",
  5102=>"111111001",
  5103=>"001000100",
  5104=>"001101111",
  5105=>"001111111",
  5106=>"000000000",
  5107=>"010000000",
  5108=>"111111111",
  5109=>"110100000",
  5110=>"000000111",
  5111=>"001001000",
  5112=>"000000011",
  5113=>"100010000",
  5114=>"000000000",
  5115=>"111111000",
  5116=>"000000000",
  5117=>"011000000",
  5118=>"001001111",
  5119=>"000000000",
  5120=>"011111011",
  5121=>"100000000",
  5122=>"000100111",
  5123=>"000001110",
  5124=>"100100001",
  5125=>"000000110",
  5126=>"000000000",
  5127=>"111111111",
  5128=>"011011001",
  5129=>"000011111",
  5130=>"000000110",
  5131=>"111111111",
  5132=>"000100100",
  5133=>"000000000",
  5134=>"000000111",
  5135=>"000000111",
  5136=>"110010001",
  5137=>"000000000",
  5138=>"000000000",
  5139=>"111001010",
  5140=>"111111111",
  5141=>"000100111",
  5142=>"100111111",
  5143=>"111111111",
  5144=>"111111000",
  5145=>"111011000",
  5146=>"011000010",
  5147=>"111110001",
  5148=>"000000100",
  5149=>"111111000",
  5150=>"111111000",
  5151=>"000000100",
  5152=>"000011011",
  5153=>"110110110",
  5154=>"000000000",
  5155=>"000000000",
  5156=>"111011011",
  5157=>"000000111",
  5158=>"111101100",
  5159=>"000000000",
  5160=>"000100101",
  5161=>"111000111",
  5162=>"000000111",
  5163=>"101000000",
  5164=>"000000000",
  5165=>"000000000",
  5166=>"000000111",
  5167=>"000000110",
  5168=>"111000111",
  5169=>"011011011",
  5170=>"000000000",
  5171=>"110110100",
  5172=>"111111101",
  5173=>"000100110",
  5174=>"000000000",
  5175=>"000111101",
  5176=>"101101111",
  5177=>"100001111",
  5178=>"001001000",
  5179=>"011000000",
  5180=>"111100101",
  5181=>"000110011",
  5182=>"110000000",
  5183=>"000000111",
  5184=>"100000001",
  5185=>"110110000",
  5186=>"000000111",
  5187=>"000000000",
  5188=>"000111110",
  5189=>"111111111",
  5190=>"000111111",
  5191=>"111111111",
  5192=>"111111110",
  5193=>"001001111",
  5194=>"111111011",
  5195=>"100000111",
  5196=>"111111000",
  5197=>"100000111",
  5198=>"000000011",
  5199=>"111110000",
  5200=>"001100001",
  5201=>"111111111",
  5202=>"000000000",
  5203=>"000000000",
  5204=>"000000000",
  5205=>"110000000",
  5206=>"111111111",
  5207=>"000110010",
  5208=>"000000111",
  5209=>"111000111",
  5210=>"111001001",
  5211=>"000000000",
  5212=>"000000111",
  5213=>"000000111",
  5214=>"000000100",
  5215=>"000000000",
  5216=>"000000000",
  5217=>"111111111",
  5218=>"000111111",
  5219=>"000000111",
  5220=>"010010000",
  5221=>"000111111",
  5222=>"111110000",
  5223=>"100000000",
  5224=>"000000000",
  5225=>"111111111",
  5226=>"000000100",
  5227=>"111111000",
  5228=>"010000100",
  5229=>"000000111",
  5230=>"111111000",
  5231=>"100100000",
  5232=>"001011011",
  5233=>"111111000",
  5234=>"111111000",
  5235=>"111110110",
  5236=>"111000111",
  5237=>"000111000",
  5238=>"001000000",
  5239=>"111111000",
  5240=>"000000011",
  5241=>"100100000",
  5242=>"000000000",
  5243=>"000000000",
  5244=>"110111110",
  5245=>"111111111",
  5246=>"111111000",
  5247=>"111111011",
  5248=>"000000111",
  5249=>"111111000",
  5250=>"111010000",
  5251=>"000001001",
  5252=>"101100000",
  5253=>"111000000",
  5254=>"100000000",
  5255=>"000000010",
  5256=>"111111000",
  5257=>"110101101",
  5258=>"000111111",
  5259=>"000000001",
  5260=>"000000000",
  5261=>"111000000",
  5262=>"100110111",
  5263=>"100000000",
  5264=>"111111111",
  5265=>"000000000",
  5266=>"111111000",
  5267=>"111001111",
  5268=>"100100101",
  5269=>"001000000",
  5270=>"110111111",
  5271=>"000010111",
  5272=>"000000111",
  5273=>"000000111",
  5274=>"111100000",
  5275=>"000000000",
  5276=>"111111111",
  5277=>"000000110",
  5278=>"111111000",
  5279=>"111000000",
  5280=>"100000111",
  5281=>"000000000",
  5282=>"000000001",
  5283=>"000000000",
  5284=>"000000001",
  5285=>"101111111",
  5286=>"000000111",
  5287=>"111111001",
  5288=>"110000001",
  5289=>"001000111",
  5290=>"111000000",
  5291=>"111000000",
  5292=>"111101000",
  5293=>"111111110",
  5294=>"111000101",
  5295=>"110111111",
  5296=>"110010000",
  5297=>"001001000",
  5298=>"111111110",
  5299=>"011111000",
  5300=>"000000000",
  5301=>"111111011",
  5302=>"000000000",
  5303=>"110010111",
  5304=>"000000111",
  5305=>"000000111",
  5306=>"000000100",
  5307=>"000000111",
  5308=>"111111000",
  5309=>"100000111",
  5310=>"111011000",
  5311=>"000100100",
  5312=>"111111111",
  5313=>"111100111",
  5314=>"110111000",
  5315=>"000000111",
  5316=>"110001111",
  5317=>"010011111",
  5318=>"000000000",
  5319=>"000001111",
  5320=>"111110000",
  5321=>"110111000",
  5322=>"000000000",
  5323=>"111111111",
  5324=>"000000000",
  5325=>"010111111",
  5326=>"000000101",
  5327=>"011000010",
  5328=>"011111111",
  5329=>"000000000",
  5330=>"000001011",
  5331=>"000000000",
  5332=>"000000000",
  5333=>"111111010",
  5334=>"000001100",
  5335=>"111000101",
  5336=>"111011111",
  5337=>"110111001",
  5338=>"000000000",
  5339=>"100111111",
  5340=>"111111111",
  5341=>"111100000",
  5342=>"000000001",
  5343=>"101000000",
  5344=>"000000010",
  5345=>"000000110",
  5346=>"111111110",
  5347=>"000000001",
  5348=>"101111111",
  5349=>"000000000",
  5350=>"111111111",
  5351=>"111111111",
  5352=>"111111011",
  5353=>"000011010",
  5354=>"111100000",
  5355=>"111100101",
  5356=>"111111111",
  5357=>"111111111",
  5358=>"000000000",
  5359=>"000000000",
  5360=>"000111000",
  5361=>"100100101",
  5362=>"010111000",
  5363=>"000000111",
  5364=>"000011100",
  5365=>"000000000",
  5366=>"100111100",
  5367=>"111111110",
  5368=>"000000000",
  5369=>"111111110",
  5370=>"100000111",
  5371=>"000000000",
  5372=>"111111000",
  5373=>"110110111",
  5374=>"100111111",
  5375=>"010111111",
  5376=>"000111000",
  5377=>"111111111",
  5378=>"010100111",
  5379=>"000000000",
  5380=>"111110111",
  5381=>"100011001",
  5382=>"000011000",
  5383=>"000001010",
  5384=>"000111111",
  5385=>"000000000",
  5386=>"000000000",
  5387=>"010111111",
  5388=>"000100110",
  5389=>"111111111",
  5390=>"111111000",
  5391=>"110110000",
  5392=>"000101111",
  5393=>"000101111",
  5394=>"110111010",
  5395=>"110100111",
  5396=>"011001001",
  5397=>"011011111",
  5398=>"111000011",
  5399=>"111111000",
  5400=>"000001111",
  5401=>"100000111",
  5402=>"111000000",
  5403=>"000000000",
  5404=>"000111111",
  5405=>"000000000",
  5406=>"000000111",
  5407=>"001100111",
  5408=>"010000111",
  5409=>"111111001",
  5410=>"000100001",
  5411=>"000000000",
  5412=>"000001001",
  5413=>"001011001",
  5414=>"000000000",
  5415=>"000000111",
  5416=>"111111111",
  5417=>"000011010",
  5418=>"000110111",
  5419=>"000000110",
  5420=>"000000111",
  5421=>"000000011",
  5422=>"000010000",
  5423=>"000000000",
  5424=>"000000000",
  5425=>"111111000",
  5426=>"111111000",
  5427=>"000111111",
  5428=>"100101111",
  5429=>"111111111",
  5430=>"111111101",
  5431=>"111111100",
  5432=>"000100100",
  5433=>"000000111",
  5434=>"000000000",
  5435=>"000110110",
  5436=>"000000000",
  5437=>"111111111",
  5438=>"111111111",
  5439=>"000000001",
  5440=>"000000110",
  5441=>"111111000",
  5442=>"111111111",
  5443=>"000000000",
  5444=>"011111111",
  5445=>"111111001",
  5446=>"111111001",
  5447=>"000000000",
  5448=>"000000000",
  5449=>"000100111",
  5450=>"100011000",
  5451=>"111110000",
  5452=>"001001001",
  5453=>"000000000",
  5454=>"000000000",
  5455=>"111111001",
  5456=>"101111100",
  5457=>"111111000",
  5458=>"111111111",
  5459=>"011111000",
  5460=>"000111111",
  5461=>"011011011",
  5462=>"000000000",
  5463=>"100000000",
  5464=>"000111111",
  5465=>"111111111",
  5466=>"111011000",
  5467=>"110111111",
  5468=>"100000000",
  5469=>"000111111",
  5470=>"000011011",
  5471=>"110001001",
  5472=>"111000111",
  5473=>"110111111",
  5474=>"111111011",
  5475=>"101100100",
  5476=>"111111000",
  5477=>"000000000",
  5478=>"000000000",
  5479=>"000000001",
  5480=>"101000011",
  5481=>"000000111",
  5482=>"000110000",
  5483=>"010111000",
  5484=>"010110111",
  5485=>"000111101",
  5486=>"000100110",
  5487=>"000000000",
  5488=>"000000000",
  5489=>"100111000",
  5490=>"000000000",
  5491=>"011000000",
  5492=>"000000000",
  5493=>"100100111",
  5494=>"000000000",
  5495=>"010111111",
  5496=>"001001001",
  5497=>"111000000",
  5498=>"000000000",
  5499=>"111111101",
  5500=>"000000000",
  5501=>"000000000",
  5502=>"111111001",
  5503=>"111111111",
  5504=>"000000001",
  5505=>"100000111",
  5506=>"111111111",
  5507=>"001111111",
  5508=>"000000000",
  5509=>"011111111",
  5510=>"100111111",
  5511=>"101000000",
  5512=>"000001111",
  5513=>"000000000",
  5514=>"000000000",
  5515=>"011000011",
  5516=>"101000111",
  5517=>"110110000",
  5518=>"100000110",
  5519=>"000111110",
  5520=>"110000000",
  5521=>"000000101",
  5522=>"000000011",
  5523=>"000000000",
  5524=>"000000000",
  5525=>"000010000",
  5526=>"111000101",
  5527=>"010100100",
  5528=>"000000000",
  5529=>"000000010",
  5530=>"111111111",
  5531=>"111111111",
  5532=>"100110111",
  5533=>"111111010",
  5534=>"110100000",
  5535=>"001001111",
  5536=>"010000000",
  5537=>"110100100",
  5538=>"100000100",
  5539=>"111111000",
  5540=>"100110110",
  5541=>"111001000",
  5542=>"111000000",
  5543=>"110000000",
  5544=>"000000000",
  5545=>"011011011",
  5546=>"010011011",
  5547=>"000100000",
  5548=>"011001000",
  5549=>"100111001",
  5550=>"110100000",
  5551=>"000001000",
  5552=>"110000101",
  5553=>"000000000",
  5554=>"111000001",
  5555=>"111000000",
  5556=>"000000111",
  5557=>"110100000",
  5558=>"100111000",
  5559=>"000111111",
  5560=>"111010111",
  5561=>"111001000",
  5562=>"011000000",
  5563=>"000000000",
  5564=>"000000111",
  5565=>"111101110",
  5566=>"000000110",
  5567=>"001100111",
  5568=>"100111000",
  5569=>"000000111",
  5570=>"000000111",
  5571=>"000000111",
  5572=>"110111111",
  5573=>"111000000",
  5574=>"001001111",
  5575=>"010000000",
  5576=>"110110101",
  5577=>"000000111",
  5578=>"000000000",
  5579=>"111111111",
  5580=>"101000000",
  5581=>"111111110",
  5582=>"000000000",
  5583=>"110111110",
  5584=>"000000000",
  5585=>"000000111",
  5586=>"111111111",
  5587=>"000000111",
  5588=>"111111011",
  5589=>"000000000",
  5590=>"000000000",
  5591=>"000000000",
  5592=>"111111111",
  5593=>"000000000",
  5594=>"000000111",
  5595=>"000011111",
  5596=>"000000111",
  5597=>"000000000",
  5598=>"011010000",
  5599=>"000010000",
  5600=>"000001111",
  5601=>"000000010",
  5602=>"111111111",
  5603=>"111111111",
  5604=>"111000000",
  5605=>"100100000",
  5606=>"111111010",
  5607=>"111101001",
  5608=>"111000101",
  5609=>"000111111",
  5610=>"000101111",
  5611=>"000100100",
  5612=>"100101000",
  5613=>"111111001",
  5614=>"000000000",
  5615=>"111111000",
  5616=>"000000000",
  5617=>"111111111",
  5618=>"111111000",
  5619=>"000000000",
  5620=>"100100111",
  5621=>"000000101",
  5622=>"000000000",
  5623=>"000000011",
  5624=>"111111111",
  5625=>"000000000",
  5626=>"000000001",
  5627=>"111111111",
  5628=>"100111111",
  5629=>"100100111",
  5630=>"100000000",
  5631=>"000000000",
  5632=>"011010000",
  5633=>"000000000",
  5634=>"000000011",
  5635=>"111011010",
  5636=>"000100110",
  5637=>"111111111",
  5638=>"000000000",
  5639=>"011000001",
  5640=>"111110110",
  5641=>"001000001",
  5642=>"000000000",
  5643=>"000000100",
  5644=>"000000010",
  5645=>"000111111",
  5646=>"111011000",
  5647=>"111111000",
  5648=>"011111111",
  5649=>"000000000",
  5650=>"000001001",
  5651=>"000000111",
  5652=>"000000000",
  5653=>"000000100",
  5654=>"011001001",
  5655=>"011011111",
  5656=>"101110000",
  5657=>"000000000",
  5658=>"011111111",
  5659=>"100000000",
  5660=>"000000111",
  5661=>"011011111",
  5662=>"100000000",
  5663=>"000000100",
  5664=>"111011000",
  5665=>"100100110",
  5666=>"101111011",
  5667=>"000100110",
  5668=>"100111111",
  5669=>"000000000",
  5670=>"100101101",
  5671=>"111111111",
  5672=>"100000001",
  5673=>"011111111",
  5674=>"111111111",
  5675=>"111011000",
  5676=>"111111101",
  5677=>"111111000",
  5678=>"001000000",
  5679=>"111001001",
  5680=>"110111011",
  5681=>"011111011",
  5682=>"000000000",
  5683=>"001101111",
  5684=>"001101001",
  5685=>"000000000",
  5686=>"110000000",
  5687=>"100011011",
  5688=>"011011000",
  5689=>"001001111",
  5690=>"110111111",
  5691=>"011111111",
  5692=>"001001001",
  5693=>"101111011",
  5694=>"111100110",
  5695=>"111111111",
  5696=>"000000110",
  5697=>"000010111",
  5698=>"111000000",
  5699=>"111011000",
  5700=>"100110110",
  5701=>"000000011",
  5702=>"010000010",
  5703=>"111111111",
  5704=>"100110010",
  5705=>"111111111",
  5706=>"000000111",
  5707=>"101000101",
  5708=>"000000000",
  5709=>"000000000",
  5710=>"110100101",
  5711=>"100111111",
  5712=>"111111111",
  5713=>"100100001",
  5714=>"000000010",
  5715=>"101100110",
  5716=>"011000111",
  5717=>"000000000",
  5718=>"111110111",
  5719=>"111111101",
  5720=>"100101000",
  5721=>"111111111",
  5722=>"111111111",
  5723=>"000001001",
  5724=>"000000100",
  5725=>"000000000",
  5726=>"000000100",
  5727=>"110110000",
  5728=>"000000111",
  5729=>"111111111",
  5730=>"000000000",
  5731=>"001000000",
  5732=>"110111100",
  5733=>"111111111",
  5734=>"000000000",
  5735=>"000000000",
  5736=>"111111111",
  5737=>"011000010",
  5738=>"001011111",
  5739=>"110111111",
  5740=>"111111111",
  5741=>"000111000",
  5742=>"111111101",
  5743=>"000001001",
  5744=>"100000111",
  5745=>"000010010",
  5746=>"000100101",
  5747=>"000010111",
  5748=>"111111111",
  5749=>"000000000",
  5750=>"000000000",
  5751=>"000000101",
  5752=>"000110110",
  5753=>"110110111",
  5754=>"011111000",
  5755=>"001000000",
  5756=>"100100100",
  5757=>"111111111",
  5758=>"001111111",
  5759=>"000000000",
  5760=>"111111111",
  5761=>"100000111",
  5762=>"111111111",
  5763=>"001001001",
  5764=>"111111111",
  5765=>"111111111",
  5766=>"111111000",
  5767=>"000000000",
  5768=>"111000011",
  5769=>"110011011",
  5770=>"000000000",
  5771=>"000000000",
  5772=>"111111111",
  5773=>"000000000",
  5774=>"000000001",
  5775=>"000000000",
  5776=>"111001011",
  5777=>"001000001",
  5778=>"000010010",
  5779=>"110111010",
  5780=>"011111110",
  5781=>"000011011",
  5782=>"111111111",
  5783=>"111111111",
  5784=>"000000001",
  5785=>"010000000",
  5786=>"000000000",
  5787=>"000000100",
  5788=>"001001111",
  5789=>"010110111",
  5790=>"111111111",
  5791=>"000000000",
  5792=>"011111100",
  5793=>"110110010",
  5794=>"000000000",
  5795=>"100000000",
  5796=>"000000000",
  5797=>"000000000",
  5798=>"111111000",
  5799=>"001101100",
  5800=>"111000000",
  5801=>"000000000",
  5802=>"111000000",
  5803=>"010100111",
  5804=>"000000000",
  5805=>"001111110",
  5806=>"000001000",
  5807=>"111111100",
  5808=>"000000000",
  5809=>"000000000",
  5810=>"010011010",
  5811=>"111111110",
  5812=>"001111000",
  5813=>"111111111",
  5814=>"001000000",
  5815=>"000001000",
  5816=>"000000000",
  5817=>"111111111",
  5818=>"010000100",
  5819=>"101111111",
  5820=>"010000000",
  5821=>"001001000",
  5822=>"001000000",
  5823=>"100111111",
  5824=>"111000001",
  5825=>"000100000",
  5826=>"111000010",
  5827=>"011111000",
  5828=>"111111110",
  5829=>"101111111",
  5830=>"000000111",
  5831=>"111111111",
  5832=>"010000000",
  5833=>"111111000",
  5834=>"000001001",
  5835=>"000101111",
  5836=>"000000011",
  5837=>"000000000",
  5838=>"100110111",
  5839=>"001001111",
  5840=>"000000000",
  5841=>"101000000",
  5842=>"000000000",
  5843=>"111111111",
  5844=>"000000000",
  5845=>"000100110",
  5846=>"011111111",
  5847=>"000000101",
  5848=>"000000000",
  5849=>"111111111",
  5850=>"000000110",
  5851=>"011111111",
  5852=>"111000000",
  5853=>"000000000",
  5854=>"000000000",
  5855=>"111011110",
  5856=>"110110010",
  5857=>"110111111",
  5858=>"000000000",
  5859=>"000000000",
  5860=>"000001000",
  5861=>"100100000",
  5862=>"111111111",
  5863=>"111111111",
  5864=>"010010000",
  5865=>"000000100",
  5866=>"000000000",
  5867=>"000000000",
  5868=>"001001000",
  5869=>"111111110",
  5870=>"100111111",
  5871=>"111111011",
  5872=>"111111111",
  5873=>"000111111",
  5874=>"111111111",
  5875=>"011011111",
  5876=>"000000000",
  5877=>"111000000",
  5878=>"000001000",
  5879=>"111110000",
  5880=>"000111001",
  5881=>"111111111",
  5882=>"110110000",
  5883=>"011010001",
  5884=>"000001011",
  5885=>"100100000",
  5886=>"000000111",
  5887=>"000010010",
  5888=>"110100100",
  5889=>"101000000",
  5890=>"000000000",
  5891=>"000000111",
  5892=>"000110100",
  5893=>"110010011",
  5894=>"101111111",
  5895=>"111010010",
  5896=>"001110110",
  5897=>"000000000",
  5898=>"111111111",
  5899=>"110111110",
  5900=>"111111111",
  5901=>"111001000",
  5902=>"001000101",
  5903=>"000000011",
  5904=>"110111111",
  5905=>"111111111",
  5906=>"011000000",
  5907=>"111111111",
  5908=>"111111111",
  5909=>"010000000",
  5910=>"100100100",
  5911=>"111111100",
  5912=>"100111000",
  5913=>"000000100",
  5914=>"000000000",
  5915=>"000111001",
  5916=>"001000000",
  5917=>"111100100",
  5918=>"000000111",
  5919=>"000111111",
  5920=>"101111111",
  5921=>"110111110",
  5922=>"111001000",
  5923=>"100110110",
  5924=>"110110010",
  5925=>"111111111",
  5926=>"100100000",
  5927=>"111111100",
  5928=>"111100111",
  5929=>"111111000",
  5930=>"111111001",
  5931=>"110100100",
  5932=>"111110011",
  5933=>"100111111",
  5934=>"100111111",
  5935=>"111111111",
  5936=>"010111111",
  5937=>"010010010",
  5938=>"111001111",
  5939=>"000000000",
  5940=>"110110111",
  5941=>"111111101",
  5942=>"001111111",
  5943=>"110000000",
  5944=>"010110000",
  5945=>"111111000",
  5946=>"111111111",
  5947=>"000100111",
  5948=>"000100001",
  5949=>"101001000",
  5950=>"000100100",
  5951=>"100111111",
  5952=>"000000000",
  5953=>"100000000",
  5954=>"001001011",
  5955=>"111111111",
  5956=>"000000001",
  5957=>"111111111",
  5958=>"000000000",
  5959=>"000000001",
  5960=>"000010000",
  5961=>"111111111",
  5962=>"000010010",
  5963=>"011011011",
  5964=>"000000011",
  5965=>"000000000",
  5966=>"000000000",
  5967=>"100100110",
  5968=>"000010000",
  5969=>"000000000",
  5970=>"111111111",
  5971=>"111111100",
  5972=>"000100110",
  5973=>"011011011",
  5974=>"111111111",
  5975=>"000000000",
  5976=>"011011011",
  5977=>"111001000",
  5978=>"000000000",
  5979=>"111110100",
  5980=>"111000001",
  5981=>"111111101",
  5982=>"011011011",
  5983=>"111100000",
  5984=>"111010000",
  5985=>"000000110",
  5986=>"001001001",
  5987=>"011000000",
  5988=>"100000001",
  5989=>"111010000",
  5990=>"000000000",
  5991=>"000111110",
  5992=>"111100110",
  5993=>"010000000",
  5994=>"000010111",
  5995=>"011011111",
  5996=>"100110111",
  5997=>"010000110",
  5998=>"010000000",
  5999=>"110000000",
  6000=>"011111010",
  6001=>"000000100",
  6002=>"111010110",
  6003=>"111111001",
  6004=>"111111111",
  6005=>"000000000",
  6006=>"111111111",
  6007=>"000000000",
  6008=>"111111001",
  6009=>"000000110",
  6010=>"000000110",
  6011=>"110010000",
  6012=>"110000000",
  6013=>"111111111",
  6014=>"111111100",
  6015=>"000000000",
  6016=>"000001000",
  6017=>"111111011",
  6018=>"001011100",
  6019=>"010110111",
  6020=>"000000110",
  6021=>"000000000",
  6022=>"111110111",
  6023=>"111111111",
  6024=>"010110011",
  6025=>"000000011",
  6026=>"111111111",
  6027=>"111111111",
  6028=>"111111111",
  6029=>"001001001",
  6030=>"100100000",
  6031=>"000000000",
  6032=>"001011110",
  6033=>"000000000",
  6034=>"111111101",
  6035=>"000000010",
  6036=>"111111010",
  6037=>"000010000",
  6038=>"101101111",
  6039=>"111111111",
  6040=>"111000101",
  6041=>"001001001",
  6042=>"111110111",
  6043=>"101001101",
  6044=>"000000001",
  6045=>"000000000",
  6046=>"111111111",
  6047=>"000000000",
  6048=>"000000000",
  6049=>"111011111",
  6050=>"111101111",
  6051=>"011010111",
  6052=>"111111111",
  6053=>"010110000",
  6054=>"000010000",
  6055=>"000000111",
  6056=>"111111111",
  6057=>"000111111",
  6058=>"111111111",
  6059=>"111110111",
  6060=>"110010000",
  6061=>"000000000",
  6062=>"110110110",
  6063=>"000001000",
  6064=>"000010000",
  6065=>"010110110",
  6066=>"001000000",
  6067=>"100010000",
  6068=>"000000001",
  6069=>"000000000",
  6070=>"000100100",
  6071=>"110111010",
  6072=>"011001111",
  6073=>"000000000",
  6074=>"111011111",
  6075=>"111100000",
  6076=>"010010010",
  6077=>"111110110",
  6078=>"111110101",
  6079=>"101101100",
  6080=>"000000100",
  6081=>"000000111",
  6082=>"101111111",
  6083=>"001000000",
  6084=>"000000000",
  6085=>"110000000",
  6086=>"101000111",
  6087=>"111101000",
  6088=>"000000000",
  6089=>"000000000",
  6090=>"111111000",
  6091=>"111111001",
  6092=>"011111111",
  6093=>"000000000",
  6094=>"000000011",
  6095=>"000000000",
  6096=>"100000111",
  6097=>"101001011",
  6098=>"000000000",
  6099=>"000000100",
  6100=>"100000000",
  6101=>"100110100",
  6102=>"000000000",
  6103=>"110111100",
  6104=>"000000000",
  6105=>"111001001",
  6106=>"110000000",
  6107=>"001011111",
  6108=>"111111111",
  6109=>"011000010",
  6110=>"111000101",
  6111=>"000100110",
  6112=>"000000000",
  6113=>"110000110",
  6114=>"111010001",
  6115=>"100100111",
  6116=>"111000010",
  6117=>"111110111",
  6118=>"100110111",
  6119=>"100110110",
  6120=>"111101111",
  6121=>"001001111",
  6122=>"110110111",
  6123=>"111100000",
  6124=>"001100110",
  6125=>"101111101",
  6126=>"111111111",
  6127=>"111111111",
  6128=>"000000000",
  6129=>"111111111",
  6130=>"110000000",
  6131=>"011000000",
  6132=>"101000000",
  6133=>"000000000",
  6134=>"000000000",
  6135=>"001100100",
  6136=>"101001001",
  6137=>"001001001",
  6138=>"111111010",
  6139=>"000000000",
  6140=>"000000011",
  6141=>"000000000",
  6142=>"111111111",
  6143=>"110110111",
  6144=>"000000000",
  6145=>"000000111",
  6146=>"000000111",
  6147=>"000000001",
  6148=>"000000000",
  6149=>"000000000",
  6150=>"000100110",
  6151=>"111111111",
  6152=>"011000000",
  6153=>"101111101",
  6154=>"000100110",
  6155=>"111111111",
  6156=>"110110100",
  6157=>"111111111",
  6158=>"111111111",
  6159=>"111100000",
  6160=>"001001000",
  6161=>"000111111",
  6162=>"000000101",
  6163=>"001000000",
  6164=>"000110111",
  6165=>"011000000",
  6166=>"000000100",
  6167=>"000001011",
  6168=>"010000000",
  6169=>"011110010",
  6170=>"011100111",
  6171=>"000110111",
  6172=>"000110001",
  6173=>"101111111",
  6174=>"100100101",
  6175=>"000010000",
  6176=>"001000000",
  6177=>"110110110",
  6178=>"111111110",
  6179=>"111111101",
  6180=>"101010000",
  6181=>"111110110",
  6182=>"000000000",
  6183=>"110000000",
  6184=>"001011111",
  6185=>"000000111",
  6186=>"000000010",
  6187=>"111111111",
  6188=>"110110111",
  6189=>"000100111",
  6190=>"000000000",
  6191=>"001000000",
  6192=>"111000000",
  6193=>"000000000",
  6194=>"000100100",
  6195=>"000000000",
  6196=>"111111001",
  6197=>"010011011",
  6198=>"111111111",
  6199=>"000000000",
  6200=>"111011111",
  6201=>"110110111",
  6202=>"111111111",
  6203=>"111111111",
  6204=>"111100000",
  6205=>"001101101",
  6206=>"001000000",
  6207=>"111111111",
  6208=>"110111110",
  6209=>"110100000",
  6210=>"000001000",
  6211=>"010010001",
  6212=>"001111111",
  6213=>"111111111",
  6214=>"000000001",
  6215=>"000111011",
  6216=>"111111110",
  6217=>"000000111",
  6218=>"111010111",
  6219=>"000000000",
  6220=>"110000001",
  6221=>"100110000",
  6222=>"111000000",
  6223=>"111111111",
  6224=>"110110110",
  6225=>"000000101",
  6226=>"100000110",
  6227=>"110111111",
  6228=>"000000000",
  6229=>"111111110",
  6230=>"111111100",
  6231=>"000000000",
  6232=>"000000110",
  6233=>"101000101",
  6234=>"001001111",
  6235=>"011000000",
  6236=>"111111111",
  6237=>"111100000",
  6238=>"000000000",
  6239=>"011000100",
  6240=>"000000000",
  6241=>"010110111",
  6242=>"000111110",
  6243=>"000000000",
  6244=>"110011000",
  6245=>"000000000",
  6246=>"010000000",
  6247=>"000000000",
  6248=>"111000000",
  6249=>"111100110",
  6250=>"010111111",
  6251=>"000000000",
  6252=>"000000000",
  6253=>"101000000",
  6254=>"111111111",
  6255=>"101111111",
  6256=>"000111100",
  6257=>"000001001",
  6258=>"111101100",
  6259=>"011010110",
  6260=>"000000000",
  6261=>"111111001",
  6262=>"001001111",
  6263=>"000000000",
  6264=>"001011000",
  6265=>"111111001",
  6266=>"000000000",
  6267=>"000000000",
  6268=>"101001011",
  6269=>"111111001",
  6270=>"001101100",
  6271=>"111111011",
  6272=>"111000000",
  6273=>"100110010",
  6274=>"110000000",
  6275=>"111111110",
  6276=>"111001001",
  6277=>"001000001",
  6278=>"000001111",
  6279=>"110110111",
  6280=>"111111111",
  6281=>"000000111",
  6282=>"011001111",
  6283=>"000111000",
  6284=>"000000001",
  6285=>"011011000",
  6286=>"111111000",
  6287=>"111110000",
  6288=>"000001011",
  6289=>"000000000",
  6290=>"000111111",
  6291=>"100100110",
  6292=>"010010010",
  6293=>"111001011",
  6294=>"000000110",
  6295=>"111111111",
  6296=>"000000111",
  6297=>"100001000",
  6298=>"000000000",
  6299=>"100100100",
  6300=>"100000000",
  6301=>"001010001",
  6302=>"011111111",
  6303=>"111010000",
  6304=>"000000000",
  6305=>"011000000",
  6306=>"011000010",
  6307=>"000000000",
  6308=>"000111001",
  6309=>"010111111",
  6310=>"000000000",
  6311=>"111111001",
  6312=>"000000000",
  6313=>"111111111",
  6314=>"000000000",
  6315=>"111111111",
  6316=>"011111000",
  6317=>"110100000",
  6318=>"111111111",
  6319=>"000000011",
  6320=>"000001111",
  6321=>"110000111",
  6322=>"110111110",
  6323=>"000000001",
  6324=>"011000101",
  6325=>"000101111",
  6326=>"000100111",
  6327=>"000110111",
  6328=>"111111111",
  6329=>"111111111",
  6330=>"000000000",
  6331=>"110110111",
  6332=>"000000111",
  6333=>"111111000",
  6334=>"111111111",
  6335=>"111110000",
  6336=>"010110111",
  6337=>"000111011",
  6338=>"000000001",
  6339=>"111011001",
  6340=>"000110111",
  6341=>"000000111",
  6342=>"111100000",
  6343=>"110010000",
  6344=>"001000011",
  6345=>"001010000",
  6346=>"011111111",
  6347=>"111111111",
  6348=>"111111011",
  6349=>"111110110",
  6350=>"111110000",
  6351=>"000010000",
  6352=>"101000000",
  6353=>"001100111",
  6354=>"111110111",
  6355=>"111110110",
  6356=>"000010111",
  6357=>"111110100",
  6358=>"000011111",
  6359=>"000111111",
  6360=>"000000000",
  6361=>"000111111",
  6362=>"111100110",
  6363=>"000000000",
  6364=>"001001011",
  6365=>"100111000",
  6366=>"000000111",
  6367=>"001110011",
  6368=>"111111111",
  6369=>"110111111",
  6370=>"000000000",
  6371=>"111111100",
  6372=>"000001000",
  6373=>"100110111",
  6374=>"000000100",
  6375=>"001001011",
  6376=>"110100011",
  6377=>"011011111",
  6378=>"111111000",
  6379=>"010010111",
  6380=>"000000000",
  6381=>"000001111",
  6382=>"000110111",
  6383=>"000000111",
  6384=>"100100000",
  6385=>"000111111",
  6386=>"111000000",
  6387=>"111111111",
  6388=>"100110110",
  6389=>"000000000",
  6390=>"000000000",
  6391=>"011001000",
  6392=>"111111111",
  6393=>"110111111",
  6394=>"000111111",
  6395=>"001000000",
  6396=>"011111110",
  6397=>"001001001",
  6398=>"110111000",
  6399=>"001001000",
  6400=>"101111000",
  6401=>"011000000",
  6402=>"000000000",
  6403=>"010100000",
  6404=>"010010010",
  6405=>"001001101",
  6406=>"000000111",
  6407=>"000001111",
  6408=>"111111111",
  6409=>"000000000",
  6410=>"000000100",
  6411=>"111011000",
  6412=>"111000000",
  6413=>"000001001",
  6414=>"000000011",
  6415=>"000101111",
  6416=>"100110110",
  6417=>"000000100",
  6418=>"111111111",
  6419=>"000000000",
  6420=>"000000111",
  6421=>"000000111",
  6422=>"011011010",
  6423=>"000000000",
  6424=>"110111010",
  6425=>"110111111",
  6426=>"110010110",
  6427=>"111001111",
  6428=>"011001000",
  6429=>"000000011",
  6430=>"000000000",
  6431=>"111110111",
  6432=>"000000000",
  6433=>"000000011",
  6434=>"111111000",
  6435=>"111100111",
  6436=>"001001000",
  6437=>"111111111",
  6438=>"111111111",
  6439=>"000100100",
  6440=>"000000111",
  6441=>"000000000",
  6442=>"000110111",
  6443=>"000000001",
  6444=>"111111111",
  6445=>"001111111",
  6446=>"000011111",
  6447=>"100111110",
  6448=>"111111111",
  6449=>"111111110",
  6450=>"000000000",
  6451=>"110000111",
  6452=>"000000000",
  6453=>"000000000",
  6454=>"111110100",
  6455=>"001000000",
  6456=>"000001111",
  6457=>"101000111",
  6458=>"001001000",
  6459=>"000101000",
  6460=>"000000000",
  6461=>"010011111",
  6462=>"000010010",
  6463=>"000000010",
  6464=>"011011001",
  6465=>"110111111",
  6466=>"000110111",
  6467=>"101000000",
  6468=>"001001000",
  6469=>"000010000",
  6470=>"000110110",
  6471=>"001000000",
  6472=>"000000000",
  6473=>"000000111",
  6474=>"111111111",
  6475=>"100000111",
  6476=>"000000110",
  6477=>"111111000",
  6478=>"111111111",
  6479=>"000011011",
  6480=>"110000000",
  6481=>"110000000",
  6482=>"111111010",
  6483=>"000110110",
  6484=>"000111111",
  6485=>"011011011",
  6486=>"000000000",
  6487=>"100110000",
  6488=>"000000000",
  6489=>"000000100",
  6490=>"110000000",
  6491=>"000000000",
  6492=>"000000000",
  6493=>"111111111",
  6494=>"001000101",
  6495=>"001111010",
  6496=>"000000000",
  6497=>"000110111",
  6498=>"011111111",
  6499=>"111000000",
  6500=>"000000000",
  6501=>"000000000",
  6502=>"000000111",
  6503=>"011111110",
  6504=>"000000000",
  6505=>"100110110",
  6506=>"111111000",
  6507=>"011111111",
  6508=>"000000110",
  6509=>"000011000",
  6510=>"000000000",
  6511=>"000000110",
  6512=>"000000111",
  6513=>"111111100",
  6514=>"000111111",
  6515=>"011111001",
  6516=>"000000000",
  6517=>"001000000",
  6518=>"000000000",
  6519=>"010010000",
  6520=>"000000011",
  6521=>"111011111",
  6522=>"111111111",
  6523=>"000000110",
  6524=>"110100111",
  6525=>"001010111",
  6526=>"111111111",
  6527=>"000000000",
  6528=>"110110100",
  6529=>"111110000",
  6530=>"001001000",
  6531=>"000000000",
  6532=>"111111010",
  6533=>"111111111",
  6534=>"110110110",
  6535=>"011111111",
  6536=>"111111111",
  6537=>"110111011",
  6538=>"000000000",
  6539=>"010000101",
  6540=>"111000111",
  6541=>"000000000",
  6542=>"100100000",
  6543=>"111111111",
  6544=>"000000000",
  6545=>"011111110",
  6546=>"001000001",
  6547=>"000000000",
  6548=>"111111111",
  6549=>"000001000",
  6550=>"011111000",
  6551=>"000000000",
  6552=>"111011111",
  6553=>"111110110",
  6554=>"100000000",
  6555=>"000000101",
  6556=>"100000000",
  6557=>"001111111",
  6558=>"000000000",
  6559=>"000000000",
  6560=>"110110000",
  6561=>"110100000",
  6562=>"000000000",
  6563=>"000000000",
  6564=>"001000001",
  6565=>"000101111",
  6566=>"111000000",
  6567=>"110110100",
  6568=>"000000000",
  6569=>"000111010",
  6570=>"000010000",
  6571=>"001000001",
  6572=>"000000000",
  6573=>"001000111",
  6574=>"000000000",
  6575=>"000000000",
  6576=>"001111111",
  6577=>"011001000",
  6578=>"001001111",
  6579=>"000111111",
  6580=>"000100000",
  6581=>"111111111",
  6582=>"000000000",
  6583=>"000000000",
  6584=>"011000000",
  6585=>"000010010",
  6586=>"000110111",
  6587=>"100000111",
  6588=>"011000011",
  6589=>"111111111",
  6590=>"111011011",
  6591=>"001000000",
  6592=>"111110110",
  6593=>"111111111",
  6594=>"111111111",
  6595=>"000000000",
  6596=>"001001000",
  6597=>"000000000",
  6598=>"000000000",
  6599=>"011011000",
  6600=>"001000100",
  6601=>"000000000",
  6602=>"000000111",
  6603=>"010111000",
  6604=>"000001011",
  6605=>"100110000",
  6606=>"001000011",
  6607=>"000000000",
  6608=>"000000011",
  6609=>"111111111",
  6610=>"110000000",
  6611=>"111111111",
  6612=>"000001111",
  6613=>"000010000",
  6614=>"000010000",
  6615=>"110011000",
  6616=>"000010010",
  6617=>"001011011",
  6618=>"000000000",
  6619=>"000111000",
  6620=>"111111111",
  6621=>"111111111",
  6622=>"000000000",
  6623=>"000000000",
  6624=>"011001000",
  6625=>"111110110",
  6626=>"010110110",
  6627=>"001011000",
  6628=>"111111000",
  6629=>"001000000",
  6630=>"000110111",
  6631=>"100100111",
  6632=>"111111011",
  6633=>"001000000",
  6634=>"100110010",
  6635=>"111111001",
  6636=>"000111111",
  6637=>"001011001",
  6638=>"111001000",
  6639=>"001111111",
  6640=>"000000000",
  6641=>"111100000",
  6642=>"100000000",
  6643=>"100111001",
  6644=>"001111000",
  6645=>"110011010",
  6646=>"111111110",
  6647=>"110100111",
  6648=>"000000000",
  6649=>"101111011",
  6650=>"001011111",
  6651=>"011001111",
  6652=>"111111111",
  6653=>"000110110",
  6654=>"000000000",
  6655=>"000000000",
  6656=>"111111110",
  6657=>"011000000",
  6658=>"000001100",
  6659=>"111111111",
  6660=>"111111111",
  6661=>"011001000",
  6662=>"000000100",
  6663=>"111011011",
  6664=>"111111000",
  6665=>"000001011",
  6666=>"100100111",
  6667=>"111111000",
  6668=>"100100100",
  6669=>"000001011",
  6670=>"001000000",
  6671=>"000000000",
  6672=>"111000000",
  6673=>"000000100",
  6674=>"000000000",
  6675=>"000000010",
  6676=>"000111111",
  6677=>"111111111",
  6678=>"111011000",
  6679=>"111110000",
  6680=>"110110000",
  6681=>"100100001",
  6682=>"111110000",
  6683=>"001000100",
  6684=>"100111100",
  6685=>"111111000",
  6686=>"110111110",
  6687=>"111111000",
  6688=>"111111111",
  6689=>"000000001",
  6690=>"111111111",
  6691=>"001001111",
  6692=>"100111111",
  6693=>"000001111",
  6694=>"000000000",
  6695=>"111111100",
  6696=>"000000111",
  6697=>"000000110",
  6698=>"000000000",
  6699=>"000000000",
  6700=>"000000000",
  6701=>"111111001",
  6702=>"000000100",
  6703=>"000111111",
  6704=>"110000110",
  6705=>"111111011",
  6706=>"000100010",
  6707=>"111111111",
  6708=>"111111111",
  6709=>"010000000",
  6710=>"111111000",
  6711=>"111111111",
  6712=>"000100110",
  6713=>"001000110",
  6714=>"100100000",
  6715=>"100110000",
  6716=>"111001000",
  6717=>"011111111",
  6718=>"111111111",
  6719=>"000111111",
  6720=>"000000000",
  6721=>"101111111",
  6722=>"111111111",
  6723=>"111111111",
  6724=>"110001001",
  6725=>"000000101",
  6726=>"000000000",
  6727=>"000000000",
  6728=>"000000000",
  6729=>"100000100",
  6730=>"111001111",
  6731=>"000000111",
  6732=>"010000000",
  6733=>"111111100",
  6734=>"000000101",
  6735=>"000000000",
  6736=>"101000000",
  6737=>"111111011",
  6738=>"000000000",
  6739=>"000000000",
  6740=>"110010000",
  6741=>"000000000",
  6742=>"111111111",
  6743=>"000000000",
  6744=>"100000000",
  6745=>"000000111",
  6746=>"111111111",
  6747=>"011111111",
  6748=>"000100100",
  6749=>"111111111",
  6750=>"000011000",
  6751=>"111111111",
  6752=>"111000000",
  6753=>"111111001",
  6754=>"111111111",
  6755=>"000000101",
  6756=>"111000110",
  6757=>"111000110",
  6758=>"111011011",
  6759=>"000000111",
  6760=>"111111100",
  6761=>"100000000",
  6762=>"111111111",
  6763=>"000000000",
  6764=>"001111111",
  6765=>"000111111",
  6766=>"000000000",
  6767=>"000000000",
  6768=>"111111111",
  6769=>"101110111",
  6770=>"111100000",
  6771=>"000000000",
  6772=>"000000000",
  6773=>"010110111",
  6774=>"000000000",
  6775=>"000111100",
  6776=>"111011000",
  6777=>"111011111",
  6778=>"000000000",
  6779=>"000101111",
  6780=>"111111110",
  6781=>"111111001",
  6782=>"000000000",
  6783=>"110110111",
  6784=>"000001000",
  6785=>"000000000",
  6786=>"111111111",
  6787=>"101111000",
  6788=>"111111111",
  6789=>"100000001",
  6790=>"100111011",
  6791=>"000000100",
  6792=>"111111100",
  6793=>"000000000",
  6794=>"111110000",
  6795=>"100110111",
  6796=>"000000111",
  6797=>"001111000",
  6798=>"010000000",
  6799=>"000000111",
  6800=>"000000000",
  6801=>"000000011",
  6802=>"011000000",
  6803=>"111111000",
  6804=>"111110100",
  6805=>"000000000",
  6806=>"101000000",
  6807=>"011011111",
  6808=>"000000010",
  6809=>"000111111",
  6810=>"010111111",
  6811=>"111111100",
  6812=>"101000111",
  6813=>"011000000",
  6814=>"000000011",
  6815=>"111111111",
  6816=>"111001111",
  6817=>"111101000",
  6818=>"001000000",
  6819=>"111000000",
  6820=>"000000000",
  6821=>"111100111",
  6822=>"111101111",
  6823=>"111110100",
  6824=>"111111111",
  6825=>"010010111",
  6826=>"100000111",
  6827=>"101101001",
  6828=>"001000000",
  6829=>"000000000",
  6830=>"111111111",
  6831=>"000000111",
  6832=>"000000000",
  6833=>"000000000",
  6834=>"111111111",
  6835=>"010100101",
  6836=>"010010000",
  6837=>"011111111",
  6838=>"000111111",
  6839=>"000000001",
  6840=>"000111111",
  6841=>"011111110",
  6842=>"000000001",
  6843=>"111000100",
  6844=>"000111111",
  6845=>"111111000",
  6846=>"111111110",
  6847=>"001111100",
  6848=>"111111100",
  6849=>"000001111",
  6850=>"111111111",
  6851=>"000111111",
  6852=>"001111111",
  6853=>"011001111",
  6854=>"100111011",
  6855=>"000000000",
  6856=>"001000100",
  6857=>"111111111",
  6858=>"100001001",
  6859=>"000000001",
  6860=>"111111001",
  6861=>"000111110",
  6862=>"111111111",
  6863=>"000000100",
  6864=>"000111100",
  6865=>"111111111",
  6866=>"100000000",
  6867=>"100111111",
  6868=>"111111101",
  6869=>"111111111",
  6870=>"000000000",
  6871=>"111111110",
  6872=>"000000111",
  6873=>"100111110",
  6874=>"111001110",
  6875=>"000000000",
  6876=>"111111110",
  6877=>"000000000",
  6878=>"000000100",
  6879=>"010000001",
  6880=>"000000000",
  6881=>"101101000",
  6882=>"111000000",
  6883=>"000100111",
  6884=>"111111101",
  6885=>"100111111",
  6886=>"111110010",
  6887=>"110110111",
  6888=>"111111111",
  6889=>"000000000",
  6890=>"001000000",
  6891=>"000100100",
  6892=>"111000011",
  6893=>"101000000",
  6894=>"111011111",
  6895=>"000011011",
  6896=>"001001000",
  6897=>"000000001",
  6898=>"111110110",
  6899=>"000000111",
  6900=>"111011000",
  6901=>"100111111",
  6902=>"000000000",
  6903=>"010110110",
  6904=>"111111111",
  6905=>"110000000",
  6906=>"010111111",
  6907=>"111010000",
  6908=>"000000001",
  6909=>"110111010",
  6910=>"000000000",
  6911=>"010000111",
  6912=>"000000000",
  6913=>"111110110",
  6914=>"111000000",
  6915=>"111110100",
  6916=>"000001000",
  6917=>"000110111",
  6918=>"110111111",
  6919=>"111101111",
  6920=>"000000000",
  6921=>"000000000",
  6922=>"111111000",
  6923=>"111101001",
  6924=>"111101111",
  6925=>"001000111",
  6926=>"001110111",
  6927=>"001000000",
  6928=>"011001000",
  6929=>"111110000",
  6930=>"000000001",
  6931=>"010001000",
  6932=>"111111111",
  6933=>"000000000",
  6934=>"010111111",
  6935=>"000000000",
  6936=>"111111001",
  6937=>"001001011",
  6938=>"111001000",
  6939=>"000001001",
  6940=>"111111100",
  6941=>"100000000",
  6942=>"000001101",
  6943=>"000100111",
  6944=>"110111000",
  6945=>"000000111",
  6946=>"001001000",
  6947=>"111000110",
  6948=>"011110110",
  6949=>"111111111",
  6950=>"011111110",
  6951=>"001111111",
  6952=>"000100111",
  6953=>"100000000",
  6954=>"001000000",
  6955=>"000000000",
  6956=>"000000000",
  6957=>"110000000",
  6958=>"101111001",
  6959=>"111111011",
  6960=>"110011000",
  6961=>"111111110",
  6962=>"111111111",
  6963=>"000000000",
  6964=>"111111111",
  6965=>"000000000",
  6966=>"000000111",
  6967=>"000000110",
  6968=>"000111111",
  6969=>"000000111",
  6970=>"111111111",
  6971=>"111111000",
  6972=>"001000000",
  6973=>"100000000",
  6974=>"000000100",
  6975=>"000000000",
  6976=>"000000000",
  6977=>"111000000",
  6978=>"100000000",
  6979=>"000111111",
  6980=>"110111111",
  6981=>"111111000",
  6982=>"111111111",
  6983=>"000000000",
  6984=>"111100010",
  6985=>"010010010",
  6986=>"000111111",
  6987=>"011111111",
  6988=>"000000000",
  6989=>"111111100",
  6990=>"100111011",
  6991=>"010000000",
  6992=>"111111101",
  6993=>"001001111",
  6994=>"000000111",
  6995=>"000000000",
  6996=>"000000000",
  6997=>"011010000",
  6998=>"111111110",
  6999=>"000000000",
  7000=>"111111111",
  7001=>"111010000",
  7002=>"111000000",
  7003=>"010001001",
  7004=>"011011111",
  7005=>"000000000",
  7006=>"011011111",
  7007=>"100001001",
  7008=>"011000101",
  7009=>"000000000",
  7010=>"110110111",
  7011=>"111111000",
  7012=>"111111000",
  7013=>"001001000",
  7014=>"011000011",
  7015=>"001111110",
  7016=>"001001101",
  7017=>"111111110",
  7018=>"000100111",
  7019=>"110110110",
  7020=>"110111011",
  7021=>"000000000",
  7022=>"000000000",
  7023=>"110000010",
  7024=>"011111000",
  7025=>"111010000",
  7026=>"000000000",
  7027=>"110111011",
  7028=>"000100110",
  7029=>"000000000",
  7030=>"111111101",
  7031=>"111110000",
  7032=>"000000111",
  7033=>"111110100",
  7034=>"000000100",
  7035=>"111111111",
  7036=>"000100111",
  7037=>"000000111",
  7038=>"111000111",
  7039=>"000001001",
  7040=>"000000100",
  7041=>"000101111",
  7042=>"000000110",
  7043=>"000111111",
  7044=>"000000111",
  7045=>"000000000",
  7046=>"001001111",
  7047=>"111010000",
  7048=>"111111101",
  7049=>"111110000",
  7050=>"000000000",
  7051=>"000000000",
  7052=>"000000111",
  7053=>"110110111",
  7054=>"111000101",
  7055=>"000000000",
  7056=>"000000000",
  7057=>"011100001",
  7058=>"110111100",
  7059=>"111111111",
  7060=>"011000010",
  7061=>"100110000",
  7062=>"001111111",
  7063=>"001111111",
  7064=>"011011000",
  7065=>"111111111",
  7066=>"000000101",
  7067=>"111111111",
  7068=>"000000111",
  7069=>"111111111",
  7070=>"011111111",
  7071=>"111111111",
  7072=>"000001111",
  7073=>"001111011",
  7074=>"111001000",
  7075=>"001111011",
  7076=>"111111101",
  7077=>"011010000",
  7078=>"000000111",
  7079=>"001000000",
  7080=>"111111111",
  7081=>"011110110",
  7082=>"000100111",
  7083=>"000000011",
  7084=>"000000000",
  7085=>"111100000",
  7086=>"000000100",
  7087=>"000000000",
  7088=>"000000100",
  7089=>"000110111",
  7090=>"011001111",
  7091=>"000000001",
  7092=>"111101000",
  7093=>"111111000",
  7094=>"000001001",
  7095=>"000110111",
  7096=>"000000110",
  7097=>"010000000",
  7098=>"100000000",
  7099=>"101000000",
  7100=>"000110111",
  7101=>"000000001",
  7102=>"111000000",
  7103=>"001111111",
  7104=>"000000000",
  7105=>"000000111",
  7106=>"111000000",
  7107=>"111111000",
  7108=>"111111111",
  7109=>"110000000",
  7110=>"000001110",
  7111=>"111001000",
  7112=>"000000111",
  7113=>"000000000",
  7114=>"000100110",
  7115=>"101000000",
  7116=>"000000000",
  7117=>"000000000",
  7118=>"000000001",
  7119=>"000001111",
  7120=>"000111111",
  7121=>"111100000",
  7122=>"001101100",
  7123=>"001000000",
  7124=>"110100000",
  7125=>"111111111",
  7126=>"001111000",
  7127=>"111111111",
  7128=>"000111111",
  7129=>"011100111",
  7130=>"111111010",
  7131=>"000000111",
  7132=>"111111111",
  7133=>"000000111",
  7134=>"110111111",
  7135=>"000000000",
  7136=>"110111110",
  7137=>"000111111",
  7138=>"000000000",
  7139=>"000000011",
  7140=>"010011111",
  7141=>"011010000",
  7142=>"111111111",
  7143=>"000000000",
  7144=>"000000000",
  7145=>"010111011",
  7146=>"111111101",
  7147=>"001000000",
  7148=>"111110100",
  7149=>"000100100",
  7150=>"000100111",
  7151=>"011010000",
  7152=>"000000001",
  7153=>"111111110",
  7154=>"111111111",
  7155=>"111111111",
  7156=>"111001000",
  7157=>"000001111",
  7158=>"111001001",
  7159=>"111111100",
  7160=>"000111111",
  7161=>"101101111",
  7162=>"100000000",
  7163=>"111111111",
  7164=>"000000100",
  7165=>"111000000",
  7166=>"000000000",
  7167=>"100000000",
  7168=>"101111111",
  7169=>"000001000",
  7170=>"000101000",
  7171=>"000000000",
  7172=>"001001001",
  7173=>"110111001",
  7174=>"111111111",
  7175=>"000101000",
  7176=>"000000000",
  7177=>"100110110",
  7178=>"000111000",
  7179=>"000000000",
  7180=>"001110010",
  7181=>"000110111",
  7182=>"010110111",
  7183=>"111111111",
  7184=>"010011111",
  7185=>"111010000",
  7186=>"111100111",
  7187=>"000111111",
  7188=>"000000000",
  7189=>"111011000",
  7190=>"111111111",
  7191=>"100100111",
  7192=>"011111110",
  7193=>"111111001",
  7194=>"000000111",
  7195=>"000000000",
  7196=>"000000000",
  7197=>"111111111",
  7198=>"001000011",
  7199=>"011110000",
  7200=>"000101000",
  7201=>"111111111",
  7202=>"001001001",
  7203=>"111011111",
  7204=>"111000111",
  7205=>"000000000",
  7206=>"000001111",
  7207=>"111100000",
  7208=>"101001111",
  7209=>"011001000",
  7210=>"011111000",
  7211=>"000111111",
  7212=>"100000111",
  7213=>"101100111",
  7214=>"010111011",
  7215=>"000101111",
  7216=>"000000000",
  7217=>"111000011",
  7218=>"000100111",
  7219=>"111111111",
  7220=>"101011111",
  7221=>"100001101",
  7222=>"000100001",
  7223=>"100101111",
  7224=>"000000111",
  7225=>"001000000",
  7226=>"001000000",
  7227=>"000000000",
  7228=>"000000111",
  7229=>"000000000",
  7230=>"111111111",
  7231=>"000111111",
  7232=>"000000000",
  7233=>"010010110",
  7234=>"110110000",
  7235=>"001000101",
  7236=>"000000000",
  7237=>"011001001",
  7238=>"111111000",
  7239=>"111111111",
  7240=>"110100110",
  7241=>"100100100",
  7242=>"111111111",
  7243=>"001001000",
  7244=>"000000000",
  7245=>"000000101",
  7246=>"100100000",
  7247=>"000000111",
  7248=>"000001000",
  7249=>"000000001",
  7250=>"000001100",
  7251=>"011101000",
  7252=>"101111111",
  7253=>"101000111",
  7254=>"000111100",
  7255=>"111001111",
  7256=>"000111011",
  7257=>"000111000",
  7258=>"000010011",
  7259=>"100100000",
  7260=>"000110000",
  7261=>"000000101",
  7262=>"111111011",
  7263=>"111111001",
  7264=>"000100000",
  7265=>"000001001",
  7266=>"111011011",
  7267=>"010010000",
  7268=>"111111111",
  7269=>"000111100",
  7270=>"000000000",
  7271=>"100000101",
  7272=>"000111111",
  7273=>"000000001",
  7274=>"010000110",
  7275=>"111111000",
  7276=>"111111111",
  7277=>"111111111",
  7278=>"110011011",
  7279=>"111000001",
  7280=>"000001001",
  7281=>"000000101",
  7282=>"101010010",
  7283=>"000001000",
  7284=>"000011111",
  7285=>"111111111",
  7286=>"000110111",
  7287=>"111111111",
  7288=>"000110000",
  7289=>"111111111",
  7290=>"111111111",
  7291=>"000000111",
  7292=>"000001001",
  7293=>"100001111",
  7294=>"110111111",
  7295=>"011000000",
  7296=>"000100111",
  7297=>"100101101",
  7298=>"000000000",
  7299=>"011110000",
  7300=>"111001011",
  7301=>"111000111",
  7302=>"111111000",
  7303=>"001001000",
  7304=>"011111111",
  7305=>"000100111",
  7306=>"000000001",
  7307=>"111111111",
  7308=>"111011000",
  7309=>"010011111",
  7310=>"111000000",
  7311=>"001100111",
  7312=>"000110110",
  7313=>"110110000",
  7314=>"001001111",
  7315=>"000000000",
  7316=>"111101001",
  7317=>"111111000",
  7318=>"000000000",
  7319=>"000111000",
  7320=>"000101111",
  7321=>"111111111",
  7322=>"100000111",
  7323=>"000000000",
  7324=>"100100000",
  7325=>"000101000",
  7326=>"000000111",
  7327=>"111111111",
  7328=>"101111111",
  7329=>"111111000",
  7330=>"000010001",
  7331=>"000001000",
  7332=>"000100101",
  7333=>"111100011",
  7334=>"111010111",
  7335=>"001000111",
  7336=>"000111000",
  7337=>"000000000",
  7338=>"001111111",
  7339=>"010111000",
  7340=>"001001111",
  7341=>"001000100",
  7342=>"110111011",
  7343=>"001001001",
  7344=>"000111000",
  7345=>"111111110",
  7346=>"110110111",
  7347=>"111000111",
  7348=>"111111000",
  7349=>"011110110",
  7350=>"111111111",
  7351=>"000000000",
  7352=>"000000001",
  7353=>"111110110",
  7354=>"110001101",
  7355=>"000101101",
  7356=>"011111111",
  7357=>"001111111",
  7358=>"000101111",
  7359=>"010010000",
  7360=>"111111000",
  7361=>"000000000",
  7362=>"111111000",
  7363=>"000101001",
  7364=>"011011001",
  7365=>"000000111",
  7366=>"111111111",
  7367=>"000011011",
  7368=>"100111111",
  7369=>"000000000",
  7370=>"111000011",
  7371=>"111111111",
  7372=>"000100000",
  7373=>"111000111",
  7374=>"001111011",
  7375=>"111101000",
  7376=>"000101000",
  7377=>"111111001",
  7378=>"110111000",
  7379=>"000000000",
  7380=>"011000011",
  7381=>"001001011",
  7382=>"000000000",
  7383=>"100101111",
  7384=>"111111001",
  7385=>"000001101",
  7386=>"000111111",
  7387=>"000111111",
  7388=>"000001000",
  7389=>"000111011",
  7390=>"010010000",
  7391=>"000000000",
  7392=>"000010000",
  7393=>"011011111",
  7394=>"111110000",
  7395=>"000000000",
  7396=>"000000110",
  7397=>"001000000",
  7398=>"111111111",
  7399=>"001111111",
  7400=>"001000000",
  7401=>"111111111",
  7402=>"111000001",
  7403=>"111111001",
  7404=>"010010010",
  7405=>"111111011",
  7406=>"001111000",
  7407=>"001111111",
  7408=>"111000111",
  7409=>"000110100",
  7410=>"001011000",
  7411=>"000101111",
  7412=>"111101111",
  7413=>"110000100",
  7414=>"110000101",
  7415=>"001001001",
  7416=>"110000000",
  7417=>"000000000",
  7418=>"000110000",
  7419=>"111111111",
  7420=>"111100110",
  7421=>"010011011",
  7422=>"001001000",
  7423=>"100111111",
  7424=>"000000111",
  7425=>"011011111",
  7426=>"000000000",
  7427=>"000001011",
  7428=>"000000001",
  7429=>"111111000",
  7430=>"000000001",
  7431=>"001100001",
  7432=>"000000100",
  7433=>"111111111",
  7434=>"000000000",
  7435=>"001111111",
  7436=>"000100110",
  7437=>"001111111",
  7438=>"101111000",
  7439=>"011111101",
  7440=>"000000110",
  7441=>"000100000",
  7442=>"110010111",
  7443=>"100111111",
  7444=>"111111000",
  7445=>"011001000",
  7446=>"111110110",
  7447=>"111101100",
  7448=>"111001001",
  7449=>"000000111",
  7450=>"000000000",
  7451=>"100110100",
  7452=>"111011111",
  7453=>"000000001",
  7454=>"111111111",
  7455=>"000111000",
  7456=>"111111101",
  7457=>"000111000",
  7458=>"110000100",
  7459=>"100100001",
  7460=>"010110110",
  7461=>"111111000",
  7462=>"000111011",
  7463=>"011011011",
  7464=>"101111111",
  7465=>"111010011",
  7466=>"001001001",
  7467=>"001101000",
  7468=>"000000100",
  7469=>"111001101",
  7470=>"010111000",
  7471=>"000000000",
  7472=>"000000000",
  7473=>"000000111",
  7474=>"100111100",
  7475=>"000000000",
  7476=>"000000000",
  7477=>"100101000",
  7478=>"001111111",
  7479=>"111111100",
  7480=>"100111111",
  7481=>"111111100",
  7482=>"110100111",
  7483=>"001000000",
  7484=>"000001000",
  7485=>"001000000",
  7486=>"000111111",
  7487=>"111111010",
  7488=>"000011001",
  7489=>"000000111",
  7490=>"000111101",
  7491=>"000000100",
  7492=>"100111111",
  7493=>"000000000",
  7494=>"110100111",
  7495=>"110110110",
  7496=>"000111110",
  7497=>"000111000",
  7498=>"011111001",
  7499=>"001000000",
  7500=>"111111000",
  7501=>"111101111",
  7502=>"001111101",
  7503=>"011011100",
  7504=>"000000111",
  7505=>"111111101",
  7506=>"000000111",
  7507=>"011011001",
  7508=>"000000111",
  7509=>"000000000",
  7510=>"111110111",
  7511=>"000000111",
  7512=>"111101000",
  7513=>"000110000",
  7514=>"011111111",
  7515=>"111110100",
  7516=>"000000000",
  7517=>"111111110",
  7518=>"111111000",
  7519=>"111111101",
  7520=>"000000000",
  7521=>"011000111",
  7522=>"000100100",
  7523=>"000000000",
  7524=>"110111111",
  7525=>"000001001",
  7526=>"000000111",
  7527=>"101101001",
  7528=>"110111000",
  7529=>"110110011",
  7530=>"111010111",
  7531=>"111100100",
  7532=>"001001000",
  7533=>"010111111",
  7534=>"111111000",
  7535=>"000000000",
  7536=>"111111000",
  7537=>"000000111",
  7538=>"000001001",
  7539=>"111110110",
  7540=>"111111001",
  7541=>"111111111",
  7542=>"000111010",
  7543=>"001001011",
  7544=>"111111111",
  7545=>"000010000",
  7546=>"111000000",
  7547=>"000111101",
  7548=>"111111010",
  7549=>"000000111",
  7550=>"110100000",
  7551=>"000000000",
  7552=>"100110000",
  7553=>"111111111",
  7554=>"100000000",
  7555=>"011111000",
  7556=>"000100000",
  7557=>"000000010",
  7558=>"000000010",
  7559=>"110110000",
  7560=>"000010000",
  7561=>"000011000",
  7562=>"001000001",
  7563=>"000010000",
  7564=>"001111111",
  7565=>"011101110",
  7566=>"111111111",
  7567=>"111111111",
  7568=>"000100110",
  7569=>"100101000",
  7570=>"100000011",
  7571=>"000000000",
  7572=>"000000000",
  7573=>"000000100",
  7574=>"111010011",
  7575=>"000101000",
  7576=>"011001001",
  7577=>"111111011",
  7578=>"111111110",
  7579=>"010011111",
  7580=>"111111110",
  7581=>"111111110",
  7582=>"110100111",
  7583=>"000000000",
  7584=>"111111111",
  7585=>"001100110",
  7586=>"001111110",
  7587=>"000011111",
  7588=>"000000000",
  7589=>"000111111",
  7590=>"000000000",
  7591=>"000111000",
  7592=>"000000000",
  7593=>"000000111",
  7594=>"000010000",
  7595=>"111111011",
  7596=>"000000011",
  7597=>"011111000",
  7598=>"000011011",
  7599=>"110100000",
  7600=>"111000011",
  7601=>"000000001",
  7602=>"011001000",
  7603=>"000000000",
  7604=>"000000000",
  7605=>"000000000",
  7606=>"000010100",
  7607=>"000000000",
  7608=>"100010111",
  7609=>"000000111",
  7610=>"001111111",
  7611=>"100101000",
  7612=>"111111010",
  7613=>"111011001",
  7614=>"111111111",
  7615=>"100101101",
  7616=>"111100011",
  7617=>"010111111",
  7618=>"000000000",
  7619=>"110110100",
  7620=>"000000100",
  7621=>"110110100",
  7622=>"111111111",
  7623=>"001111101",
  7624=>"000000111",
  7625=>"111111011",
  7626=>"000000000",
  7627=>"111000000",
  7628=>"111111000",
  7629=>"000000111",
  7630=>"000000101",
  7631=>"111011000",
  7632=>"000101000",
  7633=>"100110110",
  7634=>"000000000",
  7635=>"000000111",
  7636=>"000101111",
  7637=>"000100111",
  7638=>"111111111",
  7639=>"000110000",
  7640=>"000111110",
  7641=>"001001110",
  7642=>"111111000",
  7643=>"000100010",
  7644=>"011010010",
  7645=>"001101000",
  7646=>"000111000",
  7647=>"110100100",
  7648=>"111001001",
  7649=>"110000111",
  7650=>"111000000",
  7651=>"000000101",
  7652=>"000100111",
  7653=>"001111111",
  7654=>"111111000",
  7655=>"001111111",
  7656=>"100000000",
  7657=>"001111111",
  7658=>"000001101",
  7659=>"111111111",
  7660=>"011111000",
  7661=>"000000011",
  7662=>"000000100",
  7663=>"000000000",
  7664=>"111010111",
  7665=>"111111110",
  7666=>"100110111",
  7667=>"111111111",
  7668=>"111111111",
  7669=>"000001000",
  7670=>"000110110",
  7671=>"111001001",
  7672=>"000000000",
  7673=>"001101000",
  7674=>"111111111",
  7675=>"000011111",
  7676=>"111111111",
  7677=>"011000000",
  7678=>"111101101",
  7679=>"010011011",
  7680=>"111110110",
  7681=>"111111011",
  7682=>"111001000",
  7683=>"000000000",
  7684=>"001000000",
  7685=>"000000000",
  7686=>"111011000",
  7687=>"000000000",
  7688=>"111111000",
  7689=>"011000110",
  7690=>"000001011",
  7691=>"111000001",
  7692=>"111111111",
  7693=>"111111111",
  7694=>"111111111",
  7695=>"111111111",
  7696=>"000101111",
  7697=>"111110100",
  7698=>"000011111",
  7699=>"100000000",
  7700=>"010000011",
  7701=>"000000000",
  7702=>"000100001",
  7703=>"000101101",
  7704=>"111111011",
  7705=>"101000011",
  7706=>"100000000",
  7707=>"111111111",
  7708=>"101111111",
  7709=>"101101000",
  7710=>"000001101",
  7711=>"000000000",
  7712=>"100000001",
  7713=>"101111111",
  7714=>"111111111",
  7715=>"000000100",
  7716=>"001000001",
  7717=>"111110111",
  7718=>"111111101",
  7719=>"111010001",
  7720=>"111111111",
  7721=>"000000000",
  7722=>"000000000",
  7723=>"110110111",
  7724=>"000001000",
  7725=>"000111111",
  7726=>"101011000",
  7727=>"001111111",
  7728=>"100110111",
  7729=>"111111111",
  7730=>"001011101",
  7731=>"000000001",
  7732=>"000000000",
  7733=>"111111111",
  7734=>"001011011",
  7735=>"111101111",
  7736=>"000000111",
  7737=>"000000000",
  7738=>"000000000",
  7739=>"000000100",
  7740=>"111101000",
  7741=>"011011001",
  7742=>"100100100",
  7743=>"000000000",
  7744=>"000000000",
  7745=>"100111111",
  7746=>"000000111",
  7747=>"111111111",
  7748=>"111110011",
  7749=>"001001001",
  7750=>"001000000",
  7751=>"111111111",
  7752=>"111111111",
  7753=>"001001111",
  7754=>"001101101",
  7755=>"100000000",
  7756=>"000000000",
  7757=>"111111100",
  7758=>"101001101",
  7759=>"000000110",
  7760=>"001111100",
  7761=>"111001100",
  7762=>"111011000",
  7763=>"111111100",
  7764=>"000000000",
  7765=>"100000000",
  7766=>"000000111",
  7767=>"111011001",
  7768=>"000000000",
  7769=>"001000000",
  7770=>"000000000",
  7771=>"001000110",
  7772=>"000000000",
  7773=>"000100000",
  7774=>"000011111",
  7775=>"001011111",
  7776=>"111111111",
  7777=>"111100110",
  7778=>"000000001",
  7779=>"111111111",
  7780=>"111111111",
  7781=>"001111111",
  7782=>"111100100",
  7783=>"000000000",
  7784=>"111111110",
  7785=>"110111111",
  7786=>"001000000",
  7787=>"111000000",
  7788=>"011111111",
  7789=>"111000000",
  7790=>"010000000",
  7791=>"001001000",
  7792=>"000110000",
  7793=>"000010111",
  7794=>"110100000",
  7795=>"111011011",
  7796=>"111111111",
  7797=>"111001000",
  7798=>"000000100",
  7799=>"001010000",
  7800=>"000000010",
  7801=>"111111111",
  7802=>"001000000",
  7803=>"111000000",
  7804=>"100100110",
  7805=>"111111111",
  7806=>"000000000",
  7807=>"001000000",
  7808=>"000000000",
  7809=>"111111111",
  7810=>"000100100",
  7811=>"100111111",
  7812=>"000000000",
  7813=>"110010000",
  7814=>"111111111",
  7815=>"111111111",
  7816=>"000000111",
  7817=>"000000000",
  7818=>"110110111",
  7819=>"011011010",
  7820=>"010110110",
  7821=>"000000000",
  7822=>"111011011",
  7823=>"000000000",
  7824=>"111111111",
  7825=>"000000000",
  7826=>"111111111",
  7827=>"000000000",
  7828=>"110101111",
  7829=>"001000000",
  7830=>"000000000",
  7831=>"000000000",
  7832=>"111111101",
  7833=>"000000000",
  7834=>"111111111",
  7835=>"000000000",
  7836=>"000001101",
  7837=>"000000100",
  7838=>"001111111",
  7839=>"111001001",
  7840=>"111001111",
  7841=>"111111111",
  7842=>"111111111",
  7843=>"111011011",
  7844=>"000000000",
  7845=>"111011000",
  7846=>"111111111",
  7847=>"111011011",
  7848=>"111111111",
  7849=>"100000111",
  7850=>"000000000",
  7851=>"000111111",
  7852=>"111110000",
  7853=>"011011111",
  7854=>"000000011",
  7855=>"001000111",
  7856=>"111111111",
  7857=>"101101100",
  7858=>"010010111",
  7859=>"100000111",
  7860=>"000001001",
  7861=>"000000000",
  7862=>"000000000",
  7863=>"111111111",
  7864=>"111111111",
  7865=>"000100101",
  7866=>"111111011",
  7867=>"110000111",
  7868=>"111111000",
  7869=>"111011100",
  7870=>"111111111",
  7871=>"100000000",
  7872=>"000000000",
  7873=>"000010000",
  7874=>"000000000",
  7875=>"101101100",
  7876=>"111111010",
  7877=>"001111111",
  7878=>"111111111",
  7879=>"000000000",
  7880=>"000110110",
  7881=>"000000000",
  7882=>"000110111",
  7883=>"111011000",
  7884=>"101100100",
  7885=>"111001110",
  7886=>"001100111",
  7887=>"001000000",
  7888=>"111100000",
  7889=>"111111111",
  7890=>"111111111",
  7891=>"000000000",
  7892=>"001011000",
  7893=>"010010000",
  7894=>"000111100",
  7895=>"111111111",
  7896=>"000001011",
  7897=>"111111111",
  7898=>"111111111",
  7899=>"111111111",
  7900=>"000000000",
  7901=>"001111111",
  7902=>"000000000",
  7903=>"001010111",
  7904=>"100111111",
  7905=>"000000101",
  7906=>"111111000",
  7907=>"000000000",
  7908=>"000000011",
  7909=>"001001000",
  7910=>"111011001",
  7911=>"000011011",
  7912=>"000000000",
  7913=>"001000101",
  7914=>"000100100",
  7915=>"000000000",
  7916=>"011000000",
  7917=>"111000000",
  7918=>"111111111",
  7919=>"000000000",
  7920=>"000000001",
  7921=>"001000111",
  7922=>"000100101",
  7923=>"000000011",
  7924=>"001111111",
  7925=>"111111111",
  7926=>"000000000",
  7927=>"111111111",
  7928=>"000000000",
  7929=>"111000011",
  7930=>"111100000",
  7931=>"110111110",
  7932=>"100111111",
  7933=>"000110110",
  7934=>"000101000",
  7935=>"001000000",
  7936=>"000000000",
  7937=>"000110110",
  7938=>"101111111",
  7939=>"001000000",
  7940=>"000000001",
  7941=>"111000000",
  7942=>"111111111",
  7943=>"001000000",
  7944=>"100100000",
  7945=>"011000011",
  7946=>"110000001",
  7947=>"000000100",
  7948=>"100100000",
  7949=>"001000000",
  7950=>"110111111",
  7951=>"111001000",
  7952=>"000110111",
  7953=>"111111111",
  7954=>"001001000",
  7955=>"111011111",
  7956=>"100000000",
  7957=>"111111000",
  7958=>"111111111",
  7959=>"111111111",
  7960=>"110110100",
  7961=>"111111110",
  7962=>"111111101",
  7963=>"100000000",
  7964=>"000101111",
  7965=>"000000000",
  7966=>"010011010",
  7967=>"111111111",
  7968=>"000000011",
  7969=>"111111111",
  7970=>"000000000",
  7971=>"011111111",
  7972=>"000111111",
  7973=>"111110000",
  7974=>"101100100",
  7975=>"000000000",
  7976=>"111111111",
  7977=>"000000000",
  7978=>"011111111",
  7979=>"000000000",
  7980=>"001001000",
  7981=>"111000110",
  7982=>"111111110",
  7983=>"111111111",
  7984=>"000000000",
  7985=>"111111111",
  7986=>"000000000",
  7987=>"000000011",
  7988=>"000000100",
  7989=>"111011111",
  7990=>"100111001",
  7991=>"111110101",
  7992=>"000000111",
  7993=>"111110110",
  7994=>"110110111",
  7995=>"110000000",
  7996=>"010000000",
  7997=>"111111111",
  7998=>"000001011",
  7999=>"000000110",
  8000=>"011111111",
  8001=>"000000000",
  8002=>"111001001",
  8003=>"001111111",
  8004=>"111111011",
  8005=>"111111111",
  8006=>"000000000",
  8007=>"000000000",
  8008=>"110110100",
  8009=>"000000000",
  8010=>"001101000",
  8011=>"011011001",
  8012=>"000000000",
  8013=>"010000000",
  8014=>"000000000",
  8015=>"100000000",
  8016=>"001001000",
  8017=>"001000010",
  8018=>"111111111",
  8019=>"100000000",
  8020=>"000000000",
  8021=>"011001001",
  8022=>"000000101",
  8023=>"000000000",
  8024=>"101111111",
  8025=>"111111111",
  8026=>"111011111",
  8027=>"111111111",
  8028=>"111111111",
  8029=>"111111111",
  8030=>"000000100",
  8031=>"111110000",
  8032=>"110111111",
  8033=>"100100110",
  8034=>"000100111",
  8035=>"110000000",
  8036=>"110110110",
  8037=>"011011011",
  8038=>"000000000",
  8039=>"111111000",
  8040=>"010110000",
  8041=>"111100100",
  8042=>"001001111",
  8043=>"111101101",
  8044=>"111110110",
  8045=>"000000000",
  8046=>"111111111",
  8047=>"000111111",
  8048=>"111111111",
  8049=>"000000000",
  8050=>"000001011",
  8051=>"111111111",
  8052=>"111011000",
  8053=>"111111111",
  8054=>"011111110",
  8055=>"001001001",
  8056=>"000000011",
  8057=>"110110010",
  8058=>"000000000",
  8059=>"100101001",
  8060=>"000000001",
  8061=>"001111111",
  8062=>"111111111",
  8063=>"111111111",
  8064=>"110110111",
  8065=>"110111111",
  8066=>"000000000",
  8067=>"000000000",
  8068=>"101000000",
  8069=>"000111000",
  8070=>"001001000",
  8071=>"000000000",
  8072=>"111000111",
  8073=>"000000000",
  8074=>"111000000",
  8075=>"000000000",
  8076=>"111111111",
  8077=>"100000001",
  8078=>"100110111",
  8079=>"000000001",
  8080=>"000000000",
  8081=>"111111111",
  8082=>"111100000",
  8083=>"000010000",
  8084=>"001001000",
  8085=>"001000000",
  8086=>"011011011",
  8087=>"111111111",
  8088=>"111111111",
  8089=>"110111000",
  8090=>"001000000",
  8091=>"000000011",
  8092=>"101001001",
  8093=>"000000011",
  8094=>"110110100",
  8095=>"000000100",
  8096=>"111111111",
  8097=>"001000000",
  8098=>"111111111",
  8099=>"000000000",
  8100=>"000000000",
  8101=>"000000000",
  8102=>"000000000",
  8103=>"111111001",
  8104=>"110111110",
  8105=>"011011111",
  8106=>"000000000",
  8107=>"110110110",
  8108=>"111000000",
  8109=>"111111011",
  8110=>"000010000",
  8111=>"000000000",
  8112=>"000010111",
  8113=>"100101110",
  8114=>"111111001",
  8115=>"111100011",
  8116=>"000100100",
  8117=>"111001001",
  8118=>"000000100",
  8119=>"000000111",
  8120=>"000100001",
  8121=>"000000101",
  8122=>"111111111",
  8123=>"000000000",
  8124=>"000000111",
  8125=>"000001111",
  8126=>"111010000",
  8127=>"100111100",
  8128=>"011011011",
  8129=>"000111111",
  8130=>"000000000",
  8131=>"100000000",
  8132=>"000000000",
  8133=>"110100110",
  8134=>"000000000",
  8135=>"000000100",
  8136=>"011010000",
  8137=>"000000000",
  8138=>"111111111",
  8139=>"101100111",
  8140=>"011011111",
  8141=>"111111111",
  8142=>"111101000",
  8143=>"000000000",
  8144=>"000000000",
  8145=>"000000000",
  8146=>"111111110",
  8147=>"100111000",
  8148=>"111111111",
  8149=>"011110000",
  8150=>"111101101",
  8151=>"000100101",
  8152=>"010010011",
  8153=>"000000000",
  8154=>"000000001",
  8155=>"000000011",
  8156=>"110000111",
  8157=>"111111001",
  8158=>"000000111",
  8159=>"010000000",
  8160=>"111001001",
  8161=>"000000111",
  8162=>"011001011",
  8163=>"000000001",
  8164=>"110111111",
  8165=>"111111111",
  8166=>"011000000",
  8167=>"000000000",
  8168=>"001000000",
  8169=>"111111000",
  8170=>"000000000",
  8171=>"000000000",
  8172=>"000101101",
  8173=>"110111111",
  8174=>"111111111",
  8175=>"001000000",
  8176=>"111111111",
  8177=>"111111111",
  8178=>"000000000",
  8179=>"100110110",
  8180=>"010000011",
  8181=>"011000000",
  8182=>"111111111",
  8183=>"110110111",
  8184=>"111111000",
  8185=>"001001111",
  8186=>"011011011",
  8187=>"000000000",
  8188=>"101101001",
  8189=>"010000000",
  8190=>"110100001",
  8191=>"010111111",
  8192=>"011111001",
  8193=>"111001000",
  8194=>"111111111",
  8195=>"000000000",
  8196=>"111111110",
  8197=>"000000000",
  8198=>"111111101",
  8199=>"101000000",
  8200=>"000000000",
  8201=>"111111000",
  8202=>"111111000",
  8203=>"000001111",
  8204=>"011001001",
  8205=>"111111111",
  8206=>"111111111",
  8207=>"011111111",
  8208=>"111111111",
  8209=>"000001001",
  8210=>"000000000",
  8211=>"001000000",
  8212=>"111111111",
  8213=>"000000000",
  8214=>"111111111",
  8215=>"110110000",
  8216=>"111100110",
  8217=>"000000000",
  8218=>"000000000",
  8219=>"000000001",
  8220=>"000000000",
  8221=>"111111111",
  8222=>"011011010",
  8223=>"000000000",
  8224=>"000000011",
  8225=>"000000000",
  8226=>"100110111",
  8227=>"111110010",
  8228=>"000011111",
  8229=>"100000000",
  8230=>"001100000",
  8231=>"111111000",
  8232=>"111111111",
  8233=>"100000000",
  8234=>"111111111",
  8235=>"100100111",
  8236=>"111111111",
  8237=>"000100000",
  8238=>"111111111",
  8239=>"000000000",
  8240=>"001001111",
  8241=>"010111010",
  8242=>"000100111",
  8243=>"000000110",
  8244=>"000001111",
  8245=>"010000000",
  8246=>"101100000",
  8247=>"100110111",
  8248=>"000001111",
  8249=>"110111011",
  8250=>"000000000",
  8251=>"010111111",
  8252=>"110000010",
  8253=>"111111111",
  8254=>"110110000",
  8255=>"111111111",
  8256=>"011001001",
  8257=>"000000000",
  8258=>"111111111",
  8259=>"111000111",
  8260=>"111001000",
  8261=>"111101001",
  8262=>"010000000",
  8263=>"000000000",
  8264=>"111011111",
  8265=>"011000000",
  8266=>"111111111",
  8267=>"001001111",
  8268=>"111100100",
  8269=>"000000000",
  8270=>"111101000",
  8271=>"010111111",
  8272=>"000000010",
  8273=>"111111100",
  8274=>"000000000",
  8275=>"001001001",
  8276=>"001001011",
  8277=>"111100000",
  8278=>"000000000",
  8279=>"111100110",
  8280=>"010000111",
  8281=>"111111111",
  8282=>"000000000",
  8283=>"110110011",
  8284=>"111111111",
  8285=>"000000000",
  8286=>"111000011",
  8287=>"000000011",
  8288=>"111001000",
  8289=>"000000000",
  8290=>"111001001",
  8291=>"111100000",
  8292=>"101100111",
  8293=>"000000000",
  8294=>"111111111",
  8295=>"110100001",
  8296=>"111111111",
  8297=>"000001110",
  8298=>"111111000",
  8299=>"000000000",
  8300=>"011011001",
  8301=>"000111111",
  8302=>"011011111",
  8303=>"100101111",
  8304=>"000000000",
  8305=>"001000000",
  8306=>"111111111",
  8307=>"111011111",
  8308=>"000000000",
  8309=>"000000000",
  8310=>"000000000",
  8311=>"000000000",
  8312=>"011011111",
  8313=>"111111111",
  8314=>"001000000",
  8315=>"011000000",
  8316=>"010000001",
  8317=>"111111101",
  8318=>"111111111",
  8319=>"000001100",
  8320=>"111111100",
  8321=>"111011000",
  8322=>"000111111",
  8323=>"011000111",
  8324=>"000000001",
  8325=>"111000000",
  8326=>"110000000",
  8327=>"111111111",
  8328=>"111111111",
  8329=>"110111111",
  8330=>"111111111",
  8331=>"111111111",
  8332=>"010111111",
  8333=>"011010000",
  8334=>"111001111",
  8335=>"000000000",
  8336=>"000000000",
  8337=>"001001111",
  8338=>"000000000",
  8339=>"000000000",
  8340=>"111111000",
  8341=>"000000000",
  8342=>"000000000",
  8343=>"111111111",
  8344=>"000000000",
  8345=>"000000000",
  8346=>"000010010",
  8347=>"111111110",
  8348=>"111111111",
  8349=>"011001001",
  8350=>"000000000",
  8351=>"111111111",
  8352=>"101001000",
  8353=>"001000001",
  8354=>"000000000",
  8355=>"000000000",
  8356=>"011111110",
  8357=>"000000000",
  8358=>"111000000",
  8359=>"000110010",
  8360=>"000000000",
  8361=>"000001001",
  8362=>"111111111",
  8363=>"000000000",
  8364=>"111111000",
  8365=>"111100000",
  8366=>"000000000",
  8367=>"001011101",
  8368=>"000001111",
  8369=>"100100000",
  8370=>"111111110",
  8371=>"111000001",
  8372=>"111111111",
  8373=>"000000100",
  8374=>"000000000",
  8375=>"111111111",
  8376=>"111111111",
  8377=>"000000000",
  8378=>"000000110",
  8379=>"000101111",
  8380=>"000000000",
  8381=>"000010010",
  8382=>"111111111",
  8383=>"000000000",
  8384=>"111110111",
  8385=>"000111111",
  8386=>"111111101",
  8387=>"100000000",
  8388=>"111111111",
  8389=>"111111111",
  8390=>"111000100",
  8391=>"001000111",
  8392=>"100110110",
  8393=>"111101111",
  8394=>"011000001",
  8395=>"000001000",
  8396=>"001000000",
  8397=>"000000000",
  8398=>"000000000",
  8399=>"011011010",
  8400=>"000000001",
  8401=>"000000000",
  8402=>"011111111",
  8403=>"111100001",
  8404=>"001111110",
  8405=>"111111111",
  8406=>"100100100",
  8407=>"000000111",
  8408=>"110000111",
  8409=>"111111111",
  8410=>"000000101",
  8411=>"111111101",
  8412=>"000000000",
  8413=>"011101111",
  8414=>"000000000",
  8415=>"000000000",
  8416=>"111000000",
  8417=>"000000000",
  8418=>"110000000",
  8419=>"000000000",
  8420=>"000000011",
  8421=>"101111110",
  8422=>"110111111",
  8423=>"111111000",
  8424=>"001000001",
  8425=>"001001111",
  8426=>"000000000",
  8427=>"001100110",
  8428=>"000000000",
  8429=>"000000111",
  8430=>"000111111",
  8431=>"000000000",
  8432=>"101100000",
  8433=>"000000000",
  8434=>"000000000",
  8435=>"000100110",
  8436=>"111111111",
  8437=>"111110111",
  8438=>"000000000",
  8439=>"000000101",
  8440=>"111111111",
  8441=>"111000000",
  8442=>"000000000",
  8443=>"000000011",
  8444=>"001001000",
  8445=>"110110111",
  8446=>"111010000",
  8447=>"000000000",
  8448=>"111111111",
  8449=>"010011110",
  8450=>"000000001",
  8451=>"111111000",
  8452=>"111111111",
  8453=>"101100100",
  8454=>"000000100",
  8455=>"001000000",
  8456=>"111000000",
  8457=>"000000000",
  8458=>"111111111",
  8459=>"111000011",
  8460=>"100000000",
  8461=>"001011111",
  8462=>"000000000",
  8463=>"010000000",
  8464=>"000000000",
  8465=>"000000000",
  8466=>"111111111",
  8467=>"000000101",
  8468=>"000000111",
  8469=>"111111000",
  8470=>"111111111",
  8471=>"111111111",
  8472=>"001001101",
  8473=>"000000000",
  8474=>"101111111",
  8475=>"100000000",
  8476=>"001001011",
  8477=>"111011001",
  8478=>"111111101",
  8479=>"011011000",
  8480=>"000000000",
  8481=>"111011001",
  8482=>"111011111",
  8483=>"011011001",
  8484=>"111111111",
  8485=>"000000100",
  8486=>"111111111",
  8487=>"001001001",
  8488=>"000000111",
  8489=>"000000000",
  8490=>"001000000",
  8491=>"111111111",
  8492=>"001001000",
  8493=>"100100100",
  8494=>"000000000",
  8495=>"000000000",
  8496=>"000000000",
  8497=>"111000000",
  8498=>"111111111",
  8499=>"111111111",
  8500=>"000000000",
  8501=>"000000001",
  8502=>"000000001",
  8503=>"111100000",
  8504=>"000000000",
  8505=>"111000001",
  8506=>"111111000",
  8507=>"010010000",
  8508=>"111110100",
  8509=>"101101000",
  8510=>"111111011",
  8511=>"111111111",
  8512=>"111111111",
  8513=>"000000000",
  8514=>"000000001",
  8515=>"111111111",
  8516=>"001000111",
  8517=>"110110110",
  8518=>"011111111",
  8519=>"000000000",
  8520=>"000000000",
  8521=>"011111111",
  8522=>"011001111",
  8523=>"000000000",
  8524=>"111111111",
  8525=>"010011001",
  8526=>"101101001",
  8527=>"000000001",
  8528=>"001001001",
  8529=>"111110111",
  8530=>"000000000",
  8531=>"110111100",
  8532=>"000000100",
  8533=>"011000000",
  8534=>"000000000",
  8535=>"000000000",
  8536=>"111111111",
  8537=>"101001010",
  8538=>"110110010",
  8539=>"100100100",
  8540=>"101000000",
  8541=>"111000000",
  8542=>"001011111",
  8543=>"110110010",
  8544=>"111111111",
  8545=>"111111111",
  8546=>"000000000",
  8547=>"111011000",
  8548=>"111111000",
  8549=>"000000000",
  8550=>"000000000",
  8551=>"111111111",
  8552=>"000001011",
  8553=>"000000000",
  8554=>"010100100",
  8555=>"000011100",
  8556=>"001001011",
  8557=>"011011110",
  8558=>"111100000",
  8559=>"000111011",
  8560=>"000000000",
  8561=>"000111111",
  8562=>"001001011",
  8563=>"110110111",
  8564=>"111111111",
  8565=>"000000100",
  8566=>"011111111",
  8567=>"100100000",
  8568=>"111111111",
  8569=>"111111100",
  8570=>"000000000",
  8571=>"111100000",
  8572=>"000000001",
  8573=>"001000000",
  8574=>"111000000",
  8575=>"111111111",
  8576=>"011011111",
  8577=>"001001011",
  8578=>"000000000",
  8579=>"001001001",
  8580=>"110110100",
  8581=>"000000001",
  8582=>"110110111",
  8583=>"011000000",
  8584=>"100100000",
  8585=>"111111011",
  8586=>"111111111",
  8587=>"011111111",
  8588=>"111000000",
  8589=>"111111110",
  8590=>"000000000",
  8591=>"100000000",
  8592=>"111111111",
  8593=>"000000001",
  8594=>"000000000",
  8595=>"111111111",
  8596=>"110111111",
  8597=>"000011011",
  8598=>"010000001",
  8599=>"111111111",
  8600=>"000000000",
  8601=>"000000000",
  8602=>"001000001",
  8603=>"111111111",
  8604=>"000000000",
  8605=>"111111111",
  8606=>"001000110",
  8607=>"000000000",
  8608=>"000000000",
  8609=>"001000000",
  8610=>"000000100",
  8611=>"111111001",
  8612=>"111000111",
  8613=>"010100111",
  8614=>"000110111",
  8615=>"011111111",
  8616=>"111111011",
  8617=>"111111111",
  8618=>"000000000",
  8619=>"000000000",
  8620=>"000000000",
  8621=>"000000000",
  8622=>"111010000",
  8623=>"000000011",
  8624=>"010000000",
  8625=>"000000000",
  8626=>"000000000",
  8627=>"000111111",
  8628=>"001001111",
  8629=>"111111111",
  8630=>"111111111",
  8631=>"000000000",
  8632=>"000111111",
  8633=>"011111111",
  8634=>"001001000",
  8635=>"000100000",
  8636=>"000000000",
  8637=>"011001000",
  8638=>"000000000",
  8639=>"111111110",
  8640=>"100000000",
  8641=>"000000000",
  8642=>"000011001",
  8643=>"111111111",
  8644=>"000000000",
  8645=>"100100100",
  8646=>"111111111",
  8647=>"000000000",
  8648=>"000000000",
  8649=>"000000100",
  8650=>"001000000",
  8651=>"111111111",
  8652=>"000111000",
  8653=>"111111101",
  8654=>"011001111",
  8655=>"000111111",
  8656=>"000101111",
  8657=>"000100001",
  8658=>"111111111",
  8659=>"010110010",
  8660=>"100100111",
  8661=>"011000000",
  8662=>"111111000",
  8663=>"000000000",
  8664=>"111111111",
  8665=>"100111111",
  8666=>"111000000",
  8667=>"000000000",
  8668=>"111111110",
  8669=>"111001101",
  8670=>"000000000",
  8671=>"111111011",
  8672=>"110101000",
  8673=>"110000000",
  8674=>"000000000",
  8675=>"111111111",
  8676=>"000000000",
  8677=>"111101100",
  8678=>"111111000",
  8679=>"111111111",
  8680=>"111111111",
  8681=>"000000000",
  8682=>"000000000",
  8683=>"000000110",
  8684=>"011111111",
  8685=>"000100111",
  8686=>"000000000",
  8687=>"111010110",
  8688=>"001000000",
  8689=>"111111011",
  8690=>"101100111",
  8691=>"111110000",
  8692=>"010111001",
  8693=>"000000000",
  8694=>"001001000",
  8695=>"001011011",
  8696=>"111111011",
  8697=>"000001000",
  8698=>"111111001",
  8699=>"111111111",
  8700=>"111111111",
  8701=>"110110000",
  8702=>"001001000",
  8703=>"111100000",
  8704=>"111000001",
  8705=>"111111000",
  8706=>"001101111",
  8707=>"000000000",
  8708=>"000000000",
  8709=>"000111111",
  8710=>"000000100",
  8711=>"110111111",
  8712=>"000000000",
  8713=>"111111111",
  8714=>"101000000",
  8715=>"110000000",
  8716=>"110000000",
  8717=>"100100000",
  8718=>"000000001",
  8719=>"111111111",
  8720=>"111111111",
  8721=>"000101111",
  8722=>"000000111",
  8723=>"000100111",
  8724=>"000100111",
  8725=>"101111111",
  8726=>"000000110",
  8727=>"111111111",
  8728=>"111111001",
  8729=>"111010000",
  8730=>"111111110",
  8731=>"111001001",
  8732=>"000101000",
  8733=>"011000000",
  8734=>"001001001",
  8735=>"000000000",
  8736=>"010000110",
  8737=>"000000110",
  8738=>"000000100",
  8739=>"111111111",
  8740=>"000000000",
  8741=>"100001111",
  8742=>"000000000",
  8743=>"000000000",
  8744=>"000000000",
  8745=>"101111111",
  8746=>"110010011",
  8747=>"111001000",
  8748=>"000111000",
  8749=>"101111001",
  8750=>"000000000",
  8751=>"111111010",
  8752=>"000000000",
  8753=>"111101000",
  8754=>"111110100",
  8755=>"011111111",
  8756=>"010010000",
  8757=>"000000010",
  8758=>"001011001",
  8759=>"001000000",
  8760=>"111111111",
  8761=>"000100111",
  8762=>"000000000",
  8763=>"000000000",
  8764=>"000000000",
  8765=>"000100000",
  8766=>"000000110",
  8767=>"000000000",
  8768=>"000000001",
  8769=>"000001000",
  8770=>"100000001",
  8771=>"111111111",
  8772=>"101111111",
  8773=>"111111111",
  8774=>"100100001",
  8775=>"111111111",
  8776=>"110100100",
  8777=>"111001111",
  8778=>"011011111",
  8779=>"000000111",
  8780=>"100111111",
  8781=>"000000100",
  8782=>"000000001",
  8783=>"000000000",
  8784=>"011000000",
  8785=>"100101011",
  8786=>"100000000",
  8787=>"000000011",
  8788=>"111111000",
  8789=>"111100000",
  8790=>"111110000",
  8791=>"000000000",
  8792=>"111111111",
  8793=>"100000000",
  8794=>"001000000",
  8795=>"101000000",
  8796=>"111111111",
  8797=>"101101111",
  8798=>"101111111",
  8799=>"111000000",
  8800=>"000000001",
  8801=>"100110000",
  8802=>"100000000",
  8803=>"000000000",
  8804=>"000001101",
  8805=>"000010010",
  8806=>"101111111",
  8807=>"011010000",
  8808=>"000111111",
  8809=>"110111111",
  8810=>"111111111",
  8811=>"111101011",
  8812=>"000000001",
  8813=>"111111111",
  8814=>"100111111",
  8815=>"000000100",
  8816=>"111110111",
  8817=>"000000001",
  8818=>"111111111",
  8819=>"111111111",
  8820=>"111111110",
  8821=>"001111111",
  8822=>"111111111",
  8823=>"111001000",
  8824=>"011000000",
  8825=>"000000000",
  8826=>"111110100",
  8827=>"000000001",
  8828=>"100100000",
  8829=>"000000000",
  8830=>"000000000",
  8831=>"000011111",
  8832=>"111111111",
  8833=>"000000111",
  8834=>"010000000",
  8835=>"000000100",
  8836=>"000001000",
  8837=>"000000000",
  8838=>"000000010",
  8839=>"101111111",
  8840=>"000000000",
  8841=>"000000001",
  8842=>"100111111",
  8843=>"111111001",
  8844=>"011011000",
  8845=>"000000000",
  8846=>"110000001",
  8847=>"000000000",
  8848=>"101111111",
  8849=>"000000000",
  8850=>"111111111",
  8851=>"100000000",
  8852=>"010000011",
  8853=>"001111101",
  8854=>"000011111",
  8855=>"111000000",
  8856=>"000000111",
  8857=>"111111011",
  8858=>"100000000",
  8859=>"000001100",
  8860=>"111111111",
  8861=>"110000000",
  8862=>"000000111",
  8863=>"111000000",
  8864=>"000000111",
  8865=>"101000000",
  8866=>"100100111",
  8867=>"111111000",
  8868=>"111001000",
  8869=>"111000100",
  8870=>"001111111",
  8871=>"101100000",
  8872=>"000011000",
  8873=>"000000001",
  8874=>"000000000",
  8875=>"000000111",
  8876=>"101000000",
  8877=>"111011111",
  8878=>"100010111",
  8879=>"001001011",
  8880=>"000000000",
  8881=>"101100110",
  8882=>"100100000",
  8883=>"000000100",
  8884=>"111011000",
  8885=>"111001111",
  8886=>"000000000",
  8887=>"111111111",
  8888=>"111111011",
  8889=>"011111000",
  8890=>"111111110",
  8891=>"111111110",
  8892=>"111111000",
  8893=>"011011111",
  8894=>"111111001",
  8895=>"111111000",
  8896=>"111000000",
  8897=>"000000000",
  8898=>"110000001",
  8899=>"110000000",
  8900=>"011111111",
  8901=>"000000000",
  8902=>"111100000",
  8903=>"000001000",
  8904=>"000110111",
  8905=>"111111111",
  8906=>"000000000",
  8907=>"111111111",
  8908=>"100000000",
  8909=>"111111110",
  8910=>"111111000",
  8911=>"111000010",
  8912=>"110111000",
  8913=>"111111111",
  8914=>"101001111",
  8915=>"000111111",
  8916=>"001000001",
  8917=>"100111111",
  8918=>"000001001",
  8919=>"011111111",
  8920=>"011000111",
  8921=>"111111011",
  8922=>"000100110",
  8923=>"111111111",
  8924=>"000000000",
  8925=>"000000101",
  8926=>"111111111",
  8927=>"101100100",
  8928=>"111000000",
  8929=>"000000000",
  8930=>"010111100",
  8931=>"100110111",
  8932=>"000000000",
  8933=>"111111110",
  8934=>"111111110",
  8935=>"111011011",
  8936=>"110000000",
  8937=>"010000000",
  8938=>"111111111",
  8939=>"000100111",
  8940=>"111111111",
  8941=>"111000000",
  8942=>"111000111",
  8943=>"000000111",
  8944=>"110111111",
  8945=>"111111111",
  8946=>"000111111",
  8947=>"001000000",
  8948=>"111000000",
  8949=>"100111111",
  8950=>"100111101",
  8951=>"110000000",
  8952=>"111100100",
  8953=>"000000000",
  8954=>"000000001",
  8955=>"001101000",
  8956=>"111111010",
  8957=>"001001000",
  8958=>"111111100",
  8959=>"011111011",
  8960=>"100000000",
  8961=>"101111111",
  8962=>"111111000",
  8963=>"111111111",
  8964=>"111111111",
  8965=>"011011001",
  8966=>"010110111",
  8967=>"000000000",
  8968=>"111111111",
  8969=>"000000000",
  8970=>"000000101",
  8971=>"000111111",
  8972=>"000000000",
  8973=>"100000000",
  8974=>"000101111",
  8975=>"111001111",
  8976=>"101111101",
  8977=>"111111111",
  8978=>"111101000",
  8979=>"101001000",
  8980=>"111111111",
  8981=>"111000011",
  8982=>"000110101",
  8983=>"000000000",
  8984=>"000000000",
  8985=>"111111011",
  8986=>"000010110",
  8987=>"111111111",
  8988=>"111001000",
  8989=>"000110111",
  8990=>"000000000",
  8991=>"110111111",
  8992=>"000000100",
  8993=>"011011001",
  8994=>"100100110",
  8995=>"000000000",
  8996=>"000000110",
  8997=>"000000000",
  8998=>"011011111",
  8999=>"111000000",
  9000=>"001000000",
  9001=>"000001000",
  9002=>"000111111",
  9003=>"000000000",
  9004=>"111111000",
  9005=>"111111000",
  9006=>"100000000",
  9007=>"111000000",
  9008=>"110011111",
  9009=>"000000000",
  9010=>"000000000",
  9011=>"011000000",
  9012=>"000000000",
  9013=>"011000000",
  9014=>"010111101",
  9015=>"111100000",
  9016=>"000000111",
  9017=>"000000100",
  9018=>"100000000",
  9019=>"111111111",
  9020=>"000000000",
  9021=>"000000111",
  9022=>"110110111",
  9023=>"000000101",
  9024=>"011011011",
  9025=>"111111001",
  9026=>"100000000",
  9027=>"000000000",
  9028=>"000000101",
  9029=>"000000111",
  9030=>"111011111",
  9031=>"111111110",
  9032=>"111111000",
  9033=>"000011111",
  9034=>"000000000",
  9035=>"010110100",
  9036=>"000000001",
  9037=>"011111000",
  9038=>"111111111",
  9039=>"100100001",
  9040=>"000000010",
  9041=>"111101000",
  9042=>"111000111",
  9043=>"111111111",
  9044=>"110110111",
  9045=>"011001011",
  9046=>"110110111",
  9047=>"011111111",
  9048=>"010100111",
  9049=>"000000000",
  9050=>"100000000",
  9051=>"000000000",
  9052=>"111111011",
  9053=>"000000111",
  9054=>"111111001",
  9055=>"111001001",
  9056=>"111111111",
  9057=>"000000000",
  9058=>"000110100",
  9059=>"110110000",
  9060=>"000000000",
  9061=>"111000000",
  9062=>"000000000",
  9063=>"000000000",
  9064=>"000000001",
  9065=>"100010110",
  9066=>"000000111",
  9067=>"101111000",
  9068=>"110110110",
  9069=>"111111101",
  9070=>"111110100",
  9071=>"100110111",
  9072=>"111111111",
  9073=>"111111111",
  9074=>"100000110",
  9075=>"000111111",
  9076=>"111100000",
  9077=>"100010011",
  9078=>"000110111",
  9079=>"111111111",
  9080=>"100000000",
  9081=>"000110111",
  9082=>"000000110",
  9083=>"100100000",
  9084=>"000100100",
  9085=>"111111110",
  9086=>"000000000",
  9087=>"000000111",
  9088=>"000000000",
  9089=>"111100000",
  9090=>"111110111",
  9091=>"011011000",
  9092=>"000000000",
  9093=>"001111111",
  9094=>"110111111",
  9095=>"000000000",
  9096=>"000111111",
  9097=>"111111000",
  9098=>"001011101",
  9099=>"011011111",
  9100=>"110000111",
  9101=>"001101101",
  9102=>"100000011",
  9103=>"010000000",
  9104=>"001001101",
  9105=>"011000000",
  9106=>"000000000",
  9107=>"000000000",
  9108=>"001001111",
  9109=>"000000001",
  9110=>"111110000",
  9111=>"100000000",
  9112=>"111111111",
  9113=>"111111111",
  9114=>"000000111",
  9115=>"000000000",
  9116=>"111110100",
  9117=>"100111111",
  9118=>"110000111",
  9119=>"000110000",
  9120=>"000000000",
  9121=>"101111100",
  9122=>"000000000",
  9123=>"000111111",
  9124=>"100000000",
  9125=>"111001000",
  9126=>"111001001",
  9127=>"111001000",
  9128=>"000111111",
  9129=>"000011011",
  9130=>"100000000",
  9131=>"000010101",
  9132=>"000000000",
  9133=>"100000000",
  9134=>"110000000",
  9135=>"111000000",
  9136=>"000000011",
  9137=>"011000000",
  9138=>"000000001",
  9139=>"000000011",
  9140=>"110111111",
  9141=>"000111111",
  9142=>"001000111",
  9143=>"111101000",
  9144=>"000100111",
  9145=>"111111101",
  9146=>"110110111",
  9147=>"000000111",
  9148=>"111111111",
  9149=>"000000100",
  9150=>"111111101",
  9151=>"101101101",
  9152=>"000000101",
  9153=>"111011001",
  9154=>"111111111",
  9155=>"000000000",
  9156=>"111111111",
  9157=>"001001111",
  9158=>"001001101",
  9159=>"011111011",
  9160=>"000000001",
  9161=>"111100000",
  9162=>"000000000",
  9163=>"100000000",
  9164=>"001001000",
  9165=>"110110000",
  9166=>"001001001",
  9167=>"101100110",
  9168=>"000001011",
  9169=>"111111111",
  9170=>"111111111",
  9171=>"111111110",
  9172=>"101111111",
  9173=>"011000000",
  9174=>"111111100",
  9175=>"100100011",
  9176=>"000000000",
  9177=>"100000000",
  9178=>"000000110",
  9179=>"100100001",
  9180=>"100100101",
  9181=>"011001000",
  9182=>"000111100",
  9183=>"111101100",
  9184=>"111111011",
  9185=>"000000000",
  9186=>"000000000",
  9187=>"011001011",
  9188=>"000000000",
  9189=>"000010000",
  9190=>"011111111",
  9191=>"000000111",
  9192=>"000000001",
  9193=>"000010000",
  9194=>"000000000",
  9195=>"111111111",
  9196=>"111000000",
  9197=>"011000100",
  9198=>"000000000",
  9199=>"100000111",
  9200=>"000000100",
  9201=>"011001011",
  9202=>"111100000",
  9203=>"111111111",
  9204=>"100000111",
  9205=>"000000000",
  9206=>"111101000",
  9207=>"101100110",
  9208=>"011001000",
  9209=>"100110100",
  9210=>"100100000",
  9211=>"111111001",
  9212=>"000000111",
  9213=>"100110111",
  9214=>"100001001",
  9215=>"110100101",
  9216=>"000000000",
  9217=>"110110111",
  9218=>"111111101",
  9219=>"001111111",
  9220=>"111111111",
  9221=>"000000001",
  9222=>"001101111",
  9223=>"101000100",
  9224=>"111111000",
  9225=>"000000111",
  9226=>"101001111",
  9227=>"000000111",
  9228=>"100100000",
  9229=>"000000000",
  9230=>"111000100",
  9231=>"111111110",
  9232=>"000011000",
  9233=>"000010111",
  9234=>"000000000",
  9235=>"111111111",
  9236=>"001000000",
  9237=>"001101111",
  9238=>"011011000",
  9239=>"100110000",
  9240=>"000000000",
  9241=>"100110010",
  9242=>"111000100",
  9243=>"000000000",
  9244=>"110110000",
  9245=>"101000000",
  9246=>"000000000",
  9247=>"110111000",
  9248=>"100111111",
  9249=>"001011000",
  9250=>"101111000",
  9251=>"111111111",
  9252=>"000000111",
  9253=>"111111111",
  9254=>"000100110",
  9255=>"110000000",
  9256=>"000000001",
  9257=>"111111000",
  9258=>"000000000",
  9259=>"111110000",
  9260=>"111011011",
  9261=>"111101110",
  9262=>"101000001",
  9263=>"101001111",
  9264=>"000101101",
  9265=>"000000000",
  9266=>"000000100",
  9267=>"111111111",
  9268=>"000000000",
  9269=>"101111111",
  9270=>"111000001",
  9271=>"001000000",
  9272=>"001001100",
  9273=>"011111000",
  9274=>"001000000",
  9275=>"000000110",
  9276=>"101101111",
  9277=>"111110111",
  9278=>"100101111",
  9279=>"111111111",
  9280=>"111111110",
  9281=>"111011000",
  9282=>"000000000",
  9283=>"000000111",
  9284=>"111111111",
  9285=>"000000100",
  9286=>"000000111",
  9287=>"000110000",
  9288=>"111110000",
  9289=>"111101111",
  9290=>"000000000",
  9291=>"000000001",
  9292=>"001001010",
  9293=>"000000100",
  9294=>"100111110",
  9295=>"001000000",
  9296=>"010000000",
  9297=>"000000000",
  9298=>"111111111",
  9299=>"100111111",
  9300=>"100000111",
  9301=>"111110000",
  9302=>"111000100",
  9303=>"111100000",
  9304=>"000000000",
  9305=>"001000111",
  9306=>"011000001",
  9307=>"110111111",
  9308=>"100000000",
  9309=>"101111111",
  9310=>"111111100",
  9311=>"100111000",
  9312=>"100100000",
  9313=>"111111111",
  9314=>"000000000",
  9315=>"111111111",
  9316=>"000000000",
  9317=>"110111111",
  9318=>"101111111",
  9319=>"000000000",
  9320=>"000000000",
  9321=>"111111000",
  9322=>"000111111",
  9323=>"000000100",
  9324=>"001001111",
  9325=>"111101001",
  9326=>"000000010",
  9327=>"000000000",
  9328=>"110111111",
  9329=>"111001001",
  9330=>"100000000",
  9331=>"111101000",
  9332=>"000000000",
  9333=>"011000000",
  9334=>"000001111",
  9335=>"000101111",
  9336=>"111111011",
  9337=>"011001001",
  9338=>"001000000",
  9339=>"000000001",
  9340=>"000100000",
  9341=>"000000111",
  9342=>"000000000",
  9343=>"000110110",
  9344=>"111110000",
  9345=>"111111111",
  9346=>"000000000",
  9347=>"110111111",
  9348=>"000000000",
  9349=>"000000111",
  9350=>"111111110",
  9351=>"000111110",
  9352=>"111111111",
  9353=>"101000000",
  9354=>"111100111",
  9355=>"100000100",
  9356=>"111111101",
  9357=>"000000000",
  9358=>"010110110",
  9359=>"001000000",
  9360=>"111000001",
  9361=>"100000000",
  9362=>"000000000",
  9363=>"011011000",
  9364=>"111001000",
  9365=>"000000111",
  9366=>"001010000",
  9367=>"000000000",
  9368=>"111000111",
  9369=>"111111111",
  9370=>"111111111",
  9371=>"111111111",
  9372=>"111111000",
  9373=>"000000000",
  9374=>"001001001",
  9375=>"000000010",
  9376=>"001001000",
  9377=>"001000000",
  9378=>"111100110",
  9379=>"001101001",
  9380=>"100000000",
  9381=>"110010010",
  9382=>"101000110",
  9383=>"111111111",
  9384=>"000000100",
  9385=>"100000000",
  9386=>"111111111",
  9387=>"111111111",
  9388=>"000000000",
  9389=>"110110110",
  9390=>"000000000",
  9391=>"111100000",
  9392=>"000000000",
  9393=>"011010000",
  9394=>"110111111",
  9395=>"000000100",
  9396=>"000010011",
  9397=>"000000010",
  9398=>"111100110",
  9399=>"000000000",
  9400=>"000000110",
  9401=>"111101111",
  9402=>"010000000",
  9403=>"111101011",
  9404=>"000111110",
  9405=>"111111111",
  9406=>"111111111",
  9407=>"000000110",
  9408=>"111111111",
  9409=>"000000101",
  9410=>"111110100",
  9411=>"111111111",
  9412=>"111111111",
  9413=>"000000000",
  9414=>"000000001",
  9415=>"110000000",
  9416=>"000001011",
  9417=>"111111111",
  9418=>"000000010",
  9419=>"001000000",
  9420=>"110110110",
  9421=>"000000000",
  9422=>"000000100",
  9423=>"011010000",
  9424=>"000000000",
  9425=>"000100111",
  9426=>"010110000",
  9427=>"000000000",
  9428=>"100010010",
  9429=>"001001001",
  9430=>"111111111",
  9431=>"101101101",
  9432=>"000001000",
  9433=>"111001000",
  9434=>"110000000",
  9435=>"100110111",
  9436=>"001111100",
  9437=>"000110111",
  9438=>"111001000",
  9439=>"000001110",
  9440=>"101111111",
  9441=>"111000000",
  9442=>"111111000",
  9443=>"111010100",
  9444=>"111111111",
  9445=>"111111111",
  9446=>"100000101",
  9447=>"101111111",
  9448=>"111111111",
  9449=>"111111111",
  9450=>"001101101",
  9451=>"111111000",
  9452=>"111111000",
  9453=>"000000000",
  9454=>"000011110",
  9455=>"111000000",
  9456=>"111111111",
  9457=>"111111111",
  9458=>"110110110",
  9459=>"000100000",
  9460=>"001110111",
  9461=>"010111010",
  9462=>"000000000",
  9463=>"111001111",
  9464=>"100111111",
  9465=>"011111110",
  9466=>"111111110",
  9467=>"111111111",
  9468=>"011011001",
  9469=>"001000000",
  9470=>"111000100",
  9471=>"001001000",
  9472=>"100111100",
  9473=>"100100100",
  9474=>"000000001",
  9475=>"000000000",
  9476=>"100000000",
  9477=>"111111111",
  9478=>"000000000",
  9479=>"111111111",
  9480=>"011110001",
  9481=>"000000000",
  9482=>"000000001",
  9483=>"100100100",
  9484=>"100000100",
  9485=>"001010111",
  9486=>"110111111",
  9487=>"111110000",
  9488=>"000001011",
  9489=>"001111011",
  9490=>"000000010",
  9491=>"000000000",
  9492=>"000111000",
  9493=>"000111111",
  9494=>"011111111",
  9495=>"111111000",
  9496=>"100100000",
  9497=>"111111010",
  9498=>"100100000",
  9499=>"110000001",
  9500=>"100001000",
  9501=>"111111111",
  9502=>"101111001",
  9503=>"111000000",
  9504=>"000000000",
  9505=>"000000011",
  9506=>"101001101",
  9507=>"101001111",
  9508=>"111010001",
  9509=>"100100100",
  9510=>"110110110",
  9511=>"000000000",
  9512=>"111001001",
  9513=>"000000000",
  9514=>"101110000",
  9515=>"000000000",
  9516=>"111111110",
  9517=>"000000000",
  9518=>"000111111",
  9519=>"110000100",
  9520=>"000000000",
  9521=>"000001011",
  9522=>"111111111",
  9523=>"111111011",
  9524=>"110111001",
  9525=>"000011000",
  9526=>"000000000",
  9527=>"111100100",
  9528=>"000000010",
  9529=>"000000011",
  9530=>"011100000",
  9531=>"000010110",
  9532=>"100100111",
  9533=>"000000100",
  9534=>"000000000",
  9535=>"111100100",
  9536=>"000000000",
  9537=>"111000011",
  9538=>"000000000",
  9539=>"111000111",
  9540=>"111111110",
  9541=>"111001111",
  9542=>"111101011",
  9543=>"000000000",
  9544=>"100101000",
  9545=>"100111000",
  9546=>"111111111",
  9547=>"101000000",
  9548=>"000001001",
  9549=>"000000000",
  9550=>"101100100",
  9551=>"000000000",
  9552=>"000000100",
  9553=>"000001111",
  9554=>"000000010",
  9555=>"010110010",
  9556=>"000000111",
  9557=>"011011011",
  9558=>"000000000",
  9559=>"111111111",
  9560=>"111110111",
  9561=>"110111111",
  9562=>"000000011",
  9563=>"110110100",
  9564=>"000000000",
  9565=>"001000000",
  9566=>"000000111",
  9567=>"101111111",
  9568=>"111111111",
  9569=>"111010000",
  9570=>"001001101",
  9571=>"111111111",
  9572=>"001111000",
  9573=>"111111111",
  9574=>"000000000",
  9575=>"000000000",
  9576=>"001001001",
  9577=>"001111111",
  9578=>"111110111",
  9579=>"111111111",
  9580=>"110111011",
  9581=>"000000110",
  9582=>"000000000",
  9583=>"111111111",
  9584=>"000110100",
  9585=>"111111111",
  9586=>"100111111",
  9587=>"011110111",
  9588=>"111111100",
  9589=>"100000000",
  9590=>"000001100",
  9591=>"101101001",
  9592=>"000000000",
  9593=>"000000000",
  9594=>"111111111",
  9595=>"111111101",
  9596=>"010000000",
  9597=>"000001011",
  9598=>"001001001",
  9599=>"111000000",
  9600=>"111111111",
  9601=>"000000001",
  9602=>"001001001",
  9603=>"111001000",
  9604=>"111111111",
  9605=>"000000000",
  9606=>"000000000",
  9607=>"110111111",
  9608=>"000000000",
  9609=>"011010011",
  9610=>"111111111",
  9611=>"111111010",
  9612=>"101111111",
  9613=>"011111100",
  9614=>"111111111",
  9615=>"111111111",
  9616=>"111111111",
  9617=>"111111111",
  9618=>"000000000",
  9619=>"011001100",
  9620=>"000110000",
  9621=>"011000000",
  9622=>"000000000",
  9623=>"000000000",
  9624=>"000001011",
  9625=>"111110111",
  9626=>"111111111",
  9627=>"111111111",
  9628=>"011011111",
  9629=>"000000001",
  9630=>"000001011",
  9631=>"111111111",
  9632=>"000000000",
  9633=>"000000100",
  9634=>"100100001",
  9635=>"111111111",
  9636=>"111111111",
  9637=>"111111111",
  9638=>"100101111",
  9639=>"000000011",
  9640=>"000000000",
  9641=>"111100100",
  9642=>"000000100",
  9643=>"000000000",
  9644=>"110010000",
  9645=>"111010000",
  9646=>"110110100",
  9647=>"111111000",
  9648=>"111101111",
  9649=>"000000110",
  9650=>"111111111",
  9651=>"000000011",
  9652=>"000000110",
  9653=>"101001000",
  9654=>"111101111",
  9655=>"111111111",
  9656=>"000000100",
  9657=>"000000010",
  9658=>"000000010",
  9659=>"000100111",
  9660=>"000000000",
  9661=>"110111101",
  9662=>"001000100",
  9663=>"111111101",
  9664=>"101001111",
  9665=>"010000111",
  9666=>"000000000",
  9667=>"111111111",
  9668=>"110110100",
  9669=>"111010010",
  9670=>"000010001",
  9671=>"000000111",
  9672=>"000000100",
  9673=>"111101000",
  9674=>"101100000",
  9675=>"000000110",
  9676=>"010111001",
  9677=>"100111011",
  9678=>"110010010",
  9679=>"000100100",
  9680=>"000000000",
  9681=>"000000001",
  9682=>"000000000",
  9683=>"111111111",
  9684=>"111111000",
  9685=>"000000000",
  9686=>"000000110",
  9687=>"011010010",
  9688=>"100000001",
  9689=>"001000000",
  9690=>"110000000",
  9691=>"100100100",
  9692=>"000000000",
  9693=>"111111111",
  9694=>"000000000",
  9695=>"110110100",
  9696=>"000000000",
  9697=>"111111111",
  9698=>"111001111",
  9699=>"111111111",
  9700=>"110000011",
  9701=>"001001001",
  9702=>"011111111",
  9703=>"111110000",
  9704=>"101100101",
  9705=>"111111110",
  9706=>"000000010",
  9707=>"000010111",
  9708=>"111111111",
  9709=>"110111010",
  9710=>"000001111",
  9711=>"001111100",
  9712=>"010000000",
  9713=>"111111110",
  9714=>"111111111",
  9715=>"100000100",
  9716=>"010111111",
  9717=>"001001000",
  9718=>"111111001",
  9719=>"000000100",
  9720=>"010111110",
  9721=>"100100000",
  9722=>"000001111",
  9723=>"111111111",
  9724=>"000001000",
  9725=>"001001111",
  9726=>"110111111",
  9727=>"000000001",
  9728=>"000001001",
  9729=>"000110111",
  9730=>"000001111",
  9731=>"000000001",
  9732=>"000000011",
  9733=>"111000000",
  9734=>"110111010",
  9735=>"010111101",
  9736=>"111001011",
  9737=>"111111111",
  9738=>"111001111",
  9739=>"000111111",
  9740=>"000001001",
  9741=>"011000001",
  9742=>"000111011",
  9743=>"111110010",
  9744=>"110110110",
  9745=>"010110110",
  9746=>"000000001",
  9747=>"110000010",
  9748=>"000101111",
  9749=>"101101001",
  9750=>"000000011",
  9751=>"101111111",
  9752=>"000001001",
  9753=>"111111011",
  9754=>"000000000",
  9755=>"100000000",
  9756=>"101101111",
  9757=>"011011001",
  9758=>"000100100",
  9759=>"000000000",
  9760=>"110110000",
  9761=>"000000000",
  9762=>"111111010",
  9763=>"111010000",
  9764=>"000000111",
  9765=>"000000000",
  9766=>"011000110",
  9767=>"100100111",
  9768=>"000000000",
  9769=>"101101111",
  9770=>"100101111",
  9771=>"000001000",
  9772=>"111111111",
  9773=>"001111111",
  9774=>"000001001",
  9775=>"011011011",
  9776=>"110110010",
  9777=>"111001000",
  9778=>"001000001",
  9779=>"000000000",
  9780=>"101111001",
  9781=>"010001001",
  9782=>"111100000",
  9783=>"111111111",
  9784=>"000101111",
  9785=>"001110111",
  9786=>"001000000",
  9787=>"011000000",
  9788=>"000000000",
  9789=>"011111110",
  9790=>"001000010",
  9791=>"111111111",
  9792=>"111111111",
  9793=>"110110001",
  9794=>"000000011",
  9795=>"111111000",
  9796=>"110110111",
  9797=>"000000100",
  9798=>"000000000",
  9799=>"011000000",
  9800=>"001001001",
  9801=>"101101000",
  9802=>"000001000",
  9803=>"010000000",
  9804=>"001000001",
  9805=>"111101110",
  9806=>"111101101",
  9807=>"111110111",
  9808=>"110111110",
  9809=>"111101000",
  9810=>"000000101",
  9811=>"000010100",
  9812=>"001000000",
  9813=>"111101101",
  9814=>"000000101",
  9815=>"011000000",
  9816=>"111111111",
  9817=>"100100000",
  9818=>"111001001",
  9819=>"110110100",
  9820=>"000000111",
  9821=>"110000000",
  9822=>"000000000",
  9823=>"000111011",
  9824=>"000001000",
  9825=>"101111111",
  9826=>"000010000",
  9827=>"111100100",
  9828=>"001001111",
  9829=>"110110110",
  9830=>"111110000",
  9831=>"000000000",
  9832=>"101000101",
  9833=>"000101111",
  9834=>"110110111",
  9835=>"000000000",
  9836=>"000000100",
  9837=>"000001111",
  9838=>"000000100",
  9839=>"000000100",
  9840=>"111111111",
  9841=>"010010000",
  9842=>"111011111",
  9843=>"111111111",
  9844=>"000000000",
  9845=>"000010010",
  9846=>"111000000",
  9847=>"001101111",
  9848=>"110110000",
  9849=>"011111110",
  9850=>"000000110",
  9851=>"001001001",
  9852=>"110110100",
  9853=>"000000000",
  9854=>"000000111",
  9855=>"000001001",
  9856=>"100110110",
  9857=>"111110110",
  9858=>"000001101",
  9859=>"000000111",
  9860=>"000011111",
  9861=>"111111000",
  9862=>"000010000",
  9863=>"000000000",
  9864=>"000000000",
  9865=>"111000000",
  9866=>"110000111",
  9867=>"000000111",
  9868=>"111111000",
  9869=>"011001111",
  9870=>"000001111",
  9871=>"110110110",
  9872=>"101001101",
  9873=>"000000000",
  9874=>"111111111",
  9875=>"110111101",
  9876=>"000000110",
  9877=>"010010000",
  9878=>"000000000",
  9879=>"000000000",
  9880=>"110110000",
  9881=>"000111111",
  9882=>"010010110",
  9883=>"001001001",
  9884=>"000000000",
  9885=>"110110110",
  9886=>"011111111",
  9887=>"111111111",
  9888=>"000000000",
  9889=>"000000100",
  9890=>"001000001",
  9891=>"000000101",
  9892=>"000100100",
  9893=>"011011100",
  9894=>"001000111",
  9895=>"011001100",
  9896=>"100101100",
  9897=>"000000000",
  9898=>"110111001",
  9899=>"111000111",
  9900=>"000000110",
  9901=>"001001111",
  9902=>"000000110",
  9903=>"000110000",
  9904=>"000011111",
  9905=>"110110100",
  9906=>"000111111",
  9907=>"000000000",
  9908=>"000000000",
  9909=>"111111111",
  9910=>"000000010",
  9911=>"100111001",
  9912=>"000000000",
  9913=>"000000110",
  9914=>"000000010",
  9915=>"110110101",
  9916=>"111001001",
  9917=>"001001001",
  9918=>"111111000",
  9919=>"111110000",
  9920=>"001000111",
  9921=>"000000111",
  9922=>"111001111",
  9923=>"000010000",
  9924=>"001011001",
  9925=>"000010010",
  9926=>"000000000",
  9927=>"000000000",
  9928=>"110110110",
  9929=>"101001111",
  9930=>"111101101",
  9931=>"000000000",
  9932=>"000000000",
  9933=>"001001000",
  9934=>"000101111",
  9935=>"000001001",
  9936=>"110010010",
  9937=>"000000000",
  9938=>"011000000",
  9939=>"000000000",
  9940=>"111111000",
  9941=>"001111111",
  9942=>"111000001",
  9943=>"011100000",
  9944=>"001001001",
  9945=>"000001000",
  9946=>"101101101",
  9947=>"001111111",
  9948=>"001000000",
  9949=>"111111011",
  9950=>"000000111",
  9951=>"000000101",
  9952=>"111111111",
  9953=>"111111111",
  9954=>"111110000",
  9955=>"000000111",
  9956=>"111111110",
  9957=>"011011011",
  9958=>"001001111",
  9959=>"010110010",
  9960=>"111111100",
  9961=>"000001001",
  9962=>"111111111",
  9963=>"000000000",
  9964=>"000000101",
  9965=>"111111111",
  9966=>"110000010",
  9967=>"101000000",
  9968=>"000000000",
  9969=>"000000011",
  9970=>"111101101",
  9971=>"000000000",
  9972=>"011011000",
  9973=>"100110110",
  9974=>"100000000",
  9975=>"001000000",
  9976=>"110111111",
  9977=>"000000000",
  9978=>"111111111",
  9979=>"011000011",
  9980=>"100001011",
  9981=>"100000001",
  9982=>"001101111",
  9983=>"110111110",
  9984=>"000001111",
  9985=>"011011001",
  9986=>"000000000",
  9987=>"111101111",
  9988=>"111111001",
  9989=>"000111111",
  9990=>"110110100",
  9991=>"010010000",
  9992=>"000000100",
  9993=>"111111111",
  9994=>"111111110",
  9995=>"110110110",
  9996=>"001000000",
  9997=>"111111011",
  9998=>"010000110",
  9999=>"011000000",
  10000=>"010001101",
  10001=>"000001001",
  10002=>"101000101",
  10003=>"101101111",
  10004=>"110111000",
  10005=>"100100100",
  10006=>"001001101",
  10007=>"000000000",
  10008=>"000010011",
  10009=>"111000111",
  10010=>"000000000",
  10011=>"000010000",
  10012=>"101111001",
  10013=>"001000101",
  10014=>"111000000",
  10015=>"110010011",
  10016=>"000000011",
  10017=>"001000000",
  10018=>"000000100",
  10019=>"010110110",
  10020=>"111111111",
  10021=>"111011111",
  10022=>"001000100",
  10023=>"100000001",
  10024=>"110111011",
  10025=>"000000000",
  10026=>"000000110",
  10027=>"111111111",
  10028=>"001010010",
  10029=>"111011111",
  10030=>"011111011",
  10031=>"000000000",
  10032=>"101111111",
  10033=>"010000000",
  10034=>"111111101",
  10035=>"000111010",
  10036=>"011011010",
  10037=>"000000000",
  10038=>"111111011",
  10039=>"110110000",
  10040=>"000000010",
  10041=>"000000000",
  10042=>"011010111",
  10043=>"001111111",
  10044=>"110010001",
  10045=>"001001001",
  10046=>"000000001",
  10047=>"110010000",
  10048=>"000000000",
  10049=>"000000000",
  10050=>"110101111",
  10051=>"001000001",
  10052=>"111111111",
  10053=>"001101111",
  10054=>"000000000",
  10055=>"111111111",
  10056=>"000000111",
  10057=>"110010000",
  10058=>"110110110",
  10059=>"000000000",
  10060=>"010111000",
  10061=>"100111111",
  10062=>"111111110",
  10063=>"110110100",
  10064=>"000001001",
  10065=>"000000001",
  10066=>"111111010",
  10067=>"011000000",
  10068=>"000000000",
  10069=>"011011011",
  10070=>"010011111",
  10071=>"111001111",
  10072=>"100000000",
  10073=>"001100001",
  10074=>"000110111",
  10075=>"000000000",
  10076=>"100110100",
  10077=>"000000000",
  10078=>"000000111",
  10079=>"110000110",
  10080=>"110100110",
  10081=>"111000000",
  10082=>"000001011",
  10083=>"000000010",
  10084=>"100001001",
  10085=>"001101101",
  10086=>"111111111",
  10087=>"011011101",
  10088=>"000001111",
  10089=>"000000000",
  10090=>"001000001",
  10091=>"101100110",
  10092=>"001000100",
  10093=>"000000000",
  10094=>"100101001",
  10095=>"000000111",
  10096=>"000000000",
  10097=>"001001111",
  10098=>"000001001",
  10099=>"011011011",
  10100=>"111111000",
  10101=>"001001000",
  10102=>"111101001",
  10103=>"110000000",
  10104=>"001000100",
  10105=>"000000000",
  10106=>"110000000",
  10107=>"011111011",
  10108=>"001000111",
  10109=>"000000110",
  10110=>"000000000",
  10111=>"000111111",
  10112=>"110110110",
  10113=>"000011011",
  10114=>"000000000",
  10115=>"111000000",
  10116=>"000000111",
  10117=>"000011111",
  10118=>"001001101",
  10119=>"110111111",
  10120=>"111101101",
  10121=>"010011111",
  10122=>"101001101",
  10123=>"000110111",
  10124=>"100111111",
  10125=>"000010110",
  10126=>"100111111",
  10127=>"000000011",
  10128=>"000000000",
  10129=>"010010010",
  10130=>"000000000",
  10131=>"101001101",
  10132=>"000000000",
  10133=>"000000000",
  10134=>"011000000",
  10135=>"001001111",
  10136=>"000001001",
  10137=>"110110110",
  10138=>"011111011",
  10139=>"110111111",
  10140=>"011000001",
  10141=>"000001001",
  10142=>"000000000",
  10143=>"000111111",
  10144=>"010000000",
  10145=>"111011001",
  10146=>"011011101",
  10147=>"111111111",
  10148=>"000011111",
  10149=>"010011000",
  10150=>"001001011",
  10151=>"111111111",
  10152=>"011000111",
  10153=>"000110110",
  10154=>"011000001",
  10155=>"000010111",
  10156=>"000000000",
  10157=>"000000101",
  10158=>"000010110",
  10159=>"001000000",
  10160=>"111111111",
  10161=>"001111011",
  10162=>"011111000",
  10163=>"001001101",
  10164=>"111110111",
  10165=>"000010000",
  10166=>"110000001",
  10167=>"111111111",
  10168=>"000000000",
  10169=>"011111111",
  10170=>"110100111",
  10171=>"111111111",
  10172=>"111101001",
  10173=>"000110111",
  10174=>"001000000",
  10175=>"010001001",
  10176=>"101111111",
  10177=>"001101000",
  10178=>"111111111",
  10179=>"110111111",
  10180=>"111111110",
  10181=>"011011011",
  10182=>"000100111",
  10183=>"001001101",
  10184=>"000110111",
  10185=>"000001111",
  10186=>"000001100",
  10187=>"011000000",
  10188=>"000100110",
  10189=>"110110000",
  10190=>"000000010",
  10191=>"000000000",
  10192=>"000001111",
  10193=>"110110010",
  10194=>"001111111",
  10195=>"000000000",
  10196=>"000110111",
  10197=>"111111011",
  10198=>"111111111",
  10199=>"001001111",
  10200=>"111110010",
  10201=>"011000000",
  10202=>"111111111",
  10203=>"111000111",
  10204=>"111011111",
  10205=>"110110110",
  10206=>"000000011",
  10207=>"001000000",
  10208=>"001110110",
  10209=>"000111111",
  10210=>"100110000",
  10211=>"001000111",
  10212=>"000000000",
  10213=>"110000000",
  10214=>"100000000",
  10215=>"101101111",
  10216=>"000100110",
  10217=>"111111110",
  10218=>"111101111",
  10219=>"100110100",
  10220=>"110110010",
  10221=>"000000110",
  10222=>"000000101",
  10223=>"111110010",
  10224=>"000000001",
  10225=>"111111001",
  10226=>"111101101",
  10227=>"000000001",
  10228=>"000001111",
  10229=>"111011000",
  10230=>"011011001",
  10231=>"111111111",
  10232=>"000000000",
  10233=>"000000100",
  10234=>"000111111",
  10235=>"111111001",
  10236=>"001001111",
  10237=>"000000000",
  10238=>"000000000",
  10239=>"001000001",
  10240=>"111111111",
  10241=>"011010100",
  10242=>"111000000",
  10243=>"100111110",
  10244=>"111000100",
  10245=>"110000101",
  10246=>"111000010",
  10247=>"111111111",
  10248=>"110001111",
  10249=>"000000101",
  10250=>"111111001",
  10251=>"110111111",
  10252=>"111011011",
  10253=>"000111111",
  10254=>"000000111",
  10255=>"010000000",
  10256=>"101110111",
  10257=>"111111011",
  10258=>"111110111",
  10259=>"111111111",
  10260=>"111111111",
  10261=>"111101111",
  10262=>"100000000",
  10263=>"111100000",
  10264=>"011111011",
  10265=>"001001101",
  10266=>"100111101",
  10267=>"000000000",
  10268=>"111111111",
  10269=>"000010000",
  10270=>"111111111",
  10271=>"111111111",
  10272=>"111111111",
  10273=>"110111110",
  10274=>"110110000",
  10275=>"111011010",
  10276=>"100000000",
  10277=>"000000000",
  10278=>"111111011",
  10279=>"011000000",
  10280=>"110100100",
  10281=>"111111000",
  10282=>"011111111",
  10283=>"000000000",
  10284=>"000000000",
  10285=>"110111111",
  10286=>"011011011",
  10287=>"111111111",
  10288=>"000110000",
  10289=>"111111111",
  10290=>"111111111",
  10291=>"111111101",
  10292=>"100000000",
  10293=>"000000000",
  10294=>"010000000",
  10295=>"100111111",
  10296=>"011011011",
  10297=>"000000000",
  10298=>"000000000",
  10299=>"011001111",
  10300=>"100110111",
  10301=>"000000000",
  10302=>"000000110",
  10303=>"000000000",
  10304=>"000000000",
  10305=>"000000000",
  10306=>"110111011",
  10307=>"000001001",
  10308=>"000000011",
  10309=>"111111111",
  10310=>"001111111",
  10311=>"000000000",
  10312=>"000001001",
  10313=>"000000000",
  10314=>"111111001",
  10315=>"101111111",
  10316=>"111111111",
  10317=>"011011111",
  10318=>"111000000",
  10319=>"010111000",
  10320=>"001000000",
  10321=>"000000000",
  10322=>"111111110",
  10323=>"110100100",
  10324=>"000000100",
  10325=>"000000000",
  10326=>"000011000",
  10327=>"110100000",
  10328=>"010000000",
  10329=>"000000111",
  10330=>"100001111",
  10331=>"110001111",
  10332=>"111111111",
  10333=>"000000000",
  10334=>"101111011",
  10335=>"100111111",
  10336=>"110111111",
  10337=>"000101101",
  10338=>"111110000",
  10339=>"011001101",
  10340=>"000000011",
  10341=>"001001101",
  10342=>"111111111",
  10343=>"000000000",
  10344=>"001000000",
  10345=>"001001000",
  10346=>"000000111",
  10347=>"001000000",
  10348=>"011111111",
  10349=>"111111010",
  10350=>"111111111",
  10351=>"111110111",
  10352=>"000000000",
  10353=>"010000000",
  10354=>"000000000",
  10355=>"110111111",
  10356=>"101100100",
  10357=>"000001111",
  10358=>"101111111",
  10359=>"011111000",
  10360=>"111111111",
  10361=>"011000100",
  10362=>"111111110",
  10363=>"111111111",
  10364=>"000000110",
  10365=>"000111101",
  10366=>"011110010",
  10367=>"001000101",
  10368=>"111000111",
  10369=>"100101001",
  10370=>"000000000",
  10371=>"100110111",
  10372=>"111100101",
  10373=>"110100110",
  10374=>"111111111",
  10375=>"000111111",
  10376=>"000000000",
  10377=>"111111011",
  10378=>"011111111",
  10379=>"011111111",
  10380=>"010000001",
  10381=>"000000000",
  10382=>"010000000",
  10383=>"100000111",
  10384=>"111011011",
  10385=>"000000101",
  10386=>"111010000",
  10387=>"000000001",
  10388=>"000110100",
  10389=>"111111111",
  10390=>"110000000",
  10391=>"100101111",
  10392=>"110100000",
  10393=>"111100000",
  10394=>"000000000",
  10395=>"000000001",
  10396=>"000000000",
  10397=>"011001101",
  10398=>"000001111",
  10399=>"101111111",
  10400=>"111101000",
  10401=>"000000001",
  10402=>"111111111",
  10403=>"111111111",
  10404=>"111011011",
  10405=>"011001011",
  10406=>"111111111",
  10407=>"000110110",
  10408=>"000000000",
  10409=>"111000100",
  10410=>"110110010",
  10411=>"000000000",
  10412=>"001110011",
  10413=>"001001001",
  10414=>"111111110",
  10415=>"111111100",
  10416=>"000000000",
  10417=>"000100111",
  10418=>"111101111",
  10419=>"111111111",
  10420=>"110111111",
  10421=>"000011100",
  10422=>"110000000",
  10423=>"000000000",
  10424=>"011001000",
  10425=>"000000000",
  10426=>"110000000",
  10427=>"011010111",
  10428=>"000000000",
  10429=>"111111111",
  10430=>"111111000",
  10431=>"111111111",
  10432=>"000000000",
  10433=>"000000000",
  10434=>"110110111",
  10435=>"111111111",
  10436=>"111011000",
  10437=>"000000000",
  10438=>"011001111",
  10439=>"100100111",
  10440=>"000000000",
  10441=>"000000011",
  10442=>"011000000",
  10443=>"111111110",
  10444=>"000010110",
  10445=>"111110000",
  10446=>"001001111",
  10447=>"100111111",
  10448=>"111000100",
  10449=>"011010000",
  10450=>"000000001",
  10451=>"100100111",
  10452=>"110111011",
  10453=>"111111111",
  10454=>"000000000",
  10455=>"000000100",
  10456=>"111111111",
  10457=>"000000000",
  10458=>"000000000",
  10459=>"111111011",
  10460=>"001000000",
  10461=>"111111111",
  10462=>"111111000",
  10463=>"011111111",
  10464=>"000100111",
  10465=>"111111111",
  10466=>"000100110",
  10467=>"000000111",
  10468=>"000011111",
  10469=>"111111111",
  10470=>"000000001",
  10471=>"001000110",
  10472=>"101101111",
  10473=>"010111001",
  10474=>"110111111",
  10475=>"000000010",
  10476=>"000000000",
  10477=>"111001000",
  10478=>"111010000",
  10479=>"000000111",
  10480=>"011111111",
  10481=>"111111111",
  10482=>"100100000",
  10483=>"010110000",
  10484=>"100111111",
  10485=>"001111111",
  10486=>"111111100",
  10487=>"100010000",
  10488=>"001001001",
  10489=>"111101101",
  10490=>"011111110",
  10491=>"000000000",
  10492=>"011011011",
  10493=>"000100000",
  10494=>"111111110",
  10495=>"111111001",
  10496=>"111111000",
  10497=>"111111111",
  10498=>"111111111",
  10499=>"111101111",
  10500=>"000000000",
  10501=>"000000000",
  10502=>"010111111",
  10503=>"011011000",
  10504=>"111111011",
  10505=>"001000001",
  10506=>"111111101",
  10507=>"000001011",
  10508=>"001001111",
  10509=>"000110000",
  10510=>"000000001",
  10511=>"000000101",
  10512=>"111111111",
  10513=>"111111111",
  10514=>"000000010",
  10515=>"011011011",
  10516=>"111111100",
  10517=>"100011000",
  10518=>"011110100",
  10519=>"111111000",
  10520=>"111111111",
  10521=>"111111010",
  10522=>"000000000",
  10523=>"000100000",
  10524=>"000000000",
  10525=>"111111000",
  10526=>"000111111",
  10527=>"111111101",
  10528=>"111111011",
  10529=>"110110100",
  10530=>"011011000",
  10531=>"000000000",
  10532=>"111111011",
  10533=>"000000000",
  10534=>"011011111",
  10535=>"111111000",
  10536=>"111111111",
  10537=>"001000000",
  10538=>"000010001",
  10539=>"100111111",
  10540=>"000000111",
  10541=>"001001001",
  10542=>"111111111",
  10543=>"101111111",
  10544=>"011011000",
  10545=>"111111111",
  10546=>"100000000",
  10547=>"111110010",
  10548=>"111101101",
  10549=>"100011110",
  10550=>"110101101",
  10551=>"111111100",
  10552=>"000000001",
  10553=>"000000001",
  10554=>"111111110",
  10555=>"000000000",
  10556=>"111111111",
  10557=>"110111111",
  10558=>"000111111",
  10559=>"111000111",
  10560=>"001001111",
  10561=>"111111111",
  10562=>"111111111",
  10563=>"111111111",
  10564=>"111111111",
  10565=>"011111111",
  10566=>"110111111",
  10567=>"111111101",
  10568=>"100110100",
  10569=>"100000101",
  10570=>"000000100",
  10571=>"100100101",
  10572=>"111111100",
  10573=>"000100000",
  10574=>"111011011",
  10575=>"000001001",
  10576=>"000000110",
  10577=>"001011010",
  10578=>"100100000",
  10579=>"111111111",
  10580=>"111010011",
  10581=>"000000000",
  10582=>"111000000",
  10583=>"010110110",
  10584=>"011011011",
  10585=>"001001001",
  10586=>"011110111",
  10587=>"111111000",
  10588=>"011110110",
  10589=>"000000000",
  10590=>"010000000",
  10591=>"111010000",
  10592=>"000000000",
  10593=>"111111111",
  10594=>"110111111",
  10595=>"011000000",
  10596=>"000110000",
  10597=>"000110100",
  10598=>"000000000",
  10599=>"000000000",
  10600=>"000100100",
  10601=>"000000000",
  10602=>"000000001",
  10603=>"111111111",
  10604=>"011001000",
  10605=>"111000111",
  10606=>"000000110",
  10607=>"111111111",
  10608=>"000100100",
  10609=>"111111010",
  10610=>"000000000",
  10611=>"011001111",
  10612=>"001001000",
  10613=>"111000101",
  10614=>"111001000",
  10615=>"001101111",
  10616=>"111111011",
  10617=>"000001111",
  10618=>"000000000",
  10619=>"100111111",
  10620=>"100110111",
  10621=>"111111011",
  10622=>"000000000",
  10623=>"000000000",
  10624=>"000110010",
  10625=>"111100101",
  10626=>"011111111",
  10627=>"000000000",
  10628=>"000000111",
  10629=>"111111111",
  10630=>"111100110",
  10631=>"110111111",
  10632=>"111001101",
  10633=>"000001111",
  10634=>"010010000",
  10635=>"111101100",
  10636=>"000000000",
  10637=>"110010001",
  10638=>"011000000",
  10639=>"111001111",
  10640=>"111111111",
  10641=>"111000000",
  10642=>"111111000",
  10643=>"111011011",
  10644=>"001000101",
  10645=>"110111101",
  10646=>"111010000",
  10647=>"011111110",
  10648=>"010111111",
  10649=>"001011011",
  10650=>"010111111",
  10651=>"000000001",
  10652=>"100000101",
  10653=>"001001111",
  10654=>"000000000",
  10655=>"111111111",
  10656=>"000000000",
  10657=>"111110100",
  10658=>"000000000",
  10659=>"111111111",
  10660=>"110111111",
  10661=>"110111111",
  10662=>"100110111",
  10663=>"000000000",
  10664=>"001000000",
  10665=>"000101100",
  10666=>"111111111",
  10667=>"000000101",
  10668=>"100111111",
  10669=>"000000110",
  10670=>"000000000",
  10671=>"111111111",
  10672=>"000000000",
  10673=>"000000000",
  10674=>"000111111",
  10675=>"111111111",
  10676=>"100000111",
  10677=>"101001000",
  10678=>"011011101",
  10679=>"111001001",
  10680=>"001011011",
  10681=>"111111111",
  10682=>"001001111",
  10683=>"000001110",
  10684=>"000101111",
  10685=>"011011001",
  10686=>"000110111",
  10687=>"011011111",
  10688=>"111001100",
  10689=>"001001001",
  10690=>"111111111",
  10691=>"000000000",
  10692=>"000000000",
  10693=>"111111001",
  10694=>"010000000",
  10695=>"000101111",
  10696=>"111011111",
  10697=>"100010000",
  10698=>"110000101",
  10699=>"111111111",
  10700=>"000000111",
  10701=>"111111001",
  10702=>"110100101",
  10703=>"000000000",
  10704=>"001001101",
  10705=>"111111111",
  10706=>"111011011",
  10707=>"000000000",
  10708=>"111111110",
  10709=>"111111000",
  10710=>"111111111",
  10711=>"011111100",
  10712=>"000000000",
  10713=>"000000000",
  10714=>"111111111",
  10715=>"000000010",
  10716=>"010101111",
  10717=>"000000000",
  10718=>"101100111",
  10719=>"111111111",
  10720=>"011111100",
  10721=>"100000000",
  10722=>"111111111",
  10723=>"000000000",
  10724=>"111011010",
  10725=>"110011011",
  10726=>"011110111",
  10727=>"000000000",
  10728=>"100111001",
  10729=>"101001111",
  10730=>"000000110",
  10731=>"011000000",
  10732=>"000000100",
  10733=>"110110110",
  10734=>"111111111",
  10735=>"010000000",
  10736=>"111111111",
  10737=>"010000100",
  10738=>"000011001",
  10739=>"000001111",
  10740=>"110111111",
  10741=>"100100110",
  10742=>"011000000",
  10743=>"111111111",
  10744=>"101111111",
  10745=>"000000000",
  10746=>"000000001",
  10747=>"001111001",
  10748=>"110011111",
  10749=>"001001000",
  10750=>"001111001",
  10751=>"111000101",
  10752=>"000000100",
  10753=>"111011001",
  10754=>"111111111",
  10755=>"111011001",
  10756=>"100001101",
  10757=>"000000000",
  10758=>"101111001",
  10759=>"101101111",
  10760=>"111111111",
  10761=>"111000001",
  10762=>"111110100",
  10763=>"011011001",
  10764=>"110000000",
  10765=>"011011111",
  10766=>"111110111",
  10767=>"111111111",
  10768=>"111111111",
  10769=>"111011111",
  10770=>"000011111",
  10771=>"000000000",
  10772=>"111111111",
  10773=>"000100111",
  10774=>"000000000",
  10775=>"000000000",
  10776=>"000000000",
  10777=>"000000000",
  10778=>"000000111",
  10779=>"101000100",
  10780=>"100000000",
  10781=>"101001001",
  10782=>"100110110",
  10783=>"000100100",
  10784=>"000000000",
  10785=>"111111011",
  10786=>"111111111",
  10787=>"111000111",
  10788=>"000000110",
  10789=>"011011111",
  10790=>"110010000",
  10791=>"110100110",
  10792=>"000000111",
  10793=>"111111111",
  10794=>"110000100",
  10795=>"001000000",
  10796=>"110000100",
  10797=>"000000000",
  10798=>"011011011",
  10799=>"000100100",
  10800=>"000000000",
  10801=>"000000000",
  10802=>"110110110",
  10803=>"000000001",
  10804=>"000000000",
  10805=>"001000100",
  10806=>"100100000",
  10807=>"011000000",
  10808=>"111111110",
  10809=>"000000000",
  10810=>"000000101",
  10811=>"000000000",
  10812=>"000000100",
  10813=>"111110111",
  10814=>"100000000",
  10815=>"111011100",
  10816=>"111101111",
  10817=>"111111111",
  10818=>"111111000",
  10819=>"111101001",
  10820=>"110000000",
  10821=>"000001000",
  10822=>"110110111",
  10823=>"000000000",
  10824=>"100100100",
  10825=>"101101111",
  10826=>"000000000",
  10827=>"000111111",
  10828=>"100000000",
  10829=>"111000011",
  10830=>"000010000",
  10831=>"000000000",
  10832=>"111111111",
  10833=>"000000100",
  10834=>"000000000",
  10835=>"110111110",
  10836=>"000000000",
  10837=>"000000100",
  10838=>"000110111",
  10839=>"000000000",
  10840=>"000000000",
  10841=>"000000111",
  10842=>"111111111",
  10843=>"111111111",
  10844=>"011111111",
  10845=>"000000000",
  10846=>"111111111",
  10847=>"010111110",
  10848=>"111010000",
  10849=>"011011000",
  10850=>"000100100",
  10851=>"000000000",
  10852=>"110101101",
  10853=>"000000000",
  10854=>"011011111",
  10855=>"111111001",
  10856=>"111111000",
  10857=>"011111111",
  10858=>"000000000",
  10859=>"110111111",
  10860=>"000000001",
  10861=>"111011111",
  10862=>"111111001",
  10863=>"011111011",
  10864=>"111000000",
  10865=>"110110010",
  10866=>"010110110",
  10867=>"000000000",
  10868=>"000000000",
  10869=>"000000000",
  10870=>"000000000",
  10871=>"000001111",
  10872=>"110111110",
  10873=>"000000000",
  10874=>"011011011",
  10875=>"000000000",
  10876=>"110100110",
  10877=>"000000000",
  10878=>"000000000",
  10879=>"000000000",
  10880=>"111111111",
  10881=>"001000000",
  10882=>"101101111",
  10883=>"111001000",
  10884=>"111001011",
  10885=>"111111111",
  10886=>"000001000",
  10887=>"100000000",
  10888=>"001011111",
  10889=>"111101001",
  10890=>"000001111",
  10891=>"000000000",
  10892=>"111111111",
  10893=>"111111110",
  10894=>"000000000",
  10895=>"111111111",
  10896=>"111111111",
  10897=>"010000010",
  10898=>"111111111",
  10899=>"111111111",
  10900=>"111001000",
  10901=>"000000000",
  10902=>"000001111",
  10903=>"000000000",
  10904=>"000000000",
  10905=>"001100110",
  10906=>"111111011",
  10907=>"111111111",
  10908=>"011000000",
  10909=>"100000100",
  10910=>"111101000",
  10911=>"111111111",
  10912=>"101111111",
  10913=>"011010110",
  10914=>"000000100",
  10915=>"111111111",
  10916=>"000000011",
  10917=>"100100000",
  10918=>"000000111",
  10919=>"001000001",
  10920=>"111111111",
  10921=>"000111111",
  10922=>"111111111",
  10923=>"001100000",
  10924=>"011000011",
  10925=>"000000100",
  10926=>"000000110",
  10927=>"000000111",
  10928=>"111111110",
  10929=>"000000000",
  10930=>"110110111",
  10931=>"000000010",
  10932=>"111111111",
  10933=>"111011011",
  10934=>"000001111",
  10935=>"111101101",
  10936=>"000000000",
  10937=>"000000111",
  10938=>"100111111",
  10939=>"101000001",
  10940=>"000010111",
  10941=>"101100111",
  10942=>"000110111",
  10943=>"000111101",
  10944=>"000000000",
  10945=>"111111111",
  10946=>"000000000",
  10947=>"000000000",
  10948=>"101000100",
  10949=>"001001000",
  10950=>"000100111",
  10951=>"111111111",
  10952=>"000011011",
  10953=>"000100000",
  10954=>"000111111",
  10955=>"001011111",
  10956=>"111111100",
  10957=>"000001100",
  10958=>"100110111",
  10959=>"111111101",
  10960=>"000111111",
  10961=>"110000000",
  10962=>"000000000",
  10963=>"111111111",
  10964=>"111111111",
  10965=>"111000000",
  10966=>"000000001",
  10967=>"000110100",
  10968=>"010000000",
  10969=>"111111100",
  10970=>"111111111",
  10971=>"110110111",
  10972=>"111100100",
  10973=>"011111110",
  10974=>"101100100",
  10975=>"111111111",
  10976=>"111000100",
  10977=>"111111111",
  10978=>"000100111",
  10979=>"111111001",
  10980=>"111111111",
  10981=>"111111111",
  10982=>"101111110",
  10983=>"111111111",
  10984=>"110100011",
  10985=>"000000000",
  10986=>"111111111",
  10987=>"000000000",
  10988=>"000000000",
  10989=>"111111111",
  10990=>"000000000",
  10991=>"000000100",
  10992=>"001111111",
  10993=>"001000000",
  10994=>"000111110",
  10995=>"001001000",
  10996=>"011111011",
  10997=>"001011011",
  10998=>"000100110",
  10999=>"111111111",
  11000=>"001000000",
  11001=>"011111001",
  11002=>"111100000",
  11003=>"000000000",
  11004=>"111111111",
  11005=>"111101111",
  11006=>"000000000",
  11007=>"111111110",
  11008=>"111111111",
  11009=>"001001101",
  11010=>"111111111",
  11011=>"011001000",
  11012=>"000000000",
  11013=>"000000100",
  11014=>"000100100",
  11015=>"111110100",
  11016=>"111111111",
  11017=>"000000000",
  11018=>"111001000",
  11019=>"100000000",
  11020=>"000000000",
  11021=>"000000000",
  11022=>"000000000",
  11023=>"011001001",
  11024=>"000000001",
  11025=>"000000110",
  11026=>"111111111",
  11027=>"000000001",
  11028=>"000001001",
  11029=>"111000001",
  11030=>"110111110",
  11031=>"000000100",
  11032=>"100100100",
  11033=>"000000000",
  11034=>"100100100",
  11035=>"000000110",
  11036=>"111011111",
  11037=>"001101111",
  11038=>"111111111",
  11039=>"111111000",
  11040=>"000000110",
  11041=>"000000000",
  11042=>"111111111",
  11043=>"111111111",
  11044=>"000000000",
  11045=>"100100000",
  11046=>"001001111",
  11047=>"111111111",
  11048=>"000000000",
  11049=>"110110100",
  11050=>"011111100",
  11051=>"000111111",
  11052=>"111111100",
  11053=>"110010110",
  11054=>"000011111",
  11055=>"101101000",
  11056=>"111100100",
  11057=>"111111000",
  11058=>"111111111",
  11059=>"000110110",
  11060=>"111111111",
  11061=>"110011011",
  11062=>"111000000",
  11063=>"111111111",
  11064=>"111100000",
  11065=>"011111111",
  11066=>"000000011",
  11067=>"111111111",
  11068=>"100100100",
  11069=>"110000100",
  11070=>"100111111",
  11071=>"111111100",
  11072=>"000111000",
  11073=>"011011111",
  11074=>"111110000",
  11075=>"000111111",
  11076=>"000000100",
  11077=>"000000000",
  11078=>"111111111",
  11079=>"000000000",
  11080=>"000000000",
  11081=>"111111111",
  11082=>"000000111",
  11083=>"111111110",
  11084=>"111111111",
  11085=>"101101000",
  11086=>"111100100",
  11087=>"000000000",
  11088=>"100100000",
  11089=>"000011111",
  11090=>"110111111",
  11091=>"000000000",
  11092=>"100010011",
  11093=>"011011011",
  11094=>"011011011",
  11095=>"111111111",
  11096=>"111111111",
  11097=>"000000111",
  11098=>"111100100",
  11099=>"111111100",
  11100=>"000000010",
  11101=>"011001011",
  11102=>"011111110",
  11103=>"111111111",
  11104=>"110110100",
  11105=>"001001001",
  11106=>"001001001",
  11107=>"111001001",
  11108=>"000011110",
  11109=>"000000000",
  11110=>"111000000",
  11111=>"011001001",
  11112=>"111111111",
  11113=>"001001011",
  11114=>"000000000",
  11115=>"111101001",
  11116=>"111011001",
  11117=>"111011001",
  11118=>"011100000",
  11119=>"011011110",
  11120=>"000000000",
  11121=>"000001000",
  11122=>"001000001",
  11123=>"000000000",
  11124=>"000000000",
  11125=>"101101111",
  11126=>"110100000",
  11127=>"111111111",
  11128=>"000000001",
  11129=>"000000110",
  11130=>"111111111",
  11131=>"111110100",
  11132=>"000000000",
  11133=>"111111111",
  11134=>"101111111",
  11135=>"111111111",
  11136=>"000000000",
  11137=>"001000000",
  11138=>"110110000",
  11139=>"111111111",
  11140=>"111111111",
  11141=>"111111110",
  11142=>"111111111",
  11143=>"111011000",
  11144=>"111111001",
  11145=>"111000000",
  11146=>"000000000",
  11147=>"111000111",
  11148=>"111111111",
  11149=>"110100100",
  11150=>"111110110",
  11151=>"000000000",
  11152=>"111111111",
  11153=>"000000000",
  11154=>"100010111",
  11155=>"000000000",
  11156=>"111111011",
  11157=>"100000001",
  11158=>"111111111",
  11159=>"000000000",
  11160=>"000111000",
  11161=>"000001011",
  11162=>"001001000",
  11163=>"000000000",
  11164=>"111111101",
  11165=>"100101111",
  11166=>"011011011",
  11167=>"100100100",
  11168=>"000001011",
  11169=>"011001101",
  11170=>"111111100",
  11171=>"000000000",
  11172=>"111101001",
  11173=>"000000000",
  11174=>"111111111",
  11175=>"111111111",
  11176=>"111110110",
  11177=>"000000000",
  11178=>"111111111",
  11179=>"111011010",
  11180=>"000000001",
  11181=>"111111111",
  11182=>"001000000",
  11183=>"000000000",
  11184=>"111000111",
  11185=>"111111000",
  11186=>"111111000",
  11187=>"000000000",
  11188=>"101100001",
  11189=>"110000000",
  11190=>"111111111",
  11191=>"000000000",
  11192=>"000100111",
  11193=>"111110110",
  11194=>"111001000",
  11195=>"011000000",
  11196=>"000000000",
  11197=>"111111110",
  11198=>"011111110",
  11199=>"100000100",
  11200=>"000000000",
  11201=>"000000000",
  11202=>"001001101",
  11203=>"000000111",
  11204=>"000000000",
  11205=>"000100100",
  11206=>"011111111",
  11207=>"000000000",
  11208=>"000000000",
  11209=>"100000000",
  11210=>"011001111",
  11211=>"000000010",
  11212=>"000000000",
  11213=>"111111110",
  11214=>"001011111",
  11215=>"100000111",
  11216=>"011110100",
  11217=>"000000000",
  11218=>"111000000",
  11219=>"000000000",
  11220=>"000010010",
  11221=>"111111111",
  11222=>"110100100",
  11223=>"100100010",
  11224=>"000000000",
  11225=>"001000000",
  11226=>"111111111",
  11227=>"001110110",
  11228=>"111111111",
  11229=>"101000000",
  11230=>"110110111",
  11231=>"100100100",
  11232=>"100100000",
  11233=>"111111111",
  11234=>"101111000",
  11235=>"111001101",
  11236=>"011111001",
  11237=>"111011011",
  11238=>"110110010",
  11239=>"000000000",
  11240=>"011011000",
  11241=>"000000001",
  11242=>"011100000",
  11243=>"000010111",
  11244=>"111100111",
  11245=>"011000000",
  11246=>"111111111",
  11247=>"000111100",
  11248=>"000000001",
  11249=>"000000000",
  11250=>"000000000",
  11251=>"011000010",
  11252=>"000000000",
  11253=>"111100000",
  11254=>"110000100",
  11255=>"010000000",
  11256=>"000000000",
  11257=>"000001000",
  11258=>"111111111",
  11259=>"111111111",
  11260=>"000111111",
  11261=>"000000000",
  11262=>"011001000",
  11263=>"111111111",
  11264=>"010100100",
  11265=>"100000111",
  11266=>"100000111",
  11267=>"101101110",
  11268=>"000001101",
  11269=>"000000111",
  11270=>"110110110",
  11271=>"011111111",
  11272=>"011011011",
  11273=>"000000000",
  11274=>"010010111",
  11275=>"000100000",
  11276=>"000001000",
  11277=>"011111111",
  11278=>"111111111",
  11279=>"000010010",
  11280=>"110010110",
  11281=>"110011111",
  11282=>"101101101",
  11283=>"100100101",
  11284=>"000000000",
  11285=>"100101111",
  11286=>"100100111",
  11287=>"110111111",
  11288=>"110110110",
  11289=>"000100001",
  11290=>"101100000",
  11291=>"110100011",
  11292=>"101001000",
  11293=>"111111111",
  11294=>"001111011",
  11295=>"110010011",
  11296=>"001000100",
  11297=>"001011011",
  11298=>"011100100",
  11299=>"101000001",
  11300=>"110110011",
  11301=>"001101101",
  11302=>"010010010",
  11303=>"000000010",
  11304=>"111000000",
  11305=>"111111111",
  11306=>"010000000",
  11307=>"000000000",
  11308=>"100101101",
  11309=>"111111111",
  11310=>"110010010",
  11311=>"100000111",
  11312=>"010110110",
  11313=>"100100111",
  11314=>"101100000",
  11315=>"000010011",
  11316=>"000100000",
  11317=>"101101100",
  11318=>"011000000",
  11319=>"111111011",
  11320=>"100100101",
  11321=>"000101101",
  11322=>"101101001",
  11323=>"000000101",
  11324=>"000000000",
  11325=>"000000110",
  11326=>"011111111",
  11327=>"000000000",
  11328=>"001100100",
  11329=>"000010000",
  11330=>"111011001",
  11331=>"010010010",
  11332=>"000000010",
  11333=>"001001000",
  11334=>"111000010",
  11335=>"111001001",
  11336=>"001001001",
  11337=>"000000100",
  11338=>"100111111",
  11339=>"111101111",
  11340=>"010000000",
  11341=>"010110111",
  11342=>"000001011",
  11343=>"100100000",
  11344=>"010011111",
  11345=>"011111111",
  11346=>"000000100",
  11347=>"000000000",
  11348=>"110010000",
  11349=>"011111111",
  11350=>"001101001",
  11351=>"000000000",
  11352=>"100000100",
  11353=>"111101101",
  11354=>"000000000",
  11355=>"100111101",
  11356=>"101101101",
  11357=>"010111111",
  11358=>"111110010",
  11359=>"000001011",
  11360=>"000000000",
  11361=>"011111111",
  11362=>"001000000",
  11363=>"101001101",
  11364=>"101100101",
  11365=>"100010110",
  11366=>"111111111",
  11367=>"101101101",
  11368=>"000000000",
  11369=>"111101110",
  11370=>"111110000",
  11371=>"110110101",
  11372=>"110010000",
  11373=>"010010000",
  11374=>"000000000",
  11375=>"000011111",
  11376=>"111111110",
  11377=>"111111000",
  11378=>"000000010",
  11379=>"100101111",
  11380=>"001000000",
  11381=>"100101100",
  11382=>"101101101",
  11383=>"000100000",
  11384=>"000000101",
  11385=>"000000101",
  11386=>"100100000",
  11387=>"001111111",
  11388=>"100111111",
  11389=>"101101101",
  11390=>"101100101",
  11391=>"000000000",
  11392=>"000000000",
  11393=>"001001000",
  11394=>"100111111",
  11395=>"000010010",
  11396=>"100101101",
  11397=>"111111010",
  11398=>"110110010",
  11399=>"111100000",
  11400=>"111000000",
  11401=>"010110010",
  11402=>"111100000",
  11403=>"011011110",
  11404=>"010110111",
  11405=>"101111101",
  11406=>"101100000",
  11407=>"011011000",
  11408=>"101101111",
  11409=>"000000000",
  11410=>"111101001",
  11411=>"111100100",
  11412=>"101111011",
  11413=>"001101101",
  11414=>"110000110",
  11415=>"101001101",
  11416=>"110111110",
  11417=>"011101101",
  11418=>"010111111",
  11419=>"011010001",
  11420=>"111010111",
  11421=>"000000101",
  11422=>"010010011",
  11423=>"010011011",
  11424=>"000011110",
  11425=>"010010010",
  11426=>"101101100",
  11427=>"111111111",
  11428=>"101001001",
  11429=>"100000011",
  11430=>"011011010",
  11431=>"000011001",
  11432=>"111111000",
  11433=>"001111111",
  11434=>"000000000",
  11435=>"111111011",
  11436=>"101101101",
  11437=>"000100000",
  11438=>"100000000",
  11439=>"011010011",
  11440=>"110111101",
  11441=>"010010010",
  11442=>"011111011",
  11443=>"111101000",
  11444=>"110000000",
  11445=>"000000010",
  11446=>"000001000",
  11447=>"000111111",
  11448=>"111101001",
  11449=>"000111010",
  11450=>"101100100",
  11451=>"011110010",
  11452=>"000000000",
  11453=>"010110000",
  11454=>"110110110",
  11455=>"001100101",
  11456=>"110110111",
  11457=>"111000001",
  11458=>"000100100",
  11459=>"010110111",
  11460=>"111000001",
  11461=>"000000000",
  11462=>"110100010",
  11463=>"000010011",
  11464=>"011011111",
  11465=>"001000111",
  11466=>"111111110",
  11467=>"001100101",
  11468=>"100100001",
  11469=>"111011001",
  11470=>"000101001",
  11471=>"001001111",
  11472=>"000000011",
  11473=>"111010011",
  11474=>"000000000",
  11475=>"000000100",
  11476=>"101101101",
  11477=>"001110101",
  11478=>"000000000",
  11479=>"111000000",
  11480=>"101101001",
  11481=>"000000001",
  11482=>"001000000",
  11483=>"000100111",
  11484=>"100000000",
  11485=>"010111011",
  11486=>"000100101",
  11487=>"000001001",
  11488=>"000000000",
  11489=>"010010110",
  11490=>"010001111",
  11491=>"000000110",
  11492=>"010010110",
  11493=>"111011111",
  11494=>"110110000",
  11495=>"111111011",
  11496=>"010010010",
  11497=>"000000000",
  11498=>"000000000",
  11499=>"100101000",
  11500=>"001001000",
  11501=>"000001101",
  11502=>"000000101",
  11503=>"110111111",
  11504=>"111011000",
  11505=>"000000111",
  11506=>"111101000",
  11507=>"101100100",
  11508=>"111111111",
  11509=>"001100100",
  11510=>"000000000",
  11511=>"000110111",
  11512=>"110111111",
  11513=>"001001100",
  11514=>"000110111",
  11515=>"001101101",
  11516=>"000000010",
  11517=>"010110110",
  11518=>"001001000",
  11519=>"111101000",
  11520=>"101101000",
  11521=>"100000100",
  11522=>"100101100",
  11523=>"111010010",
  11524=>"000000011",
  11525=>"001000000",
  11526=>"001101111",
  11527=>"010110011",
  11528=>"000000100",
  11529=>"100100100",
  11530=>"010110010",
  11531=>"010110111",
  11532=>"111011001",
  11533=>"000000011",
  11534=>"000101101",
  11535=>"011011000",
  11536=>"000010111",
  11537=>"111000101",
  11538=>"000001000",
  11539=>"111001101",
  11540=>"000001110",
  11541=>"011111111",
  11542=>"000101101",
  11543=>"111111111",
  11544=>"000000001",
  11545=>"001000101",
  11546=>"101101000",
  11547=>"011000000",
  11548=>"100110100",
  11549=>"101101101",
  11550=>"111001101",
  11551=>"010000100",
  11552=>"000110110",
  11553=>"100001001",
  11554=>"000011010",
  11555=>"010010111",
  11556=>"111111111",
  11557=>"000000000",
  11558=>"000001001",
  11559=>"011111000",
  11560=>"000000111",
  11561=>"000010011",
  11562=>"111110100",
  11563=>"000000011",
  11564=>"000000000",
  11565=>"011111011",
  11566=>"000010010",
  11567=>"000000100",
  11568=>"100110110",
  11569=>"000000000",
  11570=>"001101011",
  11571=>"000111111",
  11572=>"110000000",
  11573=>"000011111",
  11574=>"001011001",
  11575=>"010000000",
  11576=>"000001000",
  11577=>"001001001",
  11578=>"101101101",
  11579=>"100101111",
  11580=>"000000101",
  11581=>"000000000",
  11582=>"011001001",
  11583=>"001001000",
  11584=>"111100111",
  11585=>"111111111",
  11586=>"000000000",
  11587=>"001001000",
  11588=>"111110010",
  11589=>"010111001",
  11590=>"110000111",
  11591=>"000000100",
  11592=>"000101101",
  11593=>"010010010",
  11594=>"110110110",
  11595=>"110111111",
  11596=>"010000011",
  11597=>"010110110",
  11598=>"110011011",
  11599=>"011111101",
  11600=>"011001001",
  11601=>"000000011",
  11602=>"111101111",
  11603=>"000110111",
  11604=>"101101101",
  11605=>"011011011",
  11606=>"101001111",
  11607=>"001001001",
  11608=>"110000000",
  11609=>"100100000",
  11610=>"111010000",
  11611=>"101100101",
  11612=>"001000000",
  11613=>"011000000",
  11614=>"001001100",
  11615=>"100001110",
  11616=>"110111101",
  11617=>"001001001",
  11618=>"101111111",
  11619=>"000111111",
  11620=>"000000011",
  11621=>"000001101",
  11622=>"111111010",
  11623=>"111110111",
  11624=>"011111101",
  11625=>"111111011",
  11626=>"111111111",
  11627=>"000000110",
  11628=>"010110111",
  11629=>"101100100",
  11630=>"010010110",
  11631=>"000000000",
  11632=>"000101111",
  11633=>"111111111",
  11634=>"000000000",
  11635=>"111011011",
  11636=>"000000000",
  11637=>"111111111",
  11638=>"111000001",
  11639=>"010010000",
  11640=>"111111111",
  11641=>"111111111",
  11642=>"101001001",
  11643=>"000000000",
  11644=>"101001001",
  11645=>"001000000",
  11646=>"110111111",
  11647=>"011011011",
  11648=>"110100110",
  11649=>"000000000",
  11650=>"000001001",
  11651=>"110110111",
  11652=>"000000000",
  11653=>"010111000",
  11654=>"111111000",
  11655=>"110111111",
  11656=>"111011001",
  11657=>"100111111",
  11658=>"000000100",
  11659=>"111110000",
  11660=>"100110111",
  11661=>"001001111",
  11662=>"010010010",
  11663=>"010010010",
  11664=>"000011011",
  11665=>"000000000",
  11666=>"110111011",
  11667=>"001000101",
  11668=>"111000010",
  11669=>"000000000",
  11670=>"101001111",
  11671=>"000001011",
  11672=>"000000101",
  11673=>"011011110",
  11674=>"010111111",
  11675=>"111110000",
  11676=>"111111010",
  11677=>"100100000",
  11678=>"101101101",
  11679=>"000000000",
  11680=>"000000000",
  11681=>"100101111",
  11682=>"000000000",
  11683=>"111101100",
  11684=>"011000000",
  11685=>"100100101",
  11686=>"000000000",
  11687=>"111111111",
  11688=>"100000000",
  11689=>"010111111",
  11690=>"111101101",
  11691=>"011111110",
  11692=>"000000101",
  11693=>"000000011",
  11694=>"000111111",
  11695=>"000010000",
  11696=>"111111010",
  11697=>"101101001",
  11698=>"100101001",
  11699=>"110110110",
  11700=>"000001101",
  11701=>"001001101",
  11702=>"101001111",
  11703=>"000001101",
  11704=>"000000000",
  11705=>"101010011",
  11706=>"100001111",
  11707=>"110001000",
  11708=>"000011111",
  11709=>"001000000",
  11710=>"001001111",
  11711=>"000000001",
  11712=>"110010000",
  11713=>"000000000",
  11714=>"001101000",
  11715=>"000011111",
  11716=>"000001101",
  11717=>"001101001",
  11718=>"110110100",
  11719=>"101101011",
  11720=>"111111100",
  11721=>"000000000",
  11722=>"000100100",
  11723=>"011011010",
  11724=>"110110010",
  11725=>"000010000",
  11726=>"000000000",
  11727=>"111111111",
  11728=>"000001011",
  11729=>"011000110",
  11730=>"010000000",
  11731=>"111011011",
  11732=>"000010000",
  11733=>"000000000",
  11734=>"000010010",
  11735=>"101001011",
  11736=>"001001000",
  11737=>"010010010",
  11738=>"101000011",
  11739=>"010011111",
  11740=>"110000000",
  11741=>"111010000",
  11742=>"010010010",
  11743=>"000000001",
  11744=>"101111010",
  11745=>"110010010",
  11746=>"001001000",
  11747=>"010110010",
  11748=>"111000001",
  11749=>"001100110",
  11750=>"001001111",
  11751=>"000000110",
  11752=>"000100000",
  11753=>"011011111",
  11754=>"111011011",
  11755=>"110110010",
  11756=>"011010010",
  11757=>"100000000",
  11758=>"000000001",
  11759=>"100000000",
  11760=>"101101101",
  11761=>"111111101",
  11762=>"101011011",
  11763=>"011111111",
  11764=>"100000101",
  11765=>"000000000",
  11766=>"101111111",
  11767=>"001001001",
  11768=>"001001001",
  11769=>"001001001",
  11770=>"000000100",
  11771=>"011111010",
  11772=>"111111111",
  11773=>"110110110",
  11774=>"000000000",
  11775=>"101101101",
  11776=>"000000111",
  11777=>"111111111",
  11778=>"111111111",
  11779=>"111000000",
  11780=>"000000001",
  11781=>"111000111",
  11782=>"111111111",
  11783=>"111111111",
  11784=>"000000000",
  11785=>"001001001",
  11786=>"000000000",
  11787=>"110111110",
  11788=>"111011011",
  11789=>"011011011",
  11790=>"000000000",
  11791=>"110111111",
  11792=>"011111111",
  11793=>"111001000",
  11794=>"011000000",
  11795=>"110110111",
  11796=>"100110111",
  11797=>"110010000",
  11798=>"010000000",
  11799=>"100110111",
  11800=>"111111110",
  11801=>"010000000",
  11802=>"110100101",
  11803=>"011000111",
  11804=>"111000001",
  11805=>"111111101",
  11806=>"011111010",
  11807=>"111111111",
  11808=>"000000000",
  11809=>"110111111",
  11810=>"000000000",
  11811=>"101111111",
  11812=>"111111111",
  11813=>"111101000",
  11814=>"000000000",
  11815=>"111110111",
  11816=>"000000000",
  11817=>"000000000",
  11818=>"000000000",
  11819=>"010111011",
  11820=>"111111111",
  11821=>"111000100",
  11822=>"101000000",
  11823=>"111010111",
  11824=>"000010000",
  11825=>"111111111",
  11826=>"000000000",
  11827=>"000000000",
  11828=>"001011100",
  11829=>"001111011",
  11830=>"000000000",
  11831=>"010010000",
  11832=>"100000000",
  11833=>"000011000",
  11834=>"101000100",
  11835=>"111111100",
  11836=>"000000000",
  11837=>"101001111",
  11838=>"101011111",
  11839=>"000000000",
  11840=>"111110111",
  11841=>"000000000",
  11842=>"000100100",
  11843=>"111111111",
  11844=>"001011111",
  11845=>"001001000",
  11846=>"111111111",
  11847=>"111111111",
  11848=>"110100100",
  11849=>"000000101",
  11850=>"111111111",
  11851=>"000000001",
  11852=>"111111100",
  11853=>"111111101",
  11854=>"111100100",
  11855=>"101000001",
  11856=>"000000000",
  11857=>"111111001",
  11858=>"111011001",
  11859=>"011011000",
  11860=>"111111101",
  11861=>"000000000",
  11862=>"111111111",
  11863=>"101110111",
  11864=>"011011111",
  11865=>"000000000",
  11866=>"111111000",
  11867=>"000000100",
  11868=>"011111111",
  11869=>"000011111",
  11870=>"111001000",
  11871=>"000000100",
  11872=>"111111111",
  11873=>"000011111",
  11874=>"000000000",
  11875=>"000000000",
  11876=>"000000000",
  11877=>"000000100",
  11878=>"000000000",
  11879=>"110110111",
  11880=>"000000000",
  11881=>"100100110",
  11882=>"111111111",
  11883=>"111111100",
  11884=>"111111000",
  11885=>"111110111",
  11886=>"111111111",
  11887=>"110111111",
  11888=>"111011111",
  11889=>"011111001",
  11890=>"000110110",
  11891=>"111111000",
  11892=>"000001010",
  11893=>"110111110",
  11894=>"000000000",
  11895=>"111111111",
  11896=>"011000000",
  11897=>"111101111",
  11898=>"111011000",
  11899=>"111011011",
  11900=>"100100100",
  11901=>"100111000",
  11902=>"111111001",
  11903=>"011000000",
  11904=>"111111111",
  11905=>"000111000",
  11906=>"000110111",
  11907=>"111110110",
  11908=>"111111111",
  11909=>"000000111",
  11910=>"110100110",
  11911=>"111111010",
  11912=>"111001000",
  11913=>"000000000",
  11914=>"001000000",
  11915=>"111111111",
  11916=>"001111111",
  11917=>"111010000",
  11918=>"111111111",
  11919=>"110111000",
  11920=>"111111111",
  11921=>"111000000",
  11922=>"000000000",
  11923=>"111111111",
  11924=>"000000001",
  11925=>"100100100",
  11926=>"111111111",
  11927=>"111000000",
  11928=>"111001001",
  11929=>"111111111",
  11930=>"100110111",
  11931=>"111111100",
  11932=>"000000111",
  11933=>"000000000",
  11934=>"111111000",
  11935=>"100000000",
  11936=>"000000100",
  11937=>"111100000",
  11938=>"000000000",
  11939=>"100100100",
  11940=>"111111001",
  11941=>"111100100",
  11942=>"111111111",
  11943=>"011111000",
  11944=>"111111011",
  11945=>"000000000",
  11946=>"100100000",
  11947=>"000001001",
  11948=>"000000101",
  11949=>"111100110",
  11950=>"000000000",
  11951=>"000000111",
  11952=>"000111000",
  11953=>"111000000",
  11954=>"111111010",
  11955=>"000000100",
  11956=>"111111011",
  11957=>"111011000",
  11958=>"000101100",
  11959=>"111111111",
  11960=>"100100000",
  11961=>"000000000",
  11962=>"111000000",
  11963=>"110000000",
  11964=>"111111111",
  11965=>"000000000",
  11966=>"111111111",
  11967=>"110111111",
  11968=>"111111111",
  11969=>"110100111",
  11970=>"001000100",
  11971=>"000000000",
  11972=>"000000000",
  11973=>"011011011",
  11974=>"000000000",
  11975=>"111110111",
  11976=>"001001000",
  11977=>"000000001",
  11978=>"100100101",
  11979=>"111111111",
  11980=>"111111000",
  11981=>"000000110",
  11982=>"110111111",
  11983=>"010000000",
  11984=>"111010010",
  11985=>"000110111",
  11986=>"111000000",
  11987=>"000100000",
  11988=>"000000000",
  11989=>"000000000",
  11990=>"000010011",
  11991=>"000000000",
  11992=>"111111111",
  11993=>"000010111",
  11994=>"000000001",
  11995=>"010000000",
  11996=>"000000111",
  11997=>"000000000",
  11998=>"000000000",
  11999=>"010000011",
  12000=>"001101000",
  12001=>"000000000",
  12002=>"001011110",
  12003=>"111011011",
  12004=>"110000100",
  12005=>"100001001",
  12006=>"111111111",
  12007=>"111000000",
  12008=>"111111111",
  12009=>"000000001",
  12010=>"100100001",
  12011=>"110110111",
  12012=>"111111111",
  12013=>"000000000",
  12014=>"000000110",
  12015=>"000000000",
  12016=>"010111000",
  12017=>"100100000",
  12018=>"111111111",
  12019=>"000000000",
  12020=>"111001001",
  12021=>"001001001",
  12022=>"001111111",
  12023=>"110110010",
  12024=>"111111111",
  12025=>"000000000",
  12026=>"111111000",
  12027=>"001111111",
  12028=>"110111111",
  12029=>"001111111",
  12030=>"000000011",
  12031=>"110111111",
  12032=>"000000011",
  12033=>"000000000",
  12034=>"111111111",
  12035=>"011111111",
  12036=>"000000001",
  12037=>"000000001",
  12038=>"000100111",
  12039=>"000000000",
  12040=>"000101111",
  12041=>"001001000",
  12042=>"000001001",
  12043=>"111111111",
  12044=>"111101111",
  12045=>"000000000",
  12046=>"111111001",
  12047=>"000000000",
  12048=>"000000001",
  12049=>"001101111",
  12050=>"000000100",
  12051=>"111000000",
  12052=>"110110111",
  12053=>"111111011",
  12054=>"001011111",
  12055=>"001000000",
  12056=>"001001100",
  12057=>"001001000",
  12058=>"000010111",
  12059=>"111111111",
  12060=>"000000010",
  12061=>"010011011",
  12062=>"000000000",
  12063=>"001000111",
  12064=>"000000100",
  12065=>"111111111",
  12066=>"000000000",
  12067=>"000000100",
  12068=>"111111111",
  12069=>"000000100",
  12070=>"111111110",
  12071=>"110100000",
  12072=>"000000000",
  12073=>"100000000",
  12074=>"000000000",
  12075=>"000000000",
  12076=>"111111001",
  12077=>"111111111",
  12078=>"111101110",
  12079=>"000000000",
  12080=>"111011011",
  12081=>"000000110",
  12082=>"111111110",
  12083=>"111111111",
  12084=>"111001000",
  12085=>"111111111",
  12086=>"000000000",
  12087=>"111001100",
  12088=>"111111000",
  12089=>"111111100",
  12090=>"110000111",
  12091=>"100000000",
  12092=>"001000000",
  12093=>"000000000",
  12094=>"111011111",
  12095=>"000010010",
  12096=>"000000000",
  12097=>"000000000",
  12098=>"111111111",
  12099=>"110100111",
  12100=>"000000100",
  12101=>"001001001",
  12102=>"110000011",
  12103=>"111111111",
  12104=>"111011000",
  12105=>"000111111",
  12106=>"000100110",
  12107=>"111111111",
  12108=>"000000000",
  12109=>"011111111",
  12110=>"000001111",
  12111=>"000010111",
  12112=>"111111111",
  12113=>"000000100",
  12114=>"001100111",
  12115=>"000111111",
  12116=>"000000000",
  12117=>"011011011",
  12118=>"000000000",
  12119=>"011111000",
  12120=>"000000000",
  12121=>"100100111",
  12122=>"011011001",
  12123=>"111001101",
  12124=>"111111111",
  12125=>"111111101",
  12126=>"001000001",
  12127=>"100010000",
  12128=>"111111110",
  12129=>"111111111",
  12130=>"111111111",
  12131=>"111000111",
  12132=>"000001000",
  12133=>"000000000",
  12134=>"000000111",
  12135=>"000000000",
  12136=>"111111111",
  12137=>"000000000",
  12138=>"011111011",
  12139=>"110010111",
  12140=>"000000000",
  12141=>"111100000",
  12142=>"000100100",
  12143=>"001000000",
  12144=>"100100110",
  12145=>"111111000",
  12146=>"000000111",
  12147=>"111111000",
  12148=>"000000000",
  12149=>"000100000",
  12150=>"100000000",
  12151=>"011011111",
  12152=>"000000000",
  12153=>"111111000",
  12154=>"000000000",
  12155=>"111000011",
  12156=>"111110000",
  12157=>"110111111",
  12158=>"000000000",
  12159=>"000000101",
  12160=>"000000000",
  12161=>"000000101",
  12162=>"000000000",
  12163=>"100101111",
  12164=>"000000001",
  12165=>"100100110",
  12166=>"000000101",
  12167=>"000000000",
  12168=>"000000000",
  12169=>"001000000",
  12170=>"001000011",
  12171=>"000000000",
  12172=>"001111111",
  12173=>"001000000",
  12174=>"000000000",
  12175=>"110111111",
  12176=>"000000000",
  12177=>"000000000",
  12178=>"110110000",
  12179=>"100100000",
  12180=>"111111100",
  12181=>"000000000",
  12182=>"111101001",
  12183=>"001001000",
  12184=>"111111111",
  12185=>"000001001",
  12186=>"111111111",
  12187=>"000000000",
  12188=>"111111111",
  12189=>"110010111",
  12190=>"111001011",
  12191=>"111110110",
  12192=>"111011000",
  12193=>"001011010",
  12194=>"111101111",
  12195=>"111101000",
  12196=>"011111111",
  12197=>"000000111",
  12198=>"000000011",
  12199=>"000110011",
  12200=>"001000100",
  12201=>"000000000",
  12202=>"001001111",
  12203=>"000000000",
  12204=>"011001001",
  12205=>"011111111",
  12206=>"111111111",
  12207=>"110111110",
  12208=>"111100000",
  12209=>"101000000",
  12210=>"111111111",
  12211=>"000000000",
  12212=>"111111111",
  12213=>"000100100",
  12214=>"000111111",
  12215=>"000000000",
  12216=>"000000100",
  12217=>"111111111",
  12218=>"111111111",
  12219=>"111111000",
  12220=>"000000000",
  12221=>"110110110",
  12222=>"111111111",
  12223=>"111111111",
  12224=>"011000111",
  12225=>"000000111",
  12226=>"011111111",
  12227=>"000100101",
  12228=>"111111111",
  12229=>"111011011",
  12230=>"111111111",
  12231=>"111111111",
  12232=>"111100000",
  12233=>"000000011",
  12234=>"000000000",
  12235=>"111111111",
  12236=>"000000000",
  12237=>"111111111",
  12238=>"000000000",
  12239=>"101011111",
  12240=>"111111111",
  12241=>"001000000",
  12242=>"111111111",
  12243=>"101000111",
  12244=>"111111111",
  12245=>"001011100",
  12246=>"000000000",
  12247=>"100110010",
  12248=>"101101111",
  12249=>"111111111",
  12250=>"000000111",
  12251=>"101001111",
  12252=>"111100100",
  12253=>"011001111",
  12254=>"010000000",
  12255=>"011011000",
  12256=>"111111111",
  12257=>"000000000",
  12258=>"000000000",
  12259=>"111111111",
  12260=>"111110011",
  12261=>"000000000",
  12262=>"000000000",
  12263=>"000000000",
  12264=>"111100000",
  12265=>"111111000",
  12266=>"000000000",
  12267=>"000011011",
  12268=>"000100111",
  12269=>"001000001",
  12270=>"111000000",
  12271=>"111111111",
  12272=>"001000001",
  12273=>"000000100",
  12274=>"000110111",
  12275=>"111111111",
  12276=>"111111001",
  12277=>"000000000",
  12278=>"011010000",
  12279=>"110110110",
  12280=>"000000000",
  12281=>"001001000",
  12282=>"000000000",
  12283=>"110110111",
  12284=>"010011010",
  12285=>"000000000",
  12286=>"000000000",
  12287=>"101111001",
  12288=>"000000000",
  12289=>"111001000",
  12290=>"000001111",
  12291=>"000000101",
  12292=>"000000111",
  12293=>"100000000",
  12294=>"111000000",
  12295=>"000000000",
  12296=>"000000111",
  12297=>"000000000",
  12298=>"000000100",
  12299=>"011011001",
  12300=>"111111000",
  12301=>"000000111",
  12302=>"011000000",
  12303=>"000000001",
  12304=>"000000000",
  12305=>"000001000",
  12306=>"111111100",
  12307=>"111111010",
  12308=>"111111110",
  12309=>"000000111",
  12310=>"110111111",
  12311=>"000000000",
  12312=>"011011011",
  12313=>"011100100",
  12314=>"000000110",
  12315=>"011000111",
  12316=>"110111111",
  12317=>"000000001",
  12318=>"110011011",
  12319=>"000001000",
  12320=>"000000000",
  12321=>"111110110",
  12322=>"011100000",
  12323=>"111111100",
  12324=>"111111111",
  12325=>"011011111",
  12326=>"000000000",
  12327=>"000000111",
  12328=>"101111111",
  12329=>"101100100",
  12330=>"000110111",
  12331=>"000000110",
  12332=>"000100111",
  12333=>"000000000",
  12334=>"111111000",
  12335=>"001011000",
  12336=>"000001001",
  12337=>"000011000",
  12338=>"000010000",
  12339=>"000000011",
  12340=>"000000000",
  12341=>"000010000",
  12342=>"000100111",
  12343=>"000111001",
  12344=>"110000111",
  12345=>"111111100",
  12346=>"001000111",
  12347=>"111111111",
  12348=>"001111111",
  12349=>"100100110",
  12350=>"001001011",
  12351=>"110000000",
  12352=>"111111111",
  12353=>"000010010",
  12354=>"001010011",
  12355=>"011111111",
  12356=>"011001000",
  12357=>"011001111",
  12358=>"111110001",
  12359=>"111111000",
  12360=>"110111110",
  12361=>"000000001",
  12362=>"111111101",
  12363=>"011000111",
  12364=>"000111111",
  12365=>"000000111",
  12366=>"111001101",
  12367=>"111111000",
  12368=>"000000100",
  12369=>"000000111",
  12370=>"000111111",
  12371=>"000100100",
  12372=>"000000000",
  12373=>"001111111",
  12374=>"110110010",
  12375=>"000111111",
  12376=>"000101111",
  12377=>"101000000",
  12378=>"110000000",
  12379=>"111100110",
  12380=>"111111010",
  12381=>"000000000",
  12382=>"000000110",
  12383=>"111001000",
  12384=>"001001001",
  12385=>"011001000",
  12386=>"001000000",
  12387=>"000000000",
  12388=>"111111111",
  12389=>"011111111",
  12390=>"000000000",
  12391=>"001000001",
  12392=>"111111111",
  12393=>"111000000",
  12394=>"111111111",
  12395=>"111111010",
  12396=>"000000010",
  12397=>"111111111",
  12398=>"111111111",
  12399=>"100000100",
  12400=>"000111110",
  12401=>"000110011",
  12402=>"001000100",
  12403=>"111000001",
  12404=>"111111100",
  12405=>"001001101",
  12406=>"000000000",
  12407=>"111000000",
  12408=>"000000000",
  12409=>"000011001",
  12410=>"000000000",
  12411=>"000000000",
  12412=>"000000000",
  12413=>"000001101",
  12414=>"000000000",
  12415=>"111110111",
  12416=>"101111111",
  12417=>"111110000",
  12418=>"111001000",
  12419=>"100110100",
  12420=>"000000001",
  12421=>"000000001",
  12422=>"100000000",
  12423=>"111111100",
  12424=>"111101100",
  12425=>"001001111",
  12426=>"000000010",
  12427=>"101101100",
  12428=>"110011000",
  12429=>"111110000",
  12430=>"000000010",
  12431=>"111011000",
  12432=>"000100111",
  12433=>"000000111",
  12434=>"000100100",
  12435=>"000011111",
  12436=>"000000110",
  12437=>"111111000",
  12438=>"111111000",
  12439=>"111011000",
  12440=>"101000101",
  12441=>"101111001",
  12442=>"111111111",
  12443=>"000000011",
  12444=>"111111111",
  12445=>"111111111",
  12446=>"111111111",
  12447=>"111111001",
  12448=>"100111110",
  12449=>"011001000",
  12450=>"011011111",
  12451=>"000000001",
  12452=>"001111111",
  12453=>"111111111",
  12454=>"000000000",
  12455=>"000011011",
  12456=>"000000010",
  12457=>"000001001",
  12458=>"000000000",
  12459=>"000001111",
  12460=>"111111111",
  12461=>"000000000",
  12462=>"111111111",
  12463=>"011001000",
  12464=>"111100000",
  12465=>"110110001",
  12466=>"000100010",
  12467=>"000000000",
  12468=>"100111111",
  12469=>"100100110",
  12470=>"101111111",
  12471=>"000111111",
  12472=>"001111111",
  12473=>"111111100",
  12474=>"000111010",
  12475=>"000000000",
  12476=>"111000000",
  12477=>"100100111",
  12478=>"001111000",
  12479=>"011111010",
  12480=>"000000000",
  12481=>"101001001",
  12482=>"000001011",
  12483=>"000000000",
  12484=>"011011111",
  12485=>"000000000",
  12486=>"000000001",
  12487=>"111000000",
  12488=>"111101111",
  12489=>"111110110",
  12490=>"000000000",
  12491=>"101100001",
  12492=>"111011011",
  12493=>"111110110",
  12494=>"111001001",
  12495=>"111000000",
  12496=>"011001111",
  12497=>"111001000",
  12498=>"111111111",
  12499=>"001001011",
  12500=>"011011111",
  12501=>"101111000",
  12502=>"111111001",
  12503=>"000001111",
  12504=>"000000000",
  12505=>"000000001",
  12506=>"111111111",
  12507=>"000000000",
  12508=>"001001111",
  12509=>"111111111",
  12510=>"000000110",
  12511=>"101100111",
  12512=>"100000000",
  12513=>"000110000",
  12514=>"110111111",
  12515=>"111111111",
  12516=>"000110000",
  12517=>"011011111",
  12518=>"111110100",
  12519=>"111111000",
  12520=>"111111000",
  12521=>"111110111",
  12522=>"001000000",
  12523=>"111001011",
  12524=>"111111000",
  12525=>"000000000",
  12526=>"110111111",
  12527=>"000000110",
  12528=>"010000000",
  12529=>"111111111",
  12530=>"100100110",
  12531=>"111111110",
  12532=>"101001111",
  12533=>"000000000",
  12534=>"010010100",
  12535=>"011000000",
  12536=>"000000000",
  12537=>"000111111",
  12538=>"000000111",
  12539=>"000001001",
  12540=>"111111111",
  12541=>"001011011",
  12542=>"111111000",
  12543=>"111111000",
  12544=>"111100000",
  12545=>"000100100",
  12546=>"001001000",
  12547=>"000111110",
  12548=>"111110100",
  12549=>"111111111",
  12550=>"111101111",
  12551=>"001111111",
  12552=>"000000111",
  12553=>"001000000",
  12554=>"111011111",
  12555=>"111111001",
  12556=>"100000000",
  12557=>"000000100",
  12558=>"000000001",
  12559=>"000000110",
  12560=>"000000000",
  12561=>"000000111",
  12562=>"000000111",
  12563=>"000001111",
  12564=>"100111111",
  12565=>"111110000",
  12566=>"001001111",
  12567=>"000000000",
  12568=>"010000000",
  12569=>"010111111",
  12570=>"111111111",
  12571=>"111001000",
  12572=>"000111111",
  12573=>"000001111",
  12574=>"000000000",
  12575=>"111111111",
  12576=>"000010110",
  12577=>"001111011",
  12578=>"111011011",
  12579=>"111100111",
  12580=>"011001001",
  12581=>"000000101",
  12582=>"111100111",
  12583=>"111111110",
  12584=>"000100100",
  12585=>"111100000",
  12586=>"000111100",
  12587=>"000000000",
  12588=>"000000010",
  12589=>"000111011",
  12590=>"000000000",
  12591=>"100100111",
  12592=>"000101011",
  12593=>"111101000",
  12594=>"111111111",
  12595=>"000111111",
  12596=>"000000000",
  12597=>"001000000",
  12598=>"000000000",
  12599=>"111000000",
  12600=>"111000000",
  12601=>"111000101",
  12602=>"101000000",
  12603=>"001011111",
  12604=>"111111110",
  12605=>"000000111",
  12606=>"001101100",
  12607=>"000000000",
  12608=>"000110111",
  12609=>"000111001",
  12610=>"111111110",
  12611=>"000000001",
  12612=>"000000000",
  12613=>"000000111",
  12614=>"111111111",
  12615=>"111111111",
  12616=>"000000000",
  12617=>"111011111",
  12618=>"001101111",
  12619=>"111100001",
  12620=>"111001101",
  12621=>"000000111",
  12622=>"111000110",
  12623=>"000000011",
  12624=>"111000000",
  12625=>"001111111",
  12626=>"000000111",
  12627=>"111111000",
  12628=>"111100100",
  12629=>"011011001",
  12630=>"111111111",
  12631=>"000011111",
  12632=>"001000111",
  12633=>"001000000",
  12634=>"110110000",
  12635=>"111111111",
  12636=>"111001001",
  12637=>"000001100",
  12638=>"111000101",
  12639=>"111000000",
  12640=>"111010000",
  12641=>"000001011",
  12642=>"000000100",
  12643=>"111111010",
  12644=>"011011111",
  12645=>"000000000",
  12646=>"111111000",
  12647=>"111111110",
  12648=>"001000000",
  12649=>"011111111",
  12650=>"011101000",
  12651=>"011011110",
  12652=>"000000000",
  12653=>"000000000",
  12654=>"011000000",
  12655=>"000110111",
  12656=>"101000001",
  12657=>"001111000",
  12658=>"000000001",
  12659=>"000111001",
  12660=>"000000000",
  12661=>"001000000",
  12662=>"111011000",
  12663=>"011110100",
  12664=>"111111111",
  12665=>"000000111",
  12666=>"100000001",
  12667=>"000000000",
  12668=>"011011011",
  12669=>"001110111",
  12670=>"000100000",
  12671=>"000111111",
  12672=>"011111111",
  12673=>"011111110",
  12674=>"111011101",
  12675=>"000000011",
  12676=>"110000000",
  12677=>"011111011",
  12678=>"001000011",
  12679=>"001000000",
  12680=>"111001001",
  12681=>"110110000",
  12682=>"000000000",
  12683=>"000000000",
  12684=>"111111111",
  12685=>"001011000",
  12686=>"000000000",
  12687=>"000111111",
  12688=>"000000000",
  12689=>"111111110",
  12690=>"001001000",
  12691=>"100111111",
  12692=>"010001111",
  12693=>"000000000",
  12694=>"100110100",
  12695=>"011110100",
  12696=>"000000000",
  12697=>"111100000",
  12698=>"111111111",
  12699=>"000000110",
  12700=>"000000000",
  12701=>"000000100",
  12702=>"001111110",
  12703=>"000100000",
  12704=>"111000000",
  12705=>"111000111",
  12706=>"000010000",
  12707=>"111000000",
  12708=>"000111100",
  12709=>"100101001",
  12710=>"000000111",
  12711=>"111111111",
  12712=>"000000000",
  12713=>"000000000",
  12714=>"000000110",
  12715=>"000000110",
  12716=>"111111000",
  12717=>"111000100",
  12718=>"111000010",
  12719=>"000010011",
  12720=>"111111011",
  12721=>"111000110",
  12722=>"011001111",
  12723=>"000000000",
  12724=>"000000111",
  12725=>"000000000",
  12726=>"000001011",
  12727=>"111110111",
  12728=>"100100111",
  12729=>"111110000",
  12730=>"111111111",
  12731=>"001001011",
  12732=>"000011111",
  12733=>"111000000",
  12734=>"000000000",
  12735=>"001100100",
  12736=>"110111011",
  12737=>"111000110",
  12738=>"000000000",
  12739=>"111111000",
  12740=>"111111000",
  12741=>"000000010",
  12742=>"000000000",
  12743=>"110000000",
  12744=>"111100000",
  12745=>"000000000",
  12746=>"111111000",
  12747=>"111111111",
  12748=>"000100100",
  12749=>"000000000",
  12750=>"000000111",
  12751=>"000000000",
  12752=>"111101111",
  12753=>"000000111",
  12754=>"011000000",
  12755=>"000111110",
  12756=>"001000001",
  12757=>"111000000",
  12758=>"010111010",
  12759=>"110110100",
  12760=>"100000100",
  12761=>"111111110",
  12762=>"111010110",
  12763=>"110000000",
  12764=>"000000111",
  12765=>"101101111",
  12766=>"000011110",
  12767=>"111111110",
  12768=>"111111000",
  12769=>"101100000",
  12770=>"000100110",
  12771=>"001001000",
  12772=>"111111010",
  12773=>"001111101",
  12774=>"000000111",
  12775=>"011000000",
  12776=>"000001101",
  12777=>"111000000",
  12778=>"111110000",
  12779=>"111111100",
  12780=>"001000110",
  12781=>"000110011",
  12782=>"111111111",
  12783=>"111111100",
  12784=>"001111111",
  12785=>"000001111",
  12786=>"111101000",
  12787=>"111001000",
  12788=>"111111000",
  12789=>"000000000",
  12790=>"000000100",
  12791=>"010010010",
  12792=>"000010000",
  12793=>"100110111",
  12794=>"001000000",
  12795=>"110000000",
  12796=>"111111111",
  12797=>"111011110",
  12798=>"000000000",
  12799=>"000000000",
  12800=>"010000000",
  12801=>"000000000",
  12802=>"111111111",
  12803=>"000000000",
  12804=>"000100111",
  12805=>"111111111",
  12806=>"011000000",
  12807=>"000000101",
  12808=>"000000000",
  12809=>"000111011",
  12810=>"101000000",
  12811=>"101111111",
  12812=>"111100111",
  12813=>"000000110",
  12814=>"010000000",
  12815=>"000111111",
  12816=>"101000001",
  12817=>"000000110",
  12818=>"001001000",
  12819=>"111101001",
  12820=>"000000101",
  12821=>"111111111",
  12822=>"000000000",
  12823=>"111111111",
  12824=>"111111100",
  12825=>"011011000",
  12826=>"101111111",
  12827=>"101011011",
  12828=>"000111111",
  12829=>"111110000",
  12830=>"000110111",
  12831=>"000000000",
  12832=>"000100100",
  12833=>"110100110",
  12834=>"000000110",
  12835=>"000000000",
  12836=>"111111111",
  12837=>"111111111",
  12838=>"111111000",
  12839=>"111111100",
  12840=>"111111011",
  12841=>"010010111",
  12842=>"000001111",
  12843=>"111111111",
  12844=>"111111111",
  12845=>"000101000",
  12846=>"001111111",
  12847=>"111111101",
  12848=>"000000101",
  12849=>"111111000",
  12850=>"011110000",
  12851=>"011011000",
  12852=>"000000000",
  12853=>"111111111",
  12854=>"111111111",
  12855=>"111111111",
  12856=>"000000000",
  12857=>"011000111",
  12858=>"101100100",
  12859=>"111111111",
  12860=>"000000000",
  12861=>"100010011",
  12862=>"100111111",
  12863=>"101100110",
  12864=>"110010111",
  12865=>"010000011",
  12866=>"010011000",
  12867=>"000000111",
  12868=>"000101111",
  12869=>"001111111",
  12870=>"000000100",
  12871=>"100100100",
  12872=>"001011011",
  12873=>"111111111",
  12874=>"000000111",
  12875=>"000000111",
  12876=>"010011111",
  12877=>"011000000",
  12878=>"001011011",
  12879=>"000000000",
  12880=>"100011000",
  12881=>"101111111",
  12882=>"111110000",
  12883=>"000110000",
  12884=>"111011111",
  12885=>"111000000",
  12886=>"000000000",
  12887=>"111111111",
  12888=>"111111111",
  12889=>"111000000",
  12890=>"000000011",
  12891=>"110111111",
  12892=>"000000000",
  12893=>"000000100",
  12894=>"000000000",
  12895=>"111111111",
  12896=>"000000000",
  12897=>"111100100",
  12898=>"100110110",
  12899=>"000000000",
  12900=>"010010110",
  12901=>"000000111",
  12902=>"000000000",
  12903=>"100100111",
  12904=>"111111111",
  12905=>"000000000",
  12906=>"111111111",
  12907=>"111111111",
  12908=>"100110100",
  12909=>"000000000",
  12910=>"111000000",
  12911=>"111111111",
  12912=>"000010010",
  12913=>"111111111",
  12914=>"011011011",
  12915=>"010010000",
  12916=>"000000000",
  12917=>"000000111",
  12918=>"111111111",
  12919=>"001110110",
  12920=>"111111111",
  12921=>"000000000",
  12922=>"000000000",
  12923=>"111111111",
  12924=>"111111110",
  12925=>"111111111",
  12926=>"011011000",
  12927=>"111011000",
  12928=>"000000100",
  12929=>"101000000",
  12930=>"000100000",
  12931=>"000001001",
  12932=>"001101111",
  12933=>"000000000",
  12934=>"000000100",
  12935=>"000000000",
  12936=>"000000000",
  12937=>"000001000",
  12938=>"000000000",
  12939=>"011111111",
  12940=>"101000111",
  12941=>"111111011",
  12942=>"000000001",
  12943=>"001000000",
  12944=>"000000000",
  12945=>"111111111",
  12946=>"100111111",
  12947=>"000000110",
  12948=>"000000000",
  12949=>"000000100",
  12950=>"001111111",
  12951=>"000000000",
  12952=>"100100000",
  12953=>"100000000",
  12954=>"000100000",
  12955=>"111001000",
  12956=>"000000101",
  12957=>"001000010",
  12958=>"111011011",
  12959=>"000111100",
  12960=>"111111111",
  12961=>"111110000",
  12962=>"011000110",
  12963=>"111111111",
  12964=>"000000000",
  12965=>"111111111",
  12966=>"111111000",
  12967=>"100110111",
  12968=>"111111011",
  12969=>"001001000",
  12970=>"111111110",
  12971=>"111011111",
  12972=>"000000101",
  12973=>"110110110",
  12974=>"001000100",
  12975=>"000000000",
  12976=>"111111111",
  12977=>"011000111",
  12978=>"111111111",
  12979=>"000000000",
  12980=>"100100001",
  12981=>"100111001",
  12982=>"001000000",
  12983=>"000110111",
  12984=>"001000100",
  12985=>"111111111",
  12986=>"000000100",
  12987=>"011000000",
  12988=>"100000100",
  12989=>"000110000",
  12990=>"000110110",
  12991=>"001001000",
  12992=>"100100101",
  12993=>"000000110",
  12994=>"001011011",
  12995=>"111111000",
  12996=>"000000000",
  12997=>"000000000",
  12998=>"000000111",
  12999=>"000000001",
  13000=>"110110110",
  13001=>"110100110",
  13002=>"111111101",
  13003=>"111110100",
  13004=>"111100111",
  13005=>"011111111",
  13006=>"111111111",
  13007=>"011011101",
  13008=>"011000000",
  13009=>"000000000",
  13010=>"000000100",
  13011=>"000000000",
  13012=>"000000000",
  13013=>"111111000",
  13014=>"010111111",
  13015=>"111110110",
  13016=>"011001111",
  13017=>"000110100",
  13018=>"000000000",
  13019=>"111111111",
  13020=>"000000000",
  13021=>"100000000",
  13022=>"110110110",
  13023=>"111111000",
  13024=>"000010011",
  13025=>"101101111",
  13026=>"111000000",
  13027=>"111111111",
  13028=>"111101000",
  13029=>"001001000",
  13030=>"000000001",
  13031=>"000000111",
  13032=>"111111000",
  13033=>"001111111",
  13034=>"000000000",
  13035=>"100100111",
  13036=>"000011111",
  13037=>"000000111",
  13038=>"000001000",
  13039=>"111111100",
  13040=>"000000001",
  13041=>"000000000",
  13042=>"100110111",
  13043=>"000000001",
  13044=>"000000000",
  13045=>"110111111",
  13046=>"011000000",
  13047=>"111111111",
  13048=>"100100100",
  13049=>"111111111",
  13050=>"100110110",
  13051=>"110000000",
  13052=>"011011011",
  13053=>"011010110",
  13054=>"000100001",
  13055=>"000000001",
  13056=>"100110100",
  13057=>"110110100",
  13058=>"111101001",
  13059=>"111111101",
  13060=>"000110111",
  13061=>"000100000",
  13062=>"000000101",
  13063=>"001001000",
  13064=>"000100111",
  13065=>"000000000",
  13066=>"111111111",
  13067=>"111111111",
  13068=>"000000110",
  13069=>"111000000",
  13070=>"111101110",
  13071=>"111111111",
  13072=>"101100111",
  13073=>"000000000",
  13074=>"100000111",
  13075=>"100100000",
  13076=>"111111111",
  13077=>"111000100",
  13078=>"100110000",
  13079=>"000111111",
  13080=>"110110110",
  13081=>"100000001",
  13082=>"111111100",
  13083=>"000000000",
  13084=>"100110100",
  13085=>"111110100",
  13086=>"101011001",
  13087=>"111111111",
  13088=>"000000100",
  13089=>"000000000",
  13090=>"000100101",
  13091=>"000000000",
  13092=>"111111110",
  13093=>"000000000",
  13094=>"000000000",
  13095=>"000101111",
  13096=>"111100000",
  13097=>"000001001",
  13098=>"110110101",
  13099=>"011111111",
  13100=>"111111101",
  13101=>"111110010",
  13102=>"000000000",
  13103=>"001010111",
  13104=>"111001001",
  13105=>"011011011",
  13106=>"000000000",
  13107=>"100110111",
  13108=>"111001000",
  13109=>"000111111",
  13110=>"111000111",
  13111=>"001000000",
  13112=>"000000000",
  13113=>"011001011",
  13114=>"000000011",
  13115=>"110111100",
  13116=>"110110011",
  13117=>"011010000",
  13118=>"000000000",
  13119=>"111111000",
  13120=>"000010000",
  13121=>"000000000",
  13122=>"110110000",
  13123=>"000000000",
  13124=>"111100000",
  13125=>"111100110",
  13126=>"011001000",
  13127=>"000011111",
  13128=>"000100100",
  13129=>"000000000",
  13130=>"011000000",
  13131=>"111111000",
  13132=>"000000000",
  13133=>"111111100",
  13134=>"101111001",
  13135=>"110111100",
  13136=>"011111001",
  13137=>"111111111",
  13138=>"111111100",
  13139=>"101000000",
  13140=>"101111000",
  13141=>"011011001",
  13142=>"100000000",
  13143=>"111111111",
  13144=>"000000000",
  13145=>"000000000",
  13146=>"010000000",
  13147=>"000110111",
  13148=>"011000000",
  13149=>"000111111",
  13150=>"000000000",
  13151=>"001111111",
  13152=>"111011011",
  13153=>"111110111",
  13154=>"001011011",
  13155=>"001001000",
  13156=>"111111111",
  13157=>"000000000",
  13158=>"000000000",
  13159=>"111111111",
  13160=>"011001101",
  13161=>"000000000",
  13162=>"000101000",
  13163=>"110010000",
  13164=>"111000100",
  13165=>"000000111",
  13166=>"000001111",
  13167=>"010011000",
  13168=>"000000000",
  13169=>"111111111",
  13170=>"011111111",
  13171=>"001011011",
  13172=>"111111001",
  13173=>"111110000",
  13174=>"010010000",
  13175=>"100111001",
  13176=>"001000000",
  13177=>"111000110",
  13178=>"000000110",
  13179=>"111000100",
  13180=>"000000010",
  13181=>"000000000",
  13182=>"111111100",
  13183=>"101000000",
  13184=>"111111111",
  13185=>"101001101",
  13186=>"111111111",
  13187=>"110111001",
  13188=>"000100111",
  13189=>"000011001",
  13190=>"000011011",
  13191=>"111111100",
  13192=>"000111111",
  13193=>"000100111",
  13194=>"101101101",
  13195=>"111000000",
  13196=>"101100101",
  13197=>"110110110",
  13198=>"001000101",
  13199=>"000000000",
  13200=>"110000000",
  13201=>"111111100",
  13202=>"000000000",
  13203=>"000000100",
  13204=>"000000000",
  13205=>"001111011",
  13206=>"000000100",
  13207=>"010110000",
  13208=>"111111000",
  13209=>"111111110",
  13210=>"011111111",
  13211=>"010011000",
  13212=>"011001001",
  13213=>"111111111",
  13214=>"011111001",
  13215=>"101100000",
  13216=>"111111111",
  13217=>"011011011",
  13218=>"111111111",
  13219=>"000001000",
  13220=>"000000110",
  13221=>"111111001",
  13222=>"000000000",
  13223=>"100100111",
  13224=>"011111000",
  13225=>"000100111",
  13226=>"001000000",
  13227=>"000010110",
  13228=>"100100100",
  13229=>"111110111",
  13230=>"000000100",
  13231=>"111110100",
  13232=>"000110000",
  13233=>"000000110",
  13234=>"111111111",
  13235=>"000111011",
  13236=>"000110111",
  13237=>"100111111",
  13238=>"111111111",
  13239=>"111110101",
  13240=>"111011100",
  13241=>"000111111",
  13242=>"111000100",
  13243=>"001111111",
  13244=>"000000111",
  13245=>"111001000",
  13246=>"000000000",
  13247=>"000100110",
  13248=>"111111111",
  13249=>"110110111",
  13250=>"000000000",
  13251=>"000000010",
  13252=>"100110111",
  13253=>"000001111",
  13254=>"000000000",
  13255=>"111111000",
  13256=>"000000000",
  13257=>"001001000",
  13258=>"001001000",
  13259=>"000000000",
  13260=>"000000000",
  13261=>"111111111",
  13262=>"000000000",
  13263=>"000010010",
  13264=>"000000000",
  13265=>"111111111",
  13266=>"111111111",
  13267=>"100000111",
  13268=>"001001001",
  13269=>"000110111",
  13270=>"101101111",
  13271=>"100000100",
  13272=>"000000000",
  13273=>"111000001",
  13274=>"010010000",
  13275=>"001110110",
  13276=>"111111111",
  13277=>"001001001",
  13278=>"000100100",
  13279=>"011111111",
  13280=>"010111111",
  13281=>"101111111",
  13282=>"100111111",
  13283=>"111111111",
  13284=>"000010111",
  13285=>"000000111",
  13286=>"000000110",
  13287=>"000000110",
  13288=>"111111111",
  13289=>"111111111",
  13290=>"110110110",
  13291=>"000000000",
  13292=>"001111111",
  13293=>"001011001",
  13294=>"000000000",
  13295=>"000010011",
  13296=>"000000000",
  13297=>"011110111",
  13298=>"111111111",
  13299=>"110000111",
  13300=>"001000000",
  13301=>"001011000",
  13302=>"111111111",
  13303=>"111000100",
  13304=>"111111000",
  13305=>"001001001",
  13306=>"101000110",
  13307=>"111111111",
  13308=>"010110111",
  13309=>"111111111",
  13310=>"000000011",
  13311=>"000000000",
  13312=>"000001011",
  13313=>"111000010",
  13314=>"100000100",
  13315=>"000000000",
  13316=>"111011101",
  13317=>"111111111",
  13318=>"011011000",
  13319=>"110110100",
  13320=>"000001000",
  13321=>"110000000",
  13322=>"001001001",
  13323=>"000000100",
  13324=>"101000000",
  13325=>"001000111",
  13326=>"010000100",
  13327=>"000010100",
  13328=>"100100001",
  13329=>"001110100",
  13330=>"111111001",
  13331=>"001001011",
  13332=>"010000000",
  13333=>"001001110",
  13334=>"010000000",
  13335=>"000110110",
  13336=>"111111110",
  13337=>"111111111",
  13338=>"001000000",
  13339=>"111111110",
  13340=>"011010011",
  13341=>"000000001",
  13342=>"011000000",
  13343=>"010111000",
  13344=>"100111011",
  13345=>"000000000",
  13346=>"100110111",
  13347=>"000000000",
  13348=>"000000000",
  13349=>"100110110",
  13350=>"000000000",
  13351=>"111100010",
  13352=>"001111000",
  13353=>"100000000",
  13354=>"010110110",
  13355=>"110100100",
  13356=>"000100111",
  13357=>"001001000",
  13358=>"111111011",
  13359=>"111111000",
  13360=>"000000000",
  13361=>"000000001",
  13362=>"000100000",
  13363=>"111011011",
  13364=>"001001001",
  13365=>"111111111",
  13366=>"111000000",
  13367=>"111111000",
  13368=>"111001001",
  13369=>"010000111",
  13370=>"111111111",
  13371=>"100000100",
  13372=>"100100101",
  13373=>"110100100",
  13374=>"000000000",
  13375=>"111111111",
  13376=>"110100100",
  13377=>"000011011",
  13378=>"000000000",
  13379=>"111100111",
  13380=>"111111111",
  13381=>"011111111",
  13382=>"000011000",
  13383=>"100000100",
  13384=>"000000001",
  13385=>"000000000",
  13386=>"111111110",
  13387=>"000000100",
  13388=>"000000000",
  13389=>"000100100",
  13390=>"100000011",
  13391=>"010101100",
  13392=>"111011011",
  13393=>"101001000",
  13394=>"110111111",
  13395=>"110110001",
  13396=>"001100001",
  13397=>"111111111",
  13398=>"100000100",
  13399=>"110111111",
  13400=>"001011011",
  13401=>"111101100",
  13402=>"111011000",
  13403=>"110100100",
  13404=>"111010011",
  13405=>"000001011",
  13406=>"110110100",
  13407=>"111111111",
  13408=>"000000000",
  13409=>"000000000",
  13410=>"001000000",
  13411=>"111111111",
  13412=>"000000001",
  13413=>"000110111",
  13414=>"111001000",
  13415=>"001101111",
  13416=>"000000010",
  13417=>"111011111",
  13418=>"111000111",
  13419=>"000110110",
  13420=>"000001011",
  13421=>"000000011",
  13422=>"110111110",
  13423=>"011101111",
  13424=>"011000000",
  13425=>"111111111",
  13426=>"111100000",
  13427=>"000000000",
  13428=>"011011000",
  13429=>"111101101",
  13430=>"011000000",
  13431=>"001000000",
  13432=>"000000111",
  13433=>"111111110",
  13434=>"001001001",
  13435=>"111111011",
  13436=>"111110111",
  13437=>"101111111",
  13438=>"001001011",
  13439=>"000000000",
  13440=>"110110011",
  13441=>"111111111",
  13442=>"000000000",
  13443=>"100100100",
  13444=>"111011101",
  13445=>"111111111",
  13446=>"000000000",
  13447=>"000000000",
  13448=>"000000111",
  13449=>"110111111",
  13450=>"000100111",
  13451=>"111111000",
  13452=>"101000001",
  13453=>"111111110",
  13454=>"111111111",
  13455=>"111110111",
  13456=>"111111111",
  13457=>"111111000",
  13458=>"000000111",
  13459=>"000000000",
  13460=>"000111111",
  13461=>"000110110",
  13462=>"111000000",
  13463=>"111111111",
  13464=>"000000001",
  13465=>"000000001",
  13466=>"000000000",
  13467=>"000110100",
  13468=>"111111110",
  13469=>"000011101",
  13470=>"111011111",
  13471=>"111111111",
  13472=>"000000000",
  13473=>"111111111",
  13474=>"111011011",
  13475=>"100100110",
  13476=>"011001001",
  13477=>"111111110",
  13478=>"000000000",
  13479=>"111111001",
  13480=>"001000000",
  13481=>"101000000",
  13482=>"001000000",
  13483=>"111111111",
  13484=>"111000011",
  13485=>"100110100",
  13486=>"111111011",
  13487=>"111101101",
  13488=>"111111111",
  13489=>"111111111",
  13490=>"111010011",
  13491=>"010000000",
  13492=>"111111011",
  13493=>"110011001",
  13494=>"000000000",
  13495=>"000000111",
  13496=>"000000000",
  13497=>"111111011",
  13498=>"001101000",
  13499=>"100100110",
  13500=>"000110000",
  13501=>"110110111",
  13502=>"000000000",
  13503=>"111110111",
  13504=>"000000101",
  13505=>"111111111",
  13506=>"000010011",
  13507=>"000000000",
  13508=>"111111010",
  13509=>"000000001",
  13510=>"011111000",
  13511=>"111111111",
  13512=>"000000000",
  13513=>"100000000",
  13514=>"010111111",
  13515=>"001011010",
  13516=>"111111101",
  13517=>"111111111",
  13518=>"000000000",
  13519=>"010000000",
  13520=>"000010000",
  13521=>"000000001",
  13522=>"000011011",
  13523=>"000000000",
  13524=>"011011111",
  13525=>"100000000",
  13526=>"000000001",
  13527=>"000000001",
  13528=>"000001001",
  13529=>"111111110",
  13530=>"000000000",
  13531=>"100000000",
  13532=>"000000000",
  13533=>"111111111",
  13534=>"111111001",
  13535=>"100111111",
  13536=>"001001111",
  13537=>"000000100",
  13538=>"100000000",
  13539=>"111111111",
  13540=>"000000000",
  13541=>"010011011",
  13542=>"000000010",
  13543=>"000000010",
  13544=>"111101110",
  13545=>"001001011",
  13546=>"111111111",
  13547=>"001000001",
  13548=>"000000000",
  13549=>"000000110",
  13550=>"111100110",
  13551=>"000000000",
  13552=>"010010011",
  13553=>"011000010",
  13554=>"111111111",
  13555=>"101101101",
  13556=>"011000011",
  13557=>"111111100",
  13558=>"110100101",
  13559=>"111111111",
  13560=>"000000000",
  13561=>"000000000",
  13562=>"111011111",
  13563=>"111111111",
  13564=>"000000000",
  13565=>"000001101",
  13566=>"100100111",
  13567=>"101001001",
  13568=>"100000111",
  13569=>"110111111",
  13570=>"111111001",
  13571=>"010010000",
  13572=>"001001101",
  13573=>"111110000",
  13574=>"101001000",
  13575=>"100000101",
  13576=>"101101111",
  13577=>"000000000",
  13578=>"000100100",
  13579=>"100000100",
  13580=>"000000000",
  13581=>"111011001",
  13582=>"111111111",
  13583=>"000000000",
  13584=>"101000000",
  13585=>"111111111",
  13586=>"000000000",
  13587=>"000101111",
  13588=>"000011011",
  13589=>"111111111",
  13590=>"100100100",
  13591=>"000000101",
  13592=>"010010111",
  13593=>"111111011",
  13594=>"111111111",
  13595=>"000111011",
  13596=>"011011101",
  13597=>"111111111",
  13598=>"111111111",
  13599=>"000011001",
  13600=>"000000001",
  13601=>"111111000",
  13602=>"111111000",
  13603=>"000000000",
  13604=>"111011000",
  13605=>"000100000",
  13606=>"011001000",
  13607=>"000011011",
  13608=>"000000000",
  13609=>"011000000",
  13610=>"100110111",
  13611=>"000000011",
  13612=>"111111111",
  13613=>"111110110",
  13614=>"000110010",
  13615=>"111000000",
  13616=>"111000001",
  13617=>"011011111",
  13618=>"000010100",
  13619=>"000000001",
  13620=>"000000000",
  13621=>"001011001",
  13622=>"111111111",
  13623=>"101101111",
  13624=>"001001111",
  13625=>"000000100",
  13626=>"011000100",
  13627=>"111100000",
  13628=>"110000110",
  13629=>"000001001",
  13630=>"010111111",
  13631=>"000010110",
  13632=>"000000101",
  13633=>"000000000",
  13634=>"110010110",
  13635=>"000101111",
  13636=>"111111111",
  13637=>"110000000",
  13638=>"000011111",
  13639=>"111100000",
  13640=>"100100111",
  13641=>"000000000",
  13642=>"111000000",
  13643=>"000000000",
  13644=>"000011011",
  13645=>"111111011",
  13646=>"100011100",
  13647=>"001001001",
  13648=>"010010011",
  13649=>"110000100",
  13650=>"111011111",
  13651=>"001000000",
  13652=>"100101001",
  13653=>"001000000",
  13654=>"110000000",
  13655=>"000000000",
  13656=>"100111111",
  13657=>"110100000",
  13658=>"110100100",
  13659=>"111100111",
  13660=>"000000000",
  13661=>"001001011",
  13662=>"111111111",
  13663=>"110111111",
  13664=>"111111110",
  13665=>"011011111",
  13666=>"101000000",
  13667=>"000000111",
  13668=>"000001001",
  13669=>"111111111",
  13670=>"000001111",
  13671=>"000000000",
  13672=>"000000000",
  13673=>"000000001",
  13674=>"000000000",
  13675=>"000000000",
  13676=>"111011001",
  13677=>"100100000",
  13678=>"000100000",
  13679=>"111111111",
  13680=>"111000001",
  13681=>"100100011",
  13682=>"111111111",
  13683=>"000000000",
  13684=>"011011000",
  13685=>"000000011",
  13686=>"110111000",
  13687=>"100111100",
  13688=>"000000111",
  13689=>"101000000",
  13690=>"001000100",
  13691=>"100100111",
  13692=>"011011111",
  13693=>"111111111",
  13694=>"110000000",
  13695=>"000000100",
  13696=>"110110000",
  13697=>"001001001",
  13698=>"110011011",
  13699=>"011011111",
  13700=>"110000000",
  13701=>"001001000",
  13702=>"000010000",
  13703=>"100000000",
  13704=>"011011010",
  13705=>"011010111",
  13706=>"111111111",
  13707=>"000000000",
  13708=>"111111111",
  13709=>"110110001",
  13710=>"101000000",
  13711=>"010110011",
  13712=>"000000000",
  13713=>"110110100",
  13714=>"000000000",
  13715=>"001000011",
  13716=>"000000000",
  13717=>"000011011",
  13718=>"100000000",
  13719=>"111100101",
  13720=>"100000101",
  13721=>"111111110",
  13722=>"000000111",
  13723=>"111111111",
  13724=>"111111111",
  13725=>"111110001",
  13726=>"111000001",
  13727=>"000000000",
  13728=>"011001000",
  13729=>"111001000",
  13730=>"100000100",
  13731=>"111001001",
  13732=>"000000000",
  13733=>"101101111",
  13734=>"001000000",
  13735=>"000110110",
  13736=>"100000000",
  13737=>"111111110",
  13738=>"111111100",
  13739=>"111111111",
  13740=>"000000000",
  13741=>"111100011",
  13742=>"000000000",
  13743=>"111010010",
  13744=>"110000000",
  13745=>"000100000",
  13746=>"101100100",
  13747=>"001111100",
  13748=>"001011000",
  13749=>"111011001",
  13750=>"101101111",
  13751=>"000000011",
  13752=>"011000000",
  13753=>"100000000",
  13754=>"111111111",
  13755=>"000110111",
  13756=>"000000000",
  13757=>"000000000",
  13758=>"100001011",
  13759=>"100000000",
  13760=>"101100011",
  13761=>"110111010",
  13762=>"111011001",
  13763=>"111000000",
  13764=>"110000000",
  13765=>"000010110",
  13766=>"110110000",
  13767=>"000101111",
  13768=>"111100111",
  13769=>"100100000",
  13770=>"001000000",
  13771=>"000011011",
  13772=>"111101000",
  13773=>"000000000",
  13774=>"100100111",
  13775=>"111111111",
  13776=>"000000000",
  13777=>"000000000",
  13778=>"000001011",
  13779=>"111111111",
  13780=>"111101001",
  13781=>"111010000",
  13782=>"111111111",
  13783=>"110000111",
  13784=>"111111111",
  13785=>"011111100",
  13786=>"111111101",
  13787=>"111111111",
  13788=>"111110100",
  13789=>"101111101",
  13790=>"000010110",
  13791=>"111111001",
  13792=>"000000001",
  13793=>"000000000",
  13794=>"010000000",
  13795=>"100001011",
  13796=>"010000000",
  13797=>"000001111",
  13798=>"000000000",
  13799=>"010000110",
  13800=>"100110000",
  13801=>"100101101",
  13802=>"111111111",
  13803=>"000000101",
  13804=>"000000111",
  13805=>"000000000",
  13806=>"011001011",
  13807=>"010010111",
  13808=>"000110111",
  13809=>"111111111",
  13810=>"111111111",
  13811=>"000001001",
  13812=>"111101111",
  13813=>"000000000",
  13814=>"111111111",
  13815=>"000000000",
  13816=>"111001111",
  13817=>"000001011",
  13818=>"111001111",
  13819=>"001001011",
  13820=>"000101101",
  13821=>"100111111",
  13822=>"111111111",
  13823=>"111011011",
  13824=>"111111111",
  13825=>"000000000",
  13826=>"111111000",
  13827=>"001011000",
  13828=>"000000000",
  13829=>"000000111",
  13830=>"111111000",
  13831=>"000000000",
  13832=>"000000000",
  13833=>"111111111",
  13834=>"111111000",
  13835=>"000000011",
  13836=>"000100101",
  13837=>"001111111",
  13838=>"111111111",
  13839=>"111111111",
  13840=>"101111111",
  13841=>"111001111",
  13842=>"000000000",
  13843=>"001000000",
  13844=>"111111111",
  13845=>"000000000",
  13846=>"000000000",
  13847=>"000000000",
  13848=>"111011101",
  13849=>"001000110",
  13850=>"000000101",
  13851=>"000000000",
  13852=>"011011000",
  13853=>"111110100",
  13854=>"001011001",
  13855=>"010111111",
  13856=>"000111111",
  13857=>"110110110",
  13858=>"000000000",
  13859=>"111111111",
  13860=>"000011111",
  13861=>"000000000",
  13862=>"111010111",
  13863=>"000000000",
  13864=>"001000000",
  13865=>"000000000",
  13866=>"111111000",
  13867=>"000000000",
  13868=>"111000001",
  13869=>"111111111",
  13870=>"101111001",
  13871=>"100000000",
  13872=>"010000000",
  13873=>"000000000",
  13874=>"111111111",
  13875=>"000101111",
  13876=>"000101101",
  13877=>"000000000",
  13878=>"000100101",
  13879=>"101100100",
  13880=>"111111111",
  13881=>"000000000",
  13882=>"001001000",
  13883=>"110111110",
  13884=>"000000000",
  13885=>"111111111",
  13886=>"110110100",
  13887=>"000000000",
  13888=>"111111100",
  13889=>"111000001",
  13890=>"111111111",
  13891=>"001001101",
  13892=>"111111111",
  13893=>"000000000",
  13894=>"000110000",
  13895=>"111111111",
  13896=>"000000000",
  13897=>"111111110",
  13898=>"101111111",
  13899=>"111111100",
  13900=>"000000000",
  13901=>"000000000",
  13902=>"000000000",
  13903=>"111110000",
  13904=>"000000111",
  13905=>"001001001",
  13906=>"111111111",
  13907=>"000110110",
  13908=>"000000000",
  13909=>"001001000",
  13910=>"111111111",
  13911=>"000000000",
  13912=>"000010010",
  13913=>"110111011",
  13914=>"111100111",
  13915=>"000100001",
  13916=>"111111111",
  13917=>"000000000",
  13918=>"010111111",
  13919=>"000000000",
  13920=>"000000000",
  13921=>"000111111",
  13922=>"011111111",
  13923=>"100100111",
  13924=>"111111111",
  13925=>"101011011",
  13926=>"000000000",
  13927=>"111000000",
  13928=>"111111110",
  13929=>"011111111",
  13930=>"001001000",
  13931=>"111101111",
  13932=>"000000101",
  13933=>"111011111",
  13934=>"111111111",
  13935=>"000000111",
  13936=>"000000100",
  13937=>"000000000",
  13938=>"001111011",
  13939=>"111000000",
  13940=>"000000111",
  13941=>"111100000",
  13942=>"100100000",
  13943=>"000000110",
  13944=>"011111000",
  13945=>"000000000",
  13946=>"000001111",
  13947=>"010000000",
  13948=>"000000000",
  13949=>"000000000",
  13950=>"000000000",
  13951=>"000000100",
  13952=>"111111111",
  13953=>"000001111",
  13954=>"000000000",
  13955=>"000111111",
  13956=>"111101111",
  13957=>"111001000",
  13958=>"011111111",
  13959=>"111000000",
  13960=>"100111111",
  13961=>"111000000",
  13962=>"111111000",
  13963=>"000000000",
  13964=>"111101100",
  13965=>"111110101",
  13966=>"000011110",
  13967=>"001001000",
  13968=>"000000000",
  13969=>"000101000",
  13970=>"000000000",
  13971=>"000000100",
  13972=>"011011111",
  13973=>"000010110",
  13974=>"111011000",
  13975=>"000000000",
  13976=>"111111100",
  13977=>"111111111",
  13978=>"111111111",
  13979=>"111111111",
  13980=>"000000000",
  13981=>"001001111",
  13982=>"000000000",
  13983=>"000000111",
  13984=>"001001111",
  13985=>"001101110",
  13986=>"111111111",
  13987=>"000000000",
  13988=>"100100110",
  13989=>"000011111",
  13990=>"111111111",
  13991=>"000001000",
  13992=>"001000000",
  13993=>"000011000",
  13994=>"111111111",
  13995=>"000011111",
  13996=>"111111000",
  13997=>"111111111",
  13998=>"000000000",
  13999=>"000000100",
  14000=>"110010111",
  14001=>"100111000",
  14002=>"111111110",
  14003=>"111111110",
  14004=>"111110000",
  14005=>"111111000",
  14006=>"000111111",
  14007=>"111111111",
  14008=>"110110000",
  14009=>"111111111",
  14010=>"000000000",
  14011=>"011001001",
  14012=>"000000000",
  14013=>"001000001",
  14014=>"100000000",
  14015=>"000001101",
  14016=>"100000111",
  14017=>"000000001",
  14018=>"000000000",
  14019=>"000000000",
  14020=>"110110000",
  14021=>"000000000",
  14022=>"111111011",
  14023=>"001111111",
  14024=>"011111110",
  14025=>"111111110",
  14026=>"110000110",
  14027=>"000000000",
  14028=>"111111111",
  14029=>"000000000",
  14030=>"000000000",
  14031=>"011011000",
  14032=>"001001111",
  14033=>"000000000",
  14034=>"111111111",
  14035=>"011011000",
  14036=>"000000000",
  14037=>"000000000",
  14038=>"111111000",
  14039=>"001000000",
  14040=>"011011111",
  14041=>"000011011",
  14042=>"111111111",
  14043=>"111001001",
  14044=>"000000000",
  14045=>"011011110",
  14046=>"111011111",
  14047=>"011011000",
  14048=>"111111111",
  14049=>"110000000",
  14050=>"111001000",
  14051=>"111100000",
  14052=>"100110110",
  14053=>"100111100",
  14054=>"111111111",
  14055=>"000000000",
  14056=>"000000000",
  14057=>"000001000",
  14058=>"111111111",
  14059=>"000010111",
  14060=>"000000000",
  14061=>"110000111",
  14062=>"111011001",
  14063=>"000010110",
  14064=>"111111111",
  14065=>"000100010",
  14066=>"111111111",
  14067=>"100000000",
  14068=>"110000000",
  14069=>"001000000",
  14070=>"101101011",
  14071=>"111000000",
  14072=>"000000000",
  14073=>"011001001",
  14074=>"000000000",
  14075=>"010000000",
  14076=>"000001001",
  14077=>"000011111",
  14078=>"000011001",
  14079=>"111111111",
  14080=>"000000000",
  14081=>"011011011",
  14082=>"000000000",
  14083=>"111111000",
  14084=>"000000000",
  14085=>"111111111",
  14086=>"111110111",
  14087=>"000000000",
  14088=>"000000011",
  14089=>"000000000",
  14090=>"000000001",
  14091=>"000111110",
  14092=>"111111000",
  14093=>"111111000",
  14094=>"111111001",
  14095=>"000000000",
  14096=>"000010010",
  14097=>"000000000",
  14098=>"101111111",
  14099=>"111111111",
  14100=>"000000000",
  14101=>"000000000",
  14102=>"000000000",
  14103=>"000000000",
  14104=>"011110110",
  14105=>"110000111",
  14106=>"000000000",
  14107=>"001001111",
  14108=>"111111111",
  14109=>"111111101",
  14110=>"000011010",
  14111=>"000000000",
  14112=>"111111111",
  14113=>"000000111",
  14114=>"001000010",
  14115=>"111111111",
  14116=>"100110101",
  14117=>"000000000",
  14118=>"001000000",
  14119=>"000000000",
  14120=>"001000000",
  14121=>"000110000",
  14122=>"000000000",
  14123=>"111111111",
  14124=>"011110110",
  14125=>"001011111",
  14126=>"110110111",
  14127=>"000010000",
  14128=>"010010110",
  14129=>"001111111",
  14130=>"011000000",
  14131=>"011010011",
  14132=>"111111111",
  14133=>"100000000",
  14134=>"000000111",
  14135=>"000000000",
  14136=>"111111110",
  14137=>"111000111",
  14138=>"111001111",
  14139=>"111000000",
  14140=>"011011011",
  14141=>"000110000",
  14142=>"111111111",
  14143=>"000000000",
  14144=>"000000000",
  14145=>"110110110",
  14146=>"110111110",
  14147=>"000000000",
  14148=>"001011011",
  14149=>"000000000",
  14150=>"000000000",
  14151=>"110111000",
  14152=>"000000111",
  14153=>"111111111",
  14154=>"001111111",
  14155=>"000101000",
  14156=>"011000000",
  14157=>"011001000",
  14158=>"000011111",
  14159=>"100110110",
  14160=>"000000000",
  14161=>"000000000",
  14162=>"000100000",
  14163=>"001000000",
  14164=>"010111111",
  14165=>"011011011",
  14166=>"110111111",
  14167=>"000000000",
  14168=>"111111111",
  14169=>"101111110",
  14170=>"111111100",
  14171=>"000111111",
  14172=>"111001001",
  14173=>"111111000",
  14174=>"000000000",
  14175=>"110100000",
  14176=>"111111111",
  14177=>"000000000",
  14178=>"100111111",
  14179=>"010011000",
  14180=>"111111111",
  14181=>"000000010",
  14182=>"000000001",
  14183=>"111111111",
  14184=>"001011000",
  14185=>"000001000",
  14186=>"001001000",
  14187=>"111111111",
  14188=>"111111111",
  14189=>"111111111",
  14190=>"000000000",
  14191=>"111111111",
  14192=>"101001001",
  14193=>"111111111",
  14194=>"000000011",
  14195=>"010001011",
  14196=>"111111110",
  14197=>"001001001",
  14198=>"111110111",
  14199=>"011010000",
  14200=>"000000000",
  14201=>"000000000",
  14202=>"000000000",
  14203=>"011111011",
  14204=>"000000010",
  14205=>"111001000",
  14206=>"000000000",
  14207=>"111111001",
  14208=>"111110111",
  14209=>"111111111",
  14210=>"000000000",
  14211=>"000000000",
  14212=>"001000011",
  14213=>"110111000",
  14214=>"011111111",
  14215=>"000000000",
  14216=>"111111111",
  14217=>"000000000",
  14218=>"111111111",
  14219=>"111111111",
  14220=>"111111111",
  14221=>"000010000",
  14222=>"000011111",
  14223=>"101000000",
  14224=>"000000001",
  14225=>"101100000",
  14226=>"111011100",
  14227=>"111111111",
  14228=>"000000000",
  14229=>"000000000",
  14230=>"111100111",
  14231=>"000000000",
  14232=>"000000000",
  14233=>"000110110",
  14234=>"110000000",
  14235=>"111111111",
  14236=>"000000000",
  14237=>"000001001",
  14238=>"111000000",
  14239=>"100111111",
  14240=>"001000000",
  14241=>"110110110",
  14242=>"000000001",
  14243=>"111111111",
  14244=>"110000000",
  14245=>"110110000",
  14246=>"000000111",
  14247=>"000000000",
  14248=>"000111111",
  14249=>"000111111",
  14250=>"110110111",
  14251=>"000000000",
  14252=>"000000000",
  14253=>"000000000",
  14254=>"010110000",
  14255=>"001111101",
  14256=>"000000000",
  14257=>"111011000",
  14258=>"000010000",
  14259=>"111011111",
  14260=>"111111111",
  14261=>"000000000",
  14262=>"100101111",
  14263=>"110111010",
  14264=>"001011111",
  14265=>"100001000",
  14266=>"000100100",
  14267=>"111111111",
  14268=>"000000000",
  14269=>"010010000",
  14270=>"000000011",
  14271=>"000000000",
  14272=>"100100000",
  14273=>"000000000",
  14274=>"000101100",
  14275=>"110100101",
  14276=>"110000100",
  14277=>"111111111",
  14278=>"101000000",
  14279=>"111111111",
  14280=>"000000000",
  14281=>"000000000",
  14282=>"100111111",
  14283=>"000001001",
  14284=>"011111111",
  14285=>"000000000",
  14286=>"111011111",
  14287=>"000000000",
  14288=>"000000000",
  14289=>"011000001",
  14290=>"000000000",
  14291=>"000000000",
  14292=>"111111111",
  14293=>"000000000",
  14294=>"001011111",
  14295=>"100100101",
  14296=>"111111111",
  14297=>"110010000",
  14298=>"111110000",
  14299=>"101000101",
  14300=>"011111111",
  14301=>"111001110",
  14302=>"000110111",
  14303=>"011010000",
  14304=>"111111111",
  14305=>"000000000",
  14306=>"000000000",
  14307=>"111001111",
  14308=>"011000000",
  14309=>"000000001",
  14310=>"000000000",
  14311=>"000000001",
  14312=>"111011111",
  14313=>"100100011",
  14314=>"111111111",
  14315=>"000011111",
  14316=>"001000000",
  14317=>"100111111",
  14318=>"110110000",
  14319=>"110100111",
  14320=>"111110000",
  14321=>"000111111",
  14322=>"111111111",
  14323=>"111111111",
  14324=>"011111111",
  14325=>"000000000",
  14326=>"011011001",
  14327=>"011001111",
  14328=>"111111000",
  14329=>"000000000",
  14330=>"101001111",
  14331=>"000000000",
  14332=>"111111111",
  14333=>"111111111",
  14334=>"101001000",
  14335=>"111111111",
  14336=>"000000001",
  14337=>"111111010",
  14338=>"111111111",
  14339=>"111111111",
  14340=>"000110111",
  14341=>"000000101",
  14342=>"000000000",
  14343=>"111001111",
  14344=>"111111111",
  14345=>"000001101",
  14346=>"100111111",
  14347=>"100111111",
  14348=>"100000000",
  14349=>"000000111",
  14350=>"001000000",
  14351=>"000000000",
  14352=>"000010111",
  14353=>"000000001",
  14354=>"000000000",
  14355=>"110000000",
  14356=>"000111000",
  14357=>"100110111",
  14358=>"011000000",
  14359=>"000000111",
  14360=>"000000000",
  14361=>"111011111",
  14362=>"111111101",
  14363=>"000001111",
  14364=>"000000000",
  14365=>"011111111",
  14366=>"011011011",
  14367=>"010010000",
  14368=>"110110001",
  14369=>"111101001",
  14370=>"000001001",
  14371=>"111111000",
  14372=>"000000000",
  14373=>"001101111",
  14374=>"101101100",
  14375=>"100101111",
  14376=>"000110100",
  14377=>"000000000",
  14378=>"110100101",
  14379=>"010111010",
  14380=>"001111111",
  14381=>"000000000",
  14382=>"100111111",
  14383=>"111111111",
  14384=>"000111001",
  14385=>"001111011",
  14386=>"001011111",
  14387=>"000110110",
  14388=>"100110101",
  14389=>"100001000",
  14390=>"111111111",
  14391=>"111111110",
  14392=>"000001001",
  14393=>"111111111",
  14394=>"000110111",
  14395=>"000000001",
  14396=>"101000100",
  14397=>"010111111",
  14398=>"000000000",
  14399=>"010101111",
  14400=>"111111110",
  14401=>"101111111",
  14402=>"000000000",
  14403=>"000001110",
  14404=>"000001011",
  14405=>"001001000",
  14406=>"000000111",
  14407=>"000101111",
  14408=>"011011011",
  14409=>"000000000",
  14410=>"001111111",
  14411=>"001111111",
  14412=>"110111110",
  14413=>"100101011",
  14414=>"111001101",
  14415=>"111111111",
  14416=>"111110100",
  14417=>"010111111",
  14418=>"000000000",
  14419=>"101000001",
  14420=>"000100111",
  14421=>"000000000",
  14422=>"111111111",
  14423=>"110110111",
  14424=>"000001000",
  14425=>"000000111",
  14426=>"001111111",
  14427=>"110100001",
  14428=>"000000000",
  14429=>"111111111",
  14430=>"110000000",
  14431=>"000001011",
  14432=>"000000001",
  14433=>"111111110",
  14434=>"000100111",
  14435=>"111111111",
  14436=>"000000001",
  14437=>"111000000",
  14438=>"001000000",
  14439=>"001001011",
  14440=>"000000000",
  14441=>"101001101",
  14442=>"001011001",
  14443=>"000000000",
  14444=>"000011000",
  14445=>"000000000",
  14446=>"000000001",
  14447=>"010000000",
  14448=>"000111111",
  14449=>"001001100",
  14450=>"100100101",
  14451=>"111110110",
  14452=>"111111000",
  14453=>"111111111",
  14454=>"011111011",
  14455=>"001000101",
  14456=>"100000010",
  14457=>"100000000",
  14458=>"001001001",
  14459=>"111111111",
  14460=>"100110100",
  14461=>"000000100",
  14462=>"011111000",
  14463=>"000000000",
  14464=>"100000000",
  14465=>"000111111",
  14466=>"000000000",
  14467=>"000000000",
  14468=>"000000000",
  14469=>"110000000",
  14470=>"110110000",
  14471=>"000000000",
  14472=>"111111011",
  14473=>"000000000",
  14474=>"111110000",
  14475=>"111100000",
  14476=>"111111111",
  14477=>"101100100",
  14478=>"000000100",
  14479=>"000001001",
  14480=>"111111101",
  14481=>"111111001",
  14482=>"010100000",
  14483=>"100110111",
  14484=>"101000010",
  14485=>"111111101",
  14486=>"000000100",
  14487=>"000100100",
  14488=>"111111001",
  14489=>"111111110",
  14490=>"001000000",
  14491=>"110111001",
  14492=>"100101011",
  14493=>"110010000",
  14494=>"000001111",
  14495=>"100000000",
  14496=>"000010000",
  14497=>"010111111",
  14498=>"011001001",
  14499=>"111110000",
  14500=>"100000000",
  14501=>"101100000",
  14502=>"001001001",
  14503=>"010010011",
  14504=>"000000100",
  14505=>"000000000",
  14506=>"000000000",
  14507=>"111000111",
  14508=>"000000111",
  14509=>"100110100",
  14510=>"000111001",
  14511=>"000101111",
  14512=>"111000000",
  14513=>"100101001",
  14514=>"011111111",
  14515=>"000000111",
  14516=>"101101100",
  14517=>"000000001",
  14518=>"000000100",
  14519=>"000000000",
  14520=>"111111111",
  14521=>"000000001",
  14522=>"110100000",
  14523=>"000000000",
  14524=>"111111111",
  14525=>"000001001",
  14526=>"111111010",
  14527=>"111101111",
  14528=>"001001111",
  14529=>"011111111",
  14530=>"111000100",
  14531=>"000111111",
  14532=>"101111111",
  14533=>"011011011",
  14534=>"100001011",
  14535=>"000000000",
  14536=>"110111111",
  14537=>"111111110",
  14538=>"000000000",
  14539=>"110111111",
  14540=>"000000111",
  14541=>"001001111",
  14542=>"000000000",
  14543=>"110111011",
  14544=>"111111111",
  14545=>"111111111",
  14546=>"111111111",
  14547=>"000000100",
  14548=>"111000000",
  14549=>"000001000",
  14550=>"000000000",
  14551=>"100000000",
  14552=>"000000000",
  14553=>"111111101",
  14554=>"111111111",
  14555=>"000000000",
  14556=>"000100100",
  14557=>"111110110",
  14558=>"000000000",
  14559=>"000101001",
  14560=>"000011001",
  14561=>"011010000",
  14562=>"000000111",
  14563=>"000000000",
  14564=>"111001000",
  14565=>"001101101",
  14566=>"001001001",
  14567=>"111111101",
  14568=>"000000000",
  14569=>"000001111",
  14570=>"111110110",
  14571=>"000000000",
  14572=>"111111111",
  14573=>"000000110",
  14574=>"111111000",
  14575=>"101000000",
  14576=>"111010000",
  14577=>"111111111",
  14578=>"000000000",
  14579=>"000101111",
  14580=>"000000000",
  14581=>"000100000",
  14582=>"100100111",
  14583=>"000000000",
  14584=>"000000100",
  14585=>"010000000",
  14586=>"001111010",
  14587=>"000111111",
  14588=>"100000001",
  14589=>"110110000",
  14590=>"001101111",
  14591=>"000111111",
  14592=>"010111000",
  14593=>"000000110",
  14594=>"000000000",
  14595=>"111110000",
  14596=>"110111000",
  14597=>"000111010",
  14598=>"000000111",
  14599=>"000001000",
  14600=>"001011100",
  14601=>"101000000",
  14602=>"000000000",
  14603=>"111111111",
  14604=>"001001000",
  14605=>"000110110",
  14606=>"111111011",
  14607=>"011001101",
  14608=>"111111101",
  14609=>"001111111",
  14610=>"011011011",
  14611=>"000000000",
  14612=>"110010000",
  14613=>"111011011",
  14614=>"111111111",
  14615=>"111111111",
  14616=>"111011111",
  14617=>"111000000",
  14618=>"000000100",
  14619=>"001000000",
  14620=>"000101001",
  14621=>"100000110",
  14622=>"111111110",
  14623=>"111000000",
  14624=>"000000000",
  14625=>"101100100",
  14626=>"111111111",
  14627=>"111111111",
  14628=>"110110110",
  14629=>"000000011",
  14630=>"000000000",
  14631=>"111000101",
  14632=>"111110000",
  14633=>"111111111",
  14634=>"000000111",
  14635=>"000011010",
  14636=>"000001101",
  14637=>"000000101",
  14638=>"000111000",
  14639=>"000000000",
  14640=>"000001001",
  14641=>"000000000",
  14642=>"110111111",
  14643=>"000000000",
  14644=>"111101001",
  14645=>"000000000",
  14646=>"000000000",
  14647=>"100111001",
  14648=>"000000000",
  14649=>"000000111",
  14650=>"111101111",
  14651=>"100111010",
  14652=>"011111111",
  14653=>"111111111",
  14654=>"011000000",
  14655=>"101100100",
  14656=>"100000011",
  14657=>"000011001",
  14658=>"110111111",
  14659=>"111111111",
  14660=>"001011111",
  14661=>"111111000",
  14662=>"000000000",
  14663=>"110111011",
  14664=>"000000000",
  14665=>"110000000",
  14666=>"011011110",
  14667=>"000000111",
  14668=>"000001000",
  14669=>"000000000",
  14670=>"000001011",
  14671=>"000100100",
  14672=>"000000100",
  14673=>"000001001",
  14674=>"111111111",
  14675=>"111000000",
  14676=>"001000000",
  14677=>"011010011",
  14678=>"100110111",
  14679=>"111111110",
  14680=>"000000100",
  14681=>"111111011",
  14682=>"100000010",
  14683=>"100111111",
  14684=>"000000000",
  14685=>"000000000",
  14686=>"111001001",
  14687=>"111111000",
  14688=>"111100111",
  14689=>"111111111",
  14690=>"110110100",
  14691=>"111111110",
  14692=>"000000110",
  14693=>"000001111",
  14694=>"111111111",
  14695=>"111111111",
  14696=>"000000100",
  14697=>"001111100",
  14698=>"001000101",
  14699=>"110110111",
  14700=>"111111001",
  14701=>"010111111",
  14702=>"111111111",
  14703=>"111111111",
  14704=>"000000000",
  14705=>"101000001",
  14706=>"011110010",
  14707=>"000001001",
  14708=>"111110111",
  14709=>"000111001",
  14710=>"111101001",
  14711=>"000000001",
  14712=>"000000101",
  14713=>"111011011",
  14714=>"000000000",
  14715=>"110111110",
  14716=>"010011011",
  14717=>"000010001",
  14718=>"111100001",
  14719=>"101100101",
  14720=>"001111010",
  14721=>"001101110",
  14722=>"110000010",
  14723=>"000000000",
  14724=>"011100000",
  14725=>"000000000",
  14726=>"110000000",
  14727=>"000000000",
  14728=>"000000000",
  14729=>"000110100",
  14730=>"111000100",
  14731=>"111100100",
  14732=>"111111111",
  14733=>"000110111",
  14734=>"111111100",
  14735=>"000000000",
  14736=>"000000000",
  14737=>"110110000",
  14738=>"000001101",
  14739=>"111100111",
  14740=>"000000000",
  14741=>"000000010",
  14742=>"000000101",
  14743=>"111011001",
  14744=>"000011001",
  14745=>"110110110",
  14746=>"000000000",
  14747=>"000110111",
  14748=>"000001111",
  14749=>"110011111",
  14750=>"110110110",
  14751=>"101111111",
  14752=>"111101001",
  14753=>"110010000",
  14754=>"001111111",
  14755=>"000000000",
  14756=>"000000000",
  14757=>"111101101",
  14758=>"001001001",
  14759=>"000000111",
  14760=>"000010110",
  14761=>"100000000",
  14762=>"000000000",
  14763=>"111111111",
  14764=>"000000010",
  14765=>"000010000",
  14766=>"111111111",
  14767=>"111100100",
  14768=>"111111111",
  14769=>"111111111",
  14770=>"111111001",
  14771=>"000000000",
  14772=>"000101000",
  14773=>"111111000",
  14774=>"101111111",
  14775=>"111111111",
  14776=>"000000000",
  14777=>"111011111",
  14778=>"000000010",
  14779=>"000000000",
  14780=>"010010000",
  14781=>"000101111",
  14782=>"000000000",
  14783=>"111111111",
  14784=>"101100000",
  14785=>"000000010",
  14786=>"000001111",
  14787=>"111110110",
  14788=>"000000000",
  14789=>"010010101",
  14790=>"101111001",
  14791=>"001111111",
  14792=>"000000000",
  14793=>"000010011",
  14794=>"001001000",
  14795=>"110110110",
  14796=>"000011111",
  14797=>"000111111",
  14798=>"110110000",
  14799=>"000001001",
  14800=>"101001000",
  14801=>"000000010",
  14802=>"111011111",
  14803=>"000110010",
  14804=>"000000000",
  14805=>"111111000",
  14806=>"000000111",
  14807=>"000000000",
  14808=>"001111111",
  14809=>"000000001",
  14810=>"000000010",
  14811=>"110101000",
  14812=>"110000000",
  14813=>"001011001",
  14814=>"111111100",
  14815=>"011010000",
  14816=>"011111111",
  14817=>"111100110",
  14818=>"000000000",
  14819=>"000100110",
  14820=>"111110000",
  14821=>"111000000",
  14822=>"000000000",
  14823=>"000000000",
  14824=>"000010110",
  14825=>"100000000",
  14826=>"111000111",
  14827=>"001000000",
  14828=>"111010110",
  14829=>"000100000",
  14830=>"000001111",
  14831=>"111111011",
  14832=>"001011011",
  14833=>"001000000",
  14834=>"011011000",
  14835=>"111101100",
  14836=>"000000111",
  14837=>"100100000",
  14838=>"011111111",
  14839=>"111101100",
  14840=>"111110110",
  14841=>"000100111",
  14842=>"011011111",
  14843=>"000001101",
  14844=>"111111000",
  14845=>"000011111",
  14846=>"110110110",
  14847=>"011111111",
  14848=>"000000000",
  14849=>"000000000",
  14850=>"111111111",
  14851=>"000000001",
  14852=>"000000001",
  14853=>"100000111",
  14854=>"011111111",
  14855=>"111000000",
  14856=>"101100111",
  14857=>"000000000",
  14858=>"000000001",
  14859=>"111000000",
  14860=>"100100100",
  14861=>"111111001",
  14862=>"111111010",
  14863=>"111111111",
  14864=>"000011000",
  14865=>"011111011",
  14866=>"010000000",
  14867=>"000000000",
  14868=>"111111100",
  14869=>"000100110",
  14870=>"000000000",
  14871=>"111111111",
  14872=>"100000010",
  14873=>"000010011",
  14874=>"001011111",
  14875=>"001011001",
  14876=>"111001000",
  14877=>"100100000",
  14878=>"111000000",
  14879=>"011111100",
  14880=>"100100000",
  14881=>"000000000",
  14882=>"110000100",
  14883=>"111111101",
  14884=>"000000111",
  14885=>"111111110",
  14886=>"000000111",
  14887=>"111111111",
  14888=>"000000111",
  14889=>"111111111",
  14890=>"011011111",
  14891=>"011011111",
  14892=>"010111111",
  14893=>"001101100",
  14894=>"000101111",
  14895=>"110010010",
  14896=>"110000111",
  14897=>"000001000",
  14898=>"000000000",
  14899=>"110110110",
  14900=>"111111001",
  14901=>"111000010",
  14902=>"010000011",
  14903=>"011011010",
  14904=>"111100111",
  14905=>"111000101",
  14906=>"010111111",
  14907=>"000000000",
  14908=>"100100100",
  14909=>"111000100",
  14910=>"000010011",
  14911=>"111100111",
  14912=>"000000100",
  14913=>"101001000",
  14914=>"000000000",
  14915=>"000000000",
  14916=>"110010010",
  14917=>"001011011",
  14918=>"000000100",
  14919=>"000000000",
  14920=>"000110110",
  14921=>"110111110",
  14922=>"011001101",
  14923=>"010001000",
  14924=>"111111111",
  14925=>"001101111",
  14926=>"110000011",
  14927=>"000000000",
  14928=>"111111101",
  14929=>"101011011",
  14930=>"000110000",
  14931=>"000000111",
  14932=>"011000011",
  14933=>"011111111",
  14934=>"010000101",
  14935=>"111111001",
  14936=>"110101011",
  14937=>"101000000",
  14938=>"111111111",
  14939=>"011001101",
  14940=>"011001000",
  14941=>"000000000",
  14942=>"000111111",
  14943=>"111101111",
  14944=>"111111111",
  14945=>"100110000",
  14946=>"000011010",
  14947=>"101000000",
  14948=>"100100110",
  14949=>"010001100",
  14950=>"111110111",
  14951=>"001101100",
  14952=>"111111000",
  14953=>"111111111",
  14954=>"000101111",
  14955=>"101111111",
  14956=>"000000000",
  14957=>"111100000",
  14958=>"000000000",
  14959=>"000000000",
  14960=>"000000000",
  14961=>"101001011",
  14962=>"011001001",
  14963=>"111111011",
  14964=>"011111110",
  14965=>"000000000",
  14966=>"000000111",
  14967=>"010000000",
  14968=>"111111111",
  14969=>"000111111",
  14970=>"111111111",
  14971=>"000000000",
  14972=>"110110010",
  14973=>"111111100",
  14974=>"010000000",
  14975=>"000000000",
  14976=>"111101100",
  14977=>"111111111",
  14978=>"111111111",
  14979=>"000001001",
  14980=>"000000000",
  14981=>"100000000",
  14982=>"110110000",
  14983=>"101011110",
  14984=>"111111111",
  14985=>"011011001",
  14986=>"111111100",
  14987=>"100100111",
  14988=>"111101101",
  14989=>"000000000",
  14990=>"101001000",
  14991=>"110000000",
  14992=>"111100000",
  14993=>"101101111",
  14994=>"110100000",
  14995=>"001111111",
  14996=>"111111111",
  14997=>"010010011",
  14998=>"001111111",
  14999=>"100100100",
  15000=>"110000001",
  15001=>"111111000",
  15002=>"000101000",
  15003=>"101001000",
  15004=>"111000000",
  15005=>"000000001",
  15006=>"110110111",
  15007=>"111111111",
  15008=>"000100110",
  15009=>"000000000",
  15010=>"111111010",
  15011=>"000000000",
  15012=>"000000000",
  15013=>"000000000",
  15014=>"111111000",
  15015=>"011111111",
  15016=>"011000110",
  15017=>"000010000",
  15018=>"110100110",
  15019=>"111111111",
  15020=>"111111110",
  15021=>"000000000",
  15022=>"000000000",
  15023=>"000101000",
  15024=>"111111111",
  15025=>"010000001",
  15026=>"111111110",
  15027=>"101000100",
  15028=>"111011111",
  15029=>"000000000",
  15030=>"110100111",
  15031=>"000000100",
  15032=>"001011001",
  15033=>"111000000",
  15034=>"010100000",
  15035=>"110101100",
  15036=>"000100110",
  15037=>"111000000",
  15038=>"011000000",
  15039=>"101111111",
  15040=>"110110011",
  15041=>"000000000",
  15042=>"111111111",
  15043=>"111111110",
  15044=>"000110110",
  15045=>"000000000",
  15046=>"111111000",
  15047=>"011000000",
  15048=>"000111111",
  15049=>"000000000",
  15050=>"000000000",
  15051=>"100000100",
  15052=>"011111110",
  15053=>"001111111",
  15054=>"001001000",
  15055=>"011101100",
  15056=>"101111111",
  15057=>"110110111",
  15058=>"000000010",
  15059=>"000000100",
  15060=>"011011111",
  15061=>"111110011",
  15062=>"000000000",
  15063=>"111111111",
  15064=>"111010111",
  15065=>"101111111",
  15066=>"111111111",
  15067=>"011110110",
  15068=>"110110000",
  15069=>"001111111",
  15070=>"111000000",
  15071=>"110010100",
  15072=>"111111111",
  15073=>"100001111",
  15074=>"100111111",
  15075=>"111111100",
  15076=>"011111111",
  15077=>"110000010",
  15078=>"001001000",
  15079=>"000000100",
  15080=>"111111111",
  15081=>"000000000",
  15082=>"000000111",
  15083=>"110011000",
  15084=>"011010000",
  15085=>"001000100",
  15086=>"001000100",
  15087=>"100100100",
  15088=>"001001111",
  15089=>"001100111",
  15090=>"110110000",
  15091=>"110100101",
  15092=>"011011111",
  15093=>"011011111",
  15094=>"110110011",
  15095=>"100000000",
  15096=>"000111111",
  15097=>"000111111",
  15098=>"000001011",
  15099=>"111111111",
  15100=>"011111111",
  15101=>"000000011",
  15102=>"110111011",
  15103=>"000110100",
  15104=>"000000100",
  15105=>"110000000",
  15106=>"011011011",
  15107=>"000000100",
  15108=>"001111110",
  15109=>"111111111",
  15110=>"011111001",
  15111=>"000100100",
  15112=>"000000000",
  15113=>"101101101",
  15114=>"011011111",
  15115=>"100101101",
  15116=>"000000000",
  15117=>"000000000",
  15118=>"000000111",
  15119=>"101001000",
  15120=>"000001101",
  15121=>"111111111",
  15122=>"111000000",
  15123=>"100000000",
  15124=>"000000001",
  15125=>"000001001",
  15126=>"010011011",
  15127=>"011010010",
  15128=>"111111111",
  15129=>"001100111",
  15130=>"000000111",
  15131=>"000011011",
  15132=>"110000010",
  15133=>"001110110",
  15134=>"000000000",
  15135=>"010000100",
  15136=>"010000111",
  15137=>"111111001",
  15138=>"000000010",
  15139=>"000000000",
  15140=>"000000000",
  15141=>"000000000",
  15142=>"000000000",
  15143=>"000001001",
  15144=>"000110111",
  15145=>"011011000",
  15146=>"111111101",
  15147=>"100000111",
  15148=>"000011111",
  15149=>"000100010",
  15150=>"000000000",
  15151=>"011111111",
  15152=>"011011111",
  15153=>"110000100",
  15154=>"011111111",
  15155=>"001111111",
  15156=>"111111111",
  15157=>"001000000",
  15158=>"111111100",
  15159=>"010000000",
  15160=>"111001000",
  15161=>"111111111",
  15162=>"110010011",
  15163=>"111001111",
  15164=>"111010000",
  15165=>"111111111",
  15166=>"000000000",
  15167=>"111011000",
  15168=>"000000001",
  15169=>"010000111",
  15170=>"000000100",
  15171=>"111111111",
  15172=>"001001000",
  15173=>"010000000",
  15174=>"011011011",
  15175=>"000000000",
  15176=>"000000000",
  15177=>"001111111",
  15178=>"100100000",
  15179=>"111110110",
  15180=>"111011000",
  15181=>"111100010",
  15182=>"000000100",
  15183=>"000110110",
  15184=>"111111111",
  15185=>"001101111",
  15186=>"010011111",
  15187=>"110110110",
  15188=>"000110100",
  15189=>"000011010",
  15190=>"111101111",
  15191=>"101111111",
  15192=>"000111100",
  15193=>"100110000",
  15194=>"000000111",
  15195=>"110100000",
  15196=>"101000000",
  15197=>"011000000",
  15198=>"110110111",
  15199=>"000000100",
  15200=>"000000000",
  15201=>"111011001",
  15202=>"000000011",
  15203=>"111111101",
  15204=>"110010010",
  15205=>"000000011",
  15206=>"000000000",
  15207=>"000000000",
  15208=>"100000001",
  15209=>"101101000",
  15210=>"000101111",
  15211=>"011011111",
  15212=>"101100111",
  15213=>"111010000",
  15214=>"000000000",
  15215=>"110110000",
  15216=>"010000000",
  15217=>"111111111",
  15218=>"000000000",
  15219=>"011000000",
  15220=>"000000000",
  15221=>"000000000",
  15222=>"001000000",
  15223=>"001111111",
  15224=>"000100111",
  15225=>"001100110",
  15226=>"111111111",
  15227=>"000000000",
  15228=>"011011000",
  15229=>"100000000",
  15230=>"000001001",
  15231=>"111111111",
  15232=>"010110000",
  15233=>"111100000",
  15234=>"000000000",
  15235=>"001011111",
  15236=>"000001000",
  15237=>"111111111",
  15238=>"111111101",
  15239=>"000000000",
  15240=>"110111111",
  15241=>"111111111",
  15242=>"100100111",
  15243=>"101101000",
  15244=>"111111101",
  15245=>"011011001",
  15246=>"000001111",
  15247=>"000011001",
  15248=>"000000000",
  15249=>"100100000",
  15250=>"111110110",
  15251=>"000000000",
  15252=>"000000000",
  15253=>"001001001",
  15254=>"110000000",
  15255=>"011011111",
  15256=>"111100000",
  15257=>"011000110",
  15258=>"111110110",
  15259=>"000001011",
  15260=>"011111111",
  15261=>"111111111",
  15262=>"011011001",
  15263=>"001011011",
  15264=>"111111111",
  15265=>"010011001",
  15266=>"010000000",
  15267=>"001000000",
  15268=>"101101000",
  15269=>"111111111",
  15270=>"110010000",
  15271=>"111111111",
  15272=>"000000011",
  15273=>"000000110",
  15274=>"000000000",
  15275=>"111011011",
  15276=>"000000011",
  15277=>"011001100",
  15278=>"000000110",
  15279=>"111111111",
  15280=>"000000000",
  15281=>"000111111",
  15282=>"111010001",
  15283=>"000000000",
  15284=>"011000000",
  15285=>"101111111",
  15286=>"100100000",
  15287=>"000110111",
  15288=>"010000110",
  15289=>"110110111",
  15290=>"001001011",
  15291=>"000111110",
  15292=>"000000000",
  15293=>"110110110",
  15294=>"111111111",
  15295=>"010011000",
  15296=>"000000000",
  15297=>"000100000",
  15298=>"111111011",
  15299=>"000000000",
  15300=>"100000111",
  15301=>"110110000",
  15302=>"100001001",
  15303=>"101000000",
  15304=>"011000000",
  15305=>"000000000",
  15306=>"000000000",
  15307=>"110111111",
  15308=>"000111000",
  15309=>"110111101",
  15310=>"110110000",
  15311=>"000000000",
  15312=>"100111111",
  15313=>"111111111",
  15314=>"001100000",
  15315=>"000000000",
  15316=>"000010000",
  15317=>"111111111",
  15318=>"111001111",
  15319=>"011001000",
  15320=>"011000111",
  15321=>"111000001",
  15322=>"000000100",
  15323=>"000000110",
  15324=>"001000000",
  15325=>"011000000",
  15326=>"000000000",
  15327=>"000001011",
  15328=>"111111011",
  15329=>"000000000",
  15330=>"000000000",
  15331=>"000001000",
  15332=>"110010000",
  15333=>"000000000",
  15334=>"101111111",
  15335=>"100110110",
  15336=>"111111100",
  15337=>"011101111",
  15338=>"011111110",
  15339=>"000000111",
  15340=>"110000000",
  15341=>"011111111",
  15342=>"111111000",
  15343=>"111011001",
  15344=>"011111111",
  15345=>"000000001",
  15346=>"001010111",
  15347=>"101001111",
  15348=>"111001000",
  15349=>"001001000",
  15350=>"111111111",
  15351=>"000100000",
  15352=>"100100100",
  15353=>"011011111",
  15354=>"100110110",
  15355=>"100111111",
  15356=>"001001000",
  15357=>"110110000",
  15358=>"010000000",
  15359=>"111101111",
  15360=>"000000000",
  15361=>"111110000",
  15362=>"100000111",
  15363=>"000000000",
  15364=>"111010010",
  15365=>"011111111",
  15366=>"011111111",
  15367=>"111111111",
  15368=>"011000111",
  15369=>"111111111",
  15370=>"000000000",
  15371=>"000000001",
  15372=>"110111111",
  15373=>"111111111",
  15374=>"000001000",
  15375=>"111111011",
  15376=>"111111001",
  15377=>"000011011",
  15378=>"011011000",
  15379=>"011000000",
  15380=>"111111111",
  15381=>"111111111",
  15382=>"000000000",
  15383=>"110100111",
  15384=>"100100000",
  15385=>"100000000",
  15386=>"111111111",
  15387=>"100100000",
  15388=>"001111111",
  15389=>"110111111",
  15390=>"001001000",
  15391=>"100000000",
  15392=>"010111111",
  15393=>"011000000",
  15394=>"000000000",
  15395=>"111111111",
  15396=>"011000000",
  15397=>"000100000",
  15398=>"000000000",
  15399=>"010000000",
  15400=>"000000000",
  15401=>"000000001",
  15402=>"000000000",
  15403=>"111111000",
  15404=>"111111101",
  15405=>"100100100",
  15406=>"000000110",
  15407=>"101100100",
  15408=>"111111111",
  15409=>"000000000",
  15410=>"011101111",
  15411=>"100111111",
  15412=>"000101101",
  15413=>"111111111",
  15414=>"000000000",
  15415=>"110111011",
  15416=>"111111111",
  15417=>"110110000",
  15418=>"111111111",
  15419=>"000000000",
  15420=>"001001111",
  15421=>"000000000",
  15422=>"101011000",
  15423=>"111111111",
  15424=>"001000011",
  15425=>"111111111",
  15426=>"000101111",
  15427=>"111000111",
  15428=>"001000101",
  15429=>"000000111",
  15430=>"110101000",
  15431=>"000001111",
  15432=>"111101111",
  15433=>"000000000",
  15434=>"000000000",
  15435=>"111010001",
  15436=>"001000111",
  15437=>"100110000",
  15438=>"000110011",
  15439=>"000000111",
  15440=>"110111000",
  15441=>"111111001",
  15442=>"000000100",
  15443=>"000000000",
  15444=>"001001001",
  15445=>"000000000",
  15446=>"010000000",
  15447=>"000000000",
  15448=>"100100010",
  15449=>"111111111",
  15450=>"010011010",
  15451=>"011111111",
  15452=>"011001001",
  15453=>"000000000",
  15454=>"000000000",
  15455=>"111111001",
  15456=>"001000000",
  15457=>"001001000",
  15458=>"111111011",
  15459=>"000000000",
  15460=>"000000000",
  15461=>"111110000",
  15462=>"100000000",
  15463=>"110111111",
  15464=>"000000000",
  15465=>"100000000",
  15466=>"011011010",
  15467=>"000000000",
  15468=>"111101000",
  15469=>"111110000",
  15470=>"011000001",
  15471=>"000100100",
  15472=>"000000111",
  15473=>"111011001",
  15474=>"010110000",
  15475=>"100000000",
  15476=>"010000000",
  15477=>"111010111",
  15478=>"000000000",
  15479=>"000000000",
  15480=>"000000000",
  15481=>"000000000",
  15482=>"001001001",
  15483=>"000001001",
  15484=>"100100111",
  15485=>"011001000",
  15486=>"111111111",
  15487=>"000010000",
  15488=>"000000000",
  15489=>"111000000",
  15490=>"110110111",
  15491=>"000000000",
  15492=>"111111111",
  15493=>"001000111",
  15494=>"111111110",
  15495=>"111111000",
  15496=>"111111111",
  15497=>"000000001",
  15498=>"001000000",
  15499=>"111011100",
  15500=>"000000000",
  15501=>"111011111",
  15502=>"001001001",
  15503=>"000011011",
  15504=>"000101111",
  15505=>"011011011",
  15506=>"110111111",
  15507=>"000011111",
  15508=>"111111111",
  15509=>"111111111",
  15510=>"000000100",
  15511=>"111111100",
  15512=>"001000000",
  15513=>"000000001",
  15514=>"111111111",
  15515=>"000000000",
  15516=>"000001111",
  15517=>"110110111",
  15518=>"111111000",
  15519=>"011111011",
  15520=>"001111111",
  15521=>"011111100",
  15522=>"000000000",
  15523=>"011111100",
  15524=>"110010010",
  15525=>"000100111",
  15526=>"000000000",
  15527=>"111111110",
  15528=>"000000000",
  15529=>"000000001",
  15530=>"111000000",
  15531=>"111111111",
  15532=>"111111111",
  15533=>"110011111",
  15534=>"111111111",
  15535=>"000010010",
  15536=>"000000000",
  15537=>"110111011",
  15538=>"011011000",
  15539=>"111111111",
  15540=>"011111111",
  15541=>"010000001",
  15542=>"000000000",
  15543=>"111111000",
  15544=>"000000000",
  15545=>"011001111",
  15546=>"000000001",
  15547=>"011001001",
  15548=>"111000000",
  15549=>"111000101",
  15550=>"000000000",
  15551=>"111001001",
  15552=>"111111011",
  15553=>"011111011",
  15554=>"011111110",
  15555=>"000000000",
  15556=>"111011001",
  15557=>"000000000",
  15558=>"010000001",
  15559=>"111111010",
  15560=>"000111111",
  15561=>"000000100",
  15562=>"011010000",
  15563=>"011111111",
  15564=>"100000101",
  15565=>"000100100",
  15566=>"101111111",
  15567=>"010000000",
  15568=>"010000000",
  15569=>"001111111",
  15570=>"111111111",
  15571=>"000101101",
  15572=>"100000000",
  15573=>"000001001",
  15574=>"000000000",
  15575=>"111111111",
  15576=>"111111000",
  15577=>"000000000",
  15578=>"000000000",
  15579=>"000000111",
  15580=>"111111010",
  15581=>"111111111",
  15582=>"000000000",
  15583=>"111111100",
  15584=>"001111000",
  15585=>"000000000",
  15586=>"000100000",
  15587=>"111111111",
  15588=>"111110000",
  15589=>"011010000",
  15590=>"000100111",
  15591=>"001000000",
  15592=>"000000000",
  15593=>"111111111",
  15594=>"111111111",
  15595=>"000000100",
  15596=>"000000000",
  15597=>"000000000",
  15598=>"000000110",
  15599=>"000110000",
  15600=>"110000000",
  15601=>"111111111",
  15602=>"111000100",
  15603=>"000010111",
  15604=>"000100111",
  15605=>"111100110",
  15606=>"110110001",
  15607=>"111111111",
  15608=>"111111111",
  15609=>"000000000",
  15610=>"111011011",
  15611=>"000000000",
  15612=>"000000001",
  15613=>"111111111",
  15614=>"111100110",
  15615=>"000000000",
  15616=>"011000000",
  15617=>"110110000",
  15618=>"111111111",
  15619=>"001001111",
  15620=>"000000000",
  15621=>"001001000",
  15622=>"111000000",
  15623=>"111111000",
  15624=>"001011000",
  15625=>"111111111",
  15626=>"111111111",
  15627=>"101111111",
  15628=>"111011111",
  15629=>"110000000",
  15630=>"011011000",
  15631=>"100000000",
  15632=>"111111110",
  15633=>"010010111",
  15634=>"111111111",
  15635=>"001001101",
  15636=>"111111001",
  15637=>"111111111",
  15638=>"111011011",
  15639=>"001000111",
  15640=>"111011011",
  15641=>"000000010",
  15642=>"110011000",
  15643=>"000000000",
  15644=>"110100100",
  15645=>"100100000",
  15646=>"000000000",
  15647=>"111111111",
  15648=>"011111111",
  15649=>"000001011",
  15650=>"111111111",
  15651=>"000000111",
  15652=>"111000000",
  15653=>"000011110",
  15654=>"100100110",
  15655=>"110010000",
  15656=>"011110110",
  15657=>"111111111",
  15658=>"111111111",
  15659=>"111111111",
  15660=>"101001111",
  15661=>"110111111",
  15662=>"000000000",
  15663=>"111111111",
  15664=>"000000000",
  15665=>"001000000",
  15666=>"000111111",
  15667=>"111111111",
  15668=>"000000000",
  15669=>"000000100",
  15670=>"000000000",
  15671=>"111111111",
  15672=>"000000000",
  15673=>"111111111",
  15674=>"000000000",
  15675=>"110000000",
  15676=>"000000000",
  15677=>"000000000",
  15678=>"111111100",
  15679=>"001000000",
  15680=>"000011111",
  15681=>"000000000",
  15682=>"111011000",
  15683=>"001000000",
  15684=>"111111111",
  15685=>"010000101",
  15686=>"000100111",
  15687=>"000000000",
  15688=>"011000000",
  15689=>"110111111",
  15690=>"111110110",
  15691=>"000000100",
  15692=>"001000000",
  15693=>"111101001",
  15694=>"000000001",
  15695=>"001001001",
  15696=>"000001001",
  15697=>"011100110",
  15698=>"000001011",
  15699=>"000110111",
  15700=>"001000000",
  15701=>"001000000",
  15702=>"111001111",
  15703=>"111111111",
  15704=>"000000000",
  15705=>"111111111",
  15706=>"000111111",
  15707=>"111111111",
  15708=>"000000000",
  15709=>"000000011",
  15710=>"111110111",
  15711=>"000000000",
  15712=>"110111100",
  15713=>"111111111",
  15714=>"110010000",
  15715=>"000000000",
  15716=>"000000001",
  15717=>"000010000",
  15718=>"100100100",
  15719=>"111111111",
  15720=>"000000001",
  15721=>"000000000",
  15722=>"100100111",
  15723=>"111110010",
  15724=>"000101000",
  15725=>"010000111",
  15726=>"111111111",
  15727=>"001000000",
  15728=>"011011001",
  15729=>"111111111",
  15730=>"001000001",
  15731=>"111111100",
  15732=>"000001000",
  15733=>"000000000",
  15734=>"010011111",
  15735=>"000000000",
  15736=>"111101111",
  15737=>"000000000",
  15738=>"111001001",
  15739=>"000111110",
  15740=>"110000100",
  15741=>"000000000",
  15742=>"000000000",
  15743=>"000000000",
  15744=>"111111001",
  15745=>"101111111",
  15746=>"100000001",
  15747=>"111111011",
  15748=>"000000111",
  15749=>"000000111",
  15750=>"110110000",
  15751=>"111111111",
  15752=>"100000000",
  15753=>"100111111",
  15754=>"001111011",
  15755=>"000001000",
  15756=>"111111111",
  15757=>"101110110",
  15758=>"000000000",
  15759=>"000010000",
  15760=>"000000100",
  15761=>"111111011",
  15762=>"000010000",
  15763=>"011001001",
  15764=>"110000000",
  15765=>"000000000",
  15766=>"001000001",
  15767=>"100000001",
  15768=>"001101111",
  15769=>"011001011",
  15770=>"000000000",
  15771=>"000111111",
  15772=>"000000000",
  15773=>"110001000",
  15774=>"010010001",
  15775=>"000000000",
  15776=>"011111111",
  15777=>"111111111",
  15778=>"000001001",
  15779=>"000011111",
  15780=>"000000100",
  15781=>"000000000",
  15782=>"000000000",
  15783=>"111111111",
  15784=>"100110000",
  15785=>"111011110",
  15786=>"111010110",
  15787=>"111111111",
  15788=>"000000000",
  15789=>"001100100",
  15790=>"100110111",
  15791=>"111011011",
  15792=>"100000110",
  15793=>"000010110",
  15794=>"111001000",
  15795=>"000000000",
  15796=>"000100110",
  15797=>"000000000",
  15798=>"101111111",
  15799=>"000000000",
  15800=>"000000000",
  15801=>"111111111",
  15802=>"000001100",
  15803=>"001001001",
  15804=>"000000111",
  15805=>"111111111",
  15806=>"001000110",
  15807=>"110000000",
  15808=>"011000101",
  15809=>"111111000",
  15810=>"111111001",
  15811=>"000000000",
  15812=>"000000101",
  15813=>"111111111",
  15814=>"111111111",
  15815=>"110111111",
  15816=>"011001001",
  15817=>"011111010",
  15818=>"001011111",
  15819=>"000011111",
  15820=>"000000000",
  15821=>"000000000",
  15822=>"001011010",
  15823=>"110100110",
  15824=>"000010010",
  15825=>"000011111",
  15826=>"000000110",
  15827=>"000000000",
  15828=>"111000100",
  15829=>"111111110",
  15830=>"000110011",
  15831=>"000000010",
  15832=>"000000000",
  15833=>"110110001",
  15834=>"010111000",
  15835=>"001000100",
  15836=>"000001001",
  15837=>"111111111",
  15838=>"111111100",
  15839=>"111111111",
  15840=>"101100111",
  15841=>"011011000",
  15842=>"000000000",
  15843=>"111111111",
  15844=>"011000000",
  15845=>"111111101",
  15846=>"110010011",
  15847=>"000100100",
  15848=>"111111111",
  15849=>"011001011",
  15850=>"111111110",
  15851=>"111001001",
  15852=>"000000111",
  15853=>"000000000",
  15854=>"111111111",
  15855=>"111111001",
  15856=>"111111111",
  15857=>"001000000",
  15858=>"011011110",
  15859=>"000000001",
  15860=>"011011110",
  15861=>"000000000",
  15862=>"000000000",
  15863=>"100100101",
  15864=>"000000000",
  15865=>"000010011",
  15866=>"000000000",
  15867=>"000000000",
  15868=>"000011010",
  15869=>"110110110",
  15870=>"111000001",
  15871=>"001000110",
  15872=>"110100100",
  15873=>"011111111",
  15874=>"000001001",
  15875=>"111000000",
  15876=>"000000110",
  15877=>"111000000",
  15878=>"000000000",
  15879=>"111111111",
  15880=>"000000100",
  15881=>"000000010",
  15882=>"000000000",
  15883=>"001001001",
  15884=>"110000001",
  15885=>"111111000",
  15886=>"111111100",
  15887=>"111101111",
  15888=>"011011111",
  15889=>"111111111",
  15890=>"110100100",
  15891=>"000000000",
  15892=>"000000000",
  15893=>"000000000",
  15894=>"000000000",
  15895=>"000000000",
  15896=>"000000111",
  15897=>"111111111",
  15898=>"001000001",
  15899=>"111111111",
  15900=>"000000111",
  15901=>"000000000",
  15902=>"111111111",
  15903=>"110111111",
  15904=>"101100100",
  15905=>"100110110",
  15906=>"111111111",
  15907=>"110111111",
  15908=>"000000101",
  15909=>"111111100",
  15910=>"000001011",
  15911=>"000000111",
  15912=>"110100100",
  15913=>"000000000",
  15914=>"000000000",
  15915=>"110000100",
  15916=>"111111111",
  15917=>"111101001",
  15918=>"111111111",
  15919=>"111111111",
  15920=>"100110111",
  15921=>"111001000",
  15922=>"000000000",
  15923=>"011011111",
  15924=>"000111111",
  15925=>"111111111",
  15926=>"000000000",
  15927=>"000011110",
  15928=>"000000000",
  15929=>"111111111",
  15930=>"000000000",
  15931=>"000000111",
  15932=>"000000001",
  15933=>"111111000",
  15934=>"000011010",
  15935=>"000000000",
  15936=>"111111111",
  15937=>"000000000",
  15938=>"111000000",
  15939=>"000000000",
  15940=>"010011011",
  15941=>"000000000",
  15942=>"100110111",
  15943=>"001101101",
  15944=>"000011011",
  15945=>"000000011",
  15946=>"110110111",
  15947=>"000101101",
  15948=>"110000000",
  15949=>"111110111",
  15950=>"000000000",
  15951=>"111001101",
  15952=>"000000000",
  15953=>"101000000",
  15954=>"110100110",
  15955=>"110111000",
  15956=>"000000000",
  15957=>"000100100",
  15958=>"000001001",
  15959=>"100000101",
  15960=>"000000100",
  15961=>"000000000",
  15962=>"111111111",
  15963=>"011111111",
  15964=>"111111111",
  15965=>"111111111",
  15966=>"000000111",
  15967=>"001011101",
  15968=>"001111111",
  15969=>"000000000",
  15970=>"000000001",
  15971=>"000000000",
  15972=>"101000000",
  15973=>"000000000",
  15974=>"011111111",
  15975=>"000001111",
  15976=>"000100111",
  15977=>"000000000",
  15978=>"000000000",
  15979=>"000111111",
  15980=>"000000000",
  15981=>"111111000",
  15982=>"111111111",
  15983=>"101100111",
  15984=>"011000110",
  15985=>"111101111",
  15986=>"111111111",
  15987=>"111100111",
  15988=>"000000000",
  15989=>"101101111",
  15990=>"000000011",
  15991=>"111111000",
  15992=>"000000001",
  15993=>"111111100",
  15994=>"000001111",
  15995=>"000000111",
  15996=>"111111110",
  15997=>"111111111",
  15998=>"000100100",
  15999=>"000000000",
  16000=>"000000000",
  16001=>"000000010",
  16002=>"011000000",
  16003=>"111111110",
  16004=>"001001001",
  16005=>"111100100",
  16006=>"000000000",
  16007=>"000000111",
  16008=>"011111111",
  16009=>"000000000",
  16010=>"000000000",
  16011=>"100000111",
  16012=>"000111001",
  16013=>"000000000",
  16014=>"000111000",
  16015=>"000000011",
  16016=>"111111111",
  16017=>"011011001",
  16018=>"001000000",
  16019=>"111111100",
  16020=>"111111111",
  16021=>"000010111",
  16022=>"000000100",
  16023=>"000000101",
  16024=>"111111111",
  16025=>"111111111",
  16026=>"111111111",
  16027=>"000000000",
  16028=>"110110110",
  16029=>"001000101",
  16030=>"000000000",
  16031=>"000000000",
  16032=>"001000100",
  16033=>"000000000",
  16034=>"000000000",
  16035=>"000000000",
  16036=>"001000111",
  16037=>"010111111",
  16038=>"000000001",
  16039=>"111111111",
  16040=>"100111100",
  16041=>"111001111",
  16042=>"111111100",
  16043=>"111111111",
  16044=>"001001000",
  16045=>"000000100",
  16046=>"101111100",
  16047=>"000001001",
  16048=>"010011000",
  16049=>"011011011",
  16050=>"111111111",
  16051=>"001011111",
  16052=>"100111110",
  16053=>"100000000",
  16054=>"111111111",
  16055=>"111110111",
  16056=>"111100101",
  16057=>"010010110",
  16058=>"110100000",
  16059=>"000000000",
  16060=>"000000110",
  16061=>"111111111",
  16062=>"000000000",
  16063=>"001001001",
  16064=>"000000000",
  16065=>"000000000",
  16066=>"111111111",
  16067=>"111111111",
  16068=>"000000110",
  16069=>"111111111",
  16070=>"000000011",
  16071=>"000000000",
  16072=>"011010010",
  16073=>"000110000",
  16074=>"000000000",
  16075=>"111100101",
  16076=>"101111111",
  16077=>"000111111",
  16078=>"010000010",
  16079=>"000000000",
  16080=>"111111001",
  16081=>"000000000",
  16082=>"000000000",
  16083=>"111111100",
  16084=>"110110111",
  16085=>"110110010",
  16086=>"001000000",
  16087=>"100110000",
  16088=>"000000010",
  16089=>"111111101",
  16090=>"000100111",
  16091=>"000000110",
  16092=>"100000000",
  16093=>"000000000",
  16094=>"011001001",
  16095=>"000001000",
  16096=>"000000000",
  16097=>"000000110",
  16098=>"111111111",
  16099=>"000000000",
  16100=>"101111101",
  16101=>"111110110",
  16102=>"110110111",
  16103=>"000000000",
  16104=>"000000001",
  16105=>"111111111",
  16106=>"111110000",
  16107=>"101111111",
  16108=>"111111111",
  16109=>"000010010",
  16110=>"000010001",
  16111=>"000000111",
  16112=>"101111111",
  16113=>"111111100",
  16114=>"111100101",
  16115=>"101100000",
  16116=>"111111111",
  16117=>"000100110",
  16118=>"101001000",
  16119=>"001101111",
  16120=>"111111111",
  16121=>"000000000",
  16122=>"000000000",
  16123=>"000000000",
  16124=>"111111111",
  16125=>"010000110",
  16126=>"110000000",
  16127=>"001111111",
  16128=>"000000000",
  16129=>"000000000",
  16130=>"111111111",
  16131=>"011111101",
  16132=>"000000000",
  16133=>"000000000",
  16134=>"000111111",
  16135=>"111011100",
  16136=>"111111000",
  16137=>"010000000",
  16138=>"100110111",
  16139=>"000100000",
  16140=>"111100000",
  16141=>"000000011",
  16142=>"000000100",
  16143=>"000000000",
  16144=>"000111111",
  16145=>"111111001",
  16146=>"000000000",
  16147=>"000000000",
  16148=>"000000000",
  16149=>"111111111",
  16150=>"111111111",
  16151=>"111111000",
  16152=>"111101001",
  16153=>"000000000",
  16154=>"111001000",
  16155=>"111111011",
  16156=>"000000011",
  16157=>"000100111",
  16158=>"000110100",
  16159=>"010100101",
  16160=>"011011000",
  16161=>"000001111",
  16162=>"000000000",
  16163=>"111111101",
  16164=>"101000000",
  16165=>"111111001",
  16166=>"000100111",
  16167=>"000000101",
  16168=>"000000000",
  16169=>"000000000",
  16170=>"000101001",
  16171=>"111111110",
  16172=>"011111111",
  16173=>"000000100",
  16174=>"000000000",
  16175=>"110000000",
  16176=>"001000000",
  16177=>"000000111",
  16178=>"111111111",
  16179=>"111100111",
  16180=>"000000000",
  16181=>"011011111",
  16182=>"111111111",
  16183=>"000100100",
  16184=>"001000000",
  16185=>"111001111",
  16186=>"000110111",
  16187=>"111111111",
  16188=>"111111111",
  16189=>"000000110",
  16190=>"000000110",
  16191=>"000000000",
  16192=>"000000000",
  16193=>"111111110",
  16194=>"000000000",
  16195=>"100000000",
  16196=>"001000000",
  16197=>"111011111",
  16198=>"000000000",
  16199=>"101101000",
  16200=>"000000011",
  16201=>"001000000",
  16202=>"011000000",
  16203=>"000000000",
  16204=>"100100110",
  16205=>"111111110",
  16206=>"111111111",
  16207=>"000001001",
  16208=>"111111000",
  16209=>"110111111",
  16210=>"111111111",
  16211=>"000000000",
  16212=>"000000110",
  16213=>"001001011",
  16214=>"001011011",
  16215=>"111011011",
  16216=>"001000000",
  16217=>"111111111",
  16218=>"111111100",
  16219=>"111111111",
  16220=>"000000111",
  16221=>"000000111",
  16222=>"111111111",
  16223=>"111011011",
  16224=>"011111111",
  16225=>"111101101",
  16226=>"111111111",
  16227=>"111111111",
  16228=>"111111111",
  16229=>"111000000",
  16230=>"000000000",
  16231=>"001001001",
  16232=>"000001000",
  16233=>"100111111",
  16234=>"000000000",
  16235=>"000000000",
  16236=>"000100001",
  16237=>"111111111",
  16238=>"110110110",
  16239=>"010001000",
  16240=>"000000011",
  16241=>"000000000",
  16242=>"000111111",
  16243=>"110000111",
  16244=>"000000000",
  16245=>"111111111",
  16246=>"000000000",
  16247=>"111111110",
  16248=>"000000111",
  16249=>"111111011",
  16250=>"000000000",
  16251=>"100110100",
  16252=>"000000000",
  16253=>"011111101",
  16254=>"100100111",
  16255=>"000000000",
  16256=>"000000000",
  16257=>"000011101",
  16258=>"001011000",
  16259=>"000000000",
  16260=>"000001011",
  16261=>"000000000",
  16262=>"000000000",
  16263=>"001000000",
  16264=>"011000001",
  16265=>"011011101",
  16266=>"111011000",
  16267=>"000000000",
  16268=>"001111111",
  16269=>"111111100",
  16270=>"111111111",
  16271=>"000000000",
  16272=>"000000000",
  16273=>"000000000",
  16274=>"111111111",
  16275=>"111111111",
  16276=>"111111111",
  16277=>"000000010",
  16278=>"100101111",
  16279=>"111111110",
  16280=>"111111111",
  16281=>"100100100",
  16282=>"000101101",
  16283=>"110000000",
  16284=>"000100000",
  16285=>"000000000",
  16286=>"110111001",
  16287=>"000000000",
  16288=>"001101111",
  16289=>"111111111",
  16290=>"000011111",
  16291=>"001000011",
  16292=>"001001101",
  16293=>"011010010",
  16294=>"000000011",
  16295=>"111111111",
  16296=>"001011111",
  16297=>"001001000",
  16298=>"000000000",
  16299=>"010001111",
  16300=>"000000000",
  16301=>"001011111",
  16302=>"000000000",
  16303=>"111111111",
  16304=>"111111000",
  16305=>"000000000",
  16306=>"001001000",
  16307=>"000000000",
  16308=>"111000111",
  16309=>"000000110",
  16310=>"000010000",
  16311=>"000000000",
  16312=>"000000000",
  16313=>"000000000",
  16314=>"001001001",
  16315=>"000000000",
  16316=>"111111111",
  16317=>"100100100",
  16318=>"011001000",
  16319=>"111000010",
  16320=>"001000001",
  16321=>"000000111",
  16322=>"111111111",
  16323=>"000000001",
  16324=>"100000000",
  16325=>"110111111",
  16326=>"101001001",
  16327=>"000000000",
  16328=>"110111100",
  16329=>"010000000",
  16330=>"101000001",
  16331=>"010111111",
  16332=>"111000000",
  16333=>"000001000",
  16334=>"000000000",
  16335=>"111111111",
  16336=>"110111000",
  16337=>"011001111",
  16338=>"000001111",
  16339=>"000111111",
  16340=>"000101111",
  16341=>"000000000",
  16342=>"011011111",
  16343=>"000000000",
  16344=>"100000000",
  16345=>"100000000",
  16346=>"111111111",
  16347=>"000111100",
  16348=>"100000000",
  16349=>"110111111",
  16350=>"000000111",
  16351=>"000000000",
  16352=>"111111111",
  16353=>"000000111",
  16354=>"111100000",
  16355=>"000000000",
  16356=>"100100111",
  16357=>"000000000",
  16358=>"001000001",
  16359=>"000000000",
  16360=>"110100100",
  16361=>"111111111",
  16362=>"000000011",
  16363=>"000000100",
  16364=>"000000000",
  16365=>"101000000",
  16366=>"000000000",
  16367=>"110111111",
  16368=>"000000100",
  16369=>"000000000",
  16370=>"111000000",
  16371=>"110111110",
  16372=>"111111111",
  16373=>"111111111",
  16374=>"110111111",
  16375=>"000010111",
  16376=>"011001111",
  16377=>"000010010",
  16378=>"011011011",
  16379=>"000000000",
  16380=>"000111111",
  16381=>"111111111",
  16382=>"000001000",
  16383=>"011001001",
  16384=>"111111111",
  16385=>"110011011",
  16386=>"111000000",
  16387=>"111111110",
  16388=>"111111011",
  16389=>"111001011",
  16390=>"111101111",
  16391=>"000000000",
  16392=>"110111000",
  16393=>"000000110",
  16394=>"101111001",
  16395=>"110110111",
  16396=>"000001111",
  16397=>"000000000",
  16398=>"100100100",
  16399=>"000000100",
  16400=>"000000111",
  16401=>"110100000",
  16402=>"000100111",
  16403=>"111111001",
  16404=>"011000011",
  16405=>"000000100",
  16406=>"000100001",
  16407=>"011010110",
  16408=>"011001100",
  16409=>"100000000",
  16410=>"000000110",
  16411=>"011011110",
  16412=>"111111111",
  16413=>"000000011",
  16414=>"000110100",
  16415=>"111101000",
  16416=>"000110111",
  16417=>"111111111",
  16418=>"111111111",
  16419=>"111000000",
  16420=>"001101111",
  16421=>"111111111",
  16422=>"000010110",
  16423=>"000000000",
  16424=>"111100110",
  16425=>"111111111",
  16426=>"000100100",
  16427=>"000000001",
  16428=>"000000110",
  16429=>"000011010",
  16430=>"111111000",
  16431=>"011011000",
  16432=>"000011001",
  16433=>"111111111",
  16434=>"111101111",
  16435=>"110110010",
  16436=>"000000000",
  16437=>"101101101",
  16438=>"111111100",
  16439=>"000000000",
  16440=>"000000111",
  16441=>"111010011",
  16442=>"000000011",
  16443=>"110111100",
  16444=>"000000101",
  16445=>"000010100",
  16446=>"111111110",
  16447=>"000100100",
  16448=>"000000000",
  16449=>"010111111",
  16450=>"000000000",
  16451=>"000001011",
  16452=>"010001011",
  16453=>"001011001",
  16454=>"111111010",
  16455=>"111111111",
  16456=>"100000000",
  16457=>"000000111",
  16458=>"000001011",
  16459=>"110111111",
  16460=>"000000000",
  16461=>"100101111",
  16462=>"000001000",
  16463=>"100111111",
  16464=>"100000000",
  16465=>"000001011",
  16466=>"101100000",
  16467=>"111100001",
  16468=>"111111111",
  16469=>"111001011",
  16470=>"001101111",
  16471=>"111111111",
  16472=>"000111111",
  16473=>"110111111",
  16474=>"000010011",
  16475=>"111000001",
  16476=>"111111111",
  16477=>"000111111",
  16478=>"000000000",
  16479=>"010010011",
  16480=>"000000000",
  16481=>"000000000",
  16482=>"001001111",
  16483=>"100101100",
  16484=>"000000000",
  16485=>"111111101",
  16486=>"000011111",
  16487=>"111101000",
  16488=>"010111111",
  16489=>"000001001",
  16490=>"010000000",
  16491=>"000001001",
  16492=>"111111001",
  16493=>"001000111",
  16494=>"111111111",
  16495=>"111111001",
  16496=>"110001001",
  16497=>"111001001",
  16498=>"000000000",
  16499=>"111111111",
  16500=>"111111111",
  16501=>"111111001",
  16502=>"000100111",
  16503=>"000001000",
  16504=>"111001011",
  16505=>"111111111",
  16506=>"001000001",
  16507=>"000000000",
  16508=>"100100100",
  16509=>"111111111",
  16510=>"111111111",
  16511=>"111111111",
  16512=>"011000000",
  16513=>"000000000",
  16514=>"000111111",
  16515=>"010110110",
  16516=>"111111111",
  16517=>"000000111",
  16518=>"111111110",
  16519=>"001111111",
  16520=>"000000000",
  16521=>"000000000",
  16522=>"111111111",
  16523=>"010100111",
  16524=>"011110110",
  16525=>"000000000",
  16526=>"010000000",
  16527=>"001000111",
  16528=>"000001111",
  16529=>"110110111",
  16530=>"000001101",
  16531=>"111111111",
  16532=>"011011011",
  16533=>"000111111",
  16534=>"000000000",
  16535=>"000000000",
  16536=>"000111111",
  16537=>"000111111",
  16538=>"111111111",
  16539=>"110110100",
  16540=>"111101100",
  16541=>"100000000",
  16542=>"000000011",
  16543=>"000000000",
  16544=>"111110111",
  16545=>"010001000",
  16546=>"101111000",
  16547=>"111111111",
  16548=>"111111111",
  16549=>"111111110",
  16550=>"000000000",
  16551=>"111011000",
  16552=>"000111010",
  16553=>"101001111",
  16554=>"001001111",
  16555=>"000011111",
  16556=>"010110110",
  16557=>"100100100",
  16558=>"000000000",
  16559=>"100111110",
  16560=>"001111000",
  16561=>"101101100",
  16562=>"100100100",
  16563=>"111110110",
  16564=>"111110111",
  16565=>"000011111",
  16566=>"100000000",
  16567=>"000000110",
  16568=>"000000000",
  16569=>"110111111",
  16570=>"001001001",
  16571=>"000000000",
  16572=>"111111101",
  16573=>"111111111",
  16574=>"001111111",
  16575=>"000100101",
  16576=>"111110110",
  16577=>"001000000",
  16578=>"000000000",
  16579=>"110111000",
  16580=>"000000000",
  16581=>"111111111",
  16582=>"011001000",
  16583=>"000000111",
  16584=>"000010011",
  16585=>"101100101",
  16586=>"011001011",
  16587=>"111111110",
  16588=>"111011111",
  16589=>"000011011",
  16590=>"010010000",
  16591=>"111111001",
  16592=>"011000000",
  16593=>"011011010",
  16594=>"111111000",
  16595=>"000000000",
  16596=>"000000000",
  16597=>"100100111",
  16598=>"000000000",
  16599=>"111111111",
  16600=>"111111111",
  16601=>"011111110",
  16602=>"000000000",
  16603=>"010010010",
  16604=>"000101111",
  16605=>"000011010",
  16606=>"100110110",
  16607=>"000000000",
  16608=>"000000111",
  16609=>"000001011",
  16610=>"000000000",
  16611=>"100100101",
  16612=>"101111111",
  16613=>"000010000",
  16614=>"011111011",
  16615=>"101100110",
  16616=>"000000000",
  16617=>"001011000",
  16618=>"111110100",
  16619=>"111100111",
  16620=>"110100000",
  16621=>"000000011",
  16622=>"111011111",
  16623=>"010110111",
  16624=>"111110010",
  16625=>"010110111",
  16626=>"001111100",
  16627=>"000110100",
  16628=>"001111111",
  16629=>"000001001",
  16630=>"111011101",
  16631=>"111111001",
  16632=>"000011111",
  16633=>"000000000",
  16634=>"011111011",
  16635=>"000000000",
  16636=>"110110110",
  16637=>"000011010",
  16638=>"111110000",
  16639=>"001111111",
  16640=>"100000001",
  16641=>"100000100",
  16642=>"110111111",
  16643=>"110100110",
  16644=>"111111111",
  16645=>"110000000",
  16646=>"000010010",
  16647=>"001111111",
  16648=>"111100110",
  16649=>"111111001",
  16650=>"000010000",
  16651=>"001000000",
  16652=>"000000000",
  16653=>"100111011",
  16654=>"111111111",
  16655=>"100100100",
  16656=>"100100100",
  16657=>"100111001",
  16658=>"000010000",
  16659=>"111101111",
  16660=>"001001101",
  16661=>"100100001",
  16662=>"011111111",
  16663=>"010111111",
  16664=>"010111111",
  16665=>"100100000",
  16666=>"000000000",
  16667=>"111111111",
  16668=>"111100000",
  16669=>"111111011",
  16670=>"001001111",
  16671=>"000111111",
  16672=>"100110111",
  16673=>"000111111",
  16674=>"101100111",
  16675=>"001111111",
  16676=>"000100100",
  16677=>"111001001",
  16678=>"010011111",
  16679=>"001101111",
  16680=>"111000000",
  16681=>"000000000",
  16682=>"000000000",
  16683=>"000000000",
  16684=>"111111010",
  16685=>"110000100",
  16686=>"011010000",
  16687=>"000100000",
  16688=>"110000111",
  16689=>"100111011",
  16690=>"000000000",
  16691=>"100000000",
  16692=>"000000000",
  16693=>"110111100",
  16694=>"110111011",
  16695=>"001011000",
  16696=>"000000000",
  16697=>"000001011",
  16698=>"101110111",
  16699=>"000000000",
  16700=>"100110111",
  16701=>"110010000",
  16702=>"111111100",
  16703=>"000000000",
  16704=>"100111000",
  16705=>"110011011",
  16706=>"000000000",
  16707=>"000000000",
  16708=>"111111111",
  16709=>"110111111",
  16710=>"111110000",
  16711=>"011110111",
  16712=>"000000000",
  16713=>"111011011",
  16714=>"001000010",
  16715=>"010000000",
  16716=>"111111111",
  16717=>"001001011",
  16718=>"111111110",
  16719=>"000000000",
  16720=>"000110000",
  16721=>"000000011",
  16722=>"111111111",
  16723=>"111111111",
  16724=>"000000000",
  16725=>"000001000",
  16726=>"100000010",
  16727=>"111111001",
  16728=>"111011000",
  16729=>"011111110",
  16730=>"100110111",
  16731=>"000000000",
  16732=>"010000000",
  16733=>"100101000",
  16734=>"000000100",
  16735=>"110110111",
  16736=>"111001011",
  16737=>"001000000",
  16738=>"111110000",
  16739=>"010000000",
  16740=>"111111111",
  16741=>"001011000",
  16742=>"111111011",
  16743=>"100000000",
  16744=>"111001000",
  16745=>"111011011",
  16746=>"111111111",
  16747=>"100110111",
  16748=>"100000000",
  16749=>"010000000",
  16750=>"000000000",
  16751=>"100111111",
  16752=>"000000101",
  16753=>"111101111",
  16754=>"000001001",
  16755=>"110100110",
  16756=>"101001001",
  16757=>"111001001",
  16758=>"111111110",
  16759=>"111111111",
  16760=>"101111111",
  16761=>"000000000",
  16762=>"000000000",
  16763=>"111111111",
  16764=>"001001101",
  16765=>"111111001",
  16766=>"100100000",
  16767=>"111111000",
  16768=>"110110111",
  16769=>"000110010",
  16770=>"111111111",
  16771=>"001000111",
  16772=>"111011001",
  16773=>"000000000",
  16774=>"010010110",
  16775=>"000000111",
  16776=>"010010000",
  16777=>"110110000",
  16778=>"000000000",
  16779=>"000111011",
  16780=>"111111111",
  16781=>"111111100",
  16782=>"110111110",
  16783=>"000001111",
  16784=>"000000000",
  16785=>"101111001",
  16786=>"000000000",
  16787=>"111011111",
  16788=>"000000101",
  16789=>"001001011",
  16790=>"001101101",
  16791=>"110011101",
  16792=>"000000101",
  16793=>"111111010",
  16794=>"001000000",
  16795=>"101100101",
  16796=>"101000100",
  16797=>"111110110",
  16798=>"100000000",
  16799=>"011111111",
  16800=>"000001001",
  16801=>"000000011",
  16802=>"010000010",
  16803=>"111111011",
  16804=>"000000001",
  16805=>"011111000",
  16806=>"111111000",
  16807=>"000111111",
  16808=>"001000000",
  16809=>"000011111",
  16810=>"001111111",
  16811=>"000100000",
  16812=>"111111111",
  16813=>"111110111",
  16814=>"000000011",
  16815=>"101011001",
  16816=>"010110111",
  16817=>"100111111",
  16818=>"111011111",
  16819=>"011100000",
  16820=>"000000101",
  16821=>"000000000",
  16822=>"000000000",
  16823=>"111110111",
  16824=>"000011111",
  16825=>"000000100",
  16826=>"100000101",
  16827=>"000001010",
  16828=>"111111111",
  16829=>"000000000",
  16830=>"000000000",
  16831=>"001000100",
  16832=>"100111000",
  16833=>"111111000",
  16834=>"001111111",
  16835=>"010110000",
  16836=>"111111001",
  16837=>"100000100",
  16838=>"000001111",
  16839=>"010111000",
  16840=>"000000111",
  16841=>"000110000",
  16842=>"000000000",
  16843=>"000000011",
  16844=>"000000000",
  16845=>"000000000",
  16846=>"110111110",
  16847=>"011000001",
  16848=>"000000000",
  16849=>"000000000",
  16850=>"001011011",
  16851=>"111111111",
  16852=>"110110100",
  16853=>"100110011",
  16854=>"010010010",
  16855=>"000000000",
  16856=>"010000000",
  16857=>"100000100",
  16858=>"101101111",
  16859=>"001001100",
  16860=>"000000100",
  16861=>"000000000",
  16862=>"111111000",
  16863=>"111100100",
  16864=>"000000000",
  16865=>"000000011",
  16866=>"000110111",
  16867=>"000000000",
  16868=>"000010000",
  16869=>"000001111",
  16870=>"000010000",
  16871=>"011111111",
  16872=>"100000000",
  16873=>"000101111",
  16874=>"011011111",
  16875=>"100101001",
  16876=>"001000000",
  16877=>"000000000",
  16878=>"000010000",
  16879=>"111111111",
  16880=>"110111111",
  16881=>"000000000",
  16882=>"111111111",
  16883=>"000000000",
  16884=>"111111111",
  16885=>"111111011",
  16886=>"000000001",
  16887=>"100000110",
  16888=>"000011011",
  16889=>"000010000",
  16890=>"001001011",
  16891=>"000011110",
  16892=>"111111111",
  16893=>"000000000",
  16894=>"110110000",
  16895=>"111001111",
  16896=>"000000000",
  16897=>"000000000",
  16898=>"111111111",
  16899=>"000111111",
  16900=>"000100100",
  16901=>"000000000",
  16902=>"000000000",
  16903=>"111111111",
  16904=>"000111111",
  16905=>"000000111",
  16906=>"111111100",
  16907=>"001000000",
  16908=>"000000000",
  16909=>"000000001",
  16910=>"011011000",
  16911=>"010001000",
  16912=>"110110000",
  16913=>"000011011",
  16914=>"001001001",
  16915=>"100000000",
  16916=>"111111111",
  16917=>"011111111",
  16918=>"111111100",
  16919=>"100000010",
  16920=>"100110111",
  16921=>"100111001",
  16922=>"111110111",
  16923=>"011011000",
  16924=>"000000100",
  16925=>"101000001",
  16926=>"111111111",
  16927=>"000000000",
  16928=>"110110110",
  16929=>"111111111",
  16930=>"000000110",
  16931=>"000000000",
  16932=>"000000000",
  16933=>"100000001",
  16934=>"000000000",
  16935=>"000010111",
  16936=>"111111111",
  16937=>"000000000",
  16938=>"000000000",
  16939=>"001000000",
  16940=>"111111111",
  16941=>"000111111",
  16942=>"000000000",
  16943=>"000000000",
  16944=>"000011011",
  16945=>"111101101",
  16946=>"100000001",
  16947=>"010000001",
  16948=>"001111001",
  16949=>"111111111",
  16950=>"000000000",
  16951=>"111011110",
  16952=>"000000000",
  16953=>"000100000",
  16954=>"100001111",
  16955=>"111111000",
  16956=>"000000010",
  16957=>"000000000",
  16958=>"001000000",
  16959=>"000000000",
  16960=>"000000000",
  16961=>"000000000",
  16962=>"000000100",
  16963=>"000000000",
  16964=>"000000000",
  16965=>"111111011",
  16966=>"111000000",
  16967=>"000100100",
  16968=>"011010110",
  16969=>"000001011",
  16970=>"111111111",
  16971=>"000000000",
  16972=>"111000000",
  16973=>"111111111",
  16974=>"111111111",
  16975=>"111111111",
  16976=>"010111111",
  16977=>"000000000",
  16978=>"100000000",
  16979=>"100000000",
  16980=>"000111111",
  16981=>"000000001",
  16982=>"001001111",
  16983=>"111111111",
  16984=>"110111111",
  16985=>"111101111",
  16986=>"110100000",
  16987=>"011010000",
  16988=>"000001111",
  16989=>"000010000",
  16990=>"111000000",
  16991=>"000100000",
  16992=>"111001000",
  16993=>"110011001",
  16994=>"110010000",
  16995=>"001000111",
  16996=>"100000100",
  16997=>"000000000",
  16998=>"111111010",
  16999=>"111111011",
  17000=>"000000100",
  17001=>"101101101",
  17002=>"111111101",
  17003=>"100000000",
  17004=>"000000000",
  17005=>"000000000",
  17006=>"011000000",
  17007=>"000000000",
  17008=>"000000000",
  17009=>"111111111",
  17010=>"000000101",
  17011=>"000000100",
  17012=>"000011011",
  17013=>"000000100",
  17014=>"000000111",
  17015=>"000000000",
  17016=>"001011111",
  17017=>"111011011",
  17018=>"101111000",
  17019=>"111111111",
  17020=>"111110110",
  17021=>"000000000",
  17022=>"100000000",
  17023=>"000000000",
  17024=>"111111111",
  17025=>"111111101",
  17026=>"111111111",
  17027=>"110100000",
  17028=>"000000011",
  17029=>"111111101",
  17030=>"110010110",
  17031=>"011000000",
  17032=>"100000000",
  17033=>"000110110",
  17034=>"000000001",
  17035=>"111111100",
  17036=>"100000000",
  17037=>"111000000",
  17038=>"110110111",
  17039=>"001001000",
  17040=>"111111111",
  17041=>"000001000",
  17042=>"111111011",
  17043=>"111111111",
  17044=>"011011001",
  17045=>"011010111",
  17046=>"000000111",
  17047=>"111111111",
  17048=>"111111111",
  17049=>"001000100",
  17050=>"110010000",
  17051=>"000000000",
  17052=>"111111111",
  17053=>"111000000",
  17054=>"100000111",
  17055=>"010010000",
  17056=>"110110000",
  17057=>"111111010",
  17058=>"000000000",
  17059=>"001001111",
  17060=>"000000000",
  17061=>"010010101",
  17062=>"111111111",
  17063=>"111111111",
  17064=>"000000000",
  17065=>"111111111",
  17066=>"000100111",
  17067=>"111111111",
  17068=>"000000011",
  17069=>"010010110",
  17070=>"111111110",
  17071=>"000000100",
  17072=>"111111111",
  17073=>"000000000",
  17074=>"111100111",
  17075=>"011000000",
  17076=>"000110010",
  17077=>"001101111",
  17078=>"111111001",
  17079=>"111111111",
  17080=>"000000000",
  17081=>"111111110",
  17082=>"001101101",
  17083=>"000000000",
  17084=>"110000000",
  17085=>"100000101",
  17086=>"111110110",
  17087=>"001110110",
  17088=>"101000000",
  17089=>"111110000",
  17090=>"111111111",
  17091=>"111111011",
  17092=>"100000001",
  17093=>"000000000",
  17094=>"101001001",
  17095=>"011010000",
  17096=>"000000000",
  17097=>"000000111",
  17098=>"100000111",
  17099=>"000100000",
  17100=>"111111111",
  17101=>"000111000",
  17102=>"110111111",
  17103=>"000000000",
  17104=>"010000000",
  17105=>"110111111",
  17106=>"111000000",
  17107=>"000010110",
  17108=>"000001111",
  17109=>"000000000",
  17110=>"111000000",
  17111=>"111001000",
  17112=>"000000000",
  17113=>"110110100",
  17114=>"111000111",
  17115=>"110100000",
  17116=>"000000111",
  17117=>"111111111",
  17118=>"000000000",
  17119=>"110110111",
  17120=>"000000000",
  17121=>"000011000",
  17122=>"000000001",
  17123=>"111111111",
  17124=>"000100000",
  17125=>"101010000",
  17126=>"000000000",
  17127=>"111000000",
  17128=>"101111111",
  17129=>"000000000",
  17130=>"111111111",
  17131=>"111111111",
  17132=>"101100110",
  17133=>"000000000",
  17134=>"111111111",
  17135=>"111111111",
  17136=>"111000100",
  17137=>"111110111",
  17138=>"100111111",
  17139=>"000100000",
  17140=>"000000000",
  17141=>"111100110",
  17142=>"011011111",
  17143=>"000000000",
  17144=>"000111111",
  17145=>"111111111",
  17146=>"111111111",
  17147=>"000000000",
  17148=>"111110111",
  17149=>"001001011",
  17150=>"011001111",
  17151=>"000000000",
  17152=>"011111111",
  17153=>"111111110",
  17154=>"111111110",
  17155=>"000111111",
  17156=>"111111111",
  17157=>"111111111",
  17158=>"110110111",
  17159=>"111111111",
  17160=>"000000000",
  17161=>"111101101",
  17162=>"111111000",
  17163=>"111011001",
  17164=>"111111000",
  17165=>"000000000",
  17166=>"111111000",
  17167=>"100111000",
  17168=>"011001001",
  17169=>"000110111",
  17170=>"111000011",
  17171=>"000000000",
  17172=>"101111111",
  17173=>"110010010",
  17174=>"001101111",
  17175=>"111011000",
  17176=>"110110110",
  17177=>"000100000",
  17178=>"111110000",
  17179=>"000000111",
  17180=>"110001001",
  17181=>"110000000",
  17182=>"111111111",
  17183=>"000011011",
  17184=>"000000000",
  17185=>"111111011",
  17186=>"111101000",
  17187=>"000000000",
  17188=>"000000011",
  17189=>"000001111",
  17190=>"011010000",
  17191=>"110110010",
  17192=>"000111111",
  17193=>"111111000",
  17194=>"100010000",
  17195=>"000000000",
  17196=>"001000000",
  17197=>"000000000",
  17198=>"000111010",
  17199=>"011000100",
  17200=>"111111111",
  17201=>"000000000",
  17202=>"000000000",
  17203=>"000000000",
  17204=>"000000110",
  17205=>"000000001",
  17206=>"000000010",
  17207=>"111111111",
  17208=>"001001000",
  17209=>"111111011",
  17210=>"001100101",
  17211=>"111111111",
  17212=>"000000000",
  17213=>"011011000",
  17214=>"011001001",
  17215=>"100000000",
  17216=>"000000000",
  17217=>"111011011",
  17218=>"110010000",
  17219=>"001111111",
  17220=>"000000000",
  17221=>"001001111",
  17222=>"000000111",
  17223=>"000010010",
  17224=>"111111111",
  17225=>"110110111",
  17226=>"000000111",
  17227=>"111111101",
  17228=>"000000000",
  17229=>"111000000",
  17230=>"111111111",
  17231=>"000000000",
  17232=>"110111101",
  17233=>"011111101",
  17234=>"110111110",
  17235=>"000110110",
  17236=>"110111111",
  17237=>"011011011",
  17238=>"111000001",
  17239=>"111111111",
  17240=>"111100000",
  17241=>"000000111",
  17242=>"111011111",
  17243=>"111111000",
  17244=>"000101101",
  17245=>"001001000",
  17246=>"100100111",
  17247=>"110111010",
  17248=>"000000000",
  17249=>"111111111",
  17250=>"111101111",
  17251=>"111111111",
  17252=>"101011011",
  17253=>"000000011",
  17254=>"111011111",
  17255=>"000110000",
  17256=>"001111111",
  17257=>"000000110",
  17258=>"001000110",
  17259=>"011011111",
  17260=>"000000000",
  17261=>"101111111",
  17262=>"110111111",
  17263=>"000000100",
  17264=>"000000001",
  17265=>"110101000",
  17266=>"000000111",
  17267=>"111100100",
  17268=>"111111111",
  17269=>"111111111",
  17270=>"001101100",
  17271=>"000000000",
  17272=>"110000010",
  17273=>"111111111",
  17274=>"110110111",
  17275=>"010010010",
  17276=>"101101111",
  17277=>"110000000",
  17278=>"111011111",
  17279=>"001001000",
  17280=>"111111111",
  17281=>"111010111",
  17282=>"110000000",
  17283=>"110111111",
  17284=>"111111111",
  17285=>"000000000",
  17286=>"000000000",
  17287=>"000000111",
  17288=>"110101111",
  17289=>"111111111",
  17290=>"000000000",
  17291=>"111111111",
  17292=>"101111111",
  17293=>"000000000",
  17294=>"011001110",
  17295=>"100000000",
  17296=>"110111111",
  17297=>"000000111",
  17298=>"111111101",
  17299=>"000000000",
  17300=>"110000000",
  17301=>"000000000",
  17302=>"011000001",
  17303=>"000000000",
  17304=>"001111111",
  17305=>"111010111",
  17306=>"010111111",
  17307=>"000000000",
  17308=>"000001011",
  17309=>"000001001",
  17310=>"011001000",
  17311=>"000000000",
  17312=>"000000000",
  17313=>"111001001",
  17314=>"000001011",
  17315=>"111111111",
  17316=>"111100100",
  17317=>"000000000",
  17318=>"001001101",
  17319=>"111111111",
  17320=>"111111010",
  17321=>"110111111",
  17322=>"000000111",
  17323=>"000001001",
  17324=>"000000000",
  17325=>"000000011",
  17326=>"110000100",
  17327=>"001000101",
  17328=>"100100111",
  17329=>"111111111",
  17330=>"111111111",
  17331=>"000011000",
  17332=>"111111111",
  17333=>"000000000",
  17334=>"111111101",
  17335=>"000000000",
  17336=>"000110111",
  17337=>"000000010",
  17338=>"001111111",
  17339=>"110110000",
  17340=>"001001001",
  17341=>"111111000",
  17342=>"111110000",
  17343=>"011111111",
  17344=>"000000000",
  17345=>"000000010",
  17346=>"000000000",
  17347=>"110111111",
  17348=>"000000000",
  17349=>"011000100",
  17350=>"000000000",
  17351=>"000011000",
  17352=>"000000000",
  17353=>"001011001",
  17354=>"000000111",
  17355=>"111111111",
  17356=>"111111000",
  17357=>"111000000",
  17358=>"000000000",
  17359=>"100111111",
  17360=>"101100100",
  17361=>"111111111",
  17362=>"111111111",
  17363=>"100000000",
  17364=>"001001000",
  17365=>"100000001",
  17366=>"000000000",
  17367=>"001001011",
  17368=>"000011000",
  17369=>"000111001",
  17370=>"011011111",
  17371=>"111111110",
  17372=>"000000111",
  17373=>"111111111",
  17374=>"000000000",
  17375=>"000000110",
  17376=>"111111100",
  17377=>"000000001",
  17378=>"100100111",
  17379=>"000000000",
  17380=>"111111111",
  17381=>"011011011",
  17382=>"000000000",
  17383=>"110111111",
  17384=>"000000000",
  17385=>"111110000",
  17386=>"000000000",
  17387=>"000000000",
  17388=>"100111011",
  17389=>"000000000",
  17390=>"011000001",
  17391=>"000000000",
  17392=>"001000000",
  17393=>"100111111",
  17394=>"111001111",
  17395=>"000100100",
  17396=>"000000000",
  17397=>"111110000",
  17398=>"111111111",
  17399=>"111110010",
  17400=>"000000000",
  17401=>"100000001",
  17402=>"001001000",
  17403=>"111000000",
  17404=>"111111000",
  17405=>"000110111",
  17406=>"111011000",
  17407=>"111111111",
  17408=>"010000010",
  17409=>"000101111",
  17410=>"111101111",
  17411=>"100000000",
  17412=>"111111000",
  17413=>"100101011",
  17414=>"010111111",
  17415=>"110111111",
  17416=>"010000001",
  17417=>"001000000",
  17418=>"111101111",
  17419=>"000000000",
  17420=>"100111111",
  17421=>"000000010",
  17422=>"000000000",
  17423=>"010111000",
  17424=>"111000100",
  17425=>"000011100",
  17426=>"000000111",
  17427=>"111011111",
  17428=>"000000110",
  17429=>"000000010",
  17430=>"101000000",
  17431=>"011001001",
  17432=>"100100000",
  17433=>"000000100",
  17434=>"000000010",
  17435=>"000011000",
  17436=>"111111111",
  17437=>"000000000",
  17438=>"111000110",
  17439=>"000110111",
  17440=>"000111111",
  17441=>"000000101",
  17442=>"100111100",
  17443=>"111111000",
  17444=>"000000001",
  17445=>"111110000",
  17446=>"111001001",
  17447=>"010000000",
  17448=>"101111111",
  17449=>"111110111",
  17450=>"000000111",
  17451=>"011111111",
  17452=>"000000111",
  17453=>"010111000",
  17454=>"000000000",
  17455=>"110100110",
  17456=>"000000001",
  17457=>"000111111",
  17458=>"111101001",
  17459=>"000000000",
  17460=>"010111110",
  17461=>"000001110",
  17462=>"111001001",
  17463=>"001000000",
  17464=>"000000001",
  17465=>"110010011",
  17466=>"000111111",
  17467=>"111111111",
  17468=>"101000000",
  17469=>"111111110",
  17470=>"000000110",
  17471=>"000101111",
  17472=>"000000100",
  17473=>"111001000",
  17474=>"111111111",
  17475=>"110000000",
  17476=>"101101000",
  17477=>"000110111",
  17478=>"000000011",
  17479=>"000000111",
  17480=>"011111000",
  17481=>"111110111",
  17482=>"111100100",
  17483=>"111001000",
  17484=>"011100100",
  17485=>"000000101",
  17486=>"000111111",
  17487=>"000000101",
  17488=>"111000000",
  17489=>"000001000",
  17490=>"111000000",
  17491=>"111111000",
  17492=>"010111000",
  17493=>"101111100",
  17494=>"111101111",
  17495=>"111111011",
  17496=>"111111011",
  17497=>"111111111",
  17498=>"111111111",
  17499=>"001000110",
  17500=>"000000010",
  17501=>"111000000",
  17502=>"111100000",
  17503=>"000110000",
  17504=>"111111111",
  17505=>"000001011",
  17506=>"000111101",
  17507=>"111111111",
  17508=>"111110000",
  17509=>"101000110",
  17510=>"000000110",
  17511=>"000000111",
  17512=>"111111111",
  17513=>"010010010",
  17514=>"011111111",
  17515=>"000000000",
  17516=>"011011001",
  17517=>"000111111",
  17518=>"111101111",
  17519=>"111111111",
  17520=>"111000000",
  17521=>"000000101",
  17522=>"000111111",
  17523=>"111000000",
  17524=>"000000100",
  17525=>"011111110",
  17526=>"000000000",
  17527=>"000000001",
  17528=>"001000000",
  17529=>"000000000",
  17530=>"111000000",
  17531=>"000101101",
  17532=>"000000000",
  17533=>"000111110",
  17534=>"000000101",
  17535=>"111111000",
  17536=>"111111100",
  17537=>"100000000",
  17538=>"000000111",
  17539=>"111111001",
  17540=>"000000100",
  17541=>"000000000",
  17542=>"100000000",
  17543=>"000000000",
  17544=>"001111111",
  17545=>"111110111",
  17546=>"111101111",
  17547=>"100000111",
  17548=>"000000000",
  17549=>"111101111",
  17550=>"111111000",
  17551=>"000000011",
  17552=>"001000101",
  17553=>"111000001",
  17554=>"100111100",
  17555=>"111111000",
  17556=>"000000000",
  17557=>"000000111",
  17558=>"111000000",
  17559=>"000000100",
  17560=>"101000101",
  17561=>"011111111",
  17562=>"000000000",
  17563=>"000000000",
  17564=>"111110000",
  17565=>"111000000",
  17566=>"111100010",
  17567=>"111110111",
  17568=>"000000000",
  17569=>"001000000",
  17570=>"111111001",
  17571=>"011001011",
  17572=>"111001001",
  17573=>"000111111",
  17574=>"000000000",
  17575=>"000100110",
  17576=>"000000001",
  17577=>"001001000",
  17578=>"000000000",
  17579=>"000000000",
  17580=>"111111001",
  17581=>"100100000",
  17582=>"000000111",
  17583=>"000111111",
  17584=>"000111111",
  17585=>"000100111",
  17586=>"010111111",
  17587=>"100000000",
  17588=>"000000001",
  17589=>"001111111",
  17590=>"000011111",
  17591=>"111111110",
  17592=>"111001111",
  17593=>"111111011",
  17594=>"101000000",
  17595=>"101000000",
  17596=>"000000100",
  17597=>"010111111",
  17598=>"110111111",
  17599=>"000000001",
  17600=>"111000110",
  17601=>"101000001",
  17602=>"011111111",
  17603=>"111011000",
  17604=>"111111000",
  17605=>"111001011",
  17606=>"111000010",
  17607=>"000000000",
  17608=>"000110010",
  17609=>"100111111",
  17610=>"000001000",
  17611=>"000000001",
  17612=>"100111111",
  17613=>"000000010",
  17614=>"111111111",
  17615=>"000000111",
  17616=>"100111111",
  17617=>"101000000",
  17618=>"100000111",
  17619=>"000000000",
  17620=>"100000101",
  17621=>"111111000",
  17622=>"000000001",
  17623=>"000000000",
  17624=>"000000111",
  17625=>"111011000",
  17626=>"000000000",
  17627=>"111001111",
  17628=>"111111000",
  17629=>"000000111",
  17630=>"111111110",
  17631=>"111111111",
  17632=>"111100000",
  17633=>"000001010",
  17634=>"111000000",
  17635=>"110110111",
  17636=>"000000000",
  17637=>"000001101",
  17638=>"000000110",
  17639=>"111111111",
  17640=>"111011010",
  17641=>"101111110",
  17642=>"000001000",
  17643=>"000000000",
  17644=>"000000000",
  17645=>"000111000",
  17646=>"111000101",
  17647=>"001011011",
  17648=>"000000000",
  17649=>"111000000",
  17650=>"000000010",
  17651=>"000000110",
  17652=>"010011011",
  17653=>"011011011",
  17654=>"000000001",
  17655=>"111011011",
  17656=>"000011011",
  17657=>"000011000",
  17658=>"111110000",
  17659=>"111111111",
  17660=>"001100011",
  17661=>"000000000",
  17662=>"100000001",
  17663=>"000100111",
  17664=>"111100010",
  17665=>"111011011",
  17666=>"011010100",
  17667=>"111011011",
  17668=>"000111111",
  17669=>"001111111",
  17670=>"111101111",
  17671=>"111111001",
  17672=>"111111111",
  17673=>"111111100",
  17674=>"000000010",
  17675=>"111111000",
  17676=>"111101111",
  17677=>"000001111",
  17678=>"101001111",
  17679=>"111000000",
  17680=>"000000011",
  17681=>"000110000",
  17682=>"000000000",
  17683=>"000001110",
  17684=>"000110000",
  17685=>"000000000",
  17686=>"001111111",
  17687=>"110111111",
  17688=>"111111110",
  17689=>"111111111",
  17690=>"100111111",
  17691=>"000111111",
  17692=>"111111111",
  17693=>"111111000",
  17694=>"000000111",
  17695=>"100111111",
  17696=>"111001000",
  17697=>"111111011",
  17698=>"111111000",
  17699=>"000111111",
  17700=>"001111111",
  17701=>"000000000",
  17702=>"000111011",
  17703=>"001000000",
  17704=>"000000000",
  17705=>"010111010",
  17706=>"111111000",
  17707=>"000000111",
  17708=>"111100000",
  17709=>"001000000",
  17710=>"000000001",
  17711=>"100000000",
  17712=>"000000000",
  17713=>"000000000",
  17714=>"001111110",
  17715=>"111000000",
  17716=>"000110001",
  17717=>"010011011",
  17718=>"000000000",
  17719=>"000000000",
  17720=>"111111111",
  17721=>"111000111",
  17722=>"010000000",
  17723=>"111001000",
  17724=>"111111111",
  17725=>"000000000",
  17726=>"111111111",
  17727=>"111000011",
  17728=>"111101100",
  17729=>"000000000",
  17730=>"111100010",
  17731=>"111000001",
  17732=>"111111000",
  17733=>"111111111",
  17734=>"111111000",
  17735=>"000000000",
  17736=>"111000000",
  17737=>"000000011",
  17738=>"000111111",
  17739=>"000000000",
  17740=>"000000000",
  17741=>"111000000",
  17742=>"100100100",
  17743=>"111001111",
  17744=>"111000000",
  17745=>"101000101",
  17746=>"111000000",
  17747=>"000000110",
  17748=>"011000000",
  17749=>"011011001",
  17750=>"110111111",
  17751=>"001000000",
  17752=>"010111111",
  17753=>"110000000",
  17754=>"111011100",
  17755=>"000000000",
  17756=>"000000110",
  17757=>"000111000",
  17758=>"000001000",
  17759=>"000000001",
  17760=>"000000000",
  17761=>"101001000",
  17762=>"111001001",
  17763=>"110111111",
  17764=>"111111110",
  17765=>"111000000",
  17766=>"000000001",
  17767=>"101101001",
  17768=>"101100000",
  17769=>"001000000",
  17770=>"000000000",
  17771=>"111001111",
  17772=>"110111111",
  17773=>"101001000",
  17774=>"010111010",
  17775=>"111111111",
  17776=>"000111111",
  17777=>"111111111",
  17778=>"000000111",
  17779=>"100111000",
  17780=>"111111111",
  17781=>"111111111",
  17782=>"011000001",
  17783=>"101101000",
  17784=>"111100111",
  17785=>"111000000",
  17786=>"001000000",
  17787=>"011000000",
  17788=>"000000000",
  17789=>"111111011",
  17790=>"111100000",
  17791=>"001111000",
  17792=>"001001100",
  17793=>"000000111",
  17794=>"000100110",
  17795=>"000000001",
  17796=>"000101111",
  17797=>"111010010",
  17798=>"000001111",
  17799=>"101110000",
  17800=>"001011111",
  17801=>"111111010",
  17802=>"000000000",
  17803=>"010111111",
  17804=>"111100111",
  17805=>"110110100",
  17806=>"111100101",
  17807=>"000000000",
  17808=>"001000000",
  17809=>"100000101",
  17810=>"101100000",
  17811=>"111111111",
  17812=>"001000111",
  17813=>"111111000",
  17814=>"111111011",
  17815=>"011111110",
  17816=>"100111111",
  17817=>"001001001",
  17818=>"111010000",
  17819=>"111111001",
  17820=>"100000000",
  17821=>"111101111",
  17822=>"101000000",
  17823=>"111111110",
  17824=>"010111101",
  17825=>"111111011",
  17826=>"111010000",
  17827=>"111111101",
  17828=>"000010000",
  17829=>"000001000",
  17830=>"000000000",
  17831=>"000000000",
  17832=>"000000101",
  17833=>"000000000",
  17834=>"000000101",
  17835=>"000001011",
  17836=>"111010010",
  17837=>"000000000",
  17838=>"111000101",
  17839=>"101101000",
  17840=>"000000011",
  17841=>"000000111",
  17842=>"111111111",
  17843=>"000000000",
  17844=>"000001000",
  17845=>"011000010",
  17846=>"000000100",
  17847=>"111010111",
  17848=>"000000111",
  17849=>"000000000",
  17850=>"000111111",
  17851=>"001000000",
  17852=>"000000001",
  17853=>"000000000",
  17854=>"111000111",
  17855=>"100111111",
  17856=>"111111011",
  17857=>"000000111",
  17858=>"111111011",
  17859=>"111000000",
  17860=>"111111000",
  17861=>"000000000",
  17862=>"010000000",
  17863=>"000000001",
  17864=>"101000001",
  17865=>"000101111",
  17866=>"001000000",
  17867=>"000000000",
  17868=>"110000000",
  17869=>"011111011",
  17870=>"000000000",
  17871=>"000000000",
  17872=>"111101001",
  17873=>"100000000",
  17874=>"001111111",
  17875=>"000000011",
  17876=>"000001101",
  17877=>"000000001",
  17878=>"000000000",
  17879=>"011111111",
  17880=>"100100110",
  17881=>"111111010",
  17882=>"111000001",
  17883=>"000000001",
  17884=>"001111000",
  17885=>"000000000",
  17886=>"011000000",
  17887=>"000000111",
  17888=>"000001000",
  17889=>"110111111",
  17890=>"000000001",
  17891=>"100000000",
  17892=>"000000000",
  17893=>"000000000",
  17894=>"111111111",
  17895=>"011010011",
  17896=>"111111010",
  17897=>"111110100",
  17898=>"011000111",
  17899=>"111000000",
  17900=>"000000110",
  17901=>"000111110",
  17902=>"000000000",
  17903=>"000000110",
  17904=>"101101000",
  17905=>"000111111",
  17906=>"101100001",
  17907=>"111010000",
  17908=>"000000000",
  17909=>"000000000",
  17910=>"111111101",
  17911=>"001110110",
  17912=>"111110010",
  17913=>"001011001",
  17914=>"111111101",
  17915=>"000000001",
  17916=>"000000111",
  17917=>"111000000",
  17918=>"100111100",
  17919=>"000000111",
  17920=>"111000000",
  17921=>"001000001",
  17922=>"111111111",
  17923=>"000000100",
  17924=>"000100000",
  17925=>"000000011",
  17926=>"111111101",
  17927=>"000111111",
  17928=>"111111111",
  17929=>"111111011",
  17930=>"100001001",
  17931=>"000111111",
  17932=>"111110111",
  17933=>"000110000",
  17934=>"111101111",
  17935=>"000000101",
  17936=>"101111110",
  17937=>"110000111",
  17938=>"100100111",
  17939=>"000000001",
  17940=>"111000110",
  17941=>"001000111",
  17942=>"000111011",
  17943=>"111111111",
  17944=>"001111000",
  17945=>"111101111",
  17946=>"101001001",
  17947=>"110111111",
  17948=>"111101111",
  17949=>"000010000",
  17950=>"100110110",
  17951=>"000100000",
  17952=>"000000111",
  17953=>"111111110",
  17954=>"001001111",
  17955=>"111001000",
  17956=>"000000011",
  17957=>"111111111",
  17958=>"111110000",
  17959=>"110100011",
  17960=>"111111111",
  17961=>"000000000",
  17962=>"100101111",
  17963=>"101001000",
  17964=>"010000111",
  17965=>"011000000",
  17966=>"101111111",
  17967=>"001000000",
  17968=>"000000010",
  17969=>"101101101",
  17970=>"000000001",
  17971=>"111111111",
  17972=>"111000000",
  17973=>"111111100",
  17974=>"100000001",
  17975=>"011011111",
  17976=>"100100000",
  17977=>"101101011",
  17978=>"001000000",
  17979=>"111001000",
  17980=>"111000000",
  17981=>"100000000",
  17982=>"111001111",
  17983=>"000000001",
  17984=>"111000000",
  17985=>"000000100",
  17986=>"111111111",
  17987=>"100111111",
  17988=>"000101111",
  17989=>"000010000",
  17990=>"111111111",
  17991=>"111111111",
  17992=>"000000000",
  17993=>"000000000",
  17994=>"000000000",
  17995=>"001011000",
  17996=>"000111011",
  17997=>"000000100",
  17998=>"000000001",
  17999=>"111111101",
  18000=>"111011011",
  18001=>"111000000",
  18002=>"111111111",
  18003=>"100011110",
  18004=>"000000000",
  18005=>"011111111",
  18006=>"000100110",
  18007=>"110111111",
  18008=>"000000000",
  18009=>"101000001",
  18010=>"111111110",
  18011=>"111111111",
  18012=>"000000001",
  18013=>"000000000",
  18014=>"111111000",
  18015=>"010000010",
  18016=>"111111111",
  18017=>"111110000",
  18018=>"000110111",
  18019=>"111110111",
  18020=>"000000101",
  18021=>"000000001",
  18022=>"111110000",
  18023=>"111111111",
  18024=>"011010000",
  18025=>"111111111",
  18026=>"111111010",
  18027=>"110111010",
  18028=>"001000100",
  18029=>"111111111",
  18030=>"000000100",
  18031=>"111111111",
  18032=>"111111110",
  18033=>"000010011",
  18034=>"000000000",
  18035=>"010110110",
  18036=>"111111111",
  18037=>"100101101",
  18038=>"001001111",
  18039=>"111001000",
  18040=>"110111111",
  18041=>"010111110",
  18042=>"111110111",
  18043=>"111111110",
  18044=>"110110110",
  18045=>"000010111",
  18046=>"111111111",
  18047=>"010111110",
  18048=>"111000111",
  18049=>"111111111",
  18050=>"000000111",
  18051=>"000100000",
  18052=>"111111111",
  18053=>"000000000",
  18054=>"011000000",
  18055=>"111111111",
  18056=>"111111110",
  18057=>"100100101",
  18058=>"000000101",
  18059=>"100110111",
  18060=>"111111111",
  18061=>"111000100",
  18062=>"001000000",
  18063=>"111111111",
  18064=>"000000000",
  18065=>"000001011",
  18066=>"111111111",
  18067=>"101000000",
  18068=>"111111000",
  18069=>"000000111",
  18070=>"111001001",
  18071=>"000000000",
  18072=>"111111010",
  18073=>"101000000",
  18074=>"111111111",
  18075=>"111111111",
  18076=>"000111111",
  18077=>"000000000",
  18078=>"100101111",
  18079=>"111000100",
  18080=>"011011111",
  18081=>"111111000",
  18082=>"000000101",
  18083=>"000011111",
  18084=>"111000000",
  18085=>"100100110",
  18086=>"111111111",
  18087=>"111111001",
  18088=>"111001011",
  18089=>"010111111",
  18090=>"000111111",
  18091=>"111111111",
  18092=>"000000000",
  18093=>"101111111",
  18094=>"111111111",
  18095=>"000000001",
  18096=>"010000000",
  18097=>"111111111",
  18098=>"011111111",
  18099=>"111111111",
  18100=>"000100111",
  18101=>"000000101",
  18102=>"101100111",
  18103=>"111111011",
  18104=>"000001011",
  18105=>"111101111",
  18106=>"111000101",
  18107=>"110110111",
  18108=>"000000000",
  18109=>"000001101",
  18110=>"111111111",
  18111=>"001000011",
  18112=>"000111111",
  18113=>"111101110",
  18114=>"000000000",
  18115=>"001101111",
  18116=>"001000000",
  18117=>"111000000",
  18118=>"000000000",
  18119=>"110000000",
  18120=>"110111110",
  18121=>"001000000",
  18122=>"101000000",
  18123=>"111011110",
  18124=>"111110100",
  18125=>"000110000",
  18126=>"000001111",
  18127=>"110000100",
  18128=>"111000000",
  18129=>"000100101",
  18130=>"111110111",
  18131=>"000000000",
  18132=>"111111001",
  18133=>"101100100",
  18134=>"000000000",
  18135=>"011000111",
  18136=>"111111111",
  18137=>"110111101",
  18138=>"010010010",
  18139=>"000000000",
  18140=>"111111110",
  18141=>"111110000",
  18142=>"000111111",
  18143=>"000000110",
  18144=>"000001101",
  18145=>"011001111",
  18146=>"111111000",
  18147=>"000000000",
  18148=>"000000000",
  18149=>"111111111",
  18150=>"111011101",
  18151=>"011011110",
  18152=>"111111011",
  18153=>"110010011",
  18154=>"100000001",
  18155=>"000000100",
  18156=>"111111000",
  18157=>"111110111",
  18158=>"000000100",
  18159=>"000111111",
  18160=>"110100000",
  18161=>"000000100",
  18162=>"000111111",
  18163=>"110110000",
  18164=>"000000000",
  18165=>"100100101",
  18166=>"111011011",
  18167=>"110110000",
  18168=>"111111111",
  18169=>"110000100",
  18170=>"001001111",
  18171=>"000000000",
  18172=>"100101000",
  18173=>"000000001",
  18174=>"100100000",
  18175=>"111000000",
  18176=>"110110110",
  18177=>"001001101",
  18178=>"100111111",
  18179=>"010000001",
  18180=>"110000000",
  18181=>"001000000",
  18182=>"000000101",
  18183=>"001001111",
  18184=>"110111000",
  18185=>"000001000",
  18186=>"111111111",
  18187=>"100001001",
  18188=>"101101111",
  18189=>"000111010",
  18190=>"100111110",
  18191=>"110110111",
  18192=>"101001111",
  18193=>"000000000",
  18194=>"000000000",
  18195=>"111110110",
  18196=>"001111111",
  18197=>"111111000",
  18198=>"011001001",
  18199=>"111111111",
  18200=>"010000000",
  18201=>"111111111",
  18202=>"000001001",
  18203=>"011011000",
  18204=>"001000100",
  18205=>"011111111",
  18206=>"110111111",
  18207=>"010110111",
  18208=>"111111111",
  18209=>"000000000",
  18210=>"000000110",
  18211=>"101111111",
  18212=>"000000000",
  18213=>"000000001",
  18214=>"110111110",
  18215=>"111111111",
  18216=>"111111000",
  18217=>"100100000",
  18218=>"000000001",
  18219=>"000001001",
  18220=>"001000010",
  18221=>"110110110",
  18222=>"111110111",
  18223=>"101001001",
  18224=>"111111111",
  18225=>"111111001",
  18226=>"111111111",
  18227=>"111111111",
  18228=>"111111010",
  18229=>"001000000",
  18230=>"100100110",
  18231=>"001000000",
  18232=>"010111010",
  18233=>"111001111",
  18234=>"000000000",
  18235=>"111111110",
  18236=>"110110010",
  18237=>"111111100",
  18238=>"001111111",
  18239=>"110000011",
  18240=>"000000000",
  18241=>"110011001",
  18242=>"001001001",
  18243=>"100101101",
  18244=>"001111001",
  18245=>"000111111",
  18246=>"000001101",
  18247=>"111101001",
  18248=>"111001101",
  18249=>"000000111",
  18250=>"000000100",
  18251=>"011001001",
  18252=>"111111111",
  18253=>"000000000",
  18254=>"000100000",
  18255=>"110110111",
  18256=>"111111011",
  18257=>"110110110",
  18258=>"100000000",
  18259=>"100000000",
  18260=>"101001101",
  18261=>"111111111",
  18262=>"111000000",
  18263=>"000000000",
  18264=>"001001000",
  18265=>"111111111",
  18266=>"011111111",
  18267=>"011000010",
  18268=>"111010010",
  18269=>"001000000",
  18270=>"000000101",
  18271=>"110110100",
  18272=>"111111010",
  18273=>"010111110",
  18274=>"001001011",
  18275=>"001001000",
  18276=>"000001001",
  18277=>"111000000",
  18278=>"011111111",
  18279=>"111011001",
  18280=>"100000000",
  18281=>"000000100",
  18282=>"000000100",
  18283=>"001001011",
  18284=>"000110110",
  18285=>"111011000",
  18286=>"111101111",
  18287=>"000000100",
  18288=>"111110111",
  18289=>"010110110",
  18290=>"000111111",
  18291=>"111111101",
  18292=>"101001111",
  18293=>"100100111",
  18294=>"000000000",
  18295=>"000000111",
  18296=>"111111100",
  18297=>"111111111",
  18298=>"000000000",
  18299=>"111111111",
  18300=>"101100110",
  18301=>"111111111",
  18302=>"110111011",
  18303=>"111000101",
  18304=>"001001011",
  18305=>"111111111",
  18306=>"011110110",
  18307=>"000000000",
  18308=>"001000100",
  18309=>"111110100",
  18310=>"001000000",
  18311=>"111000000",
  18312=>"111111111",
  18313=>"110110111",
  18314=>"111110111",
  18315=>"111111110",
  18316=>"000000000",
  18317=>"110110000",
  18318=>"000000110",
  18319=>"000111001",
  18320=>"000100000",
  18321=>"000000000",
  18322=>"111111110",
  18323=>"010111111",
  18324=>"111111111",
  18325=>"000010000",
  18326=>"101100111",
  18327=>"100000011",
  18328=>"000000111",
  18329=>"111111111",
  18330=>"111111111",
  18331=>"011111111",
  18332=>"000000000",
  18333=>"010000101",
  18334=>"000001000",
  18335=>"000000001",
  18336=>"111111111",
  18337=>"011111011",
  18338=>"000000000",
  18339=>"001111000",
  18340=>"000000000",
  18341=>"111111111",
  18342=>"111110111",
  18343=>"110111110",
  18344=>"111110000",
  18345=>"000010011",
  18346=>"000000111",
  18347=>"110110111",
  18348=>"100111111",
  18349=>"000000110",
  18350=>"000110000",
  18351=>"111111101",
  18352=>"110010010",
  18353=>"101001000",
  18354=>"000100101",
  18355=>"011111111",
  18356=>"011111011",
  18357=>"111001001",
  18358=>"100111111",
  18359=>"100000101",
  18360=>"110111000",
  18361=>"000000010",
  18362=>"100011111",
  18363=>"000011010",
  18364=>"000000111",
  18365=>"111111111",
  18366=>"001000110",
  18367=>"111101001",
  18368=>"110001001",
  18369=>"001001101",
  18370=>"011000001",
  18371=>"001000000",
  18372=>"011000001",
  18373=>"011011100",
  18374=>"001000000",
  18375=>"011001001",
  18376=>"111100001",
  18377=>"000000000",
  18378=>"101000000",
  18379=>"000110111",
  18380=>"111111100",
  18381=>"000010000",
  18382=>"111001000",
  18383=>"000110111",
  18384=>"011110100",
  18385=>"111111111",
  18386=>"101000001",
  18387=>"101001111",
  18388=>"110111111",
  18389=>"000010011",
  18390=>"111100110",
  18391=>"000000000",
  18392=>"000000000",
  18393=>"101000000",
  18394=>"000000111",
  18395=>"110100000",
  18396=>"111000110",
  18397=>"111111001",
  18398=>"111111111",
  18399=>"100100110",
  18400=>"001000000",
  18401=>"111111111",
  18402=>"111111101",
  18403=>"001000000",
  18404=>"000000000",
  18405=>"000000111",
  18406=>"110011011",
  18407=>"100000000",
  18408=>"000000000",
  18409=>"000110110",
  18410=>"011000000",
  18411=>"100111000",
  18412=>"000000111",
  18413=>"111111110",
  18414=>"111111111",
  18415=>"000000111",
  18416=>"111111111",
  18417=>"000000001",
  18418=>"111110111",
  18419=>"111011001",
  18420=>"111111111",
  18421=>"000010000",
  18422=>"010111111",
  18423=>"110110110",
  18424=>"111111011",
  18425=>"111111001",
  18426=>"100000111",
  18427=>"101111111",
  18428=>"000000101",
  18429=>"000000000",
  18430=>"100000000",
  18431=>"000000011",
  18432=>"000000110",
  18433=>"110111111",
  18434=>"111111111",
  18435=>"101000110",
  18436=>"000000000",
  18437=>"111011000",
  18438=>"000000000",
  18439=>"111111111",
  18440=>"111111111",
  18441=>"000000111",
  18442=>"001001111",
  18443=>"000111111",
  18444=>"000000110",
  18445=>"000011111",
  18446=>"000000000",
  18447=>"000000000",
  18448=>"111111111",
  18449=>"000000110",
  18450=>"000000000",
  18451=>"111011000",
  18452=>"110000000",
  18453=>"000000101",
  18454=>"011000000",
  18455=>"000001111",
  18456=>"100000100",
  18457=>"101101111",
  18458=>"111111111",
  18459=>"001111111",
  18460=>"111111111",
  18461=>"001011001",
  18462=>"001000000",
  18463=>"100111111",
  18464=>"100111111",
  18465=>"101000000",
  18466=>"000011111",
  18467=>"000000000",
  18468=>"000000110",
  18469=>"111111000",
  18470=>"101000000",
  18471=>"011001111",
  18472=>"000100111",
  18473=>"000000000",
  18474=>"111000000",
  18475=>"110100111",
  18476=>"000010111",
  18477=>"000000000",
  18478=>"110110100",
  18479=>"000000010",
  18480=>"100000110",
  18481=>"000000000",
  18482=>"100000110",
  18483=>"000000000",
  18484=>"110111110",
  18485=>"001101000",
  18486=>"111111111",
  18487=>"111111111",
  18488=>"000000111",
  18489=>"111111111",
  18490=>"000000000",
  18491=>"111100000",
  18492=>"000000000",
  18493=>"101000000",
  18494=>"111111001",
  18495=>"111111000",
  18496=>"110000001",
  18497=>"100001000",
  18498=>"000110111",
  18499=>"100111111",
  18500=>"000000000",
  18501=>"000000000",
  18502=>"111101101",
  18503=>"101000000",
  18504=>"100000011",
  18505=>"000000000",
  18506=>"111111111",
  18507=>"100000111",
  18508=>"111100111",
  18509=>"000010111",
  18510=>"111000001",
  18511=>"111111000",
  18512=>"000000000",
  18513=>"000000000",
  18514=>"111110100",
  18515=>"000000000",
  18516=>"000000000",
  18517=>"000000000",
  18518=>"001000000",
  18519=>"111011011",
  18520=>"000000101",
  18521=>"000000110",
  18522=>"000000011",
  18523=>"111111001",
  18524=>"111010000",
  18525=>"000000000",
  18526=>"000000001",
  18527=>"111110111",
  18528=>"101111100",
  18529=>"000000000",
  18530=>"111000000",
  18531=>"000100111",
  18532=>"000111111",
  18533=>"000000000",
  18534=>"000000000",
  18535=>"010110010",
  18536=>"100110000",
  18537=>"000100111",
  18538=>"000000010",
  18539=>"000000000",
  18540=>"011000000",
  18541=>"111111111",
  18542=>"111111111",
  18543=>"011111011",
  18544=>"000000111",
  18545=>"000000111",
  18546=>"111111111",
  18547=>"111111111",
  18548=>"111010111",
  18549=>"010110000",
  18550=>"111111111",
  18551=>"000000001",
  18552=>"000000110",
  18553=>"000000111",
  18554=>"000000000",
  18555=>"111111111",
  18556=>"000001111",
  18557=>"111001001",
  18558=>"000000000",
  18559=>"000000111",
  18560=>"111011000",
  18561=>"100000110",
  18562=>"000000000",
  18563=>"000000000",
  18564=>"110111110",
  18565=>"000000000",
  18566=>"001000000",
  18567=>"111111110",
  18568=>"000000000",
  18569=>"000000000",
  18570=>"111100000",
  18571=>"000000000",
  18572=>"110000000",
  18573=>"000000000",
  18574=>"111111000",
  18575=>"100100111",
  18576=>"100000000",
  18577=>"000000000",
  18578=>"000000000",
  18579=>"111111101",
  18580=>"110111011",
  18581=>"000000000",
  18582=>"111111111",
  18583=>"000000000",
  18584=>"000000000",
  18585=>"111111111",
  18586=>"111000001",
  18587=>"000000000",
  18588=>"000000000",
  18589=>"001000000",
  18590=>"000000000",
  18591=>"101001000",
  18592=>"111111111",
  18593=>"111100000",
  18594=>"000011011",
  18595=>"000000011",
  18596=>"000000100",
  18597=>"111001001",
  18598=>"110111110",
  18599=>"000000000",
  18600=>"000000000",
  18601=>"110111111",
  18602=>"000000000",
  18603=>"111111000",
  18604=>"000000001",
  18605=>"011001000",
  18606=>"000000000",
  18607=>"000000000",
  18608=>"000011000",
  18609=>"111111111",
  18610=>"111111111",
  18611=>"111111111",
  18612=>"110110000",
  18613=>"000011111",
  18614=>"000000010",
  18615=>"000000000",
  18616=>"100000000",
  18617=>"100000110",
  18618=>"000000000",
  18619=>"110001111",
  18620=>"000000110",
  18621=>"111111111",
  18622=>"111111111",
  18623=>"001011110",
  18624=>"000011110",
  18625=>"000000000",
  18626=>"000000000",
  18627=>"000000000",
  18628=>"111111111",
  18629=>"110110110",
  18630=>"001110111",
  18631=>"100000100",
  18632=>"110110111",
  18633=>"000000111",
  18634=>"000000000",
  18635=>"111111111",
  18636=>"000000000",
  18637=>"111111111",
  18638=>"001011111",
  18639=>"000000000",
  18640=>"000000000",
  18641=>"000110011",
  18642=>"000000000",
  18643=>"000000001",
  18644=>"001001011",
  18645=>"000111111",
  18646=>"000000000",
  18647=>"000000000",
  18648=>"110111111",
  18649=>"110110111",
  18650=>"000000000",
  18651=>"000000011",
  18652=>"111111110",
  18653=>"100001111",
  18654=>"110000000",
  18655=>"110010000",
  18656=>"000000000",
  18657=>"000101111",
  18658=>"010000000",
  18659=>"000101111",
  18660=>"001000000",
  18661=>"100110111",
  18662=>"111111111",
  18663=>"000000000",
  18664=>"000011011",
  18665=>"111111001",
  18666=>"111000000",
  18667=>"000000000",
  18668=>"000000000",
  18669=>"011011111",
  18670=>"111110110",
  18671=>"111111001",
  18672=>"000101111",
  18673=>"111000000",
  18674=>"000000000",
  18675=>"000000000",
  18676=>"101011011",
  18677=>"111110110",
  18678=>"000000101",
  18679=>"000000100",
  18680=>"111111111",
  18681=>"000000000",
  18682=>"000000001",
  18683=>"000000000",
  18684=>"000000101",
  18685=>"111000001",
  18686=>"011000011",
  18687=>"001000001",
  18688=>"000000000",
  18689=>"001000000",
  18690=>"111111110",
  18691=>"000000001",
  18692=>"111111111",
  18693=>"100100111",
  18694=>"000000000",
  18695=>"000000101",
  18696=>"000000000",
  18697=>"111111111",
  18698=>"001001001",
  18699=>"000000000",
  18700=>"101001000",
  18701=>"000000101",
  18702=>"001101111",
  18703=>"000100111",
  18704=>"001000000",
  18705=>"000111111",
  18706=>"000000000",
  18707=>"000000110",
  18708=>"011011000",
  18709=>"111011000",
  18710=>"110111010",
  18711=>"111111000",
  18712=>"110100010",
  18713=>"001111111",
  18714=>"000000000",
  18715=>"000000000",
  18716=>"100110111",
  18717=>"111111110",
  18718=>"000000000",
  18719=>"010110110",
  18720=>"000000011",
  18721=>"110110100",
  18722=>"000000111",
  18723=>"010000000",
  18724=>"000000000",
  18725=>"000000000",
  18726=>"000000011",
  18727=>"111111111",
  18728=>"001001000",
  18729=>"000000000",
  18730=>"100100000",
  18731=>"111111010",
  18732=>"000111111",
  18733=>"000000000",
  18734=>"101000001",
  18735=>"000001001",
  18736=>"111000000",
  18737=>"000011111",
  18738=>"000000000",
  18739=>"000001000",
  18740=>"000000000",
  18741=>"001100110",
  18742=>"000000111",
  18743=>"000000000",
  18744=>"000000000",
  18745=>"111111000",
  18746=>"111111111",
  18747=>"111111111",
  18748=>"111111111",
  18749=>"000000000",
  18750=>"111111111",
  18751=>"111000000",
  18752=>"000000000",
  18753=>"000000000",
  18754=>"001111101",
  18755=>"000000000",
  18756=>"100000000",
  18757=>"000001011",
  18758=>"010011111",
  18759=>"001000000",
  18760=>"111111111",
  18761=>"111111111",
  18762=>"111100111",
  18763=>"111111000",
  18764=>"000111111",
  18765=>"000000000",
  18766=>"111111111",
  18767=>"110101100",
  18768=>"111111111",
  18769=>"000001111",
  18770=>"000111111",
  18771=>"110111111",
  18772=>"000000000",
  18773=>"001011011",
  18774=>"111111111",
  18775=>"111111111",
  18776=>"111110000",
  18777=>"111000000",
  18778=>"110111010",
  18779=>"111101100",
  18780=>"000000001",
  18781=>"111111111",
  18782=>"111111000",
  18783=>"000000100",
  18784=>"111111111",
  18785=>"010100000",
  18786=>"000000000",
  18787=>"111111111",
  18788=>"111111110",
  18789=>"000100111",
  18790=>"000000000",
  18791=>"000000100",
  18792=>"111111000",
  18793=>"000000000",
  18794=>"111101111",
  18795=>"111111111",
  18796=>"001000000",
  18797=>"000000000",
  18798=>"000010000",
  18799=>"000000000",
  18800=>"111111111",
  18801=>"111111111",
  18802=>"000000000",
  18803=>"000000000",
  18804=>"000000000",
  18805=>"111111111",
  18806=>"000000101",
  18807=>"000000000",
  18808=>"111111111",
  18809=>"111111111",
  18810=>"000000000",
  18811=>"111000011",
  18812=>"000110110",
  18813=>"110110111",
  18814=>"000000000",
  18815=>"111111111",
  18816=>"000000000",
  18817=>"110010000",
  18818=>"011000011",
  18819=>"011000000",
  18820=>"000000011",
  18821=>"000000000",
  18822=>"100001111",
  18823=>"111101001",
  18824=>"000000000",
  18825=>"111111111",
  18826=>"110111111",
  18827=>"110110111",
  18828=>"111111111",
  18829=>"000000000",
  18830=>"011000000",
  18831=>"111111000",
  18832=>"000000000",
  18833=>"011111111",
  18834=>"111111111",
  18835=>"111111111",
  18836=>"000000000",
  18837=>"000000000",
  18838=>"000000000",
  18839=>"000000100",
  18840=>"100000000",
  18841=>"111111111",
  18842=>"000000111",
  18843=>"000111111",
  18844=>"000111111",
  18845=>"000000111",
  18846=>"000000000",
  18847=>"111111111",
  18848=>"000000000",
  18849=>"111111001",
  18850=>"110100101",
  18851=>"111111111",
  18852=>"111111111",
  18853=>"111111111",
  18854=>"000000000",
  18855=>"111000111",
  18856=>"000000000",
  18857=>"000000000",
  18858=>"001001000",
  18859=>"000110010",
  18860=>"000000000",
  18861=>"000000000",
  18862=>"110100101",
  18863=>"011011111",
  18864=>"000000011",
  18865=>"000000000",
  18866=>"100000101",
  18867=>"000000111",
  18868=>"111111111",
  18869=>"111111111",
  18870=>"111111111",
  18871=>"000110110",
  18872=>"000111000",
  18873=>"110110111",
  18874=>"000110110",
  18875=>"111111001",
  18876=>"111000000",
  18877=>"000000110",
  18878=>"011000000",
  18879=>"110110010",
  18880=>"000001011",
  18881=>"001000011",
  18882=>"000000000",
  18883=>"000000000",
  18884=>"000000000",
  18885=>"000000111",
  18886=>"010001111",
  18887=>"000000000",
  18888=>"000000000",
  18889=>"000111011",
  18890=>"000000111",
  18891=>"000000111",
  18892=>"000000000",
  18893=>"000010000",
  18894=>"000000000",
  18895=>"100110111",
  18896=>"000000000",
  18897=>"111111111",
  18898=>"000001111",
  18899=>"111111111",
  18900=>"000000000",
  18901=>"111111111",
  18902=>"111111111",
  18903=>"111010011",
  18904=>"100000111",
  18905=>"111101001",
  18906=>"111111111",
  18907=>"111100111",
  18908=>"111011011",
  18909=>"111111111",
  18910=>"001000000",
  18911=>"111111111",
  18912=>"011010001",
  18913=>"000000000",
  18914=>"000000000",
  18915=>"111111000",
  18916=>"111111111",
  18917=>"000000001",
  18918=>"111111110",
  18919=>"111000000",
  18920=>"000000110",
  18921=>"101001101",
  18922=>"111111111",
  18923=>"000000001",
  18924=>"111000000",
  18925=>"000000000",
  18926=>"011011000",
  18927=>"000000000",
  18928=>"111111111",
  18929=>"000000000",
  18930=>"111111111",
  18931=>"000000111",
  18932=>"111100000",
  18933=>"000000000",
  18934=>"111111111",
  18935=>"000111111",
  18936=>"000000111",
  18937=>"000000001",
  18938=>"000100111",
  18939=>"000000000",
  18940=>"001101111",
  18941=>"111111111",
  18942=>"111111000",
  18943=>"000000000",
  18944=>"110000000",
  18945=>"000111110",
  18946=>"000000000",
  18947=>"111111000",
  18948=>"000010000",
  18949=>"111110000",
  18950=>"000000000",
  18951=>"000000000",
  18952=>"110000000",
  18953=>"110010000",
  18954=>"111000000",
  18955=>"000001111",
  18956=>"011111111",
  18957=>"000000000",
  18958=>"000000000",
  18959=>"000100100",
  18960=>"000000000",
  18961=>"000000000",
  18962=>"000000000",
  18963=>"010000110",
  18964=>"111000000",
  18965=>"110111111",
  18966=>"001000001",
  18967=>"100110111",
  18968=>"000001000",
  18969=>"000011010",
  18970=>"000000111",
  18971=>"111110110",
  18972=>"111111111",
  18973=>"000000000",
  18974=>"010111001",
  18975=>"010000100",
  18976=>"010110000",
  18977=>"000000000",
  18978=>"111111111",
  18979=>"111111111",
  18980=>"111111111",
  18981=>"000001111",
  18982=>"111111001",
  18983=>"000010111",
  18984=>"111001010",
  18985=>"011111000",
  18986=>"111111010",
  18987=>"100100000",
  18988=>"001000000",
  18989=>"101101000",
  18990=>"011111101",
  18991=>"111101111",
  18992=>"001111011",
  18993=>"000000000",
  18994=>"000000110",
  18995=>"000000000",
  18996=>"000000001",
  18997=>"000000001",
  18998=>"111111111",
  18999=>"000000000",
  19000=>"111111111",
  19001=>"001011111",
  19002=>"111111110",
  19003=>"000000000",
  19004=>"111010000",
  19005=>"111111111",
  19006=>"011000111",
  19007=>"111111110",
  19008=>"011111111",
  19009=>"110101111",
  19010=>"111001000",
  19011=>"111111111",
  19012=>"110011000",
  19013=>"111110110",
  19014=>"011001111",
  19015=>"000000000",
  19016=>"110100100",
  19017=>"111111111",
  19018=>"110000000",
  19019=>"000000111",
  19020=>"000000000",
  19021=>"000000000",
  19022=>"000000000",
  19023=>"011010111",
  19024=>"000000000",
  19025=>"111101000",
  19026=>"111111111",
  19027=>"011011000",
  19028=>"000000000",
  19029=>"000110100",
  19030=>"110110110",
  19031=>"111100000",
  19032=>"011110000",
  19033=>"100000000",
  19034=>"001101111",
  19035=>"001101011",
  19036=>"111111000",
  19037=>"111001101",
  19038=>"111111111",
  19039=>"111100110",
  19040=>"111111111",
  19041=>"100000000",
  19042=>"011111011",
  19043=>"000000000",
  19044=>"000000000",
  19045=>"000000000",
  19046=>"111111111",
  19047=>"000000011",
  19048=>"111111111",
  19049=>"111111111",
  19050=>"000000001",
  19051=>"000000000",
  19052=>"111111111",
  19053=>"000000100",
  19054=>"100000000",
  19055=>"010000000",
  19056=>"001111111",
  19057=>"000000001",
  19058=>"000001001",
  19059=>"000100000",
  19060=>"000000000",
  19061=>"111111001",
  19062=>"111110111",
  19063=>"101111111",
  19064=>"010111111",
  19065=>"111111100",
  19066=>"000000000",
  19067=>"100000010",
  19068=>"011000000",
  19069=>"000000000",
  19070=>"000000000",
  19071=>"111110111",
  19072=>"000000000",
  19073=>"000010000",
  19074=>"101000000",
  19075=>"011100000",
  19076=>"000011011",
  19077=>"110100111",
  19078=>"111111111",
  19079=>"010110111",
  19080=>"000000000",
  19081=>"111111011",
  19082=>"000101000",
  19083=>"001000100",
  19084=>"111111000",
  19085=>"000000000",
  19086=>"000000000",
  19087=>"111111111",
  19088=>"000001001",
  19089=>"100000000",
  19090=>"111111110",
  19091=>"000111110",
  19092=>"001111111",
  19093=>"100111011",
  19094=>"000000000",
  19095=>"111001000",
  19096=>"111001001",
  19097=>"111111000",
  19098=>"010000000",
  19099=>"000100110",
  19100=>"111111000",
  19101=>"001000000",
  19102=>"000000000",
  19103=>"000000000",
  19104=>"000000000",
  19105=>"000100000",
  19106=>"111111111",
  19107=>"111001001",
  19108=>"000000011",
  19109=>"001001101",
  19110=>"111000000",
  19111=>"100100100",
  19112=>"110011000",
  19113=>"111011000",
  19114=>"110110100",
  19115=>"111111111",
  19116=>"001001011",
  19117=>"011011011",
  19118=>"110110111",
  19119=>"000100001",
  19120=>"111111110",
  19121=>"010000100",
  19122=>"111100000",
  19123=>"000000000",
  19124=>"111111111",
  19125=>"000000000",
  19126=>"010011111",
  19127=>"111111111",
  19128=>"000110110",
  19129=>"000000000",
  19130=>"000000000",
  19131=>"101111111",
  19132=>"000000111",
  19133=>"111001111",
  19134=>"111111000",
  19135=>"111011111",
  19136=>"111011111",
  19137=>"111111111",
  19138=>"001000000",
  19139=>"011111111",
  19140=>"110110110",
  19141=>"100000000",
  19142=>"011000001",
  19143=>"000111111",
  19144=>"000000111",
  19145=>"100111101",
  19146=>"001001000",
  19147=>"011000000",
  19148=>"111101111",
  19149=>"000000011",
  19150=>"111011111",
  19151=>"000000010",
  19152=>"000000110",
  19153=>"000000000",
  19154=>"000011000",
  19155=>"100000111",
  19156=>"111111010",
  19157=>"111111111",
  19158=>"000000000",
  19159=>"000000000",
  19160=>"010010110",
  19161=>"111111011",
  19162=>"000000000",
  19163=>"011011000",
  19164=>"111111111",
  19165=>"100000001",
  19166=>"101111111",
  19167=>"000010001",
  19168=>"111011001",
  19169=>"111011111",
  19170=>"100000100",
  19171=>"000110110",
  19172=>"000000000",
  19173=>"111111111",
  19174=>"000000000",
  19175=>"111111111",
  19176=>"101111111",
  19177=>"000000000",
  19178=>"111111001",
  19179=>"000000000",
  19180=>"001001000",
  19181=>"111111110",
  19182=>"000110111",
  19183=>"000000000",
  19184=>"000000010",
  19185=>"000000000",
  19186=>"011001101",
  19187=>"011111000",
  19188=>"111111111",
  19189=>"111111111",
  19190=>"111011011",
  19191=>"111011000",
  19192=>"000000000",
  19193=>"000011011",
  19194=>"111111000",
  19195=>"111111111",
  19196=>"000011001",
  19197=>"000000011",
  19198=>"100000100",
  19199=>"111000000",
  19200=>"111111111",
  19201=>"111011011",
  19202=>"000000001",
  19203=>"100100000",
  19204=>"000000100",
  19205=>"011000000",
  19206=>"011000000",
  19207=>"100110001",
  19208=>"000001000",
  19209=>"000000111",
  19210=>"000000000",
  19211=>"110111111",
  19212=>"111101000",
  19213=>"100100110",
  19214=>"111111111",
  19215=>"111111001",
  19216=>"111111111",
  19217=>"000010100",
  19218=>"000000000",
  19219=>"000000000",
  19220=>"000000000",
  19221=>"111111111",
  19222=>"011100100",
  19223=>"000000001",
  19224=>"110111011",
  19225=>"000000000",
  19226=>"111101111",
  19227=>"110110000",
  19228=>"000111010",
  19229=>"000010000",
  19230=>"100100100",
  19231=>"100100000",
  19232=>"011111110",
  19233=>"000011000",
  19234=>"111111111",
  19235=>"001001001",
  19236=>"000000000",
  19237=>"111111111",
  19238=>"001000000",
  19239=>"110110000",
  19240=>"011000111",
  19241=>"000000000",
  19242=>"111111111",
  19243=>"111111111",
  19244=>"111110110",
  19245=>"101001001",
  19246=>"100000001",
  19247=>"010111111",
  19248=>"000100010",
  19249=>"000000000",
  19250=>"111111111",
  19251=>"111000000",
  19252=>"000000000",
  19253=>"111000100",
  19254=>"111000001",
  19255=>"111111111",
  19256=>"000000000",
  19257=>"000000000",
  19258=>"000000001",
  19259=>"101111110",
  19260=>"000000000",
  19261=>"001000100",
  19262=>"000111110",
  19263=>"111111000",
  19264=>"000000000",
  19265=>"000000000",
  19266=>"011111001",
  19267=>"000000011",
  19268=>"000001011",
  19269=>"111000000",
  19270=>"111111010",
  19271=>"000000000",
  19272=>"000000000",
  19273=>"000111111",
  19274=>"010100100",
  19275=>"100000000",
  19276=>"111111111",
  19277=>"111000001",
  19278=>"111111111",
  19279=>"000000000",
  19280=>"010000010",
  19281=>"110111101",
  19282=>"111111000",
  19283=>"011111111",
  19284=>"000000000",
  19285=>"000000000",
  19286=>"111111000",
  19287=>"001000101",
  19288=>"000111111",
  19289=>"000000000",
  19290=>"111111111",
  19291=>"111101111",
  19292=>"111011000",
  19293=>"000000001",
  19294=>"010111000",
  19295=>"111011011",
  19296=>"010010000",
  19297=>"000000000",
  19298=>"000000001",
  19299=>"000111111",
  19300=>"111011011",
  19301=>"000000000",
  19302=>"111111111",
  19303=>"110110011",
  19304=>"001011111",
  19305=>"000000111",
  19306=>"000100111",
  19307=>"000111111",
  19308=>"100000000",
  19309=>"001011010",
  19310=>"000000000",
  19311=>"111111111",
  19312=>"000000001",
  19313=>"000000000",
  19314=>"000000111",
  19315=>"111111111",
  19316=>"111111111",
  19317=>"000000010",
  19318=>"000011010",
  19319=>"111111111",
  19320=>"000000000",
  19321=>"001000000",
  19322=>"111111111",
  19323=>"000000000",
  19324=>"110000000",
  19325=>"000000000",
  19326=>"100111111",
  19327=>"111111111",
  19328=>"000000000",
  19329=>"000000111",
  19330=>"000011010",
  19331=>"111111111",
  19332=>"111111111",
  19333=>"111000001",
  19334=>"011000000",
  19335=>"111111000",
  19336=>"111111111",
  19337=>"011000000",
  19338=>"111111111",
  19339=>"111111111",
  19340=>"110110000",
  19341=>"000000000",
  19342=>"111111111",
  19343=>"011111100",
  19344=>"001000111",
  19345=>"000110110",
  19346=>"111111000",
  19347=>"000110010",
  19348=>"111000000",
  19349=>"111111101",
  19350=>"000110000",
  19351=>"010010000",
  19352=>"011001000",
  19353=>"111111111",
  19354=>"011000110",
  19355=>"000000000",
  19356=>"111111110",
  19357=>"001000000",
  19358=>"100111111",
  19359=>"111000000",
  19360=>"000000111",
  19361=>"001001001",
  19362=>"111111110",
  19363=>"111111111",
  19364=>"111111111",
  19365=>"000000000",
  19366=>"111111111",
  19367=>"000110000",
  19368=>"001111111",
  19369=>"010010000",
  19370=>"001001000",
  19371=>"111000000",
  19372=>"111111000",
  19373=>"111111111",
  19374=>"011011111",
  19375=>"000000100",
  19376=>"100000100",
  19377=>"111111111",
  19378=>"010000110",
  19379=>"111111111",
  19380=>"001000000",
  19381=>"111101000",
  19382=>"110100110",
  19383=>"010011011",
  19384=>"000001111",
  19385=>"010111000",
  19386=>"101111110",
  19387=>"100100111",
  19388=>"000000000",
  19389=>"001011011",
  19390=>"000000000",
  19391=>"001001001",
  19392=>"111001000",
  19393=>"111111111",
  19394=>"000001111",
  19395=>"000000111",
  19396=>"110000000",
  19397=>"011111011",
  19398=>"000011111",
  19399=>"011011000",
  19400=>"001000000",
  19401=>"111111111",
  19402=>"011111111",
  19403=>"011000111",
  19404=>"000110110",
  19405=>"111111111",
  19406=>"111111111",
  19407=>"111111111",
  19408=>"000000000",
  19409=>"100100100",
  19410=>"000000000",
  19411=>"011011010",
  19412=>"001001001",
  19413=>"000011111",
  19414=>"000000111",
  19415=>"100110100",
  19416=>"101111111",
  19417=>"000100000",
  19418=>"110111111",
  19419=>"110111111",
  19420=>"000000000",
  19421=>"111111100",
  19422=>"000110110",
  19423=>"010011011",
  19424=>"000010111",
  19425=>"010000010",
  19426=>"000000000",
  19427=>"111111111",
  19428=>"000000000",
  19429=>"111000100",
  19430=>"000000000",
  19431=>"110110000",
  19432=>"111111111",
  19433=>"000000111",
  19434=>"000010111",
  19435=>"001101000",
  19436=>"111110111",
  19437=>"111111110",
  19438=>"000000000",
  19439=>"000000100",
  19440=>"000001010",
  19441=>"111111111",
  19442=>"000000000",
  19443=>"110000000",
  19444=>"001001001",
  19445=>"111111101",
  19446=>"101111111",
  19447=>"000010011",
  19448=>"111111111",
  19449=>"111111110",
  19450=>"000000000",
  19451=>"111111111",
  19452=>"111011101",
  19453=>"100100100",
  19454=>"001101111",
  19455=>"000000000",
  19456=>"111110111",
  19457=>"111000001",
  19458=>"010000100",
  19459=>"111010111",
  19460=>"000000001",
  19461=>"000000100",
  19462=>"000000000",
  19463=>"111111111",
  19464=>"111111111",
  19465=>"111111100",
  19466=>"111111101",
  19467=>"011000000",
  19468=>"000110111",
  19469=>"111011111",
  19470=>"001000000",
  19471=>"111111111",
  19472=>"111111111",
  19473=>"111111111",
  19474=>"010000111",
  19475=>"000000000",
  19476=>"010100100",
  19477=>"011011011",
  19478=>"000000000",
  19479=>"100110111",
  19480=>"111111111",
  19481=>"111000000",
  19482=>"000000000",
  19483=>"111110110",
  19484=>"111000000",
  19485=>"001000101",
  19486=>"111111110",
  19487=>"001000011",
  19488=>"000000101",
  19489=>"000000000",
  19490=>"111111101",
  19491=>"111000000",
  19492=>"111111011",
  19493=>"100000100",
  19494=>"010011101",
  19495=>"001000000",
  19496=>"111000000",
  19497=>"010011000",
  19498=>"011001111",
  19499=>"111111111",
  19500=>"010000111",
  19501=>"100000010",
  19502=>"100111001",
  19503=>"010011001",
  19504=>"110100111",
  19505=>"110010000",
  19506=>"111101101",
  19507=>"000100100",
  19508=>"000000000",
  19509=>"000110110",
  19510=>"010010000",
  19511=>"100001101",
  19512=>"011011000",
  19513=>"000010000",
  19514=>"000000000",
  19515=>"111111111",
  19516=>"101000000",
  19517=>"011000101",
  19518=>"001001111",
  19519=>"111111111",
  19520=>"000011011",
  19521=>"111111111",
  19522=>"111000000",
  19523=>"000000000",
  19524=>"000000011",
  19525=>"111111011",
  19526=>"111000000",
  19527=>"111111111",
  19528=>"000000000",
  19529=>"000000111",
  19530=>"000000000",
  19531=>"000101100",
  19532=>"000011111",
  19533=>"000000000",
  19534=>"111101100",
  19535=>"011111000",
  19536=>"110111000",
  19537=>"111111111",
  19538=>"000100100",
  19539=>"110110000",
  19540=>"000000111",
  19541=>"000000000",
  19542=>"000000001",
  19543=>"111111111",
  19544=>"111111011",
  19545=>"000100100",
  19546=>"000011000",
  19547=>"000000101",
  19548=>"000000000",
  19549=>"111111111",
  19550=>"000111111",
  19551=>"000000000",
  19552=>"000000000",
  19553=>"111000000",
  19554=>"111111101",
  19555=>"000000000",
  19556=>"110110000",
  19557=>"111111111",
  19558=>"111111000",
  19559=>"111111111",
  19560=>"000010111",
  19561=>"000110000",
  19562=>"000110010",
  19563=>"000000000",
  19564=>"010100111",
  19565=>"000000100",
  19566=>"111111101",
  19567=>"111110000",
  19568=>"000000000",
  19569=>"000011011",
  19570=>"111101100",
  19571=>"111111111",
  19572=>"111111111",
  19573=>"000000000",
  19574=>"111111111",
  19575=>"000100000",
  19576=>"001000000",
  19577=>"110111111",
  19578=>"000100000",
  19579=>"101101101",
  19580=>"000000110",
  19581=>"111101001",
  19582=>"000000000",
  19583=>"111111111",
  19584=>"000000111",
  19585=>"000000000",
  19586=>"111111001",
  19587=>"011111111",
  19588=>"100100000",
  19589=>"111111111",
  19590=>"000000000",
  19591=>"000000000",
  19592=>"111011011",
  19593=>"110000100",
  19594=>"110000000",
  19595=>"111111111",
  19596=>"111111111",
  19597=>"111111111",
  19598=>"111111111",
  19599=>"000111111",
  19600=>"000000000",
  19601=>"101000101",
  19602=>"000011111",
  19603=>"111111110",
  19604=>"000110000",
  19605=>"111111111",
  19606=>"110111111",
  19607=>"111111111",
  19608=>"111111110",
  19609=>"111011001",
  19610=>"111111111",
  19611=>"000000000",
  19612=>"111111100",
  19613=>"000000001",
  19614=>"011111111",
  19615=>"111111111",
  19616=>"000010000",
  19617=>"000000100",
  19618=>"000000000",
  19619=>"111111111",
  19620=>"000000000",
  19621=>"111111111",
  19622=>"111111010",
  19623=>"111111011",
  19624=>"011010111",
  19625=>"000000000",
  19626=>"000000000",
  19627=>"000000000",
  19628=>"111001001",
  19629=>"011101101",
  19630=>"000000000",
  19631=>"010001000",
  19632=>"111111010",
  19633=>"101100101",
  19634=>"010111111",
  19635=>"111111111",
  19636=>"111111111",
  19637=>"111111110",
  19638=>"000000000",
  19639=>"110000000",
  19640=>"111111111",
  19641=>"000000000",
  19642=>"000111111",
  19643=>"000000110",
  19644=>"110110110",
  19645=>"111011000",
  19646=>"001000000",
  19647=>"111111011",
  19648=>"001111111",
  19649=>"101001001",
  19650=>"110100000",
  19651=>"000000001",
  19652=>"011011000",
  19653=>"111011110",
  19654=>"010000110",
  19655=>"010000101",
  19656=>"111111110",
  19657=>"111101111",
  19658=>"111101001",
  19659=>"000000000",
  19660=>"001000000",
  19661=>"000011011",
  19662=>"100100010",
  19663=>"111110111",
  19664=>"001011111",
  19665=>"000000000",
  19666=>"001001111",
  19667=>"101000100",
  19668=>"000000000",
  19669=>"000000001",
  19670=>"110110110",
  19671=>"111111100",
  19672=>"000111100",
  19673=>"011111000",
  19674=>"111100100",
  19675=>"111111111",
  19676=>"111111111",
  19677=>"000000001",
  19678=>"000000000",
  19679=>"111011100",
  19680=>"000000000",
  19681=>"000000010",
  19682=>"111111111",
  19683=>"011111111",
  19684=>"001001000",
  19685=>"111111111",
  19686=>"000000000",
  19687=>"000000000",
  19688=>"000011111",
  19689=>"000000000",
  19690=>"111111111",
  19691=>"000101111",
  19692=>"110111111",
  19693=>"111011000",
  19694=>"100000000",
  19695=>"100100110",
  19696=>"110000010",
  19697=>"000000000",
  19698=>"111111111",
  19699=>"011011000",
  19700=>"011011000",
  19701=>"000000000",
  19702=>"111111111",
  19703=>"000010011",
  19704=>"000000000",
  19705=>"100000000",
  19706=>"111111111",
  19707=>"110100111",
  19708=>"001001001",
  19709=>"000000000",
  19710=>"111111110",
  19711=>"000001010",
  19712=>"111011001",
  19713=>"111111100",
  19714=>"111001111",
  19715=>"000000110",
  19716=>"111100100",
  19717=>"111000000",
  19718=>"000000000",
  19719=>"000100111",
  19720=>"111111111",
  19721=>"000001000",
  19722=>"000000000",
  19723=>"001101111",
  19724=>"010011111",
  19725=>"000111111",
  19726=>"000000000",
  19727=>"111011000",
  19728=>"111111111",
  19729=>"000000000",
  19730=>"111100111",
  19731=>"101010000",
  19732=>"110100000",
  19733=>"000101111",
  19734=>"011110110",
  19735=>"000000000",
  19736=>"111000000",
  19737=>"000010000",
  19738=>"111111111",
  19739=>"111111111",
  19740=>"111111111",
  19741=>"111111111",
  19742=>"111111000",
  19743=>"011101101",
  19744=>"001011000",
  19745=>"000000000",
  19746=>"000000111",
  19747=>"111111111",
  19748=>"111111111",
  19749=>"001001001",
  19750=>"000111111",
  19751=>"000000000",
  19752=>"000110111",
  19753=>"100111110",
  19754=>"111111101",
  19755=>"000110110",
  19756=>"000000000",
  19757=>"011011001",
  19758=>"111111111",
  19759=>"000000000",
  19760=>"111111111",
  19761=>"000000000",
  19762=>"111111111",
  19763=>"000000000",
  19764=>"001000110",
  19765=>"111111111",
  19766=>"000000000",
  19767=>"111111111",
  19768=>"000001001",
  19769=>"011111111",
  19770=>"000000010",
  19771=>"000010111",
  19772=>"111111111",
  19773=>"000111000",
  19774=>"000000001",
  19775=>"001101101",
  19776=>"000000000",
  19777=>"111111111",
  19778=>"111111111",
  19779=>"000101111",
  19780=>"111111000",
  19781=>"110110100",
  19782=>"000000000",
  19783=>"111111111",
  19784=>"000000000",
  19785=>"111100100",
  19786=>"111111101",
  19787=>"000001101",
  19788=>"111011000",
  19789=>"011001000",
  19790=>"000000000",
  19791=>"011011011",
  19792=>"100111110",
  19793=>"000000000",
  19794=>"100100001",
  19795=>"101001111",
  19796=>"000110111",
  19797=>"000000011",
  19798=>"000000000",
  19799=>"000000000",
  19800=>"000101111",
  19801=>"111111000",
  19802=>"111111111",
  19803=>"110010111",
  19804=>"111111111",
  19805=>"000000000",
  19806=>"000000101",
  19807=>"011111000",
  19808=>"000000000",
  19809=>"010010000",
  19810=>"111001001",
  19811=>"111111111",
  19812=>"110111111",
  19813=>"011011001",
  19814=>"111111111",
  19815=>"000001001",
  19816=>"000000001",
  19817=>"110110111",
  19818=>"000000000",
  19819=>"011111111",
  19820=>"111111111",
  19821=>"111111111",
  19822=>"000000000",
  19823=>"000000000",
  19824=>"011000100",
  19825=>"100000000",
  19826=>"001000000",
  19827=>"011011011",
  19828=>"010000000",
  19829=>"000100000",
  19830=>"111111001",
  19831=>"000000000",
  19832=>"000000000",
  19833=>"000000000",
  19834=>"111101111",
  19835=>"000000000",
  19836=>"001000000",
  19837=>"000000100",
  19838=>"111101111",
  19839=>"000000111",
  19840=>"111110110",
  19841=>"010010101",
  19842=>"111010100",
  19843=>"111111111",
  19844=>"100100111",
  19845=>"000000000",
  19846=>"001011111",
  19847=>"100100111",
  19848=>"000000001",
  19849=>"011011011",
  19850=>"110110111",
  19851=>"000000000",
  19852=>"111111111",
  19853=>"111010000",
  19854=>"010010110",
  19855=>"000000000",
  19856=>"111111111",
  19857=>"111000000",
  19858=>"111111111",
  19859=>"111111111",
  19860=>"000000000",
  19861=>"000000110",
  19862=>"111101111",
  19863=>"111111011",
  19864=>"110111000",
  19865=>"111000111",
  19866=>"000000000",
  19867=>"100000101",
  19868=>"111111111",
  19869=>"111111011",
  19870=>"011111010",
  19871=>"000000000",
  19872=>"000000010",
  19873=>"110110110",
  19874=>"011000011",
  19875=>"010110111",
  19876=>"000100110",
  19877=>"111011011",
  19878=>"000000000",
  19879=>"111111111",
  19880=>"010000100",
  19881=>"000000000",
  19882=>"111111010",
  19883=>"000000000",
  19884=>"100101111",
  19885=>"011111010",
  19886=>"000000111",
  19887=>"000100101",
  19888=>"111111000",
  19889=>"001101111",
  19890=>"010001001",
  19891=>"000000000",
  19892=>"111111000",
  19893=>"111011001",
  19894=>"000100111",
  19895=>"111000000",
  19896=>"000110111",
  19897=>"010011001",
  19898=>"000000010",
  19899=>"111111111",
  19900=>"000111111",
  19901=>"111111101",
  19902=>"000000100",
  19903=>"010010000",
  19904=>"011110000",
  19905=>"111111111",
  19906=>"010010010",
  19907=>"000111110",
  19908=>"000011001",
  19909=>"010111011",
  19910=>"011011010",
  19911=>"000011000",
  19912=>"000000000",
  19913=>"011111010",
  19914=>"111000001",
  19915=>"001111111",
  19916=>"010001000",
  19917=>"000110100",
  19918=>"001001001",
  19919=>"010000100",
  19920=>"110100100",
  19921=>"011011010",
  19922=>"110000010",
  19923=>"000000000",
  19924=>"000000001",
  19925=>"000000100",
  19926=>"000100100",
  19927=>"011000000",
  19928=>"001111101",
  19929=>"000000000",
  19930=>"000000000",
  19931=>"011111111",
  19932=>"111111111",
  19933=>"000000000",
  19934=>"111111111",
  19935=>"111111101",
  19936=>"000000000",
  19937=>"011000101",
  19938=>"111111000",
  19939=>"000000100",
  19940=>"000000000",
  19941=>"100000010",
  19942=>"000100111",
  19943=>"001111111",
  19944=>"011001101",
  19945=>"000001011",
  19946=>"111111111",
  19947=>"110110100",
  19948=>"010001011",
  19949=>"101100101",
  19950=>"111011000",
  19951=>"111011000",
  19952=>"011000000",
  19953=>"101111111",
  19954=>"111111111",
  19955=>"000000000",
  19956=>"000001111",
  19957=>"111000111",
  19958=>"000000111",
  19959=>"000000000",
  19960=>"000000000",
  19961=>"000000000",
  19962=>"000000000",
  19963=>"000000000",
  19964=>"111001001",
  19965=>"100010111",
  19966=>"000010001",
  19967=>"110110111",
  19968=>"111111111",
  19969=>"111110000",
  19970=>"101100000",
  19971=>"110010000",
  19972=>"111011110",
  19973=>"000100111",
  19974=>"111111111",
  19975=>"111111111",
  19976=>"111010000",
  19977=>"010010001",
  19978=>"000000011",
  19979=>"111101101",
  19980=>"011011011",
  19981=>"001111111",
  19982=>"000000001",
  19983=>"000000000",
  19984=>"000100101",
  19985=>"001001000",
  19986=>"000000000",
  19987=>"001001111",
  19988=>"111101111",
  19989=>"111000001",
  19990=>"111111000",
  19991=>"110111111",
  19992=>"000000000",
  19993=>"110110111",
  19994=>"101101111",
  19995=>"111111111",
  19996=>"101001001",
  19997=>"000000010",
  19998=>"001111011",
  19999=>"000011011",
  20000=>"111111111",
  20001=>"110111110",
  20002=>"000001111",
  20003=>"111111111",
  20004=>"111000000",
  20005=>"000000000",
  20006=>"000000000",
  20007=>"000000000",
  20008=>"111111111",
  20009=>"111111111",
  20010=>"001001111",
  20011=>"110111110",
  20012=>"010000000",
  20013=>"000000110",
  20014=>"110010000",
  20015=>"011111111",
  20016=>"111111111",
  20017=>"100100100",
  20018=>"100100100",
  20019=>"000000011",
  20020=>"000000000",
  20021=>"110110110",
  20022=>"111111111",
  20023=>"011111110",
  20024=>"000000000",
  20025=>"000000000",
  20026=>"111111000",
  20027=>"000000111",
  20028=>"000000111",
  20029=>"000000000",
  20030=>"111111111",
  20031=>"000000111",
  20032=>"111101100",
  20033=>"000000100",
  20034=>"000011111",
  20035=>"111111111",
  20036=>"011111111",
  20037=>"001001101",
  20038=>"000000000",
  20039=>"111111000",
  20040=>"111111011",
  20041=>"111111111",
  20042=>"111111111",
  20043=>"001001000",
  20044=>"111100000",
  20045=>"110110000",
  20046=>"001011001",
  20047=>"000000111",
  20048=>"000111111",
  20049=>"110111111",
  20050=>"000000100",
  20051=>"000000000",
  20052=>"000000000",
  20053=>"101111111",
  20054=>"100000000",
  20055=>"111111110",
  20056=>"100000000",
  20057=>"101000001",
  20058=>"000000100",
  20059=>"000000001",
  20060=>"111111100",
  20061=>"011111111",
  20062=>"111111000",
  20063=>"000000000",
  20064=>"101111100",
  20065=>"000000111",
  20066=>"111101101",
  20067=>"000000011",
  20068=>"000000000",
  20069=>"110000000",
  20070=>"000111111",
  20071=>"100000000",
  20072=>"000000000",
  20073=>"111111011",
  20074=>"000111011",
  20075=>"111111111",
  20076=>"000101111",
  20077=>"111111111",
  20078=>"000000101",
  20079=>"000000000",
  20080=>"111101100",
  20081=>"001101111",
  20082=>"111111111",
  20083=>"100110100",
  20084=>"000000000",
  20085=>"000010000",
  20086=>"111111111",
  20087=>"100110110",
  20088=>"001101111",
  20089=>"101101101",
  20090=>"111000000",
  20091=>"000000000",
  20092=>"111110000",
  20093=>"000100100",
  20094=>"111111010",
  20095=>"000111110",
  20096=>"000110110",
  20097=>"001001111",
  20098=>"000100100",
  20099=>"000000000",
  20100=>"000000000",
  20101=>"111101111",
  20102=>"111111111",
  20103=>"000110110",
  20104=>"111111000",
  20105=>"000100111",
  20106=>"111111111",
  20107=>"111111111",
  20108=>"001000100",
  20109=>"000000101",
  20110=>"111110111",
  20111=>"011111111",
  20112=>"001001111",
  20113=>"000000000",
  20114=>"111101001",
  20115=>"000000101",
  20116=>"111111000",
  20117=>"001000011",
  20118=>"000000111",
  20119=>"000000000",
  20120=>"010000101",
  20121=>"111111111",
  20122=>"000010111",
  20123=>"000000000",
  20124=>"000100000",
  20125=>"001000000",
  20126=>"101111111",
  20127=>"000000000",
  20128=>"111111111",
  20129=>"011111011",
  20130=>"000011111",
  20131=>"011111111",
  20132=>"011001000",
  20133=>"011011100",
  20134=>"111111111",
  20135=>"000001000",
  20136=>"000001111",
  20137=>"100000100",
  20138=>"111111111",
  20139=>"000000000",
  20140=>"000100000",
  20141=>"110111111",
  20142=>"000001111",
  20143=>"010110000",
  20144=>"000000000",
  20145=>"011011011",
  20146=>"110111000",
  20147=>"111111111",
  20148=>"111100000",
  20149=>"000111111",
  20150=>"000000000",
  20151=>"110111010",
  20152=>"000000011",
  20153=>"111111111",
  20154=>"111001000",
  20155=>"111100000",
  20156=>"000000000",
  20157=>"111001000",
  20158=>"111110111",
  20159=>"110000000",
  20160=>"100000111",
  20161=>"000000010",
  20162=>"111111100",
  20163=>"100000011",
  20164=>"000000110",
  20165=>"000000111",
  20166=>"000001111",
  20167=>"111110000",
  20168=>"111111111",
  20169=>"111111011",
  20170=>"111000001",
  20171=>"000111111",
  20172=>"000000010",
  20173=>"100000100",
  20174=>"110110001",
  20175=>"100111111",
  20176=>"000000111",
  20177=>"100100111",
  20178=>"111111100",
  20179=>"111111001",
  20180=>"001110010",
  20181=>"110110000",
  20182=>"000000000",
  20183=>"000000000",
  20184=>"111111000",
  20185=>"000000000",
  20186=>"111111111",
  20187=>"000000111",
  20188=>"000010111",
  20189=>"000001001",
  20190=>"000000000",
  20191=>"000000000",
  20192=>"000000000",
  20193=>"000110110",
  20194=>"000000000",
  20195=>"000000000",
  20196=>"111101000",
  20197=>"000000000",
  20198=>"111111111",
  20199=>"000000001",
  20200=>"000111111",
  20201=>"111111111",
  20202=>"111111111",
  20203=>"111100111",
  20204=>"000000001",
  20205=>"111111111",
  20206=>"111111111",
  20207=>"011011011",
  20208=>"001111000",
  20209=>"111011000",
  20210=>"111101101",
  20211=>"000000000",
  20212=>"111101111",
  20213=>"000000000",
  20214=>"000000000",
  20215=>"110111111",
  20216=>"111111111",
  20217=>"111110000",
  20218=>"000000000",
  20219=>"111111111",
  20220=>"111111100",
  20221=>"111000100",
  20222=>"011111111",
  20223=>"000000000",
  20224=>"000000001",
  20225=>"001001000",
  20226=>"000000000",
  20227=>"111111000",
  20228=>"001101111",
  20229=>"011011000",
  20230=>"111111111",
  20231=>"111110000",
  20232=>"000000000",
  20233=>"000000000",
  20234=>"000000000",
  20235=>"011011010",
  20236=>"110110110",
  20237=>"000001011",
  20238=>"000000000",
  20239=>"010111111",
  20240=>"111111111",
  20241=>"001000000",
  20242=>"000000000",
  20243=>"001001001",
  20244=>"111101111",
  20245=>"101000000",
  20246=>"000000000",
  20247=>"000000000",
  20248=>"111111111",
  20249=>"111111111",
  20250=>"111010000",
  20251=>"110110110",
  20252=>"010000000",
  20253=>"000000001",
  20254=>"000000000",
  20255=>"001111111",
  20256=>"100100011",
  20257=>"010111111",
  20258=>"111111111",
  20259=>"001100111",
  20260=>"001001100",
  20261=>"001000111",
  20262=>"000000001",
  20263=>"100001000",
  20264=>"001111010",
  20265=>"111000000",
  20266=>"000001111",
  20267=>"111101111",
  20268=>"000110110",
  20269=>"001000000",
  20270=>"111011010",
  20271=>"000000000",
  20272=>"111011000",
  20273=>"000101111",
  20274=>"010111111",
  20275=>"101101000",
  20276=>"000000000",
  20277=>"111111111",
  20278=>"111100100",
  20279=>"001000001",
  20280=>"100110100",
  20281=>"111100111",
  20282=>"111111010",
  20283=>"000000101",
  20284=>"000000111",
  20285=>"111111111",
  20286=>"111001000",
  20287=>"000000000",
  20288=>"111000010",
  20289=>"000000000",
  20290=>"000000000",
  20291=>"111111111",
  20292=>"001111111",
  20293=>"000000100",
  20294=>"000000000",
  20295=>"000000111",
  20296=>"000000000",
  20297=>"000001101",
  20298=>"001000000",
  20299=>"000000000",
  20300=>"001000000",
  20301=>"111111111",
  20302=>"111111111",
  20303=>"110100100",
  20304=>"111111100",
  20305=>"111111011",
  20306=>"000000000",
  20307=>"000000111",
  20308=>"111000001",
  20309=>"011001001",
  20310=>"000000000",
  20311=>"000000000",
  20312=>"100111111",
  20313=>"000000000",
  20314=>"000001111",
  20315=>"111111001",
  20316=>"111110111",
  20317=>"000000100",
  20318=>"111000000",
  20319=>"000110110",
  20320=>"000000111",
  20321=>"011000000",
  20322=>"000110110",
  20323=>"000000100",
  20324=>"111001000",
  20325=>"000111111",
  20326=>"000000000",
  20327=>"110110000",
  20328=>"001001001",
  20329=>"001111110",
  20330=>"001111111",
  20331=>"111110000",
  20332=>"110100000",
  20333=>"000010110",
  20334=>"001000000",
  20335=>"010111011",
  20336=>"000001011",
  20337=>"110010000",
  20338=>"111101000",
  20339=>"111111111",
  20340=>"110111110",
  20341=>"000000000",
  20342=>"000000000",
  20343=>"110000000",
  20344=>"111111000",
  20345=>"101000000",
  20346=>"000000000",
  20347=>"000000010",
  20348=>"111111111",
  20349=>"000000101",
  20350=>"011111111",
  20351=>"000111011",
  20352=>"011001011",
  20353=>"011011011",
  20354=>"100110111",
  20355=>"111111111",
  20356=>"000000001",
  20357=>"010000000",
  20358=>"001101111",
  20359=>"000000000",
  20360=>"000000000",
  20361=>"000000000",
  20362=>"111111000",
  20363=>"110000000",
  20364=>"001101111",
  20365=>"010001001",
  20366=>"010011011",
  20367=>"000000111",
  20368=>"000100100",
  20369=>"001001111",
  20370=>"000000000",
  20371=>"111100100",
  20372=>"101000111",
  20373=>"000110000",
  20374=>"111111000",
  20375=>"111111000",
  20376=>"000001111",
  20377=>"100111011",
  20378=>"000000000",
  20379=>"000001011",
  20380=>"000000000",
  20381=>"111111000",
  20382=>"011011111",
  20383=>"111110111",
  20384=>"110110000",
  20385=>"011000001",
  20386=>"111111111",
  20387=>"000000101",
  20388=>"000100101",
  20389=>"111110000",
  20390=>"001101111",
  20391=>"111111111",
  20392=>"000000000",
  20393=>"100100000",
  20394=>"111101111",
  20395=>"010110111",
  20396=>"111111111",
  20397=>"111111000",
  20398=>"001000001",
  20399=>"100100100",
  20400=>"000111111",
  20401=>"000000000",
  20402=>"111111111",
  20403=>"111111111",
  20404=>"011000111",
  20405=>"000111110",
  20406=>"000000111",
  20407=>"111111111",
  20408=>"111111000",
  20409=>"111000000",
  20410=>"000000000",
  20411=>"000000000",
  20412=>"100000011",
  20413=>"111110010",
  20414=>"000111111",
  20415=>"000000011",
  20416=>"111111111",
  20417=>"000000011",
  20418=>"111111011",
  20419=>"100000000",
  20420=>"000000101",
  20421=>"000111111",
  20422=>"110110111",
  20423=>"100001111",
  20424=>"001000000",
  20425=>"000000000",
  20426=>"101000010",
  20427=>"110110110",
  20428=>"111011111",
  20429=>"000000000",
  20430=>"001000100",
  20431=>"000111111",
  20432=>"101001011",
  20433=>"011000000",
  20434=>"001000000",
  20435=>"111000101",
  20436=>"000111111",
  20437=>"001000000",
  20438=>"111100111",
  20439=>"111111111",
  20440=>"001111111",
  20441=>"001011111",
  20442=>"000100001",
  20443=>"000000000",
  20444=>"111111111",
  20445=>"111111111",
  20446=>"000100111",
  20447=>"100111000",
  20448=>"110100111",
  20449=>"000000000",
  20450=>"000111001",
  20451=>"111011000",
  20452=>"111111111",
  20453=>"000000000",
  20454=>"111111111",
  20455=>"110110100",
  20456=>"000000000",
  20457=>"111110101",
  20458=>"000100100",
  20459=>"110110001",
  20460=>"111000101",
  20461=>"111111111",
  20462=>"111001111",
  20463=>"110111110",
  20464=>"010000000",
  20465=>"111110110",
  20466=>"000000101",
  20467=>"000000110",
  20468=>"111111111",
  20469=>"000010000",
  20470=>"111111111",
  20471=>"011001000",
  20472=>"011111000",
  20473=>"000000000",
  20474=>"011011011",
  20475=>"001000000",
  20476=>"100111000",
  20477=>"101100001",
  20478=>"111111111",
  20479=>"000110110",
  20480=>"111111110",
  20481=>"111111000",
  20482=>"000000001",
  20483=>"000000000",
  20484=>"111111011",
  20485=>"000000100",
  20486=>"000000000",
  20487=>"011010111",
  20488=>"111001111",
  20489=>"111111111",
  20490=>"111111111",
  20491=>"110111110",
  20492=>"000100010",
  20493=>"111111111",
  20494=>"000001001",
  20495=>"111111111",
  20496=>"111111111",
  20497=>"000001001",
  20498=>"000000011",
  20499=>"000111111",
  20500=>"111111111",
  20501=>"111111111",
  20502=>"110000000",
  20503=>"111100100",
  20504=>"110000000",
  20505=>"000010000",
  20506=>"000000000",
  20507=>"110110110",
  20508=>"111111111",
  20509=>"111111111",
  20510=>"011100100",
  20511=>"000010000",
  20512=>"001001000",
  20513=>"110010010",
  20514=>"100100000",
  20515=>"111110111",
  20516=>"111000001",
  20517=>"111111110",
  20518=>"000000011",
  20519=>"111001000",
  20520=>"111111111",
  20521=>"111111111",
  20522=>"111011011",
  20523=>"000000000",
  20524=>"111111111",
  20525=>"111101100",
  20526=>"000000000",
  20527=>"001100111",
  20528=>"001000000",
  20529=>"110111111",
  20530=>"111111110",
  20531=>"010111011",
  20532=>"100000000",
  20533=>"001001000",
  20534=>"000000000",
  20535=>"001101111",
  20536=>"111111111",
  20537=>"001000100",
  20538=>"000000000",
  20539=>"111111011",
  20540=>"111111111",
  20541=>"111111111",
  20542=>"000000011",
  20543=>"111111111",
  20544=>"111111000",
  20545=>"111111111",
  20546=>"101000000",
  20547=>"111111111",
  20548=>"000100000",
  20549=>"111111111",
  20550=>"111100000",
  20551=>"111011011",
  20552=>"000000000",
  20553=>"111111111",
  20554=>"111111111",
  20555=>"011001000",
  20556=>"000001011",
  20557=>"000011111",
  20558=>"111101000",
  20559=>"000000000",
  20560=>"111111111",
  20561=>"010010111",
  20562=>"000000000",
  20563=>"001000000",
  20564=>"111111111",
  20565=>"010000000",
  20566=>"111111001",
  20567=>"111111111",
  20568=>"111011001",
  20569=>"101000100",
  20570=>"000100110",
  20571=>"111011111",
  20572=>"111111111",
  20573=>"001100110",
  20574=>"011111111",
  20575=>"000111111",
  20576=>"100000000",
  20577=>"111111111",
  20578=>"111111111",
  20579=>"000000000",
  20580=>"111110110",
  20581=>"101001111",
  20582=>"111111111",
  20583=>"101000111",
  20584=>"111110110",
  20585=>"000000000",
  20586=>"111111111",
  20587=>"111111111",
  20588=>"000000111",
  20589=>"111111111",
  20590=>"111001111",
  20591=>"110110110",
  20592=>"111101001",
  20593=>"000000100",
  20594=>"100110111",
  20595=>"001111111",
  20596=>"000000000",
  20597=>"000111111",
  20598=>"111111111",
  20599=>"000000110",
  20600=>"001001001",
  20601=>"000010000",
  20602=>"000000000",
  20603=>"001101001",
  20604=>"000000000",
  20605=>"101101000",
  20606=>"000000000",
  20607=>"110010001",
  20608=>"111111111",
  20609=>"001000000",
  20610=>"101000110",
  20611=>"011001000",
  20612=>"001111111",
  20613=>"000000000",
  20614=>"010011111",
  20615=>"111111111",
  20616=>"110110010",
  20617=>"111111000",
  20618=>"111111001",
  20619=>"000000000",
  20620=>"110111111",
  20621=>"111111111",
  20622=>"000001111",
  20623=>"111101111",
  20624=>"001011111",
  20625=>"101111111",
  20626=>"111111111",
  20627=>"111111011",
  20628=>"111111111",
  20629=>"111101101",
  20630=>"111111000",
  20631=>"000000000",
  20632=>"110100101",
  20633=>"100000000",
  20634=>"111111111",
  20635=>"111111101",
  20636=>"100110110",
  20637=>"101000000",
  20638=>"111111111",
  20639=>"111100100",
  20640=>"111111111",
  20641=>"110110110",
  20642=>"000000000",
  20643=>"111111110",
  20644=>"000111111",
  20645=>"000000000",
  20646=>"111111111",
  20647=>"000000000",
  20648=>"111111111",
  20649=>"000000000",
  20650=>"000000000",
  20651=>"111111101",
  20652=>"111111110",
  20653=>"011011011",
  20654=>"111111000",
  20655=>"111011000",
  20656=>"010110110",
  20657=>"001000001",
  20658=>"000111101",
  20659=>"111111111",
  20660=>"000000000",
  20661=>"100100000",
  20662=>"111111111",
  20663=>"000000000",
  20664=>"111111111",
  20665=>"011010000",
  20666=>"001111100",
  20667=>"000000000",
  20668=>"111101000",
  20669=>"101110110",
  20670=>"110000000",
  20671=>"001001011",
  20672=>"000000000",
  20673=>"000000000",
  20674=>"111111111",
  20675=>"111111110",
  20676=>"100000000",
  20677=>"001011001",
  20678=>"001000111",
  20679=>"000001111",
  20680=>"111111111",
  20681=>"000000011",
  20682=>"001000001",
  20683=>"011111000",
  20684=>"000110110",
  20685=>"111111000",
  20686=>"111111111",
  20687=>"111111011",
  20688=>"000000100",
  20689=>"011111110",
  20690=>"000000000",
  20691=>"001000111",
  20692=>"111111111",
  20693=>"000000000",
  20694=>"111111111",
  20695=>"000111111",
  20696=>"000000000",
  20697=>"111011011",
  20698=>"111111111",
  20699=>"000000000",
  20700=>"111111111",
  20701=>"100110111",
  20702=>"111111111",
  20703=>"111111011",
  20704=>"111111111",
  20705=>"111111111",
  20706=>"001111111",
  20707=>"000000010",
  20708=>"000001000",
  20709=>"111111111",
  20710=>"000000000",
  20711=>"100111001",
  20712=>"111011000",
  20713=>"001001011",
  20714=>"111111111",
  20715=>"111101001",
  20716=>"000000000",
  20717=>"111111110",
  20718=>"111111111",
  20719=>"000000000",
  20720=>"000000000",
  20721=>"011010111",
  20722=>"000000010",
  20723=>"111111100",
  20724=>"001000000",
  20725=>"100111111",
  20726=>"111110100",
  20727=>"000000000",
  20728=>"111100100",
  20729=>"111111111",
  20730=>"100111101",
  20731=>"111111111",
  20732=>"111011111",
  20733=>"001001001",
  20734=>"111011011",
  20735=>"111111111",
  20736=>"000111000",
  20737=>"011010010",
  20738=>"001111011",
  20739=>"000000111",
  20740=>"111111110",
  20741=>"100000100",
  20742=>"000100000",
  20743=>"011001001",
  20744=>"000000111",
  20745=>"000000000",
  20746=>"110110100",
  20747=>"110000111",
  20748=>"110110110",
  20749=>"111111111",
  20750=>"000000010",
  20751=>"111111000",
  20752=>"100001001",
  20753=>"111111000",
  20754=>"101111111",
  20755=>"100110000",
  20756=>"000111111",
  20757=>"111111111",
  20758=>"001001000",
  20759=>"000000000",
  20760=>"000000100",
  20761=>"000000011",
  20762=>"000000000",
  20763=>"111111111",
  20764=>"001100000",
  20765=>"111010000",
  20766=>"111111111",
  20767=>"110111000",
  20768=>"000011011",
  20769=>"000000000",
  20770=>"000111111",
  20771=>"111111011",
  20772=>"001101111",
  20773=>"000001111",
  20774=>"000011001",
  20775=>"111111011",
  20776=>"111111111",
  20777=>"111111111",
  20778=>"111111111",
  20779=>"111111111",
  20780=>"101111111",
  20781=>"011011011",
  20782=>"011110111",
  20783=>"000000000",
  20784=>"001011011",
  20785=>"111101111",
  20786=>"000100000",
  20787=>"111101001",
  20788=>"111011000",
  20789=>"000000111",
  20790=>"100101101",
  20791=>"000000000",
  20792=>"111111110",
  20793=>"111000001",
  20794=>"001001011",
  20795=>"110010000",
  20796=>"000000000",
  20797=>"000000000",
  20798=>"000000010",
  20799=>"111111101",
  20800=>"111110000",
  20801=>"111000000",
  20802=>"111111110",
  20803=>"111000000",
  20804=>"000000000",
  20805=>"110010000",
  20806=>"000000000",
  20807=>"111111111",
  20808=>"111111111",
  20809=>"111111111",
  20810=>"111001011",
  20811=>"100100110",
  20812=>"000100100",
  20813=>"111111000",
  20814=>"100001111",
  20815=>"000000001",
  20816=>"000110000",
  20817=>"000000000",
  20818=>"111110100",
  20819=>"111111111",
  20820=>"010000000",
  20821=>"001011011",
  20822=>"000000011",
  20823=>"000000000",
  20824=>"111111111",
  20825=>"000111111",
  20826=>"111011000",
  20827=>"111111000",
  20828=>"111111111",
  20829=>"000000000",
  20830=>"111111111",
  20831=>"001001101",
  20832=>"110110111",
  20833=>"001111000",
  20834=>"101011011",
  20835=>"000000111",
  20836=>"111000100",
  20837=>"111111111",
  20838=>"111111111",
  20839=>"101001111",
  20840=>"010110111",
  20841=>"000000000",
  20842=>"100111000",
  20843=>"101011011",
  20844=>"011011011",
  20845=>"000000000",
  20846=>"000000000",
  20847=>"000000110",
  20848=>"000000000",
  20849=>"000000000",
  20850=>"111111110",
  20851=>"000000000",
  20852=>"000001000",
  20853=>"111110011",
  20854=>"110110000",
  20855=>"000000110",
  20856=>"111111111",
  20857=>"000000000",
  20858=>"110111111",
  20859=>"111111111",
  20860=>"000000000",
  20861=>"000001001",
  20862=>"111001000",
  20863=>"000000000",
  20864=>"111111100",
  20865=>"111101001",
  20866=>"111111111",
  20867=>"111111111",
  20868=>"000000000",
  20869=>"000100000",
  20870=>"111000000",
  20871=>"111111011",
  20872=>"111111111",
  20873=>"111111111",
  20874=>"000000000",
  20875=>"011000000",
  20876=>"111111111",
  20877=>"000011011",
  20878=>"111110000",
  20879=>"000111000",
  20880=>"111111111",
  20881=>"111110100",
  20882=>"001000000",
  20883=>"000000000",
  20884=>"000000000",
  20885=>"001000010",
  20886=>"100000000",
  20887=>"000000000",
  20888=>"001001000",
  20889=>"111111101",
  20890=>"000000001",
  20891=>"000001111",
  20892=>"000000000",
  20893=>"000000000",
  20894=>"001000000",
  20895=>"111111111",
  20896=>"111111111",
  20897=>"011001001",
  20898=>"110111111",
  20899=>"111111111",
  20900=>"000000001",
  20901=>"111111111",
  20902=>"111111111",
  20903=>"111001001",
  20904=>"111110110",
  20905=>"000011111",
  20906=>"000000000",
  20907=>"011111111",
  20908=>"111111111",
  20909=>"000001111",
  20910=>"001101100",
  20911=>"110111111",
  20912=>"100100000",
  20913=>"100100000",
  20914=>"000000000",
  20915=>"000000000",
  20916=>"111000000",
  20917=>"111110000",
  20918=>"111111000",
  20919=>"110100001",
  20920=>"111111110",
  20921=>"111111111",
  20922=>"000000000",
  20923=>"111110111",
  20924=>"001101000",
  20925=>"111101111",
  20926=>"111111000",
  20927=>"000000000",
  20928=>"000000000",
  20929=>"111111001",
  20930=>"111111110",
  20931=>"111011011",
  20932=>"110110110",
  20933=>"000000010",
  20934=>"000000000",
  20935=>"000001111",
  20936=>"010000000",
  20937=>"000000000",
  20938=>"011001000",
  20939=>"000000000",
  20940=>"111111000",
  20941=>"000011000",
  20942=>"111000100",
  20943=>"000110001",
  20944=>"010010000",
  20945=>"001001011",
  20946=>"111111111",
  20947=>"000000000",
  20948=>"111111111",
  20949=>"111111111",
  20950=>"000101111",
  20951=>"011011001",
  20952=>"000000000",
  20953=>"001001000",
  20954=>"111110100",
  20955=>"000011111",
  20956=>"111100111",
  20957=>"110000000",
  20958=>"101100100",
  20959=>"011111011",
  20960=>"000000000",
  20961=>"111111111",
  20962=>"000000000",
  20963=>"011111111",
  20964=>"000000000",
  20965=>"100000000",
  20966=>"010000000",
  20967=>"100100101",
  20968=>"111111000",
  20969=>"000000011",
  20970=>"000000000",
  20971=>"100010011",
  20972=>"000000000",
  20973=>"100100110",
  20974=>"001000000",
  20975=>"000000100",
  20976=>"000000000",
  20977=>"101111111",
  20978=>"100110111",
  20979=>"111111111",
  20980=>"100000000",
  20981=>"100100100",
  20982=>"111000011",
  20983=>"000011011",
  20984=>"000000000",
  20985=>"010110010",
  20986=>"100000001",
  20987=>"100111111",
  20988=>"011110111",
  20989=>"000101111",
  20990=>"000000000",
  20991=>"000000100",
  20992=>"000000000",
  20993=>"000000000",
  20994=>"110100000",
  20995=>"000111111",
  20996=>"010001000",
  20997=>"111001001",
  20998=>"000000000",
  20999=>"111111111",
  21000=>"000100000",
  21001=>"111111111",
  21002=>"001000000",
  21003=>"111111111",
  21004=>"000000000",
  21005=>"111111111",
  21006=>"111111100",
  21007=>"111111111",
  21008=>"111111111",
  21009=>"000011000",
  21010=>"010000000",
  21011=>"000100100",
  21012=>"101101000",
  21013=>"111110110",
  21014=>"000000010",
  21015=>"111111111",
  21016=>"111000000",
  21017=>"011000001",
  21018=>"111111111",
  21019=>"000100100",
  21020=>"111111111",
  21021=>"111111110",
  21022=>"110110010",
  21023=>"000000111",
  21024=>"001011111",
  21025=>"111011000",
  21026=>"111110111",
  21027=>"111111111",
  21028=>"111111100",
  21029=>"000000000",
  21030=>"100100101",
  21031=>"000000110",
  21032=>"111111111",
  21033=>"000110010",
  21034=>"111111111",
  21035=>"101000000",
  21036=>"111111111",
  21037=>"000100000",
  21038=>"000000110",
  21039=>"111111111",
  21040=>"000000000",
  21041=>"000000000",
  21042=>"110110110",
  21043=>"000000000",
  21044=>"000000000",
  21045=>"000000100",
  21046=>"111111111",
  21047=>"111111111",
  21048=>"000000100",
  21049=>"010110111",
  21050=>"010011000",
  21051=>"111111111",
  21052=>"000000100",
  21053=>"111111111",
  21054=>"000000100",
  21055=>"101001111",
  21056=>"111001000",
  21057=>"111111100",
  21058=>"110011010",
  21059=>"111111111",
  21060=>"110110110",
  21061=>"000000000",
  21062=>"000000001",
  21063=>"000000000",
  21064=>"100100111",
  21065=>"111111111",
  21066=>"000000000",
  21067=>"000000000",
  21068=>"011110000",
  21069=>"111111000",
  21070=>"111000001",
  21071=>"111111111",
  21072=>"100111001",
  21073=>"111011011",
  21074=>"111111010",
  21075=>"111111111",
  21076=>"011001000",
  21077=>"000100111",
  21078=>"000000000",
  21079=>"000000000",
  21080=>"000000100",
  21081=>"000000000",
  21082=>"000000000",
  21083=>"100100111",
  21084=>"111001000",
  21085=>"000010111",
  21086=>"111111101",
  21087=>"010110111",
  21088=>"111111111",
  21089=>"001000000",
  21090=>"000000000",
  21091=>"000000000",
  21092=>"110000000",
  21093=>"111111111",
  21094=>"111111111",
  21095=>"000000000",
  21096=>"000111111",
  21097=>"000111111",
  21098=>"000000000",
  21099=>"000000000",
  21100=>"000000110",
  21101=>"111110100",
  21102=>"100110110",
  21103=>"000000000",
  21104=>"111001100",
  21105=>"000111111",
  21106=>"001001111",
  21107=>"011011101",
  21108=>"111111111",
  21109=>"001000000",
  21110=>"000000000",
  21111=>"111111111",
  21112=>"000001001",
  21113=>"011011001",
  21114=>"110011011",
  21115=>"110111110",
  21116=>"110110110",
  21117=>"111111111",
  21118=>"000000000",
  21119=>"111001000",
  21120=>"111111111",
  21121=>"000000000",
  21122=>"111111000",
  21123=>"111111111",
  21124=>"000000001",
  21125=>"111100000",
  21126=>"110000000",
  21127=>"001001011",
  21128=>"000100100",
  21129=>"000000000",
  21130=>"111111111",
  21131=>"000000111",
  21132=>"111101101",
  21133=>"000000000",
  21134=>"000000000",
  21135=>"100000000",
  21136=>"000000000",
  21137=>"111111111",
  21138=>"111111111",
  21139=>"111111011",
  21140=>"001011111",
  21141=>"000000000",
  21142=>"000000000",
  21143=>"000000000",
  21144=>"111111111",
  21145=>"110101111",
  21146=>"010110111",
  21147=>"111111111",
  21148=>"111111111",
  21149=>"111000001",
  21150=>"111011000",
  21151=>"000000000",
  21152=>"000000000",
  21153=>"001000000",
  21154=>"011000110",
  21155=>"111111111",
  21156=>"000011001",
  21157=>"000000111",
  21158=>"111111111",
  21159=>"001001000",
  21160=>"111111111",
  21161=>"100100111",
  21162=>"111111111",
  21163=>"111111111",
  21164=>"000000000",
  21165=>"110110110",
  21166=>"000000100",
  21167=>"101000000",
  21168=>"000111111",
  21169=>"000000000",
  21170=>"001101000",
  21171=>"111111111",
  21172=>"111111111",
  21173=>"000000000",
  21174=>"000000000",
  21175=>"001001000",
  21176=>"000000000",
  21177=>"001111111",
  21178=>"000000000",
  21179=>"000000000",
  21180=>"010000110",
  21181=>"000000000",
  21182=>"100101101",
  21183=>"101111111",
  21184=>"100100110",
  21185=>"100000100",
  21186=>"000000001",
  21187=>"111111111",
  21188=>"111111111",
  21189=>"010000110",
  21190=>"000000000",
  21191=>"000000000",
  21192=>"000000000",
  21193=>"000000000",
  21194=>"111000000",
  21195=>"000000000",
  21196=>"111111100",
  21197=>"111111111",
  21198=>"000000000",
  21199=>"110000000",
  21200=>"000000000",
  21201=>"000000000",
  21202=>"111000000",
  21203=>"000000000",
  21204=>"111111111",
  21205=>"000001000",
  21206=>"011111111",
  21207=>"000000001",
  21208=>"101111111",
  21209=>"001100100",
  21210=>"000000101",
  21211=>"111111111",
  21212=>"000000100",
  21213=>"111111100",
  21214=>"001000001",
  21215=>"110111111",
  21216=>"111100110",
  21217=>"000010000",
  21218=>"111111000",
  21219=>"111111100",
  21220=>"111000000",
  21221=>"111110110",
  21222=>"111111111",
  21223=>"111111111",
  21224=>"111111000",
  21225=>"000000000",
  21226=>"011111111",
  21227=>"000000000",
  21228=>"000000000",
  21229=>"000010011",
  21230=>"011111111",
  21231=>"111000011",
  21232=>"111111111",
  21233=>"000111111",
  21234=>"000010000",
  21235=>"001000000",
  21236=>"111111111",
  21237=>"000110110",
  21238=>"100000110",
  21239=>"111111111",
  21240=>"111111111",
  21241=>"011011011",
  21242=>"000000000",
  21243=>"000000000",
  21244=>"000111111",
  21245=>"011011111",
  21246=>"000011011",
  21247=>"010110110",
  21248=>"110110110",
  21249=>"000000000",
  21250=>"000000000",
  21251=>"111111111",
  21252=>"000000111",
  21253=>"000000000",
  21254=>"111111111",
  21255=>"111111101",
  21256=>"001001100",
  21257=>"000000000",
  21258=>"001001011",
  21259=>"111111111",
  21260=>"111111011",
  21261=>"001011111",
  21262=>"000000000",
  21263=>"000000000",
  21264=>"110100000",
  21265=>"000000000",
  21266=>"000000000",
  21267=>"000000000",
  21268=>"111111111",
  21269=>"011000000",
  21270=>"100100000",
  21271=>"000000000",
  21272=>"111101001",
  21273=>"000000000",
  21274=>"000000000",
  21275=>"011000011",
  21276=>"111111111",
  21277=>"000000000",
  21278=>"000110111",
  21279=>"111001001",
  21280=>"100100111",
  21281=>"000100110",
  21282=>"111111111",
  21283=>"000000111",
  21284=>"100000000",
  21285=>"111111000",
  21286=>"111000000",
  21287=>"111111111",
  21288=>"000000000",
  21289=>"000000000",
  21290=>"010000010",
  21291=>"111111111",
  21292=>"011001000",
  21293=>"000010110",
  21294=>"111111111",
  21295=>"000000000",
  21296=>"111111110",
  21297=>"000000000",
  21298=>"110010001",
  21299=>"000000000",
  21300=>"000001001",
  21301=>"000000000",
  21302=>"111000001",
  21303=>"111111111",
  21304=>"000110000",
  21305=>"111101100",
  21306=>"000000000",
  21307=>"000000000",
  21308=>"000000000",
  21309=>"000000000",
  21310=>"000000000",
  21311=>"011011111",
  21312=>"000000000",
  21313=>"001100000",
  21314=>"111111111",
  21315=>"010000011",
  21316=>"011000111",
  21317=>"110011011",
  21318=>"011111111",
  21319=>"000000000",
  21320=>"000000011",
  21321=>"011011000",
  21322=>"000000000",
  21323=>"011001001",
  21324=>"110111111",
  21325=>"111111100",
  21326=>"111110111",
  21327=>"000000000",
  21328=>"010011010",
  21329=>"000000110",
  21330=>"000000000",
  21331=>"000001001",
  21332=>"100111111",
  21333=>"011000011",
  21334=>"000000000",
  21335=>"000000000",
  21336=>"000000011",
  21337=>"111111111",
  21338=>"111111111",
  21339=>"011000100",
  21340=>"111000000",
  21341=>"011001000",
  21342=>"111111111",
  21343=>"000000000",
  21344=>"111000001",
  21345=>"001011000",
  21346=>"011000000",
  21347=>"110000000",
  21348=>"000001000",
  21349=>"000000000",
  21350=>"000000000",
  21351=>"000000000",
  21352=>"100110100",
  21353=>"011011000",
  21354=>"000000000",
  21355=>"000000000",
  21356=>"110110111",
  21357=>"001011001",
  21358=>"111111000",
  21359=>"111000000",
  21360=>"000000000",
  21361=>"111111000",
  21362=>"111111111",
  21363=>"111111111",
  21364=>"111111111",
  21365=>"000000000",
  21366=>"100000000",
  21367=>"000000000",
  21368=>"000000000",
  21369=>"111111011",
  21370=>"000000001",
  21371=>"000000000",
  21372=>"111111111",
  21373=>"111100110",
  21374=>"000000000",
  21375=>"111111111",
  21376=>"001000000",
  21377=>"000000000",
  21378=>"000000000",
  21379=>"111111111",
  21380=>"111111111",
  21381=>"010011000",
  21382=>"111100000",
  21383=>"001011111",
  21384=>"000000000",
  21385=>"111111000",
  21386=>"001000010",
  21387=>"010010111",
  21388=>"110111111",
  21389=>"111111111",
  21390=>"000000110",
  21391=>"000000010",
  21392=>"000000000",
  21393=>"111100000",
  21394=>"011000111",
  21395=>"000000000",
  21396=>"111111111",
  21397=>"000000000",
  21398=>"000000010",
  21399=>"011011001",
  21400=>"000000000",
  21401=>"111111111",
  21402=>"111111111",
  21403=>"111111000",
  21404=>"000000000",
  21405=>"111111111",
  21406=>"111000000",
  21407=>"001111111",
  21408=>"000000000",
  21409=>"010000001",
  21410=>"000000100",
  21411=>"000101111",
  21412=>"111111111",
  21413=>"000000000",
  21414=>"111111111",
  21415=>"000000000",
  21416=>"111111100",
  21417=>"000000000",
  21418=>"111001101",
  21419=>"111001000",
  21420=>"000000000",
  21421=>"000000011",
  21422=>"110111111",
  21423=>"000000000",
  21424=>"111111011",
  21425=>"001000000",
  21426=>"111111111",
  21427=>"000001001",
  21428=>"111111111",
  21429=>"000000000",
  21430=>"111111111",
  21431=>"000011000",
  21432=>"000110111",
  21433=>"111111111",
  21434=>"111111111",
  21435=>"111011110",
  21436=>"011001001",
  21437=>"111110100",
  21438=>"001111111",
  21439=>"000010011",
  21440=>"111111101",
  21441=>"000000000",
  21442=>"111111111",
  21443=>"000000000",
  21444=>"111100100",
  21445=>"000010111",
  21446=>"000000000",
  21447=>"110110100",
  21448=>"000000000",
  21449=>"000000111",
  21450=>"111111111",
  21451=>"000000000",
  21452=>"000000000",
  21453=>"111001010",
  21454=>"111111111",
  21455=>"111111111",
  21456=>"111111111",
  21457=>"000000000",
  21458=>"101001001",
  21459=>"000000100",
  21460=>"111111111",
  21461=>"110110110",
  21462=>"000000000",
  21463=>"000000100",
  21464=>"000000000",
  21465=>"000111111",
  21466=>"000000000",
  21467=>"000000000",
  21468=>"101001111",
  21469=>"000001101",
  21470=>"000000000",
  21471=>"000000000",
  21472=>"000000111",
  21473=>"000000000",
  21474=>"111111111",
  21475=>"000000000",
  21476=>"000000000",
  21477=>"000000000",
  21478=>"000000000",
  21479=>"100011011",
  21480=>"110000000",
  21481=>"000000000",
  21482=>"000000001",
  21483=>"001000000",
  21484=>"111100000",
  21485=>"011001101",
  21486=>"000101111",
  21487=>"111111111",
  21488=>"000000000",
  21489=>"000000000",
  21490=>"111011111",
  21491=>"011110010",
  21492=>"000000000",
  21493=>"000000000",
  21494=>"111111111",
  21495=>"110000000",
  21496=>"011000000",
  21497=>"111001001",
  21498=>"000000000",
  21499=>"111001000",
  21500=>"000000000",
  21501=>"000000100",
  21502=>"111111111",
  21503=>"111111111",
  21504=>"000000111",
  21505=>"000000000",
  21506=>"000000111",
  21507=>"000111010",
  21508=>"000100110",
  21509=>"000000001",
  21510=>"100100000",
  21511=>"111100101",
  21512=>"000000000",
  21513=>"100111111",
  21514=>"001000000",
  21515=>"000000000",
  21516=>"000000000",
  21517=>"011000000",
  21518=>"000000000",
  21519=>"111111111",
  21520=>"000100100",
  21521=>"111100000",
  21522=>"111111111",
  21523=>"001000000",
  21524=>"001000000",
  21525=>"011011011",
  21526=>"000011000",
  21527=>"000000000",
  21528=>"111111110",
  21529=>"000000000",
  21530=>"111001111",
  21531=>"111111011",
  21532=>"000000000",
  21533=>"011111001",
  21534=>"110100000",
  21535=>"110000000",
  21536=>"000000000",
  21537=>"111111010",
  21538=>"000000000",
  21539=>"001000000",
  21540=>"000111110",
  21541=>"111111111",
  21542=>"001001001",
  21543=>"111101000",
  21544=>"011111001",
  21545=>"000000000",
  21546=>"000000000",
  21547=>"110000000",
  21548=>"001101000",
  21549=>"111111111",
  21550=>"100000000",
  21551=>"111111000",
  21552=>"000000010",
  21553=>"010000000",
  21554=>"111000000",
  21555=>"000000000",
  21556=>"000000010",
  21557=>"000110110",
  21558=>"000010111",
  21559=>"111000100",
  21560=>"111111000",
  21561=>"001111111",
  21562=>"000000000",
  21563=>"000000000",
  21564=>"101001101",
  21565=>"000000100",
  21566=>"111011111",
  21567=>"111000000",
  21568=>"111111001",
  21569=>"101001001",
  21570=>"000000000",
  21571=>"001000000",
  21572=>"000110110",
  21573=>"110110000",
  21574=>"111000000",
  21575=>"111111111",
  21576=>"111111000",
  21577=>"111000000",
  21578=>"101111111",
  21579=>"001000000",
  21580=>"100101000",
  21581=>"111111100",
  21582=>"000111111",
  21583=>"010000000",
  21584=>"000000101",
  21585=>"001011011",
  21586=>"000000000",
  21587=>"000000000",
  21588=>"101000000",
  21589=>"000110111",
  21590=>"000001111",
  21591=>"111111000",
  21592=>"000000000",
  21593=>"101000101",
  21594=>"111111001",
  21595=>"001000000",
  21596=>"000000000",
  21597=>"110000000",
  21598=>"000000101",
  21599=>"111111100",
  21600=>"000000000",
  21601=>"111111000",
  21602=>"000000000",
  21603=>"000000000",
  21604=>"000010010",
  21605=>"001001111",
  21606=>"111111111",
  21607=>"000011111",
  21608=>"100000000",
  21609=>"111111111",
  21610=>"000000000",
  21611=>"000011111",
  21612=>"001000000",
  21613=>"001001000",
  21614=>"100000011",
  21615=>"110111111",
  21616=>"111111111",
  21617=>"001000000",
  21618=>"111111110",
  21619=>"000000001",
  21620=>"000000000",
  21621=>"100110110",
  21622=>"000000000",
  21623=>"000110111",
  21624=>"000000000",
  21625=>"110111111",
  21626=>"111001000",
  21627=>"111000000",
  21628=>"110110110",
  21629=>"111111111",
  21630=>"011001000",
  21631=>"011000000",
  21632=>"000000111",
  21633=>"111111100",
  21634=>"111011000",
  21635=>"011011000",
  21636=>"000001111",
  21637=>"111000000",
  21638=>"000100100",
  21639=>"111111111",
  21640=>"111000000",
  21641=>"111111111",
  21642=>"000000000",
  21643=>"110101000",
  21644=>"000101111",
  21645=>"000100111",
  21646=>"001001111",
  21647=>"000001000",
  21648=>"111000000",
  21649=>"000000000",
  21650=>"001111111",
  21651=>"100000110",
  21652=>"011111001",
  21653=>"010000111",
  21654=>"011000000",
  21655=>"001000101",
  21656=>"111111111",
  21657=>"111111001",
  21658=>"011000000",
  21659=>"000000100",
  21660=>"011010010",
  21661=>"000000000",
  21662=>"000000000",
  21663=>"000111100",
  21664=>"111101100",
  21665=>"111111111",
  21666=>"101110010",
  21667=>"111111000",
  21668=>"001000000",
  21669=>"000010111",
  21670=>"111111100",
  21671=>"001111111",
  21672=>"111111111",
  21673=>"111111111",
  21674=>"111111111",
  21675=>"000001001",
  21676=>"101111001",
  21677=>"100100000",
  21678=>"000000000",
  21679=>"111101011",
  21680=>"111111110",
  21681=>"011001000",
  21682=>"110111110",
  21683=>"111101000",
  21684=>"000111111",
  21685=>"111001000",
  21686=>"000000100",
  21687=>"000001111",
  21688=>"000000001",
  21689=>"101111101",
  21690=>"111100000",
  21691=>"000000000",
  21692=>"111000111",
  21693=>"101000000",
  21694=>"111111111",
  21695=>"000111111",
  21696=>"000000000",
  21697=>"000000000",
  21698=>"000001000",
  21699=>"111111111",
  21700=>"100000111",
  21701=>"100000000",
  21702=>"011011000",
  21703=>"001000000",
  21704=>"110111111",
  21705=>"000001000",
  21706=>"110111110",
  21707=>"111000100",
  21708=>"101111111",
  21709=>"111111110",
  21710=>"000100110",
  21711=>"111111111",
  21712=>"000000000",
  21713=>"111111111",
  21714=>"111111011",
  21715=>"000001000",
  21716=>"000001011",
  21717=>"100000000",
  21718=>"000000001",
  21719=>"100110111",
  21720=>"000000111",
  21721=>"111100001",
  21722=>"000010111",
  21723=>"000000000",
  21724=>"100100100",
  21725=>"001001111",
  21726=>"000001111",
  21727=>"000001111",
  21728=>"111000000",
  21729=>"000111111",
  21730=>"000000111",
  21731=>"000000000",
  21732=>"111111111",
  21733=>"110000000",
  21734=>"110000111",
  21735=>"100000101",
  21736=>"000000000",
  21737=>"000000011",
  21738=>"111011001",
  21739=>"001000000",
  21740=>"110111111",
  21741=>"000000000",
  21742=>"000000000",
  21743=>"000111111",
  21744=>"001000101",
  21745=>"111111001",
  21746=>"111111011",
  21747=>"000000000",
  21748=>"010111111",
  21749=>"110111110",
  21750=>"100000111",
  21751=>"000111111",
  21752=>"110111111",
  21753=>"011000000",
  21754=>"000000100",
  21755=>"110111010",
  21756=>"110110110",
  21757=>"000000000",
  21758=>"000000101",
  21759=>"110100110",
  21760=>"000000101",
  21761=>"000000100",
  21762=>"111111001",
  21763=>"111111101",
  21764=>"111111111",
  21765=>"010111111",
  21766=>"000000101",
  21767=>"111111000",
  21768=>"000111010",
  21769=>"000000000",
  21770=>"001001101",
  21771=>"000000101",
  21772=>"111101111",
  21773=>"000011110",
  21774=>"000000000",
  21775=>"111111000",
  21776=>"011011111",
  21777=>"000111111",
  21778=>"011100111",
  21779=>"000000101",
  21780=>"111111111",
  21781=>"111111000",
  21782=>"111111100",
  21783=>"111000000",
  21784=>"110111111",
  21785=>"000110010",
  21786=>"111111111",
  21787=>"100000000",
  21788=>"100110000",
  21789=>"000111100",
  21790=>"000000111",
  21791=>"000000000",
  21792=>"000011001",
  21793=>"100000000",
  21794=>"011001000",
  21795=>"111111000",
  21796=>"011000000",
  21797=>"000110111",
  21798=>"111111110",
  21799=>"000000000",
  21800=>"111110000",
  21801=>"010111010",
  21802=>"000000000",
  21803=>"100000011",
  21804=>"110000000",
  21805=>"000011000",
  21806=>"111011111",
  21807=>"111101000",
  21808=>"111111111",
  21809=>"000000000",
  21810=>"110000000",
  21811=>"010011001",
  21812=>"111111111",
  21813=>"001010011",
  21814=>"001111111",
  21815=>"111000001",
  21816=>"001001000",
  21817=>"101100100",
  21818=>"000000000",
  21819=>"111111000",
  21820=>"000000000",
  21821=>"001111111",
  21822=>"000000100",
  21823=>"000000000",
  21824=>"100000111",
  21825=>"111111000",
  21826=>"111111000",
  21827=>"011000000",
  21828=>"000000000",
  21829=>"000000000",
  21830=>"000110111",
  21831=>"001111110",
  21832=>"000000010",
  21833=>"101000000",
  21834=>"000000000",
  21835=>"111000000",
  21836=>"111101111",
  21837=>"010111010",
  21838=>"000111011",
  21839=>"111111111",
  21840=>"000000000",
  21841=>"000100111",
  21842=>"111111111",
  21843=>"000000001",
  21844=>"011001000",
  21845=>"001011001",
  21846=>"111111000",
  21847=>"111111011",
  21848=>"111111111",
  21849=>"111000111",
  21850=>"100000000",
  21851=>"000000101",
  21852=>"000000000",
  21853=>"111000000",
  21854=>"001101110",
  21855=>"000000110",
  21856=>"000000001",
  21857=>"111111111",
  21858=>"001011011",
  21859=>"111000100",
  21860=>"000000000",
  21861=>"000111111",
  21862=>"111000000",
  21863=>"000101100",
  21864=>"100000000",
  21865=>"111111011",
  21866=>"101111010",
  21867=>"000000010",
  21868=>"000000000",
  21869=>"000000111",
  21870=>"000100111",
  21871=>"000000000",
  21872=>"000000000",
  21873=>"000000100",
  21874=>"111111000",
  21875=>"111111110",
  21876=>"110110000",
  21877=>"100000110",
  21878=>"100100111",
  21879=>"000000000",
  21880=>"111000000",
  21881=>"111000000",
  21882=>"000000000",
  21883=>"000011111",
  21884=>"111011000",
  21885=>"110111111",
  21886=>"111001000",
  21887=>"111000000",
  21888=>"100000100",
  21889=>"111110000",
  21890=>"111001000",
  21891=>"000000000",
  21892=>"111111111",
  21893=>"000101000",
  21894=>"000000000",
  21895=>"000000111",
  21896=>"010000110",
  21897=>"000000000",
  21898=>"000000000",
  21899=>"000100000",
  21900=>"111101111",
  21901=>"000110100",
  21902=>"000001011",
  21903=>"111111111",
  21904=>"011101100",
  21905=>"110111111",
  21906=>"111000000",
  21907=>"001000000",
  21908=>"111111111",
  21909=>"000010000",
  21910=>"000000111",
  21911=>"001001001",
  21912=>"000000101",
  21913=>"000000100",
  21914=>"111111100",
  21915=>"111000111",
  21916=>"000000000",
  21917=>"000000011",
  21918=>"001000000",
  21919=>"100111000",
  21920=>"000000000",
  21921=>"111111111",
  21922=>"100100000",
  21923=>"000111111",
  21924=>"100001001",
  21925=>"111101001",
  21926=>"111111111",
  21927=>"000111111",
  21928=>"011001000",
  21929=>"000001000",
  21930=>"111000000",
  21931=>"001001100",
  21932=>"000000000",
  21933=>"000110110",
  21934=>"000000111",
  21935=>"000000000",
  21936=>"111111111",
  21937=>"000001001",
  21938=>"111111111",
  21939=>"111111111",
  21940=>"111111111",
  21941=>"111000000",
  21942=>"001111111",
  21943=>"111001001",
  21944=>"000000111",
  21945=>"000000110",
  21946=>"111110000",
  21947=>"111000000",
  21948=>"111111111",
  21949=>"111100100",
  21950=>"001111111",
  21951=>"000000100",
  21952=>"000000011",
  21953=>"111111000",
  21954=>"111111111",
  21955=>"111111000",
  21956=>"000000001",
  21957=>"111001000",
  21958=>"000000001",
  21959=>"110111111",
  21960=>"000000000",
  21961=>"000000000",
  21962=>"111001000",
  21963=>"000111000",
  21964=>"001000000",
  21965=>"000000000",
  21966=>"101101000",
  21967=>"000111111",
  21968=>"111000000",
  21969=>"011111111",
  21970=>"000000100",
  21971=>"000000000",
  21972=>"000001001",
  21973=>"111111110",
  21974=>"000000000",
  21975=>"000000000",
  21976=>"000100100",
  21977=>"000000111",
  21978=>"000000000",
  21979=>"000000001",
  21980=>"111111001",
  21981=>"000100110",
  21982=>"011011011",
  21983=>"001011111",
  21984=>"000000000",
  21985=>"011000000",
  21986=>"000000000",
  21987=>"000101111",
  21988=>"111111111",
  21989=>"111111110",
  21990=>"111111111",
  21991=>"011011000",
  21992=>"000000001",
  21993=>"000100110",
  21994=>"000011111",
  21995=>"000000000",
  21996=>"001101001",
  21997=>"000000000",
  21998=>"000000000",
  21999=>"011011111",
  22000=>"111111100",
  22001=>"110111111",
  22002=>"011111111",
  22003=>"001000000",
  22004=>"010000000",
  22005=>"111000000",
  22006=>"000001111",
  22007=>"001100000",
  22008=>"001111111",
  22009=>"011001001",
  22010=>"111000000",
  22011=>"111111111",
  22012=>"011001011",
  22013=>"111110110",
  22014=>"000111110",
  22015=>"111111111",
  22016=>"111011000",
  22017=>"001000000",
  22018=>"000110111",
  22019=>"111110111",
  22020=>"111000000",
  22021=>"010000000",
  22022=>"000000000",
  22023=>"001000000",
  22024=>"000000000",
  22025=>"001000000",
  22026=>"111110000",
  22027=>"111110110",
  22028=>"111111111",
  22029=>"000000000",
  22030=>"000000000",
  22031=>"000000111",
  22032=>"100000100",
  22033=>"000011001",
  22034=>"000000000",
  22035=>"000000110",
  22036=>"101101101",
  22037=>"111111111",
  22038=>"111111111",
  22039=>"000000100",
  22040=>"000000111",
  22041=>"001000000",
  22042=>"000000000",
  22043=>"111100100",
  22044=>"111111000",
  22045=>"111011111",
  22046=>"000000001",
  22047=>"001001000",
  22048=>"000010000",
  22049=>"000000000",
  22050=>"000001000",
  22051=>"000000111",
  22052=>"111111111",
  22053=>"001000000",
  22054=>"010111111",
  22055=>"000000000",
  22056=>"111001110",
  22057=>"000000000",
  22058=>"111000000",
  22059=>"011011000",
  22060=>"000000000",
  22061=>"000000000",
  22062=>"010001011",
  22063=>"111111111",
  22064=>"011011000",
  22065=>"000000000",
  22066=>"111101000",
  22067=>"111111111",
  22068=>"000100101",
  22069=>"111011011",
  22070=>"111101100",
  22071=>"011000000",
  22072=>"111001000",
  22073=>"011001011",
  22074=>"000000000",
  22075=>"000110111",
  22076=>"111011111",
  22077=>"011111111",
  22078=>"011111111",
  22079=>"111111101",
  22080=>"011000000",
  22081=>"000000110",
  22082=>"111111111",
  22083=>"111110111",
  22084=>"111000000",
  22085=>"011111111",
  22086=>"111111111",
  22087=>"111111111",
  22088=>"111001000",
  22089=>"000010010",
  22090=>"111101101",
  22091=>"111000000",
  22092=>"110111111",
  22093=>"110000000",
  22094=>"000000000",
  22095=>"000111000",
  22096=>"111101100",
  22097=>"111111111",
  22098=>"111111000",
  22099=>"111111101",
  22100=>"111000000",
  22101=>"011000000",
  22102=>"111000001",
  22103=>"111100000",
  22104=>"011000000",
  22105=>"111111111",
  22106=>"100000000",
  22107=>"000100100",
  22108=>"000000000",
  22109=>"000000100",
  22110=>"000000000",
  22111=>"111111111",
  22112=>"010000000",
  22113=>"000000000",
  22114=>"111111111",
  22115=>"000111111",
  22116=>"111000111",
  22117=>"110100001",
  22118=>"111111111",
  22119=>"111111111",
  22120=>"111011000",
  22121=>"100001111",
  22122=>"100000000",
  22123=>"000000000",
  22124=>"001001000",
  22125=>"001001111",
  22126=>"011000001",
  22127=>"000000000",
  22128=>"000000000",
  22129=>"001000111",
  22130=>"001000000",
  22131=>"000000001",
  22132=>"111111111",
  22133=>"000100110",
  22134=>"100100000",
  22135=>"000000000",
  22136=>"000000001",
  22137=>"000000011",
  22138=>"000000000",
  22139=>"000000111",
  22140=>"111111001",
  22141=>"000100100",
  22142=>"000000000",
  22143=>"000000010",
  22144=>"000000000",
  22145=>"000000111",
  22146=>"000000000",
  22147=>"111100000",
  22148=>"111111100",
  22149=>"000000000",
  22150=>"111000110",
  22151=>"000000000",
  22152=>"111111111",
  22153=>"000000000",
  22154=>"000000000",
  22155=>"111111011",
  22156=>"111111111",
  22157=>"111111010",
  22158=>"111111111",
  22159=>"001111011",
  22160=>"110111111",
  22161=>"111111111",
  22162=>"000111111",
  22163=>"111011111",
  22164=>"011011010",
  22165=>"000000001",
  22166=>"001011011",
  22167=>"001000000",
  22168=>"100000001",
  22169=>"110000000",
  22170=>"000000000",
  22171=>"110110000",
  22172=>"001000000",
  22173=>"011001001",
  22174=>"000000111",
  22175=>"000000111",
  22176=>"000000111",
  22177=>"111000001",
  22178=>"111011000",
  22179=>"000000000",
  22180=>"000000000",
  22181=>"111111110",
  22182=>"111111111",
  22183=>"111111101",
  22184=>"101111000",
  22185=>"000001010",
  22186=>"111000000",
  22187=>"000011111",
  22188=>"000111110",
  22189=>"010000001",
  22190=>"001000000",
  22191=>"011111011",
  22192=>"111011111",
  22193=>"110010000",
  22194=>"110111000",
  22195=>"111111100",
  22196=>"111111111",
  22197=>"111111100",
  22198=>"000000000",
  22199=>"111010000",
  22200=>"111000000",
  22201=>"111111111",
  22202=>"000100000",
  22203=>"111111111",
  22204=>"100000111",
  22205=>"111110110",
  22206=>"000111111",
  22207=>"000000000",
  22208=>"001000000",
  22209=>"000000001",
  22210=>"001001000",
  22211=>"010000000",
  22212=>"000110010",
  22213=>"111111110",
  22214=>"011001101",
  22215=>"111011011",
  22216=>"111111010",
  22217=>"100111111",
  22218=>"001011011",
  22219=>"111111110",
  22220=>"111111000",
  22221=>"000000010",
  22222=>"111110000",
  22223=>"000000000",
  22224=>"010010001",
  22225=>"011000110",
  22226=>"111011011",
  22227=>"111111111",
  22228=>"111111000",
  22229=>"000001000",
  22230=>"111111110",
  22231=>"001011110",
  22232=>"011000011",
  22233=>"000000000",
  22234=>"000000000",
  22235=>"000000000",
  22236=>"111111010",
  22237=>"001000000",
  22238=>"011011111",
  22239=>"000000111",
  22240=>"111000000",
  22241=>"010010010",
  22242=>"111011011",
  22243=>"000000000",
  22244=>"010101011",
  22245=>"000100111",
  22246=>"000100110",
  22247=>"111111111",
  22248=>"111001111",
  22249=>"011001001",
  22250=>"111111101",
  22251=>"111000111",
  22252=>"000000000",
  22253=>"111111000",
  22254=>"111111111",
  22255=>"111111111",
  22256=>"001000100",
  22257=>"111111111",
  22258=>"101000000",
  22259=>"101000001",
  22260=>"111010000",
  22261=>"111110111",
  22262=>"001000000",
  22263=>"111111001",
  22264=>"000000110",
  22265=>"100000000",
  22266=>"111111011",
  22267=>"111111111",
  22268=>"000001011",
  22269=>"111111111",
  22270=>"010011000",
  22271=>"110000000",
  22272=>"000100111",
  22273=>"000000111",
  22274=>"111000111",
  22275=>"111111111",
  22276=>"111111111",
  22277=>"111001111",
  22278=>"111111111",
  22279=>"001001110",
  22280=>"000000000",
  22281=>"000000000",
  22282=>"001010000",
  22283=>"101000000",
  22284=>"001000000",
  22285=>"111101111",
  22286=>"110111111",
  22287=>"000111100",
  22288=>"111111000",
  22289=>"000000000",
  22290=>"000000001",
  22291=>"000000011",
  22292=>"011111111",
  22293=>"000000111",
  22294=>"000000001",
  22295=>"111110100",
  22296=>"000000000",
  22297=>"000000000",
  22298=>"111111111",
  22299=>"000000000",
  22300=>"111111110",
  22301=>"000000000",
  22302=>"000111111",
  22303=>"011010000",
  22304=>"001101001",
  22305=>"000000000",
  22306=>"111110111",
  22307=>"111111111",
  22308=>"111111110",
  22309=>"111001111",
  22310=>"000001001",
  22311=>"001011000",
  22312=>"011010011",
  22313=>"111111111",
  22314=>"111111111",
  22315=>"000001111",
  22316=>"111111110",
  22317=>"000000000",
  22318=>"111111000",
  22319=>"111111000",
  22320=>"001001101",
  22321=>"000100100",
  22322=>"000000000",
  22323=>"111111111",
  22324=>"000000000",
  22325=>"000000011",
  22326=>"001001000",
  22327=>"111111111",
  22328=>"011011111",
  22329=>"111000000",
  22330=>"000010010",
  22331=>"001001111",
  22332=>"011001001",
  22333=>"011000000",
  22334=>"000011011",
  22335=>"000000000",
  22336=>"111000000",
  22337=>"000000000",
  22338=>"011111010",
  22339=>"100000000",
  22340=>"000000000",
  22341=>"000000000",
  22342=>"000000000",
  22343=>"000000000",
  22344=>"111111111",
  22345=>"000111110",
  22346=>"011011101",
  22347=>"100111100",
  22348=>"010110111",
  22349=>"000000000",
  22350=>"111111111",
  22351=>"111111111",
  22352=>"000001000",
  22353=>"000000000",
  22354=>"000000000",
  22355=>"100111111",
  22356=>"000010110",
  22357=>"011011111",
  22358=>"011111111",
  22359=>"111101001",
  22360=>"000100111",
  22361=>"011000000",
  22362=>"000000111",
  22363=>"000000000",
  22364=>"000011010",
  22365=>"000000000",
  22366=>"001000000",
  22367=>"000000000",
  22368=>"111111111",
  22369=>"000000000",
  22370=>"011011011",
  22371=>"011111111",
  22372=>"000000000",
  22373=>"111111111",
  22374=>"111111111",
  22375=>"100110110",
  22376=>"001001001",
  22377=>"111100001",
  22378=>"111111110",
  22379=>"000000000",
  22380=>"011111111",
  22381=>"111000000",
  22382=>"000000000",
  22383=>"000011011",
  22384=>"011111111",
  22385=>"000001000",
  22386=>"111111111",
  22387=>"001000000",
  22388=>"111111000",
  22389=>"111111111",
  22390=>"111111100",
  22391=>"110111111",
  22392=>"000000000",
  22393=>"000000000",
  22394=>"111111111",
  22395=>"000000000",
  22396=>"111111111",
  22397=>"100000000",
  22398=>"000000000",
  22399=>"000000011",
  22400=>"110100111",
  22401=>"011011001",
  22402=>"110111001",
  22403=>"000000011",
  22404=>"111111111",
  22405=>"000100000",
  22406=>"000110100",
  22407=>"110011101",
  22408=>"000000100",
  22409=>"111111111",
  22410=>"111111111",
  22411=>"111111111",
  22412=>"000000001",
  22413=>"111111111",
  22414=>"111111111",
  22415=>"000000000",
  22416=>"111111111",
  22417=>"000000000",
  22418=>"111011011",
  22419=>"110110110",
  22420=>"000000000",
  22421=>"000000010",
  22422=>"111011000",
  22423=>"100000001",
  22424=>"011000000",
  22425=>"011111111",
  22426=>"000011111",
  22427=>"100000111",
  22428=>"000000000",
  22429=>"100000000",
  22430=>"111110000",
  22431=>"000000000",
  22432=>"000000000",
  22433=>"011011111",
  22434=>"111000000",
  22435=>"001011000",
  22436=>"111100100",
  22437=>"111111000",
  22438=>"111001000",
  22439=>"000000000",
  22440=>"110110110",
  22441=>"000000000",
  22442=>"000100000",
  22443=>"001000101",
  22444=>"000000000",
  22445=>"111011000",
  22446=>"110111011",
  22447=>"011011111",
  22448=>"111111110",
  22449=>"000000000",
  22450=>"111111111",
  22451=>"000100100",
  22452=>"111111111",
  22453=>"000000111",
  22454=>"111001001",
  22455=>"000000000",
  22456=>"111111111",
  22457=>"111010010",
  22458=>"000000000",
  22459=>"101101101",
  22460=>"111111000",
  22461=>"111001000",
  22462=>"011111110",
  22463=>"100000000",
  22464=>"111111111",
  22465=>"000000000",
  22466=>"000010000",
  22467=>"111111000",
  22468=>"000000000",
  22469=>"111011001",
  22470=>"001001000",
  22471=>"100111001",
  22472=>"000000000",
  22473=>"000000110",
  22474=>"011011011",
  22475=>"011011111",
  22476=>"111000000",
  22477=>"111111111",
  22478=>"000000000",
  22479=>"111111111",
  22480=>"000010111",
  22481=>"111111111",
  22482=>"101100110",
  22483=>"000111111",
  22484=>"011000001",
  22485=>"000000000",
  22486=>"100111111",
  22487=>"011011011",
  22488=>"111111111",
  22489=>"000000001",
  22490=>"110111111",
  22491=>"111111111",
  22492=>"001000000",
  22493=>"111011111",
  22494=>"000000000",
  22495=>"100100110",
  22496=>"000000110",
  22497=>"111111100",
  22498=>"100000000",
  22499=>"111011000",
  22500=>"111111101",
  22501=>"000000000",
  22502=>"111111000",
  22503=>"000001001",
  22504=>"011011000",
  22505=>"000011000",
  22506=>"110000111",
  22507=>"000000000",
  22508=>"000000000",
  22509=>"011100000",
  22510=>"101000000",
  22511=>"111111111",
  22512=>"000100000",
  22513=>"010011100",
  22514=>"000000000",
  22515=>"110111001",
  22516=>"011111111",
  22517=>"010000000",
  22518=>"000000000",
  22519=>"110111111",
  22520=>"000000000",
  22521=>"111100100",
  22522=>"000000000",
  22523=>"111111111",
  22524=>"111110011",
  22525=>"000000000",
  22526=>"111111111",
  22527=>"010100000",
  22528=>"000000110",
  22529=>"111111011",
  22530=>"000000111",
  22531=>"000000000",
  22532=>"111111000",
  22533=>"000001011",
  22534=>"000000001",
  22535=>"101111111",
  22536=>"000000000",
  22537=>"000000000",
  22538=>"000011000",
  22539=>"111111111",
  22540=>"100111011",
  22541=>"011000000",
  22542=>"000110100",
  22543=>"111001001",
  22544=>"000000000",
  22545=>"111010000",
  22546=>"000001111",
  22547=>"111111111",
  22548=>"100111111",
  22549=>"111111000",
  22550=>"101111111",
  22551=>"000111110",
  22552=>"111101111",
  22553=>"001011111",
  22554=>"100100100",
  22555=>"100000000",
  22556=>"001111111",
  22557=>"000111110",
  22558=>"001001001",
  22559=>"110100000",
  22560=>"111111001",
  22561=>"000000000",
  22562=>"111111010",
  22563=>"000000000",
  22564=>"111001000",
  22565=>"010000000",
  22566=>"000000101",
  22567=>"000011011",
  22568=>"000000000",
  22569=>"000000000",
  22570=>"001111111",
  22571=>"000001001",
  22572=>"000000001",
  22573=>"111111111",
  22574=>"000000000",
  22575=>"001101111",
  22576=>"111001000",
  22577=>"000000000",
  22578=>"000011111",
  22579=>"000000000",
  22580=>"111111111",
  22581=>"111111000",
  22582=>"111001000",
  22583=>"111000000",
  22584=>"001001000",
  22585=>"000000000",
  22586=>"000000111",
  22587=>"000110111",
  22588=>"000111111",
  22589=>"000000000",
  22590=>"010000000",
  22591=>"101000001",
  22592=>"011011000",
  22593=>"111000000",
  22594=>"000111111",
  22595=>"111111111",
  22596=>"000100010",
  22597=>"000000000",
  22598=>"111111000",
  22599=>"000111011",
  22600=>"111111111",
  22601=>"000000111",
  22602=>"111111001",
  22603=>"111111111",
  22604=>"001111111",
  22605=>"000111111",
  22606=>"110000001",
  22607=>"000000011",
  22608=>"111110000",
  22609=>"111111000",
  22610=>"111110000",
  22611=>"111110110",
  22612=>"000000000",
  22613=>"000000000",
  22614=>"000000000",
  22615=>"111111000",
  22616=>"011011111",
  22617=>"000000111",
  22618=>"000110111",
  22619=>"000000000",
  22620=>"010000000",
  22621=>"111111010",
  22622=>"000000101",
  22623=>"000000000",
  22624=>"000000001",
  22625=>"110111001",
  22626=>"000000100",
  22627=>"111111111",
  22628=>"111111000",
  22629=>"111000000",
  22630=>"000100100",
  22631=>"111000000",
  22632=>"000000110",
  22633=>"111111111",
  22634=>"000000000",
  22635=>"100111000",
  22636=>"000000000",
  22637=>"000100111",
  22638=>"000000000",
  22639=>"000000000",
  22640=>"000000001",
  22641=>"111001000",
  22642=>"111111000",
  22643=>"111111111",
  22644=>"000000111",
  22645=>"010110000",
  22646=>"000000111",
  22647=>"011000000",
  22648=>"000111011",
  22649=>"000000000",
  22650=>"000000000",
  22651=>"111111100",
  22652=>"111110000",
  22653=>"000000000",
  22654=>"111010000",
  22655=>"000000000",
  22656=>"111111000",
  22657=>"111101000",
  22658=>"001000100",
  22659=>"111111111",
  22660=>"111011010",
  22661=>"111111101",
  22662=>"101100000",
  22663=>"000000001",
  22664=>"100000000",
  22665=>"000011000",
  22666=>"000000000",
  22667=>"111000000",
  22668=>"000000000",
  22669=>"111111110",
  22670=>"111011111",
  22671=>"000110100",
  22672=>"000010000",
  22673=>"000000001",
  22674=>"000000000",
  22675=>"001011111",
  22676=>"100101100",
  22677=>"000000000",
  22678=>"111111001",
  22679=>"111111100",
  22680=>"001101101",
  22681=>"111111111",
  22682=>"111011000",
  22683=>"011000001",
  22684=>"111000000",
  22685=>"000011011",
  22686=>"111111001",
  22687=>"111111111",
  22688=>"000000110",
  22689=>"111110000",
  22690=>"000000111",
  22691=>"000000011",
  22692=>"000000001",
  22693=>"111000000",
  22694=>"110111000",
  22695=>"111111000",
  22696=>"000000100",
  22697=>"010111111",
  22698=>"000000111",
  22699=>"000000000",
  22700=>"111011000",
  22701=>"000100110",
  22702=>"111001001",
  22703=>"100111011",
  22704=>"011000001",
  22705=>"100000010",
  22706=>"110111010",
  22707=>"111111011",
  22708=>"000000000",
  22709=>"000000010",
  22710=>"000000000",
  22711=>"111111111",
  22712=>"000000011",
  22713=>"111111111",
  22714=>"000000100",
  22715=>"001000000",
  22716=>"000000000",
  22717=>"111010110",
  22718=>"111110111",
  22719=>"110110000",
  22720=>"111111110",
  22721=>"111101001",
  22722=>"111000000",
  22723=>"100111111",
  22724=>"000010111",
  22725=>"000111111",
  22726=>"111111000",
  22727=>"111111111",
  22728=>"010111111",
  22729=>"111111000",
  22730=>"111100000",
  22731=>"111000000",
  22732=>"100101111",
  22733=>"001111111",
  22734=>"000000111",
  22735=>"000000000",
  22736=>"000000000",
  22737=>"110111111",
  22738=>"000000000",
  22739=>"001001011",
  22740=>"100110000",
  22741=>"111001000",
  22742=>"000000000",
  22743=>"111001000",
  22744=>"111110101",
  22745=>"010110101",
  22746=>"000000000",
  22747=>"000010111",
  22748=>"111101111",
  22749=>"110110111",
  22750=>"111100000",
  22751=>"111111001",
  22752=>"000000000",
  22753=>"111110000",
  22754=>"110111111",
  22755=>"111111011",
  22756=>"011111001",
  22757=>"000000000",
  22758=>"000000000",
  22759=>"000000001",
  22760=>"000000000",
  22761=>"111111111",
  22762=>"011111111",
  22763=>"111111111",
  22764=>"010011111",
  22765=>"111111000",
  22766=>"111111111",
  22767=>"000111100",
  22768=>"000000101",
  22769=>"000000000",
  22770=>"100111111",
  22771=>"000110111",
  22772=>"000000000",
  22773=>"111000000",
  22774=>"001011111",
  22775=>"111111011",
  22776=>"000010011",
  22777=>"010000000",
  22778=>"110100111",
  22779=>"110111111",
  22780=>"111111111",
  22781=>"001001011",
  22782=>"111111111",
  22783=>"000000000",
  22784=>"000000000",
  22785=>"101111011",
  22786=>"001111111",
  22787=>"000001111",
  22788=>"111111110",
  22789=>"000000000",
  22790=>"111110101",
  22791=>"101000111",
  22792=>"000000000",
  22793=>"111111101",
  22794=>"111111111",
  22795=>"001001111",
  22796=>"000000111",
  22797=>"111111111",
  22798=>"111101000",
  22799=>"100110111",
  22800=>"011111111",
  22801=>"000000001",
  22802=>"000000000",
  22803=>"111111110",
  22804=>"000000000",
  22805=>"110111000",
  22806=>"001111011",
  22807=>"111000000",
  22808=>"000000000",
  22809=>"000111000",
  22810=>"001001000",
  22811=>"100000100",
  22812=>"101111111",
  22813=>"111000111",
  22814=>"000000000",
  22815=>"111111111",
  22816=>"001001000",
  22817=>"111111111",
  22818=>"100000000",
  22819=>"000000011",
  22820=>"111111011",
  22821=>"111111001",
  22822=>"100111111",
  22823=>"111111001",
  22824=>"110000000",
  22825=>"011101001",
  22826=>"110110011",
  22827=>"111111111",
  22828=>"000000000",
  22829=>"000000000",
  22830=>"110000111",
  22831=>"000000000",
  22832=>"111111110",
  22833=>"100000110",
  22834=>"100111101",
  22835=>"111111000",
  22836=>"000000000",
  22837=>"111000000",
  22838=>"111100111",
  22839=>"111111000",
  22840=>"101000000",
  22841=>"111000000",
  22842=>"111100100",
  22843=>"000000000",
  22844=>"110111111",
  22845=>"110111110",
  22846=>"111101000",
  22847=>"000110110",
  22848=>"000111111",
  22849=>"000100111",
  22850=>"111001011",
  22851=>"000110111",
  22852=>"000111001",
  22853=>"111111111",
  22854=>"001111111",
  22855=>"000000001",
  22856=>"000000000",
  22857=>"000111111",
  22858=>"100000111",
  22859=>"011111111",
  22860=>"000000111",
  22861=>"000000001",
  22862=>"000000000",
  22863=>"101111110",
  22864=>"001001000",
  22865=>"000000000",
  22866=>"111111000",
  22867=>"100111000",
  22868=>"111111111",
  22869=>"000001000",
  22870=>"000000000",
  22871=>"001101001",
  22872=>"111000111",
  22873=>"000000000",
  22874=>"111111001",
  22875=>"110101111",
  22876=>"000010010",
  22877=>"000001001",
  22878=>"000000000",
  22879=>"000000000",
  22880=>"000000000",
  22881=>"100111100",
  22882=>"000000000",
  22883=>"000111111",
  22884=>"110111110",
  22885=>"111111000",
  22886=>"111000000",
  22887=>"011000000",
  22888=>"100111111",
  22889=>"110111111",
  22890=>"011001000",
  22891=>"000000011",
  22892=>"010000000",
  22893=>"000111111",
  22894=>"111111111",
  22895=>"000000000",
  22896=>"111111001",
  22897=>"111010011",
  22898=>"100000000",
  22899=>"000000000",
  22900=>"100000000",
  22901=>"001001111",
  22902=>"010110111",
  22903=>"000111111",
  22904=>"000100111",
  22905=>"000000000",
  22906=>"111000001",
  22907=>"001001000",
  22908=>"000000111",
  22909=>"000100111",
  22910=>"000000000",
  22911=>"000000000",
  22912=>"000110111",
  22913=>"000000000",
  22914=>"000000000",
  22915=>"100000111",
  22916=>"111111111",
  22917=>"000000111",
  22918=>"000001001",
  22919=>"011111011",
  22920=>"000000000",
  22921=>"000000110",
  22922=>"000111111",
  22923=>"111110000",
  22924=>"000101111",
  22925=>"000000100",
  22926=>"111000000",
  22927=>"111111111",
  22928=>"001000000",
  22929=>"110000111",
  22930=>"111100000",
  22931=>"111111111",
  22932=>"000100000",
  22933=>"000000000",
  22934=>"111110111",
  22935=>"000000110",
  22936=>"000000000",
  22937=>"111111111",
  22938=>"000000001",
  22939=>"000000001",
  22940=>"000000001",
  22941=>"000000011",
  22942=>"000000000",
  22943=>"000000000",
  22944=>"111111000",
  22945=>"010000000",
  22946=>"111111111",
  22947=>"000000110",
  22948=>"001000110",
  22949=>"000100111",
  22950=>"000000000",
  22951=>"111111111",
  22952=>"000111111",
  22953=>"000000111",
  22954=>"111001011",
  22955=>"000000000",
  22956=>"000000000",
  22957=>"000000000",
  22958=>"111111110",
  22959=>"111111111",
  22960=>"111111000",
  22961=>"000000111",
  22962=>"011011111",
  22963=>"111111111",
  22964=>"000000000",
  22965=>"000001111",
  22966=>"010111111",
  22967=>"000000000",
  22968=>"110111111",
  22969=>"111111111",
  22970=>"111111000",
  22971=>"111111000",
  22972=>"000001011",
  22973=>"000111111",
  22974=>"111111111",
  22975=>"000000000",
  22976=>"000000000",
  22977=>"111111000",
  22978=>"111111111",
  22979=>"111000000",
  22980=>"111111111",
  22981=>"001001111",
  22982=>"100000110",
  22983=>"000010111",
  22984=>"000000000",
  22985=>"011000010",
  22986=>"001001011",
  22987=>"110111110",
  22988=>"100111000",
  22989=>"110111000",
  22990=>"001000000",
  22991=>"011001000",
  22992=>"010111111",
  22993=>"000111111",
  22994=>"111000000",
  22995=>"000010010",
  22996=>"111001001",
  22997=>"000000111",
  22998=>"001000001",
  22999=>"011000000",
  23000=>"000000111",
  23001=>"111111111",
  23002=>"000111111",
  23003=>"111001000",
  23004=>"111000111",
  23005=>"111110111",
  23006=>"111111000",
  23007=>"000110111",
  23008=>"000001010",
  23009=>"011110000",
  23010=>"000000000",
  23011=>"111000001",
  23012=>"111000000",
  23013=>"000110110",
  23014=>"000001100",
  23015=>"000000000",
  23016=>"000000000",
  23017=>"110111011",
  23018=>"111011000",
  23019=>"110111001",
  23020=>"111111111",
  23021=>"000000101",
  23022=>"111111111",
  23023=>"000101000",
  23024=>"000000000",
  23025=>"111010000",
  23026=>"100010010",
  23027=>"010111000",
  23028=>"111111111",
  23029=>"110111111",
  23030=>"111001111",
  23031=>"111000000",
  23032=>"000000100",
  23033=>"001000000",
  23034=>"100000100",
  23035=>"110000000",
  23036=>"111111101",
  23037=>"111111011",
  23038=>"110000000",
  23039=>"000000000",
  23040=>"111111111",
  23041=>"111101111",
  23042=>"000111111",
  23043=>"111000100",
  23044=>"111111111",
  23045=>"011010110",
  23046=>"111111001",
  23047=>"111111111",
  23048=>"111111111",
  23049=>"000000001",
  23050=>"111001000",
  23051=>"100111111",
  23052=>"000000000",
  23053=>"111111111",
  23054=>"000111111",
  23055=>"111111111",
  23056=>"000010010",
  23057=>"111111000",
  23058=>"100000000",
  23059=>"111110000",
  23060=>"111111111",
  23061=>"000110111",
  23062=>"111001000",
  23063=>"001000000",
  23064=>"111111111",
  23065=>"000010000",
  23066=>"000101000",
  23067=>"000100101",
  23068=>"111100000",
  23069=>"000100100",
  23070=>"010000011",
  23071=>"111000000",
  23072=>"111111111",
  23073=>"111111110",
  23074=>"000000000",
  23075=>"111111011",
  23076=>"011111111",
  23077=>"000000000",
  23078=>"111011011",
  23079=>"111001000",
  23080=>"111111111",
  23081=>"111111111",
  23082=>"111111111",
  23083=>"111010011",
  23084=>"101001000",
  23085=>"100110100",
  23086=>"000000001",
  23087=>"001001111",
  23088=>"011110111",
  23089=>"000000000",
  23090=>"000000000",
  23091=>"000000011",
  23092=>"100110000",
  23093=>"000000000",
  23094=>"000101111",
  23095=>"110101111",
  23096=>"111111111",
  23097=>"111111110",
  23098=>"101101111",
  23099=>"000000110",
  23100=>"001000000",
  23101=>"101101001",
  23102=>"110110110",
  23103=>"000000000",
  23104=>"100111110",
  23105=>"000000001",
  23106=>"000010000",
  23107=>"111111111",
  23108=>"110101111",
  23109=>"000000000",
  23110=>"111111111",
  23111=>"111001000",
  23112=>"111111110",
  23113=>"111001111",
  23114=>"011011000",
  23115=>"111111000",
  23116=>"111111111",
  23117=>"000110111",
  23118=>"000001000",
  23119=>"111111111",
  23120=>"000001001",
  23121=>"111111111",
  23122=>"111000111",
  23123=>"111111111",
  23124=>"000000000",
  23125=>"011000000",
  23126=>"111111111",
  23127=>"000000000",
  23128=>"000000000",
  23129=>"111101111",
  23130=>"000001111",
  23131=>"000010000",
  23132=>"111111111",
  23133=>"111111111",
  23134=>"000000000",
  23135=>"000000100",
  23136=>"000000000",
  23137=>"000000000",
  23138=>"110100100",
  23139=>"111111111",
  23140=>"111111111",
  23141=>"011000000",
  23142=>"000000000",
  23143=>"111111100",
  23144=>"000000000",
  23145=>"000000000",
  23146=>"111011011",
  23147=>"110111110",
  23148=>"111111010",
  23149=>"000000000",
  23150=>"000000000",
  23151=>"111111111",
  23152=>"001111111",
  23153=>"000000010",
  23154=>"111111011",
  23155=>"100101100",
  23156=>"101000000",
  23157=>"111111111",
  23158=>"100000000",
  23159=>"111111001",
  23160=>"111111111",
  23161=>"111000000",
  23162=>"100100101",
  23163=>"000000000",
  23164=>"010111110",
  23165=>"111110000",
  23166=>"001001011",
  23167=>"111111111",
  23168=>"011011111",
  23169=>"000100110",
  23170=>"000000100",
  23171=>"011110111",
  23172=>"000001000",
  23173=>"000000000",
  23174=>"111111111",
  23175=>"000000000",
  23176=>"111111010",
  23177=>"111110000",
  23178=>"000001001",
  23179=>"010000000",
  23180=>"111111111",
  23181=>"110111110",
  23182=>"000000000",
  23183=>"011011000",
  23184=>"111111000",
  23185=>"101101111",
  23186=>"000000111",
  23187=>"111100000",
  23188=>"111111111",
  23189=>"100110000",
  23190=>"111111111",
  23191=>"011011011",
  23192=>"000000000",
  23193=>"111001100",
  23194=>"001000110",
  23195=>"101101111",
  23196=>"111111111",
  23197=>"001000111",
  23198=>"000000000",
  23199=>"111111111",
  23200=>"000000110",
  23201=>"110100000",
  23202=>"000000000",
  23203=>"111111111",
  23204=>"001000000",
  23205=>"000000000",
  23206=>"010111000",
  23207=>"100000000",
  23208=>"111001011",
  23209=>"111111111",
  23210=>"111111111",
  23211=>"111111111",
  23212=>"111111100",
  23213=>"000011011",
  23214=>"001101001",
  23215=>"000000000",
  23216=>"111111111",
  23217=>"010010010",
  23218=>"111111111",
  23219=>"111111100",
  23220=>"000000000",
  23221=>"000000000",
  23222=>"000000000",
  23223=>"000000000",
  23224=>"111101110",
  23225=>"000000000",
  23226=>"101000000",
  23227=>"110000000",
  23228=>"000000010",
  23229=>"111111111",
  23230=>"000000000",
  23231=>"111011111",
  23232=>"111111111",
  23233=>"001001001",
  23234=>"000000100",
  23235=>"011011111",
  23236=>"111111111",
  23237=>"111011000",
  23238=>"111111100",
  23239=>"111111111",
  23240=>"000000000",
  23241=>"000110110",
  23242=>"101000000",
  23243=>"110110101",
  23244=>"000011111",
  23245=>"111111101",
  23246=>"110110000",
  23247=>"001000000",
  23248=>"000000100",
  23249=>"111111111",
  23250=>"111111011",
  23251=>"010011000",
  23252=>"100000000",
  23253=>"111111111",
  23254=>"000000000",
  23255=>"000000111",
  23256=>"000000000",
  23257=>"001000110",
  23258=>"111011010",
  23259=>"010111000",
  23260=>"100111111",
  23261=>"100000000",
  23262=>"000100000",
  23263=>"000000000",
  23264=>"000111111",
  23265=>"000001111",
  23266=>"111110000",
  23267=>"101101111",
  23268=>"001000000",
  23269=>"000010000",
  23270=>"111111111",
  23271=>"000000000",
  23272=>"000000000",
  23273=>"111111111",
  23274=>"011111111",
  23275=>"000000000",
  23276=>"110000000",
  23277=>"111111000",
  23278=>"000001000",
  23279=>"000000110",
  23280=>"000000000",
  23281=>"110111111",
  23282=>"111111111",
  23283=>"000000000",
  23284=>"001111111",
  23285=>"000000000",
  23286=>"101100101",
  23287=>"000000000",
  23288=>"111111111",
  23289=>"000000000",
  23290=>"000000000",
  23291=>"000111111",
  23292=>"000000000",
  23293=>"111111111",
  23294=>"011000000",
  23295=>"000000000",
  23296=>"000000000",
  23297=>"100000000",
  23298=>"111111111",
  23299=>"000100111",
  23300=>"001000000",
  23301=>"000000000",
  23302=>"111110110",
  23303=>"011111101",
  23304=>"001111111",
  23305=>"000000000",
  23306=>"000111111",
  23307=>"010111111",
  23308=>"101001000",
  23309=>"101000000",
  23310=>"000000000",
  23311=>"100000000",
  23312=>"000000000",
  23313=>"100101000",
  23314=>"111001000",
  23315=>"000000000",
  23316=>"000000000",
  23317=>"000010000",
  23318=>"001000000",
  23319=>"111111111",
  23320=>"010001000",
  23321=>"101101111",
  23322=>"000000001",
  23323=>"111111000",
  23324=>"111111001",
  23325=>"000000000",
  23326=>"011011111",
  23327=>"110100110",
  23328=>"111101001",
  23329=>"111101111",
  23330=>"000000000",
  23331=>"111111111",
  23332=>"001100000",
  23333=>"000000111",
  23334=>"000000000",
  23335=>"111001111",
  23336=>"100110110",
  23337=>"000000011",
  23338=>"000000000",
  23339=>"110100000",
  23340=>"000000110",
  23341=>"110110111",
  23342=>"111111111",
  23343=>"001001111",
  23344=>"011011011",
  23345=>"000000000",
  23346=>"111000001",
  23347=>"111111111",
  23348=>"111111111",
  23349=>"000000100",
  23350=>"000000000",
  23351=>"111000000",
  23352=>"000010010",
  23353=>"000000110",
  23354=>"001011010",
  23355=>"111111100",
  23356=>"111111111",
  23357=>"000000000",
  23358=>"101101101",
  23359=>"011011000",
  23360=>"100100100",
  23361=>"011000000",
  23362=>"100100100",
  23363=>"111111000",
  23364=>"110000001",
  23365=>"000001111",
  23366=>"100101100",
  23367=>"010111011",
  23368=>"000011000",
  23369=>"111111111",
  23370=>"000000100",
  23371=>"000000000",
  23372=>"111000000",
  23373=>"111111111",
  23374=>"000000000",
  23375=>"011011000",
  23376=>"000000000",
  23377=>"100000000",
  23378=>"000111111",
  23379=>"111111111",
  23380=>"110000000",
  23381=>"011011011",
  23382=>"001000000",
  23383=>"111101100",
  23384=>"111111111",
  23385=>"000000000",
  23386=>"100111110",
  23387=>"111111111",
  23388=>"000000000",
  23389=>"100000000",
  23390=>"000000000",
  23391=>"000010111",
  23392=>"111111111",
  23393=>"111111000",
  23394=>"001101111",
  23395=>"011111111",
  23396=>"001011011",
  23397=>"100000000",
  23398=>"001001011",
  23399=>"111111001",
  23400=>"000010000",
  23401=>"001111111",
  23402=>"000101100",
  23403=>"101111111",
  23404=>"000001001",
  23405=>"111111111",
  23406=>"111111000",
  23407=>"111111100",
  23408=>"110100000",
  23409=>"100000000",
  23410=>"111111111",
  23411=>"000000000",
  23412=>"111011110",
  23413=>"011010000",
  23414=>"100000101",
  23415=>"100111111",
  23416=>"000001011",
  23417=>"111111000",
  23418=>"111000000",
  23419=>"000111111",
  23420=>"000000000",
  23421=>"000000011",
  23422=>"101001101",
  23423=>"000000001",
  23424=>"110111111",
  23425=>"000001101",
  23426=>"000000000",
  23427=>"111111101",
  23428=>"111001000",
  23429=>"000000000",
  23430=>"000100000",
  23431=>"100000000",
  23432=>"000000000",
  23433=>"011111111",
  23434=>"111111010",
  23435=>"000000000",
  23436=>"101101111",
  23437=>"100100110",
  23438=>"000000100",
  23439=>"100100111",
  23440=>"000000000",
  23441=>"111100111",
  23442=>"001000000",
  23443=>"111111111",
  23444=>"001001000",
  23445=>"000000000",
  23446=>"000000000",
  23447=>"000010011",
  23448=>"101101111",
  23449=>"000100111",
  23450=>"000000000",
  23451=>"100111110",
  23452=>"111111111",
  23453=>"111111111",
  23454=>"000001000",
  23455=>"111111111",
  23456=>"011111111",
  23457=>"111111111",
  23458=>"001111001",
  23459=>"111000000",
  23460=>"111111111",
  23461=>"010000000",
  23462=>"111111111",
  23463=>"000111111",
  23464=>"000000110",
  23465=>"000000000",
  23466=>"000000101",
  23467=>"000000000",
  23468=>"000000000",
  23469=>"111111101",
  23470=>"011000000",
  23471=>"111111111",
  23472=>"011000010",
  23473=>"000000000",
  23474=>"000000000",
  23475=>"111000000",
  23476=>"101100001",
  23477=>"000000100",
  23478=>"001000000",
  23479=>"000000111",
  23480=>"000000111",
  23481=>"111110000",
  23482=>"000000000",
  23483=>"111100100",
  23484=>"000110111",
  23485=>"000000000",
  23486=>"000000000",
  23487=>"110010000",
  23488=>"110111111",
  23489=>"111111111",
  23490=>"111011001",
  23491=>"000000000",
  23492=>"000110111",
  23493=>"010000011",
  23494=>"111111111",
  23495=>"111100000",
  23496=>"000000000",
  23497=>"101101000",
  23498=>"000010011",
  23499=>"001001000",
  23500=>"000000000",
  23501=>"111111111",
  23502=>"000000000",
  23503=>"000110111",
  23504=>"111111001",
  23505=>"000000000",
  23506=>"111111111",
  23507=>"111111001",
  23508=>"111000111",
  23509=>"111000100",
  23510=>"001001010",
  23511=>"000000010",
  23512=>"000000000",
  23513=>"111110010",
  23514=>"000000000",
  23515=>"111111011",
  23516=>"111111111",
  23517=>"111111111",
  23518=>"111111111",
  23519=>"001000000",
  23520=>"000100000",
  23521=>"111111001",
  23522=>"111111001",
  23523=>"101101100",
  23524=>"000000000",
  23525=>"111111111",
  23526=>"111111000",
  23527=>"111111111",
  23528=>"111000000",
  23529=>"111000000",
  23530=>"000110000",
  23531=>"111111111",
  23532=>"111110100",
  23533=>"100100010",
  23534=>"000100111",
  23535=>"100110110",
  23536=>"001000000",
  23537=>"000000011",
  23538=>"000000000",
  23539=>"111111111",
  23540=>"000111111",
  23541=>"111111111",
  23542=>"011011001",
  23543=>"110011011",
  23544=>"000000010",
  23545=>"111111011",
  23546=>"000000110",
  23547=>"000000000",
  23548=>"111000111",
  23549=>"111111101",
  23550=>"111111000",
  23551=>"110110000",
  23552=>"000000001",
  23553=>"110000000",
  23554=>"111111111",
  23555=>"000000000",
  23556=>"111111000",
  23557=>"000000000",
  23558=>"100111111",
  23559=>"011111111",
  23560=>"111111111",
  23561=>"001001111",
  23562=>"001000111",
  23563=>"011111001",
  23564=>"111011000",
  23565=>"110000000",
  23566=>"110100100",
  23567=>"000001011",
  23568=>"110110110",
  23569=>"111111000",
  23570=>"101000001",
  23571=>"111011010",
  23572=>"000100111",
  23573=>"111111111",
  23574=>"000000000",
  23575=>"101000000",
  23576=>"000100110",
  23577=>"110110110",
  23578=>"111100000",
  23579=>"110000000",
  23580=>"111111111",
  23581=>"001001111",
  23582=>"000001000",
  23583=>"111110000",
  23584=>"111111001",
  23585=>"000001001",
  23586=>"011000000",
  23587=>"011111111",
  23588=>"000001000",
  23589=>"111111101",
  23590=>"000000011",
  23591=>"000000000",
  23592=>"000111111",
  23593=>"111111000",
  23594=>"000000010",
  23595=>"111011001",
  23596=>"000000000",
  23597=>"000000000",
  23598=>"110000000",
  23599=>"111111111",
  23600=>"111111000",
  23601=>"100110110",
  23602=>"000011001",
  23603=>"100100101",
  23604=>"000001001",
  23605=>"111000000",
  23606=>"001000000",
  23607=>"010111000",
  23608=>"111110000",
  23609=>"000110111",
  23610=>"111111111",
  23611=>"111001110",
  23612=>"111111111",
  23613=>"111011000",
  23614=>"111111101",
  23615=>"000000000",
  23616=>"000110110",
  23617=>"100001000",
  23618=>"111111000",
  23619=>"000000111",
  23620=>"111111000",
  23621=>"000000010",
  23622=>"111010000",
  23623=>"111111000",
  23624=>"110000000",
  23625=>"000101101",
  23626=>"000000000",
  23627=>"100111110",
  23628=>"001001001",
  23629=>"111111111",
  23630=>"110000000",
  23631=>"111111000",
  23632=>"111000000",
  23633=>"000000110",
  23634=>"000011010",
  23635=>"111111110",
  23636=>"000111000",
  23637=>"000001111",
  23638=>"000000100",
  23639=>"111011000",
  23640=>"111111111",
  23641=>"101101101",
  23642=>"011000111",
  23643=>"101101111",
  23644=>"000000001",
  23645=>"000000000",
  23646=>"000000000",
  23647=>"111110000",
  23648=>"111111111",
  23649=>"000000000",
  23650=>"000000000",
  23651=>"000000000",
  23652=>"000000111",
  23653=>"110110100",
  23654=>"111001111",
  23655=>"111111110",
  23656=>"000001100",
  23657=>"111111111",
  23658=>"100111111",
  23659=>"111111011",
  23660=>"100000000",
  23661=>"011110110",
  23662=>"001000000",
  23663=>"000001111",
  23664=>"000000000",
  23665=>"111100000",
  23666=>"000000001",
  23667=>"011000000",
  23668=>"000111101",
  23669=>"100111110",
  23670=>"111111111",
  23671=>"111111111",
  23672=>"000110111",
  23673=>"010001111",
  23674=>"111000000",
  23675=>"000000001",
  23676=>"110100100",
  23677=>"111111000",
  23678=>"110000000",
  23679=>"111110110",
  23680=>"111111111",
  23681=>"110111000",
  23682=>"000010010",
  23683=>"110110111",
  23684=>"111000000",
  23685=>"000000000",
  23686=>"000000000",
  23687=>"111100111",
  23688=>"111111111",
  23689=>"111001001",
  23690=>"111111111",
  23691=>"000111110",
  23692=>"000111111",
  23693=>"011011011",
  23694=>"100110111",
  23695=>"111111000",
  23696=>"000000000",
  23697=>"100000000",
  23698=>"111111111",
  23699=>"111111000",
  23700=>"100111100",
  23701=>"110110100",
  23702=>"111111001",
  23703=>"111011000",
  23704=>"001000111",
  23705=>"111000000",
  23706=>"111111111",
  23707=>"000111000",
  23708=>"000000000",
  23709=>"110110111",
  23710=>"011010111",
  23711=>"111111111",
  23712=>"111100100",
  23713=>"011011000",
  23714=>"000000111",
  23715=>"111110111",
  23716=>"111001011",
  23717=>"111110110",
  23718=>"011000000",
  23719=>"000000000",
  23720=>"001101111",
  23721=>"100111111",
  23722=>"000010000",
  23723=>"000001001",
  23724=>"000000000",
  23725=>"000111111",
  23726=>"111001101",
  23727=>"111000000",
  23728=>"000000010",
  23729=>"111111100",
  23730=>"000011010",
  23731=>"000001111",
  23732=>"111101101",
  23733=>"111111111",
  23734=>"111110000",
  23735=>"000101000",
  23736=>"001000001",
  23737=>"000001111",
  23738=>"101100000",
  23739=>"110110111",
  23740=>"101000000",
  23741=>"000111111",
  23742=>"100110101",
  23743=>"110111111",
  23744=>"000100111",
  23745=>"111001001",
  23746=>"110111111",
  23747=>"110000111",
  23748=>"000000111",
  23749=>"000000111",
  23750=>"001011011",
  23751=>"010000000",
  23752=>"000000011",
  23753=>"011000000",
  23754=>"000000110",
  23755=>"100111111",
  23756=>"000111111",
  23757=>"000111111",
  23758=>"110110111",
  23759=>"100110010",
  23760=>"111100100",
  23761=>"100100000",
  23762=>"111111001",
  23763=>"110000000",
  23764=>"000000000",
  23765=>"000000111",
  23766=>"111000000",
  23767=>"111111111",
  23768=>"111111000",
  23769=>"111000001",
  23770=>"000111111",
  23771=>"111100000",
  23772=>"111111011",
  23773=>"000100100",
  23774=>"000101111",
  23775=>"111000010",
  23776=>"000000111",
  23777=>"001001000",
  23778=>"111100000",
  23779=>"111000000",
  23780=>"000100000",
  23781=>"000010110",
  23782=>"111000000",
  23783=>"111111111",
  23784=>"011000000",
  23785=>"100000000",
  23786=>"111000000",
  23787=>"111101000",
  23788=>"010000000",
  23789=>"111000000",
  23790=>"001000011",
  23791=>"111111111",
  23792=>"011011111",
  23793=>"111110111",
  23794=>"000000000",
  23795=>"110001000",
  23796=>"000100110",
  23797=>"101000001",
  23798=>"000111001",
  23799=>"000000000",
  23800=>"000001000",
  23801=>"111000000",
  23802=>"111000000",
  23803=>"111000000",
  23804=>"011111111",
  23805=>"111110010",
  23806=>"111110000",
  23807=>"001011111",
  23808=>"111000000",
  23809=>"011000000",
  23810=>"000000000",
  23811=>"000100101",
  23812=>"000000000",
  23813=>"100101111",
  23814=>"000000100",
  23815=>"000000111",
  23816=>"111010000",
  23817=>"000000000",
  23818=>"000011111",
  23819=>"111000101",
  23820=>"111111001",
  23821=>"111101111",
  23822=>"111111111",
  23823=>"000001100",
  23824=>"111000110",
  23825=>"001000000",
  23826=>"000000111",
  23827=>"011111111",
  23828=>"000000111",
  23829=>"000000000",
  23830=>"111011000",
  23831=>"111111100",
  23832=>"000000100",
  23833=>"000000000",
  23834=>"111011011",
  23835=>"000000000",
  23836=>"000111011",
  23837=>"110111111",
  23838=>"111110000",
  23839=>"100000100",
  23840=>"111111000",
  23841=>"100000000",
  23842=>"000101000",
  23843=>"010000111",
  23844=>"000011000",
  23845=>"000111011",
  23846=>"111111001",
  23847=>"111111111",
  23848=>"000000000",
  23849=>"111000000",
  23850=>"011001000",
  23851=>"000000011",
  23852=>"110110111",
  23853=>"100000000",
  23854=>"111000011",
  23855=>"000000111",
  23856=>"000000001",
  23857=>"111011000",
  23858=>"100111001",
  23859=>"111110000",
  23860=>"111111100",
  23861=>"110000000",
  23862=>"111100110",
  23863=>"100111000",
  23864=>"000000000",
  23865=>"001000001",
  23866=>"101100000",
  23867=>"000111111",
  23868=>"001000000",
  23869=>"000001111",
  23870=>"001011111",
  23871=>"111011101",
  23872=>"000010100",
  23873=>"011001000",
  23874=>"001001000",
  23875=>"000000011",
  23876=>"000101111",
  23877=>"111111111",
  23878=>"111100100",
  23879=>"011000000",
  23880=>"000000011",
  23881=>"111100000",
  23882=>"111000000",
  23883=>"000001001",
  23884=>"110111111",
  23885=>"000100111",
  23886=>"111010000",
  23887=>"100100100",
  23888=>"111001000",
  23889=>"100100100",
  23890=>"000010000",
  23891=>"111111110",
  23892=>"111001000",
  23893=>"001011001",
  23894=>"100101000",
  23895=>"001001011",
  23896=>"011111111",
  23897=>"111110000",
  23898=>"110110110",
  23899=>"111000000",
  23900=>"000000111",
  23901=>"111111000",
  23902=>"110111110",
  23903=>"001111111",
  23904=>"100101111",
  23905=>"001001111",
  23906=>"000000000",
  23907=>"001111111",
  23908=>"000111110",
  23909=>"111111000",
  23910=>"111111001",
  23911=>"000111111",
  23912=>"000000000",
  23913=>"000000110",
  23914=>"111111000",
  23915=>"011111111",
  23916=>"011000100",
  23917=>"100111101",
  23918=>"000001111",
  23919=>"000000000",
  23920=>"111011000",
  23921=>"100111000",
  23922=>"111111000",
  23923=>"110111111",
  23924=>"111111111",
  23925=>"000111111",
  23926=>"100000000",
  23927=>"100000000",
  23928=>"111111111",
  23929=>"100000000",
  23930=>"110111110",
  23931=>"100000000",
  23932=>"111111100",
  23933=>"110000000",
  23934=>"110100000",
  23935=>"000111111",
  23936=>"000111111",
  23937=>"110110100",
  23938=>"000000000",
  23939=>"110100111",
  23940=>"111111110",
  23941=>"110100000",
  23942=>"000000000",
  23943=>"110000000",
  23944=>"000000000",
  23945=>"000000111",
  23946=>"000100110",
  23947=>"000111111",
  23948=>"001011111",
  23949=>"001000000",
  23950=>"001111111",
  23951=>"000111111",
  23952=>"110000000",
  23953=>"000000000",
  23954=>"000111111",
  23955=>"111001100",
  23956=>"101101101",
  23957=>"111000000",
  23958=>"000000111",
  23959=>"110000000",
  23960=>"111111000",
  23961=>"111110110",
  23962=>"111001111",
  23963=>"100100100",
  23964=>"011011000",
  23965=>"000000111",
  23966=>"000000011",
  23967=>"000111111",
  23968=>"111001111",
  23969=>"110110000",
  23970=>"001000100",
  23971=>"111000000",
  23972=>"001000101",
  23973=>"111111001",
  23974=>"111111111",
  23975=>"011111111",
  23976=>"101111111",
  23977=>"110111001",
  23978=>"110000100",
  23979=>"100100000",
  23980=>"111111000",
  23981=>"000000110",
  23982=>"000000111",
  23983=>"111111000",
  23984=>"001110100",
  23985=>"111101000",
  23986=>"001001000",
  23987=>"000100111",
  23988=>"110111111",
  23989=>"111111000",
  23990=>"000110101",
  23991=>"010110000",
  23992=>"000000111",
  23993=>"110111111",
  23994=>"000000000",
  23995=>"111111111",
  23996=>"000000011",
  23997=>"111111111",
  23998=>"111111111",
  23999=>"001001010",
  24000=>"001011100",
  24001=>"011101111",
  24002=>"000111000",
  24003=>"011111111",
  24004=>"010000111",
  24005=>"001111111",
  24006=>"000000000",
  24007=>"000001111",
  24008=>"111001000",
  24009=>"000110111",
  24010=>"111110000",
  24011=>"111111111",
  24012=>"111111000",
  24013=>"000001111",
  24014=>"101101111",
  24015=>"111100000",
  24016=>"000000100",
  24017=>"000000000",
  24018=>"100110000",
  24019=>"000000111",
  24020=>"101011011",
  24021=>"111111100",
  24022=>"110110000",
  24023=>"001011011",
  24024=>"110000000",
  24025=>"011010011",
  24026=>"111110010",
  24027=>"000000000",
  24028=>"000000000",
  24029=>"111111111",
  24030=>"011111000",
  24031=>"010000000",
  24032=>"000000000",
  24033=>"111100000",
  24034=>"110111111",
  24035=>"000000111",
  24036=>"111000000",
  24037=>"000000000",
  24038=>"110111001",
  24039=>"111100111",
  24040=>"011000000",
  24041=>"100111111",
  24042=>"100000000",
  24043=>"111111011",
  24044=>"000000000",
  24045=>"110010000",
  24046=>"000000000",
  24047=>"111111111",
  24048=>"100001010",
  24049=>"000000111",
  24050=>"111110000",
  24051=>"000011011",
  24052=>"110111111",
  24053=>"001111111",
  24054=>"100111111",
  24055=>"000000011",
  24056=>"111111000",
  24057=>"101100111",
  24058=>"111001000",
  24059=>"011011011",
  24060=>"011001101",
  24061=>"000000111",
  24062=>"110000000",
  24063=>"000010110",
  24064=>"101111001",
  24065=>"000000100",
  24066=>"000101101",
  24067=>"111111111",
  24068=>"000000001",
  24069=>"100110100",
  24070=>"111111101",
  24071=>"000000000",
  24072=>"000000111",
  24073=>"111101000",
  24074=>"000000000",
  24075=>"000110111",
  24076=>"000000000",
  24077=>"000000000",
  24078=>"000000111",
  24079=>"111111111",
  24080=>"110000000",
  24081=>"101001000",
  24082=>"000110110",
  24083=>"111100001",
  24084=>"111111111",
  24085=>"111111111",
  24086=>"000010010",
  24087=>"000000000",
  24088=>"011001001",
  24089=>"000000001",
  24090=>"000000101",
  24091=>"100101111",
  24092=>"111100000",
  24093=>"000011000",
  24094=>"001000000",
  24095=>"110110111",
  24096=>"001111111",
  24097=>"000000001",
  24098=>"000000001",
  24099=>"011000111",
  24100=>"001111111",
  24101=>"000000001",
  24102=>"110111111",
  24103=>"111111111",
  24104=>"000101011",
  24105=>"111111111",
  24106=>"111010110",
  24107=>"111111000",
  24108=>"000111111",
  24109=>"111000000",
  24110=>"111111111",
  24111=>"101101111",
  24112=>"111111111",
  24113=>"001001011",
  24114=>"100100100",
  24115=>"111111111",
  24116=>"000000000",
  24117=>"001001001",
  24118=>"111010000",
  24119=>"111101111",
  24120=>"101111100",
  24121=>"100111101",
  24122=>"111111111",
  24123=>"000000000",
  24124=>"000000111",
  24125=>"101011010",
  24126=>"011011011",
  24127=>"111111111",
  24128=>"000011000",
  24129=>"011011001",
  24130=>"000000000",
  24131=>"110111101",
  24132=>"000000000",
  24133=>"111111000",
  24134=>"110000100",
  24135=>"111111111",
  24136=>"000000000",
  24137=>"111001001",
  24138=>"100011111",
  24139=>"111111111",
  24140=>"010111111",
  24141=>"111001101",
  24142=>"000000100",
  24143=>"000000000",
  24144=>"111001111",
  24145=>"000000000",
  24146=>"000000000",
  24147=>"001010000",
  24148=>"000000000",
  24149=>"000000000",
  24150=>"000110110",
  24151=>"011111111",
  24152=>"111000000",
  24153=>"000000000",
  24154=>"000010111",
  24155=>"011111111",
  24156=>"111000000",
  24157=>"111111111",
  24158=>"111001111",
  24159=>"110110110",
  24160=>"000000101",
  24161=>"111110000",
  24162=>"000000000",
  24163=>"000000011",
  24164=>"100000011",
  24165=>"111111111",
  24166=>"110110010",
  24167=>"111111001",
  24168=>"000000000",
  24169=>"001111001",
  24170=>"111001111",
  24171=>"111111111",
  24172=>"110100000",
  24173=>"111111110",
  24174=>"110100000",
  24175=>"111001000",
  24176=>"111111011",
  24177=>"000000000",
  24178=>"111111100",
  24179=>"000110111",
  24180=>"110111111",
  24181=>"001001111",
  24182=>"000110000",
  24183=>"111111111",
  24184=>"000000000",
  24185=>"100000000",
  24186=>"111011001",
  24187=>"111111111",
  24188=>"110100000",
  24189=>"000000000",
  24190=>"000000000",
  24191=>"000111100",
  24192=>"111001001",
  24193=>"101111111",
  24194=>"000000000",
  24195=>"110110100",
  24196=>"110110111",
  24197=>"000000101",
  24198=>"001000000",
  24199=>"000000000",
  24200=>"111111101",
  24201=>"011000000",
  24202=>"000000000",
  24203=>"000000111",
  24204=>"000001001",
  24205=>"000010011",
  24206=>"000000000",
  24207=>"111111111",
  24208=>"111111111",
  24209=>"111111111",
  24210=>"101111011",
  24211=>"000000000",
  24212=>"111101100",
  24213=>"000000000",
  24214=>"111111110",
  24215=>"000000111",
  24216=>"111001000",
  24217=>"111111111",
  24218=>"000000000",
  24219=>"111111111",
  24220=>"111001001",
  24221=>"011010000",
  24222=>"000000000",
  24223=>"111111111",
  24224=>"111111111",
  24225=>"111000001",
  24226=>"111111111",
  24227=>"000000000",
  24228=>"000110100",
  24229=>"111111111",
  24230=>"111111111",
  24231=>"000000000",
  24232=>"111000000",
  24233=>"000001000",
  24234=>"001011011",
  24235=>"111101111",
  24236=>"100000000",
  24237=>"011011011",
  24238=>"000000000",
  24239=>"110110111",
  24240=>"111111100",
  24241=>"100100100",
  24242=>"111111111",
  24243=>"000000000",
  24244=>"111101000",
  24245=>"000010110",
  24246=>"111111111",
  24247=>"001000000",
  24248=>"110111111",
  24249=>"111100110",
  24250=>"001010001",
  24251=>"001011111",
  24252=>"111100110",
  24253=>"001001001",
  24254=>"111110111",
  24255=>"111111111",
  24256=>"111110110",
  24257=>"111001111",
  24258=>"011000000",
  24259=>"001000000",
  24260=>"111111111",
  24261=>"111111001",
  24262=>"111111111",
  24263=>"000100111",
  24264=>"010010111",
  24265=>"111111111",
  24266=>"111111111",
  24267=>"111111111",
  24268=>"111111111",
  24269=>"111111111",
  24270=>"000000111",
  24271=>"111011001",
  24272=>"111111100",
  24273=>"010111111",
  24274=>"010010000",
  24275=>"000001111",
  24276=>"100111111",
  24277=>"110110111",
  24278=>"000000000",
  24279=>"111110000",
  24280=>"100110000",
  24281=>"011001001",
  24282=>"000000000",
  24283=>"100000000",
  24284=>"000000000",
  24285=>"000000100",
  24286=>"110111111",
  24287=>"001111011",
  24288=>"000000000",
  24289=>"111101100",
  24290=>"000000000",
  24291=>"000000000",
  24292=>"111111011",
  24293=>"110100111",
  24294=>"111111100",
  24295=>"111111101",
  24296=>"111000000",
  24297=>"000000000",
  24298=>"000000000",
  24299=>"000011011",
  24300=>"111011111",
  24301=>"010111110",
  24302=>"000001001",
  24303=>"000100110",
  24304=>"111111111",
  24305=>"000100111",
  24306=>"000000110",
  24307=>"001001001",
  24308=>"111111111",
  24309=>"000000000",
  24310=>"100000000",
  24311=>"111111111",
  24312=>"111000000",
  24313=>"111111110",
  24314=>"111101001",
  24315=>"000000000",
  24316=>"100000000",
  24317=>"000000000",
  24318=>"000000000",
  24319=>"111110100",
  24320=>"000000000",
  24321=>"000000000",
  24322=>"000000111",
  24323=>"111001000",
  24324=>"100110110",
  24325=>"111111111",
  24326=>"000000000",
  24327=>"111111001",
  24328=>"100100000",
  24329=>"100110000",
  24330=>"010010000",
  24331=>"111111111",
  24332=>"000000110",
  24333=>"000000000",
  24334=>"111111111",
  24335=>"000100110",
  24336=>"000000100",
  24337=>"000111000",
  24338=>"111111111",
  24339=>"111111111",
  24340=>"011000011",
  24341=>"000000000",
  24342=>"000000000",
  24343=>"111111111",
  24344=>"111000001",
  24345=>"110100011",
  24346=>"100100000",
  24347=>"001111110",
  24348=>"001001001",
  24349=>"000000111",
  24350=>"111001001",
  24351=>"000000110",
  24352=>"110010000",
  24353=>"111100000",
  24354=>"110111111",
  24355=>"111011000",
  24356=>"001000000",
  24357=>"011111111",
  24358=>"000000000",
  24359=>"111111111",
  24360=>"110110111",
  24361=>"001111111",
  24362=>"111110000",
  24363=>"000010010",
  24364=>"000000000",
  24365=>"000000000",
  24366=>"000101000",
  24367=>"110100100",
  24368=>"000001001",
  24369=>"111111000",
  24370=>"000000000",
  24371=>"111111111",
  24372=>"000000000",
  24373=>"000000000",
  24374=>"110100111",
  24375=>"000010111",
  24376=>"111111000",
  24377=>"110000100",
  24378=>"000110111",
  24379=>"111111111",
  24380=>"111011011",
  24381=>"111110000",
  24382=>"111110011",
  24383=>"111001001",
  24384=>"000010000",
  24385=>"000000000",
  24386=>"000000000",
  24387=>"111111001",
  24388=>"000000001",
  24389=>"111111100",
  24390=>"111000000",
  24391=>"000000010",
  24392=>"110000000",
  24393=>"111111111",
  24394=>"011011000",
  24395=>"000100100",
  24396=>"011011011",
  24397=>"010011111",
  24398=>"100101101",
  24399=>"000000000",
  24400=>"111110110",
  24401=>"100100111",
  24402=>"110000100",
  24403=>"111111111",
  24404=>"001001000",
  24405=>"111111111",
  24406=>"000000000",
  24407=>"111111111",
  24408=>"101100000",
  24409=>"111111111",
  24410=>"111001000",
  24411=>"000111001",
  24412=>"111111111",
  24413=>"000000111",
  24414=>"111111101",
  24415=>"111111111",
  24416=>"100111111",
  24417=>"000000000",
  24418=>"000000000",
  24419=>"000000000",
  24420=>"000100100",
  24421=>"111111100",
  24422=>"111111111",
  24423=>"111111000",
  24424=>"000000000",
  24425=>"111110000",
  24426=>"000000000",
  24427=>"010111000",
  24428=>"011001101",
  24429=>"111101100",
  24430=>"111111101",
  24431=>"111111111",
  24432=>"000111111",
  24433=>"000000000",
  24434=>"000000000",
  24435=>"000000000",
  24436=>"011001101",
  24437=>"101001111",
  24438=>"111000100",
  24439=>"000000001",
  24440=>"111111111",
  24441=>"000000000",
  24442=>"000000000",
  24443=>"111011000",
  24444=>"000011001",
  24445=>"110000000",
  24446=>"100000000",
  24447=>"111000000",
  24448=>"000000111",
  24449=>"000111111",
  24450=>"111111010",
  24451=>"111111111",
  24452=>"000000000",
  24453=>"000001001",
  24454=>"111111001",
  24455=>"011000000",
  24456=>"111111111",
  24457=>"111000000",
  24458=>"000111111",
  24459=>"011000000",
  24460=>"111111111",
  24461=>"100000000",
  24462=>"111111111",
  24463=>"000000111",
  24464=>"000000000",
  24465=>"000111111",
  24466=>"100000000",
  24467=>"110111111",
  24468=>"000000000",
  24469=>"001111111",
  24470=>"110110000",
  24471=>"001000000",
  24472=>"001011000",
  24473=>"111111111",
  24474=>"100000001",
  24475=>"111001000",
  24476=>"100000000",
  24477=>"000000111",
  24478=>"000000011",
  24479=>"111111111",
  24480=>"001101111",
  24481=>"000100100",
  24482=>"000100111",
  24483=>"000000000",
  24484=>"111110111",
  24485=>"100000000",
  24486=>"111011111",
  24487=>"000000001",
  24488=>"011111111",
  24489=>"011011011",
  24490=>"111111111",
  24491=>"000111111",
  24492=>"000111111",
  24493=>"000001101",
  24494=>"011110111",
  24495=>"000110000",
  24496=>"010110000",
  24497=>"000000000",
  24498=>"000000110",
  24499=>"111100000",
  24500=>"000000000",
  24501=>"110100100",
  24502=>"001001111",
  24503=>"111111111",
  24504=>"100000010",
  24505=>"000000000",
  24506=>"100010111",
  24507=>"110010011",
  24508=>"111111010",
  24509=>"111100100",
  24510=>"111111111",
  24511=>"111001011",
  24512=>"000011011",
  24513=>"000000110",
  24514=>"000010000",
  24515=>"000011011",
  24516=>"111111111",
  24517=>"000000000",
  24518=>"000000000",
  24519=>"000000000",
  24520=>"000000000",
  24521=>"101001000",
  24522=>"111111000",
  24523=>"000110000",
  24524=>"111111001",
  24525=>"100101001",
  24526=>"000010111",
  24527=>"000111101",
  24528=>"000011001",
  24529=>"111110000",
  24530=>"111101101",
  24531=>"000000011",
  24532=>"011001011",
  24533=>"110111001",
  24534=>"100100100",
  24535=>"000100110",
  24536=>"111111101",
  24537=>"101111111",
  24538=>"000000000",
  24539=>"000000110",
  24540=>"001000000",
  24541=>"000000000",
  24542=>"110110110",
  24543=>"000001011",
  24544=>"000000000",
  24545=>"111111111",
  24546=>"100000000",
  24547=>"111001011",
  24548=>"101011011",
  24549=>"111111111",
  24550=>"000000000",
  24551=>"111110000",
  24552=>"000000000",
  24553=>"001000000",
  24554=>"000000000",
  24555=>"100100000",
  24556=>"000000000",
  24557=>"100110000",
  24558=>"000000000",
  24559=>"000000000",
  24560=>"000000001",
  24561=>"000000111",
  24562=>"111000000",
  24563=>"111111111",
  24564=>"000011001",
  24565=>"000101111",
  24566=>"111111011",
  24567=>"000001011",
  24568=>"000000111",
  24569=>"000000000",
  24570=>"111110000",
  24571=>"100110000",
  24572=>"000000100",
  24573=>"000000100",
  24574=>"001000000",
  24575=>"111110111",
  24576=>"110100000",
  24577=>"000000110",
  24578=>"111111111",
  24579=>"000000000",
  24580=>"000000000",
  24581=>"010000000",
  24582=>"101000000",
  24583=>"000000111",
  24584=>"000111111",
  24585=>"000000101",
  24586=>"000000000",
  24587=>"111011011",
  24588=>"100100000",
  24589=>"111111101",
  24590=>"111111111",
  24591=>"000100000",
  24592=>"111000001",
  24593=>"100111111",
  24594=>"111111111",
  24595=>"111111000",
  24596=>"000110110",
  24597=>"000000111",
  24598=>"000000000",
  24599=>"111100110",
  24600=>"111111001",
  24601=>"000001001",
  24602=>"000001011",
  24603=>"001001001",
  24604=>"000000111",
  24605=>"111001001",
  24606=>"000000011",
  24607=>"001000101",
  24608=>"111110000",
  24609=>"000000110",
  24610=>"100000100",
  24611=>"000000001",
  24612=>"111111011",
  24613=>"111111010",
  24614=>"111010000",
  24615=>"110111011",
  24616=>"111111111",
  24617=>"000000000",
  24618=>"011000001",
  24619=>"000001011",
  24620=>"101111111",
  24621=>"100000111",
  24622=>"110000001",
  24623=>"111111111",
  24624=>"000000000",
  24625=>"111111000",
  24626=>"000000000",
  24627=>"111111110",
  24628=>"110111100",
  24629=>"000100000",
  24630=>"000000000",
  24631=>"000000000",
  24632=>"000000000",
  24633=>"000000000",
  24634=>"000000000",
  24635=>"111111111",
  24636=>"111100110",
  24637=>"000110110",
  24638=>"000001011",
  24639=>"000100000",
  24640=>"000001001",
  24641=>"111111111",
  24642=>"000001000",
  24643=>"110110111",
  24644=>"100100000",
  24645=>"000011011",
  24646=>"111001111",
  24647=>"111111111",
  24648=>"001001000",
  24649=>"001000111",
  24650=>"111111111",
  24651=>"111111111",
  24652=>"110110110",
  24653=>"000000110",
  24654=>"111101100",
  24655=>"111111111",
  24656=>"000010111",
  24657=>"000000000",
  24658=>"111111101",
  24659=>"111001001",
  24660=>"110111111",
  24661=>"111111111",
  24662=>"000000000",
  24663=>"111101101",
  24664=>"000000000",
  24665=>"111101111",
  24666=>"000000000",
  24667=>"001000000",
  24668=>"000000000",
  24669=>"111011010",
  24670=>"111111111",
  24671=>"000000000",
  24672=>"110100111",
  24673=>"111111111",
  24674=>"111111111",
  24675=>"111111101",
  24676=>"101111000",
  24677=>"000000000",
  24678=>"111111111",
  24679=>"111111111",
  24680=>"000000000",
  24681=>"000100110",
  24682=>"000000001",
  24683=>"000000010",
  24684=>"000000000",
  24685=>"111111111",
  24686=>"111111000",
  24687=>"000110110",
  24688=>"111111111",
  24689=>"110111111",
  24690=>"000000000",
  24691=>"111000000",
  24692=>"111111111",
  24693=>"111111000",
  24694=>"111111111",
  24695=>"111111000",
  24696=>"011011011",
  24697=>"000000011",
  24698=>"111111111",
  24699=>"111000000",
  24700=>"101101100",
  24701=>"010010011",
  24702=>"111000000",
  24703=>"000000000",
  24704=>"111001111",
  24705=>"111111111",
  24706=>"000000000",
  24707=>"100100000",
  24708=>"100000001",
  24709=>"111111111",
  24710=>"000100000",
  24711=>"000000000",
  24712=>"111111111",
  24713=>"000000100",
  24714=>"110000000",
  24715=>"000111111",
  24716=>"110111111",
  24717=>"100111111",
  24718=>"000010110",
  24719=>"000000000",
  24720=>"111111111",
  24721=>"101001000",
  24722=>"000000000",
  24723=>"111111011",
  24724=>"111111000",
  24725=>"111001001",
  24726=>"000010111",
  24727=>"111111111",
  24728=>"000000000",
  24729=>"000000100",
  24730=>"000000000",
  24731=>"111111101",
  24732=>"111111011",
  24733=>"000000000",
  24734=>"000000000",
  24735=>"111111111",
  24736=>"000000000",
  24737=>"110011000",
  24738=>"000001111",
  24739=>"011011110",
  24740=>"000000000",
  24741=>"000000000",
  24742=>"010111111",
  24743=>"010010000",
  24744=>"000100000",
  24745=>"111111101",
  24746=>"111111111",
  24747=>"111000100",
  24748=>"000000000",
  24749=>"111111100",
  24750=>"101101111",
  24751=>"111111010",
  24752=>"111111100",
  24753=>"000100100",
  24754=>"110111010",
  24755=>"000000000",
  24756=>"000000100",
  24757=>"111111111",
  24758=>"000000000",
  24759=>"000111111",
  24760=>"011111111",
  24761=>"000001111",
  24762=>"000100111",
  24763=>"000100110",
  24764=>"111111001",
  24765=>"000111111",
  24766=>"000000000",
  24767=>"111111111",
  24768=>"000011111",
  24769=>"000000110",
  24770=>"000000000",
  24771=>"000000000",
  24772=>"000010011",
  24773=>"111111111",
  24774=>"111111111",
  24775=>"011111111",
  24776=>"000010111",
  24777=>"000000000",
  24778=>"111100100",
  24779=>"111111111",
  24780=>"110111101",
  24781=>"000000000",
  24782=>"000000000",
  24783=>"000001001",
  24784=>"111001000",
  24785=>"111110010",
  24786=>"001000000",
  24787=>"000000000",
  24788=>"000000000",
  24789=>"000000000",
  24790=>"111111111",
  24791=>"000001000",
  24792=>"000010111",
  24793=>"111001111",
  24794=>"000000110",
  24795=>"000000000",
  24796=>"000000110",
  24797=>"000000111",
  24798=>"000000000",
  24799=>"111110110",
  24800=>"000100110",
  24801=>"000000000",
  24802=>"000000000",
  24803=>"111111111",
  24804=>"111000111",
  24805=>"100000000",
  24806=>"110110111",
  24807=>"111111111",
  24808=>"000100000",
  24809=>"000000000",
  24810=>"100000100",
  24811=>"000000111",
  24812=>"000000000",
  24813=>"001011011",
  24814=>"100110111",
  24815=>"111111111",
  24816=>"000000000",
  24817=>"111011000",
  24818=>"111111111",
  24819=>"110101111",
  24820=>"000010111",
  24821=>"110100000",
  24822=>"000001001",
  24823=>"000111111",
  24824=>"111111111",
  24825=>"000000000",
  24826=>"000000000",
  24827=>"000001001",
  24828=>"001011000",
  24829=>"111111111",
  24830=>"100110110",
  24831=>"111111101",
  24832=>"001111110",
  24833=>"010010000",
  24834=>"111011011",
  24835=>"000000000",
  24836=>"111111111",
  24837=>"011011000",
  24838=>"000000000",
  24839=>"000000000",
  24840=>"100100100",
  24841=>"000000111",
  24842=>"111111111",
  24843=>"000000000",
  24844=>"111111110",
  24845=>"010000000",
  24846=>"000110111",
  24847=>"110111010",
  24848=>"111111101",
  24849=>"100000111",
  24850=>"111111111",
  24851=>"111110111",
  24852=>"011100111",
  24853=>"000000000",
  24854=>"011001101",
  24855=>"111111111",
  24856=>"000000101",
  24857=>"110111111",
  24858=>"110111111",
  24859=>"000111000",
  24860=>"000000000",
  24861=>"010111011",
  24862=>"111111100",
  24863=>"011000100",
  24864=>"110011011",
  24865=>"000000000",
  24866=>"111111100",
  24867=>"111111111",
  24868=>"000000100",
  24869=>"111111111",
  24870=>"011111111",
  24871=>"111111111",
  24872=>"110111111",
  24873=>"001000000",
  24874=>"111000000",
  24875=>"000000000",
  24876=>"111111000",
  24877=>"111111001",
  24878=>"111101101",
  24879=>"111011011",
  24880=>"001001101",
  24881=>"000000000",
  24882=>"000000000",
  24883=>"111111010",
  24884=>"000000000",
  24885=>"000010000",
  24886=>"111111000",
  24887=>"110111111",
  24888=>"000000000",
  24889=>"111111111",
  24890=>"010000000",
  24891=>"111111111",
  24892=>"000001111",
  24893=>"111111111",
  24894=>"010111111",
  24895=>"111111111",
  24896=>"110100110",
  24897=>"000000000",
  24898=>"000001001",
  24899=>"011000000",
  24900=>"111111111",
  24901=>"000111111",
  24902=>"010000000",
  24903=>"111111110",
  24904=>"000000000",
  24905=>"000000000",
  24906=>"011000000",
  24907=>"000000000",
  24908=>"000000010",
  24909=>"111000000",
  24910=>"111111111",
  24911=>"111011001",
  24912=>"101001000",
  24913=>"111111111",
  24914=>"000000110",
  24915=>"000000000",
  24916=>"111111110",
  24917=>"111111011",
  24918=>"000000000",
  24919=>"111111111",
  24920=>"111111111",
  24921=>"111001000",
  24922=>"100000100",
  24923=>"001100100",
  24924=>"011011111",
  24925=>"111111111",
  24926=>"111111101",
  24927=>"110111110",
  24928=>"000000000",
  24929=>"111000100",
  24930=>"100111111",
  24931=>"111111011",
  24932=>"101000000",
  24933=>"000000000",
  24934=>"000111111",
  24935=>"101000000",
  24936=>"000000000",
  24937=>"000010110",
  24938=>"111111110",
  24939=>"000000011",
  24940=>"111110110",
  24941=>"111111111",
  24942=>"111111111",
  24943=>"000000000",
  24944=>"110000000",
  24945=>"111011000",
  24946=>"010011100",
  24947=>"000000000",
  24948=>"000001001",
  24949=>"111011001",
  24950=>"000000111",
  24951=>"110110111",
  24952=>"111101111",
  24953=>"001000000",
  24954=>"111111111",
  24955=>"011111111",
  24956=>"010000000",
  24957=>"111111111",
  24958=>"111111111",
  24959=>"111111111",
  24960=>"010011011",
  24961=>"000000000",
  24962=>"111010000",
  24963=>"111111111",
  24964=>"000000000",
  24965=>"111111111",
  24966=>"001000000",
  24967=>"000010110",
  24968=>"111111111",
  24969=>"111111111",
  24970=>"111000000",
  24971=>"111111111",
  24972=>"111101111",
  24973=>"011011010",
  24974=>"000001001",
  24975=>"111111111",
  24976=>"111111111",
  24977=>"000000100",
  24978=>"110111101",
  24979=>"000110110",
  24980=>"000000000",
  24981=>"010010010",
  24982=>"000000101",
  24983=>"111111100",
  24984=>"110111111",
  24985=>"000000100",
  24986=>"111111111",
  24987=>"001001000",
  24988=>"000110111",
  24989=>"011000000",
  24990=>"111111110",
  24991=>"011000000",
  24992=>"000111111",
  24993=>"111111110",
  24994=>"110111111",
  24995=>"111111111",
  24996=>"000000001",
  24997=>"001000000",
  24998=>"111111111",
  24999=>"000000101",
  25000=>"101111000",
  25001=>"011010010",
  25002=>"110111111",
  25003=>"011010000",
  25004=>"111000000",
  25005=>"111111111",
  25006=>"000000000",
  25007=>"000000000",
  25008=>"000000011",
  25009=>"000000000",
  25010=>"000000000",
  25011=>"000000000",
  25012=>"000000010",
  25013=>"000000100",
  25014=>"111111111",
  25015=>"110110000",
  25016=>"000111101",
  25017=>"000000010",
  25018=>"111111111",
  25019=>"111111111",
  25020=>"100011111",
  25021=>"111110111",
  25022=>"111111011",
  25023=>"011111111",
  25024=>"000000000",
  25025=>"111111111",
  25026=>"000000000",
  25027=>"000000000",
  25028=>"000101111",
  25029=>"000000010",
  25030=>"111110000",
  25031=>"000000000",
  25032=>"000000000",
  25033=>"111111100",
  25034=>"000000111",
  25035=>"111111111",
  25036=>"100000000",
  25037=>"100000000",
  25038=>"000001100",
  25039=>"011111111",
  25040=>"111101111",
  25041=>"010011110",
  25042=>"100110111",
  25043=>"000000000",
  25044=>"000000000",
  25045=>"000000110",
  25046=>"110111000",
  25047=>"010010010",
  25048=>"011111111",
  25049=>"111111111",
  25050=>"111111111",
  25051=>"100111111",
  25052=>"000000000",
  25053=>"111111111",
  25054=>"000101111",
  25055=>"011111111",
  25056=>"000000111",
  25057=>"000000000",
  25058=>"011000111",
  25059=>"111011001",
  25060=>"100000111",
  25061=>"111111111",
  25062=>"000000010",
  25063=>"000000010",
  25064=>"101001101",
  25065=>"000000010",
  25066=>"000000000",
  25067=>"000001111",
  25068=>"111001000",
  25069=>"111101000",
  25070=>"110000000",
  25071=>"111111111",
  25072=>"111111111",
  25073=>"000101111",
  25074=>"111100100",
  25075=>"110110000",
  25076=>"110110100",
  25077=>"111111000",
  25078=>"111111110",
  25079=>"111111111",
  25080=>"010100111",
  25081=>"100110100",
  25082=>"111001000",
  25083=>"110011000",
  25084=>"011001000",
  25085=>"101000000",
  25086=>"111111111",
  25087=>"000000000",
  25088=>"110111111",
  25089=>"110110000",
  25090=>"101111111",
  25091=>"000000000",
  25092=>"011001000",
  25093=>"000000000",
  25094=>"000111111",
  25095=>"000000100",
  25096=>"000111111",
  25097=>"000110111",
  25098=>"111111111",
  25099=>"101011001",
  25100=>"100011000",
  25101=>"000000000",
  25102=>"111111111",
  25103=>"000111010",
  25104=>"000000000",
  25105=>"000000000",
  25106=>"100111011",
  25107=>"111111111",
  25108=>"111111111",
  25109=>"111111111",
  25110=>"000011011",
  25111=>"000000000",
  25112=>"000000000",
  25113=>"111111111",
  25114=>"000000000",
  25115=>"000000011",
  25116=>"000000000",
  25117=>"101001001",
  25118=>"000000000",
  25119=>"111111110",
  25120=>"111101111",
  25121=>"000000000",
  25122=>"000100111",
  25123=>"000000000",
  25124=>"111100111",
  25125=>"000000000",
  25126=>"000000000",
  25127=>"000000000",
  25128=>"110100111",
  25129=>"000000110",
  25130=>"111010010",
  25131=>"000000011",
  25132=>"000000011",
  25133=>"000000000",
  25134=>"111111111",
  25135=>"100101001",
  25136=>"000010011",
  25137=>"000000000",
  25138=>"000000000",
  25139=>"000000000",
  25140=>"101101000",
  25141=>"111111110",
  25142=>"111101111",
  25143=>"111110110",
  25144=>"011111111",
  25145=>"001000000",
  25146=>"000000100",
  25147=>"000000000",
  25148=>"000000000",
  25149=>"100100111",
  25150=>"111110111",
  25151=>"000000000",
  25152=>"001001100",
  25153=>"000000000",
  25154=>"000110110",
  25155=>"000000111",
  25156=>"000000110",
  25157=>"111111111",
  25158=>"000000000",
  25159=>"000111111",
  25160=>"000000010",
  25161=>"111111111",
  25162=>"111111110",
  25163=>"000100000",
  25164=>"000000000",
  25165=>"100000110",
  25166=>"111111111",
  25167=>"000000000",
  25168=>"100000111",
  25169=>"111111111",
  25170=>"110110110",
  25171=>"000000000",
  25172=>"000000000",
  25173=>"000000000",
  25174=>"001001000",
  25175=>"110010010",
  25176=>"001000000",
  25177=>"000000000",
  25178=>"001111111",
  25179=>"111100100",
  25180=>"110110111",
  25181=>"001111011",
  25182=>"100100110",
  25183=>"011111010",
  25184=>"111111011",
  25185=>"000000000",
  25186=>"011001111",
  25187=>"111010000",
  25188=>"111110110",
  25189=>"111111010",
  25190=>"001000111",
  25191=>"111111000",
  25192=>"000000000",
  25193=>"111111110",
  25194=>"111110110",
  25195=>"111111111",
  25196=>"111111100",
  25197=>"111111111",
  25198=>"000000000",
  25199=>"000000000",
  25200=>"000000000",
  25201=>"000000000",
  25202=>"110110111",
  25203=>"000000000",
  25204=>"111111110",
  25205=>"000000111",
  25206=>"111111111",
  25207=>"110111111",
  25208=>"010000000",
  25209=>"000000000",
  25210=>"001000000",
  25211=>"111000111",
  25212=>"000000000",
  25213=>"111100110",
  25214=>"111111111",
  25215=>"000000000",
  25216=>"111011011",
  25217=>"000000000",
  25218=>"110100000",
  25219=>"001001000",
  25220=>"000000000",
  25221=>"111111111",
  25222=>"110111110",
  25223=>"000000011",
  25224=>"100000001",
  25225=>"000000000",
  25226=>"000110111",
  25227=>"111111111",
  25228=>"000000001",
  25229=>"110111111",
  25230=>"100000011",
  25231=>"000000111",
  25232=>"111100111",
  25233=>"111101001",
  25234=>"111111111",
  25235=>"000000000",
  25236=>"100101011",
  25237=>"100100100",
  25238=>"000000000",
  25239=>"000000011",
  25240=>"000111111",
  25241=>"111111001",
  25242=>"000000000",
  25243=>"000100100",
  25244=>"000001111",
  25245=>"110100000",
  25246=>"000000000",
  25247=>"000000000",
  25248=>"110111000",
  25249=>"000000100",
  25250=>"011111111",
  25251=>"111111111",
  25252=>"000000000",
  25253=>"111100110",
  25254=>"101000000",
  25255=>"011011011",
  25256=>"000000000",
  25257=>"111000111",
  25258=>"100000000",
  25259=>"111011111",
  25260=>"111110110",
  25261=>"000000000",
  25262=>"011011010",
  25263=>"101111101",
  25264=>"010111111",
  25265=>"111111111",
  25266=>"110111111",
  25267=>"000000000",
  25268=>"111111111",
  25269=>"000000000",
  25270=>"000000000",
  25271=>"000010110",
  25272=>"111011111",
  25273=>"100000111",
  25274=>"000000000",
  25275=>"000000001",
  25276=>"111100111",
  25277=>"000000100",
  25278=>"110001110",
  25279=>"000111101",
  25280=>"001101111",
  25281=>"011001111",
  25282=>"000000000",
  25283=>"111111000",
  25284=>"000100011",
  25285=>"000000011",
  25286=>"100000000",
  25287=>"000000000",
  25288=>"001111111",
  25289=>"000000100",
  25290=>"100100001",
  25291=>"000000000",
  25292=>"000000000",
  25293=>"000001000",
  25294=>"000000000",
  25295=>"000000010",
  25296=>"000000001",
  25297=>"001000000",
  25298=>"111111100",
  25299=>"000000000",
  25300=>"111111111",
  25301=>"010011111",
  25302=>"000110110",
  25303=>"111111000",
  25304=>"000000111",
  25305=>"000000111",
  25306=>"111111111",
  25307=>"001010010",
  25308=>"000010100",
  25309=>"111111111",
  25310=>"111001000",
  25311=>"100000110",
  25312=>"011111111",
  25313=>"000000011",
  25314=>"111000000",
  25315=>"000000000",
  25316=>"101101000",
  25317=>"100100111",
  25318=>"000000000",
  25319=>"000000001",
  25320=>"000000000",
  25321=>"000000000",
  25322=>"111001111",
  25323=>"000000000",
  25324=>"000000000",
  25325=>"111111111",
  25326=>"110111111",
  25327=>"000110110",
  25328=>"111111111",
  25329=>"000000001",
  25330=>"111111111",
  25331=>"000000000",
  25332=>"110111111",
  25333=>"000000000",
  25334=>"111111111",
  25335=>"000110111",
  25336=>"110111111",
  25337=>"000000000",
  25338=>"110111111",
  25339=>"111111111",
  25340=>"100000000",
  25341=>"101100000",
  25342=>"111110110",
  25343=>"000110110",
  25344=>"111111111",
  25345=>"000000000",
  25346=>"100111111",
  25347=>"000000110",
  25348=>"110100100",
  25349=>"111111111",
  25350=>"101111111",
  25351=>"000000000",
  25352=>"111111111",
  25353=>"000000000",
  25354=>"100111111",
  25355=>"001111111",
  25356=>"100101000",
  25357=>"111111111",
  25358=>"000000000",
  25359=>"111111000",
  25360=>"100000111",
  25361=>"111111111",
  25362=>"000000000",
  25363=>"001011011",
  25364=>"111111111",
  25365=>"000000001",
  25366=>"100100100",
  25367=>"000000000",
  25368=>"111111110",
  25369=>"000000000",
  25370=>"000000000",
  25371=>"000000000",
  25372=>"000000000",
  25373=>"000000001",
  25374=>"111001000",
  25375=>"111111111",
  25376=>"100100000",
  25377=>"111111111",
  25378=>"111111111",
  25379=>"111111111",
  25380=>"000000000",
  25381=>"111111110",
  25382=>"000000001",
  25383=>"110110111",
  25384=>"111111111",
  25385=>"000000000",
  25386=>"100000000",
  25387=>"011000000",
  25388=>"011011111",
  25389=>"000000000",
  25390=>"111110010",
  25391=>"000110111",
  25392=>"001000011",
  25393=>"000000000",
  25394=>"110100100",
  25395=>"111111111",
  25396=>"000000010",
  25397=>"111111111",
  25398=>"111101001",
  25399=>"110110111",
  25400=>"000000000",
  25401=>"000000111",
  25402=>"111111111",
  25403=>"111111000",
  25404=>"011000000",
  25405=>"001000000",
  25406=>"111111111",
  25407=>"000100100",
  25408=>"000000000",
  25409=>"000000000",
  25410=>"000000110",
  25411=>"111010010",
  25412=>"001000000",
  25413=>"111111110",
  25414=>"000000000",
  25415=>"111111111",
  25416=>"000000000",
  25417=>"000000000",
  25418=>"110111111",
  25419=>"000000000",
  25420=>"000000000",
  25421=>"000000001",
  25422=>"100000000",
  25423=>"111111000",
  25424=>"000001001",
  25425=>"111111111",
  25426=>"001010000",
  25427=>"000110110",
  25428=>"000000011",
  25429=>"000000001",
  25430=>"000000000",
  25431=>"100000000",
  25432=>"000000000",
  25433=>"000000000",
  25434=>"111111111",
  25435=>"000000000",
  25436=>"001000001",
  25437=>"111111110",
  25438=>"111111111",
  25439=>"000011110",
  25440=>"111111111",
  25441=>"111111000",
  25442=>"000000000",
  25443=>"000111111",
  25444=>"001011111",
  25445=>"110000000",
  25446=>"111000111",
  25447=>"111111111",
  25448=>"000000000",
  25449=>"111111010",
  25450=>"111111000",
  25451=>"111111111",
  25452=>"000000110",
  25453=>"111111111",
  25454=>"100100000",
  25455=>"000000000",
  25456=>"111011111",
  25457=>"001001000",
  25458=>"000000000",
  25459=>"000000011",
  25460=>"000000001",
  25461=>"000101111",
  25462=>"000011001",
  25463=>"000100110",
  25464=>"000000000",
  25465=>"000000000",
  25466=>"111101111",
  25467=>"100100100",
  25468=>"111111111",
  25469=>"111111111",
  25470=>"111111100",
  25471=>"000101111",
  25472=>"111111110",
  25473=>"000000000",
  25474=>"111111111",
  25475=>"000000000",
  25476=>"100000000",
  25477=>"000000000",
  25478=>"100000000",
  25479=>"000000001",
  25480=>"111111111",
  25481=>"000101111",
  25482=>"111111111",
  25483=>"111111000",
  25484=>"111111111",
  25485=>"111111100",
  25486=>"110111111",
  25487=>"000000000",
  25488=>"000010010",
  25489=>"000000001",
  25490=>"111111111",
  25491=>"011111111",
  25492=>"111111011",
  25493=>"000001111",
  25494=>"000011111",
  25495=>"001000111",
  25496=>"111011111",
  25497=>"111110000",
  25498=>"000000101",
  25499=>"111111111",
  25500=>"000000000",
  25501=>"101111111",
  25502=>"110100000",
  25503=>"111111000",
  25504=>"000100111",
  25505=>"111100011",
  25506=>"001000000",
  25507=>"111111111",
  25508=>"000000000",
  25509=>"111111111",
  25510=>"111000000",
  25511=>"001111100",
  25512=>"100100000",
  25513=>"000000110",
  25514=>"111111111",
  25515=>"000000100",
  25516=>"000000000",
  25517=>"001111100",
  25518=>"000000110",
  25519=>"000000100",
  25520=>"000001000",
  25521=>"001011111",
  25522=>"000000000",
  25523=>"111111111",
  25524=>"000000000",
  25525=>"001010110",
  25526=>"111111111",
  25527=>"000101000",
  25528=>"000000000",
  25529=>"000000000",
  25530=>"110010000",
  25531=>"111111111",
  25532=>"011100000",
  25533=>"111111111",
  25534=>"000000000",
  25535=>"111111011",
  25536=>"000010111",
  25537=>"000000000",
  25538=>"111111111",
  25539=>"111111111",
  25540=>"000000000",
  25541=>"100000100",
  25542=>"001000000",
  25543=>"111011011",
  25544=>"000100001",
  25545=>"000111111",
  25546=>"000000111",
  25547=>"111100000",
  25548=>"100000000",
  25549=>"000000000",
  25550=>"000000000",
  25551=>"111111111",
  25552=>"110000000",
  25553=>"111110100",
  25554=>"000000000",
  25555=>"111010010",
  25556=>"000101001",
  25557=>"000000000",
  25558=>"111111111",
  25559=>"011011011",
  25560=>"000000000",
  25561=>"000000000",
  25562=>"010010000",
  25563=>"111111111",
  25564=>"000000000",
  25565=>"111111000",
  25566=>"000000000",
  25567=>"100110011",
  25568=>"000010111",
  25569=>"000010110",
  25570=>"000000000",
  25571=>"111111111",
  25572=>"000000000",
  25573=>"000000111",
  25574=>"000000000",
  25575=>"000000011",
  25576=>"000000000",
  25577=>"101101000",
  25578=>"011111011",
  25579=>"000000000",
  25580=>"111111111",
  25581=>"000000111",
  25582=>"101001111",
  25583=>"111111111",
  25584=>"000000000",
  25585=>"110100100",
  25586=>"111111111",
  25587=>"000000000",
  25588=>"000000111",
  25589=>"111100110",
  25590=>"000000000",
  25591=>"101000000",
  25592=>"110111111",
  25593=>"010011011",
  25594=>"111100100",
  25595=>"101111101",
  25596=>"111111111",
  25597=>"110110110",
  25598=>"000000000",
  25599=>"000111111",
  25600=>"000000100",
  25601=>"000000001",
  25602=>"111111111",
  25603=>"000110110",
  25604=>"100110001",
  25605=>"000000000",
  25606=>"001101101",
  25607=>"111101111",
  25608=>"000000110",
  25609=>"011111000",
  25610=>"101000001",
  25611=>"000011111",
  25612=>"000010000",
  25613=>"100000101",
  25614=>"000011111",
  25615=>"000000000",
  25616=>"100001111",
  25617=>"000000000",
  25618=>"100101000",
  25619=>"000001001",
  25620=>"001001011",
  25621=>"000000111",
  25622=>"111101111",
  25623=>"001011011",
  25624=>"000000111",
  25625=>"000001011",
  25626=>"110000000",
  25627=>"000010100",
  25628=>"001000111",
  25629=>"111100111",
  25630=>"111101111",
  25631=>"111111111",
  25632=>"000110111",
  25633=>"000000000",
  25634=>"110110000",
  25635=>"101111111",
  25636=>"000000000",
  25637=>"001000000",
  25638=>"000000000",
  25639=>"000000001",
  25640=>"001000001",
  25641=>"110111111",
  25642=>"001001111",
  25643=>"000001000",
  25644=>"001001001",
  25645=>"111111000",
  25646=>"000000000",
  25647=>"110111111",
  25648=>"001001101",
  25649=>"111111000",
  25650=>"000110110",
  25651=>"000000000",
  25652=>"111000100",
  25653=>"110110000",
  25654=>"110111111",
  25655=>"001101101",
  25656=>"000010010",
  25657=>"111111110",
  25658=>"110110100",
  25659=>"111001111",
  25660=>"111111111",
  25661=>"000001001",
  25662=>"000011011",
  25663=>"001000001",
  25664=>"001011011",
  25665=>"111100101",
  25666=>"100100100",
  25667=>"111000000",
  25668=>"110110110",
  25669=>"000001011",
  25670=>"000000000",
  25671=>"100111111",
  25672=>"111111100",
  25673=>"101101111",
  25674=>"011011011",
  25675=>"000001111",
  25676=>"011000000",
  25677=>"001001111",
  25678=>"010010000",
  25679=>"000000000",
  25680=>"101111100",
  25681=>"000010011",
  25682=>"000111111",
  25683=>"100110110",
  25684=>"000100000",
  25685=>"000000111",
  25686=>"011011001",
  25687=>"001011010",
  25688=>"110110000",
  25689=>"111101111",
  25690=>"100100010",
  25691=>"011111111",
  25692=>"111111000",
  25693=>"111001111",
  25694=>"101111111",
  25695=>"111111011",
  25696=>"000010000",
  25697=>"000101000",
  25698=>"000011011",
  25699=>"111111100",
  25700=>"111010100",
  25701=>"011111111",
  25702=>"100000100",
  25703=>"110000000",
  25704=>"001001001",
  25705=>"000100111",
  25706=>"110000100",
  25707=>"000001110",
  25708=>"100100000",
  25709=>"000010111",
  25710=>"111101111",
  25711=>"111111111",
  25712=>"000010010",
  25713=>"110110111",
  25714=>"111111111",
  25715=>"000000110",
  25716=>"001001111",
  25717=>"001000000",
  25718=>"000000000",
  25719=>"111100111",
  25720=>"101111111",
  25721=>"101001111",
  25722=>"111001000",
  25723=>"111111001",
  25724=>"111111100",
  25725=>"111111011",
  25726=>"101000001",
  25727=>"000000000",
  25728=>"000000000",
  25729=>"111101110",
  25730=>"111010000",
  25731=>"011111011",
  25732=>"001000000",
  25733=>"000000001",
  25734=>"110110110",
  25735=>"010101111",
  25736=>"000000110",
  25737=>"001001111",
  25738=>"101111111",
  25739=>"000001110",
  25740=>"000000111",
  25741=>"000000100",
  25742=>"000001011",
  25743=>"011001000",
  25744=>"111111111",
  25745=>"000110001",
  25746=>"111111110",
  25747=>"100110110",
  25748=>"001000000",
  25749=>"111000000",
  25750=>"111001001",
  25751=>"001001101",
  25752=>"001001111",
  25753=>"011110111",
  25754=>"110110010",
  25755=>"101000000",
  25756=>"000000110",
  25757=>"111100000",
  25758=>"110011001",
  25759=>"111111111",
  25760=>"011000000",
  25761=>"111110111",
  25762=>"000000000",
  25763=>"101000001",
  25764=>"000111111",
  25765=>"101000000",
  25766=>"000010111",
  25767=>"011111110",
  25768=>"001111111",
  25769=>"100111111",
  25770=>"111111111",
  25771=>"001100111",
  25772=>"111000001",
  25773=>"100110100",
  25774=>"000000111",
  25775=>"110110000",
  25776=>"000010110",
  25777=>"000000101",
  25778=>"010111010",
  25779=>"101100100",
  25780=>"101000000",
  25781=>"000000101",
  25782=>"100100000",
  25783=>"111011000",
  25784=>"111111111",
  25785=>"111111111",
  25786=>"101001001",
  25787=>"001001100",
  25788=>"101101001",
  25789=>"001000100",
  25790=>"001111111",
  25791=>"000000000",
  25792=>"000000000",
  25793=>"001001001",
  25794=>"000000000",
  25795=>"111100110",
  25796=>"000111101",
  25797=>"000011110",
  25798=>"001000110",
  25799=>"000101111",
  25800=>"101100010",
  25801=>"001111111",
  25802=>"001001001",
  25803=>"101000000",
  25804=>"111111011",
  25805=>"000000000",
  25806=>"111100101",
  25807=>"111011000",
  25808=>"001001111",
  25809=>"111001111",
  25810=>"000110100",
  25811=>"100101101",
  25812=>"111111100",
  25813=>"111111010",
  25814=>"111100111",
  25815=>"010110001",
  25816=>"111001111",
  25817=>"000110110",
  25818=>"101101110",
  25819=>"111011111",
  25820=>"000000111",
  25821=>"111111111",
  25822=>"000000011",
  25823=>"001111001",
  25824=>"001011011",
  25825=>"000000111",
  25826=>"010000000",
  25827=>"111101000",
  25828=>"111001000",
  25829=>"000010011",
  25830=>"000010010",
  25831=>"111111111",
  25832=>"100100100",
  25833=>"110100011",
  25834=>"110110111",
  25835=>"000000000",
  25836=>"011111011",
  25837=>"000000000",
  25838=>"110110111",
  25839=>"111010010",
  25840=>"000000100",
  25841=>"111111100",
  25842=>"000110111",
  25843=>"000010010",
  25844=>"000110111",
  25845=>"110110110",
  25846=>"111100000",
  25847=>"111111111",
  25848=>"101000100",
  25849=>"011111111",
  25850=>"100000100",
  25851=>"001110000",
  25852=>"111111111",
  25853=>"001000011",
  25854=>"011000001",
  25855=>"101110000",
  25856=>"001001001",
  25857=>"011001011",
  25858=>"001000000",
  25859=>"111101111",
  25860=>"110110000",
  25861=>"111101111",
  25862=>"110110000",
  25863=>"000000001",
  25864=>"110110111",
  25865=>"011111111",
  25866=>"000000001",
  25867=>"110111010",
  25868=>"000100000",
  25869=>"000000000",
  25870=>"101100110",
  25871=>"111111111",
  25872=>"111111000",
  25873=>"011111111",
  25874=>"000111111",
  25875=>"000110110",
  25876=>"111110010",
  25877=>"000000100",
  25878=>"000001001",
  25879=>"000000011",
  25880=>"100100011",
  25881=>"001001001",
  25882=>"110111111",
  25883=>"100100111",
  25884=>"000000000",
  25885=>"000000000",
  25886=>"000000011",
  25887=>"111111111",
  25888=>"011010000",
  25889=>"101000001",
  25890=>"000111111",
  25891=>"110111111",
  25892=>"100110110",
  25893=>"001001111",
  25894=>"111111100",
  25895=>"110110000",
  25896=>"111101000",
  25897=>"010001000",
  25898=>"000110010",
  25899=>"011011001",
  25900=>"000000011",
  25901=>"111110110",
  25902=>"111111111",
  25903=>"110010000",
  25904=>"100100100",
  25905=>"001001011",
  25906=>"111111111",
  25907=>"111100110",
  25908=>"001101000",
  25909=>"100000110",
  25910=>"000111111",
  25911=>"111111000",
  25912=>"111111111",
  25913=>"111101101",
  25914=>"101001111",
  25915=>"001000011",
  25916=>"000000000",
  25917=>"110110000",
  25918=>"011000111",
  25919=>"110111110",
  25920=>"000011010",
  25921=>"001000111",
  25922=>"101000000",
  25923=>"001011111",
  25924=>"000000111",
  25925=>"111101000",
  25926=>"000001011",
  25927=>"000000111",
  25928=>"000110110",
  25929=>"000000111",
  25930=>"110110010",
  25931=>"010011011",
  25932=>"001000101",
  25933=>"100100111",
  25934=>"111111001",
  25935=>"100000100",
  25936=>"101111111",
  25937=>"101000110",
  25938=>"111111000",
  25939=>"000111101",
  25940=>"101111111",
  25941=>"011011001",
  25942=>"011001000",
  25943=>"101000100",
  25944=>"110110000",
  25945=>"100100111",
  25946=>"111110110",
  25947=>"000000111",
  25948=>"000110100",
  25949=>"111100100",
  25950=>"101000110",
  25951=>"110100000",
  25952=>"110001001",
  25953=>"001000001",
  25954=>"100110111",
  25955=>"011001000",
  25956=>"111110100",
  25957=>"111111001",
  25958=>"111001011",
  25959=>"001101111",
  25960=>"000111111",
  25961=>"011100111",
  25962=>"010011001",
  25963=>"101110111",
  25964=>"110110111",
  25965=>"111100000",
  25966=>"011111111",
  25967=>"100100111",
  25968=>"000000111",
  25969=>"111100000",
  25970=>"000000000",
  25971=>"001100100",
  25972=>"101111111",
  25973=>"000000110",
  25974=>"001000000",
  25975=>"110111111",
  25976=>"000000000",
  25977=>"000000000",
  25978=>"111111111",
  25979=>"000000000",
  25980=>"100100110",
  25981=>"001000001",
  25982=>"111111111",
  25983=>"001000000",
  25984=>"111111000",
  25985=>"110110010",
  25986=>"000000100",
  25987=>"000000001",
  25988=>"000000000",
  25989=>"111101111",
  25990=>"001111111",
  25991=>"111110110",
  25992=>"101100110",
  25993=>"000000010",
  25994=>"001000001",
  25995=>"111111111",
  25996=>"001000001",
  25997=>"100010100",
  25998=>"101001001",
  25999=>"111101111",
  26000=>"000000001",
  26001=>"001000001",
  26002=>"111111000",
  26003=>"000000000",
  26004=>"000001011",
  26005=>"000000001",
  26006=>"101110000",
  26007=>"000001001",
  26008=>"000000000",
  26009=>"101101100",
  26010=>"111111001",
  26011=>"111111111",
  26012=>"001001001",
  26013=>"001110000",
  26014=>"001000000",
  26015=>"001011111",
  26016=>"000000111",
  26017=>"011011001",
  26018=>"010111111",
  26019=>"100000000",
  26020=>"110110111",
  26021=>"000001000",
  26022=>"111111010",
  26023=>"111100110",
  26024=>"001001111",
  26025=>"000000111",
  26026=>"100000000",
  26027=>"111001001",
  26028=>"100100111",
  26029=>"110110001",
  26030=>"101110110",
  26031=>"001000101",
  26032=>"111110110",
  26033=>"111111101",
  26034=>"111110110",
  26035=>"001001011",
  26036=>"111000000",
  26037=>"001111111",
  26038=>"000000111",
  26039=>"111001001",
  26040=>"001000000",
  26041=>"000000000",
  26042=>"001000100",
  26043=>"001001000",
  26044=>"000000000",
  26045=>"000001111",
  26046=>"000000000",
  26047=>"001111111",
  26048=>"111111001",
  26049=>"001000000",
  26050=>"111111010",
  26051=>"001000000",
  26052=>"010000001",
  26053=>"010000111",
  26054=>"110000000",
  26055=>"001000000",
  26056=>"000011000",
  26057=>"000000111",
  26058=>"101111101",
  26059=>"111111110",
  26060=>"110000000",
  26061=>"110110111",
  26062=>"111100101",
  26063=>"100000010",
  26064=>"011011000",
  26065=>"111100100",
  26066=>"111111111",
  26067=>"111000000",
  26068=>"011111100",
  26069=>"100000000",
  26070=>"111000001",
  26071=>"000110010",
  26072=>"111111001",
  26073=>"001010011",
  26074=>"100010000",
  26075=>"000000010",
  26076=>"001001111",
  26077=>"110110010",
  26078=>"111011000",
  26079=>"001001111",
  26080=>"001001111",
  26081=>"000000110",
  26082=>"011111111",
  26083=>"001001000",
  26084=>"000111111",
  26085=>"111001001",
  26086=>"110110100",
  26087=>"101001001",
  26088=>"110110000",
  26089=>"000000000",
  26090=>"110110111",
  26091=>"110111100",
  26092=>"001000000",
  26093=>"111111000",
  26094=>"101111111",
  26095=>"000001101",
  26096=>"000000110",
  26097=>"110010000",
  26098=>"000011111",
  26099=>"001011001",
  26100=>"110110101",
  26101=>"111111101",
  26102=>"111111111",
  26103=>"110110110",
  26104=>"110001011",
  26105=>"100110111",
  26106=>"000000110",
  26107=>"111111111",
  26108=>"111000101",
  26109=>"111011001",
  26110=>"111111111",
  26111=>"001001101",
  26112=>"001011000",
  26113=>"000000000",
  26114=>"001000001",
  26115=>"000001000",
  26116=>"110111101",
  26117=>"001001001",
  26118=>"111110100",
  26119=>"111111111",
  26120=>"000000001",
  26121=>"000111111",
  26122=>"111111110",
  26123=>"101001000",
  26124=>"100111111",
  26125=>"001000000",
  26126=>"111111111",
  26127=>"000001000",
  26128=>"111100111",
  26129=>"000111011",
  26130=>"110110110",
  26131=>"000001111",
  26132=>"000000011",
  26133=>"111111111",
  26134=>"111101101",
  26135=>"110110111",
  26136=>"110110110",
  26137=>"111011110",
  26138=>"111111111",
  26139=>"010000001",
  26140=>"000000000",
  26141=>"111111111",
  26142=>"011001001",
  26143=>"000001001",
  26144=>"110110100",
  26145=>"110100100",
  26146=>"110110110",
  26147=>"010010110",
  26148=>"000000000",
  26149=>"000000000",
  26150=>"001101000",
  26151=>"110111000",
  26152=>"001001001",
  26153=>"000000000",
  26154=>"000011011",
  26155=>"000000000",
  26156=>"001000000",
  26157=>"011111000",
  26158=>"000001000",
  26159=>"111111111",
  26160=>"000101001",
  26161=>"000100000",
  26162=>"011011111",
  26163=>"000000010",
  26164=>"011111111",
  26165=>"000000100",
  26166=>"000001001",
  26167=>"111000000",
  26168=>"111000110",
  26169=>"111111111",
  26170=>"000000000",
  26171=>"101111111",
  26172=>"000000001",
  26173=>"110111111",
  26174=>"111100100",
  26175=>"111110110",
  26176=>"111001001",
  26177=>"111111111",
  26178=>"000000111",
  26179=>"111110001",
  26180=>"110110110",
  26181=>"101100100",
  26182=>"111001000",
  26183=>"100100100",
  26184=>"111111111",
  26185=>"000000000",
  26186=>"000000001",
  26187=>"111011111",
  26188=>"100100110",
  26189=>"111001001",
  26190=>"001000000",
  26191=>"011110110",
  26192=>"111110010",
  26193=>"100100011",
  26194=>"111000000",
  26195=>"001000000",
  26196=>"000100111",
  26197=>"000000111",
  26198=>"111101100",
  26199=>"000101100",
  26200=>"001001101",
  26201=>"001001111",
  26202=>"011011000",
  26203=>"100110011",
  26204=>"111101000",
  26205=>"000000101",
  26206=>"000000000",
  26207=>"001110100",
  26208=>"110010010",
  26209=>"011010111",
  26210=>"000000000",
  26211=>"000000000",
  26212=>"110011010",
  26213=>"101100000",
  26214=>"111011011",
  26215=>"000010000",
  26216=>"000110110",
  26217=>"111111000",
  26218=>"111100000",
  26219=>"000010111",
  26220=>"111111111",
  26221=>"111010000",
  26222=>"110000000",
  26223=>"100111111",
  26224=>"110110110",
  26225=>"101100110",
  26226=>"001001001",
  26227=>"000000100",
  26228=>"000111111",
  26229=>"110110111",
  26230=>"010111111",
  26231=>"110110110",
  26232=>"000001000",
  26233=>"000000011",
  26234=>"100100110",
  26235=>"100100000",
  26236=>"100000100",
  26237=>"001111111",
  26238=>"100000000",
  26239=>"111111111",
  26240=>"000000000",
  26241=>"110000000",
  26242=>"000000000",
  26243=>"000000000",
  26244=>"000000000",
  26245=>"111010000",
  26246=>"001011011",
  26247=>"111111000",
  26248=>"001000000",
  26249=>"111111111",
  26250=>"000000000",
  26251=>"000000111",
  26252=>"001001001",
  26253=>"110110110",
  26254=>"110000000",
  26255=>"010010010",
  26256=>"001001001",
  26257=>"111001011",
  26258=>"111111001",
  26259=>"011000111",
  26260=>"011000000",
  26261=>"111001000",
  26262=>"001001001",
  26263=>"001100000",
  26264=>"001001001",
  26265=>"111111111",
  26266=>"010000000",
  26267=>"111101001",
  26268=>"100000001",
  26269=>"001111110",
  26270=>"000000000",
  26271=>"000000000",
  26272=>"000000000",
  26273=>"000110010",
  26274=>"111111111",
  26275=>"000111010",
  26276=>"000101001",
  26277=>"110110011",
  26278=>"001000101",
  26279=>"100000000",
  26280=>"101001101",
  26281=>"000000000",
  26282=>"000000000",
  26283=>"111101110",
  26284=>"001000101",
  26285=>"000110111",
  26286=>"111101110",
  26287=>"001001000",
  26288=>"111111110",
  26289=>"000011000",
  26290=>"111110110",
  26291=>"000000000",
  26292=>"000000000",
  26293=>"111110111",
  26294=>"000100000",
  26295=>"111111001",
  26296=>"101001000",
  26297=>"111111111",
  26298=>"100111101",
  26299=>"101111000",
  26300=>"000111111",
  26301=>"111111111",
  26302=>"100000000",
  26303=>"111110000",
  26304=>"000000000",
  26305=>"110110000",
  26306=>"000000000",
  26307=>"110110010",
  26308=>"100000000",
  26309=>"000100110",
  26310=>"000100100",
  26311=>"000000100",
  26312=>"110110000",
  26313=>"000000000",
  26314=>"000010111",
  26315=>"110111111",
  26316=>"111001011",
  26317=>"111010000",
  26318=>"101100100",
  26319=>"001101110",
  26320=>"000011000",
  26321=>"100000000",
  26322=>"111011000",
  26323=>"000000000",
  26324=>"001000001",
  26325=>"100100000",
  26326=>"000000110",
  26327=>"001011001",
  26328=>"010100000",
  26329=>"110110110",
  26330=>"001000101",
  26331=>"110111111",
  26332=>"000000000",
  26333=>"001000000",
  26334=>"000000001",
  26335=>"000010111",
  26336=>"011000010",
  26337=>"010000001",
  26338=>"000001000",
  26339=>"000000000",
  26340=>"011000111",
  26341=>"111011011",
  26342=>"000000000",
  26343=>"111111111",
  26344=>"100110000",
  26345=>"011001100",
  26346=>"110110110",
  26347=>"000000000",
  26348=>"000000000",
  26349=>"000000111",
  26350=>"011011110",
  26351=>"111111000",
  26352=>"111111000",
  26353=>"111111110",
  26354=>"110010010",
  26355=>"001001000",
  26356=>"100100101",
  26357=>"100001011",
  26358=>"101100100",
  26359=>"000000111",
  26360=>"111111110",
  26361=>"000000001",
  26362=>"101111111",
  26363=>"111001001",
  26364=>"111110111",
  26365=>"000100110",
  26366=>"111111111",
  26367=>"110100000",
  26368=>"110000010",
  26369=>"001101101",
  26370=>"110110000",
  26371=>"000001100",
  26372=>"000000000",
  26373=>"111011001",
  26374=>"001000110",
  26375=>"001000110",
  26376=>"111111111",
  26377=>"111111111",
  26378=>"001000000",
  26379=>"000110000",
  26380=>"100000000",
  26381=>"011100110",
  26382=>"000000000",
  26383=>"111111100",
  26384=>"111100000",
  26385=>"101111110",
  26386=>"001001011",
  26387=>"000001111",
  26388=>"000000000",
  26389=>"001111111",
  26390=>"110111111",
  26391=>"110000000",
  26392=>"101100000",
  26393=>"111101001",
  26394=>"000000000",
  26395=>"110000100",
  26396=>"110110110",
  26397=>"111111001",
  26398=>"010001000",
  26399=>"111111111",
  26400=>"001000001",
  26401=>"111111000",
  26402=>"000000000",
  26403=>"000000000",
  26404=>"000000000",
  26405=>"000000000",
  26406=>"111111111",
  26407=>"001011111",
  26408=>"110110110",
  26409=>"110111110",
  26410=>"001111111",
  26411=>"001000000",
  26412=>"110100111",
  26413=>"110111111",
  26414=>"000000000",
  26415=>"001000000",
  26416=>"111111101",
  26417=>"111110111",
  26418=>"001001001",
  26419=>"000000000",
  26420=>"000000000",
  26421=>"000000100",
  26422=>"001001011",
  26423=>"001001001",
  26424=>"011011111",
  26425=>"000000111",
  26426=>"110110110",
  26427=>"110000000",
  26428=>"011111111",
  26429=>"001100001",
  26430=>"001001101",
  26431=>"001001000",
  26432=>"111101111",
  26433=>"101001000",
  26434=>"001000000",
  26435=>"000011111",
  26436=>"111111110",
  26437=>"111001001",
  26438=>"100101101",
  26439=>"111001111",
  26440=>"000001101",
  26441=>"000001001",
  26442=>"000001000",
  26443=>"000000100",
  26444=>"000000000",
  26445=>"000000000",
  26446=>"111101001",
  26447=>"000000000",
  26448=>"111101101",
  26449=>"111111001",
  26450=>"000000000",
  26451=>"111111100",
  26452=>"011111000",
  26453=>"011011011",
  26454=>"111111111",
  26455=>"111111011",
  26456=>"001001101",
  26457=>"110110000",
  26458=>"000000001",
  26459=>"111111100",
  26460=>"011011011",
  26461=>"000000000",
  26462=>"010110010",
  26463=>"000000001",
  26464=>"001111101",
  26465=>"111111111",
  26466=>"100100100",
  26467=>"101101001",
  26468=>"001000001",
  26469=>"001001001",
  26470=>"011111001",
  26471=>"100000111",
  26472=>"001000101",
  26473=>"110111100",
  26474=>"001000000",
  26475=>"111000000",
  26476=>"000001001",
  26477=>"101001001",
  26478=>"000000000",
  26479=>"101000000",
  26480=>"110110110",
  26481=>"110101101",
  26482=>"000100000",
  26483=>"111111111",
  26484=>"110111111",
  26485=>"000110010",
  26486=>"111110000",
  26487=>"001101111",
  26488=>"000000000",
  26489=>"111001000",
  26490=>"001011111",
  26491=>"000000000",
  26492=>"000110110",
  26493=>"110110110",
  26494=>"011011111",
  26495=>"001000000",
  26496=>"111101111",
  26497=>"001000110",
  26498=>"100000001",
  26499=>"000000000",
  26500=>"001000000",
  26501=>"000000000",
  26502=>"000000000",
  26503=>"110111110",
  26504=>"000000000",
  26505=>"000111000",
  26506=>"000000010",
  26507=>"111110000",
  26508=>"001000001",
  26509=>"100111010",
  26510=>"001000000",
  26511=>"000000000",
  26512=>"101100110",
  26513=>"110110110",
  26514=>"001001011",
  26515=>"101001001",
  26516=>"000010010",
  26517=>"000000000",
  26518=>"000000000",
  26519=>"011111111",
  26520=>"000000110",
  26521=>"000110111",
  26522=>"101101001",
  26523=>"001000001",
  26524=>"111101100",
  26525=>"110110100",
  26526=>"000000000",
  26527=>"001111111",
  26528=>"110110100",
  26529=>"011011111",
  26530=>"110011110",
  26531=>"001000001",
  26532=>"110111110",
  26533=>"111111011",
  26534=>"111011000",
  26535=>"000000001",
  26536=>"010111110",
  26537=>"110111011",
  26538=>"110000001",
  26539=>"111000000",
  26540=>"111000100",
  26541=>"111111000",
  26542=>"110111111",
  26543=>"111100100",
  26544=>"111101101",
  26545=>"010010110",
  26546=>"000001001",
  26547=>"011000000",
  26548=>"011110010",
  26549=>"001001101",
  26550=>"001001101",
  26551=>"111111111",
  26552=>"001000000",
  26553=>"111111111",
  26554=>"000001011",
  26555=>"111111101",
  26556=>"001001111",
  26557=>"000000000",
  26558=>"101101100",
  26559=>"111111101",
  26560=>"110110110",
  26561=>"111110011",
  26562=>"111111000",
  26563=>"000000000",
  26564=>"111111111",
  26565=>"001100100",
  26566=>"111111111",
  26567=>"011011000",
  26568=>"001000001",
  26569=>"111001011",
  26570=>"011011011",
  26571=>"001000111",
  26572=>"111000111",
  26573=>"001001001",
  26574=>"000000000",
  26575=>"011001000",
  26576=>"000000000",
  26577=>"111111111",
  26578=>"000001001",
  26579=>"111111111",
  26580=>"101100101",
  26581=>"111111111",
  26582=>"010000000",
  26583=>"011010111",
  26584=>"100100110",
  26585=>"110011011",
  26586=>"001101000",
  26587=>"000000000",
  26588=>"000000000",
  26589=>"111111001",
  26590=>"111111000",
  26591=>"100100000",
  26592=>"111111000",
  26593=>"000110110",
  26594=>"000000100",
  26595=>"100100100",
  26596=>"001001111",
  26597=>"100000001",
  26598=>"000000100",
  26599=>"000000001",
  26600=>"111000000",
  26601=>"110110010",
  26602=>"111111101",
  26603=>"111110010",
  26604=>"110110110",
  26605=>"101101111",
  26606=>"000100101",
  26607=>"111111110",
  26608=>"100100100",
  26609=>"111001000",
  26610=>"111111111",
  26611=>"111101100",
  26612=>"110110110",
  26613=>"111101000",
  26614=>"111100000",
  26615=>"111100111",
  26616=>"110010010",
  26617=>"010110110",
  26618=>"110111001",
  26619=>"111111111",
  26620=>"111101111",
  26621=>"111111111",
  26622=>"111111111",
  26623=>"001000000",
  26624=>"111111000",
  26625=>"110000100",
  26626=>"100100110",
  26627=>"000001011",
  26628=>"111111011",
  26629=>"111111111",
  26630=>"111111111",
  26631=>"000000111",
  26632=>"000000000",
  26633=>"000011011",
  26634=>"111101111",
  26635=>"001000011",
  26636=>"100100110",
  26637=>"011111111",
  26638=>"110000000",
  26639=>"111111111",
  26640=>"000110100",
  26641=>"000000111",
  26642=>"011000000",
  26643=>"111111111",
  26644=>"000000000",
  26645=>"001111110",
  26646=>"100111111",
  26647=>"111001101",
  26648=>"100100101",
  26649=>"001001000",
  26650=>"111111111",
  26651=>"000010111",
  26652=>"000000000",
  26653=>"111111111",
  26654=>"100000000",
  26655=>"100000000",
  26656=>"010000000",
  26657=>"000000000",
  26658=>"111111101",
  26659=>"110000000",
  26660=>"111011111",
  26661=>"011110111",
  26662=>"000000111",
  26663=>"111000000",
  26664=>"001000000",
  26665=>"111111111",
  26666=>"000000100",
  26667=>"111111111",
  26668=>"000000000",
  26669=>"000000000",
  26670=>"111000011",
  26671=>"111011001",
  26672=>"000000000",
  26673=>"111010010",
  26674=>"000000000",
  26675=>"000000001",
  26676=>"111111111",
  26677=>"110111111",
  26678=>"111111111",
  26679=>"001011111",
  26680=>"000000000",
  26681=>"110111000",
  26682=>"111111111",
  26683=>"111111111",
  26684=>"111111001",
  26685=>"110100110",
  26686=>"000000000",
  26687=>"111111111",
  26688=>"011000000",
  26689=>"011011011",
  26690=>"111000100",
  26691=>"110000001",
  26692=>"110100100",
  26693=>"011011111",
  26694=>"111111110",
  26695=>"111011011",
  26696=>"001001000",
  26697=>"000011011",
  26698=>"000000111",
  26699=>"111011010",
  26700=>"111101111",
  26701=>"000000000",
  26702=>"111111111",
  26703=>"000000000",
  26704=>"000000000",
  26705=>"111111111",
  26706=>"000000000",
  26707=>"100111111",
  26708=>"000000000",
  26709=>"111111000",
  26710=>"111100100",
  26711=>"000000000",
  26712=>"000000000",
  26713=>"111101100",
  26714=>"000000000",
  26715=>"100000000",
  26716=>"000110111",
  26717=>"000111111",
  26718=>"000000000",
  26719=>"000001000",
  26720=>"010000000",
  26721=>"000000000",
  26722=>"111111111",
  26723=>"000000000",
  26724=>"100000000",
  26725=>"111111111",
  26726=>"111111111",
  26727=>"111111110",
  26728=>"000000000",
  26729=>"000000001",
  26730=>"111110110",
  26731=>"000000111",
  26732=>"111010000",
  26733=>"001111000",
  26734=>"111111111",
  26735=>"000010010",
  26736=>"111111111",
  26737=>"000000000",
  26738=>"101101101",
  26739=>"100111000",
  26740=>"111111111",
  26741=>"000000110",
  26742=>"000110111",
  26743=>"111111111",
  26744=>"000000000",
  26745=>"110110111",
  26746=>"110000000",
  26747=>"000000100",
  26748=>"110100100",
  26749=>"011000000",
  26750=>"110000000",
  26751=>"111111111",
  26752=>"111111111",
  26753=>"000001000",
  26754=>"011111111",
  26755=>"101111111",
  26756=>"111111111",
  26757=>"100111111",
  26758=>"101001111",
  26759=>"000000000",
  26760=>"111011111",
  26761=>"011111111",
  26762=>"000000000",
  26763=>"000000001",
  26764=>"000100111",
  26765=>"111101111",
  26766=>"111000000",
  26767=>"010000000",
  26768=>"000000000",
  26769=>"100110111",
  26770=>"000000111",
  26771=>"110000011",
  26772=>"111000001",
  26773=>"010010001",
  26774=>"000000110",
  26775=>"111111111",
  26776=>"000100011",
  26777=>"011001111",
  26778=>"111111111",
  26779=>"000000000",
  26780=>"111111111",
  26781=>"000010111",
  26782=>"100000111",
  26783=>"000011111",
  26784=>"000000000",
  26785=>"111111111",
  26786=>"000000000",
  26787=>"100110111",
  26788=>"000000000",
  26789=>"111111110",
  26790=>"000000000",
  26791=>"000110111",
  26792=>"110110111",
  26793=>"000000000",
  26794=>"000000110",
  26795=>"111011011",
  26796=>"000010111",
  26797=>"111111111",
  26798=>"111000100",
  26799=>"111111101",
  26800=>"000001001",
  26801=>"000000000",
  26802=>"111111111",
  26803=>"001111111",
  26804=>"000000000",
  26805=>"111111000",
  26806=>"111101111",
  26807=>"000000000",
  26808=>"000000000",
  26809=>"101100111",
  26810=>"010000000",
  26811=>"010000100",
  26812=>"111000011",
  26813=>"010000000",
  26814=>"001111111",
  26815=>"010111010",
  26816=>"111111111",
  26817=>"000000111",
  26818=>"000000000",
  26819=>"000000110",
  26820=>"000000000",
  26821=>"100101111",
  26822=>"101111111",
  26823=>"000000001",
  26824=>"111111110",
  26825=>"011000000",
  26826=>"111000000",
  26827=>"000000000",
  26828=>"111101000",
  26829=>"000111111",
  26830=>"011011111",
  26831=>"000000000",
  26832=>"111000111",
  26833=>"000000000",
  26834=>"111111100",
  26835=>"000000000",
  26836=>"111111111",
  26837=>"111111111",
  26838=>"000000000",
  26839=>"111111101",
  26840=>"111111100",
  26841=>"111111111",
  26842=>"000000000",
  26843=>"111111111",
  26844=>"000000100",
  26845=>"001000001",
  26846=>"001011111",
  26847=>"001000000",
  26848=>"000111111",
  26849=>"001100000",
  26850=>"000000000",
  26851=>"111100000",
  26852=>"111000011",
  26853=>"001001001",
  26854=>"000000000",
  26855=>"111111111",
  26856=>"111111001",
  26857=>"000000000",
  26858=>"001101111",
  26859=>"000000000",
  26860=>"111111111",
  26861=>"111111111",
  26862=>"000010111",
  26863=>"000110100",
  26864=>"101100111",
  26865=>"000011000",
  26866=>"000000000",
  26867=>"000000000",
  26868=>"000010110",
  26869=>"111100000",
  26870=>"111111100",
  26871=>"111111111",
  26872=>"000000000",
  26873=>"111111111",
  26874=>"111110111",
  26875=>"000100110",
  26876=>"011011001",
  26877=>"111111111",
  26878=>"011001001",
  26879=>"011111111",
  26880=>"111111100",
  26881=>"111111111",
  26882=>"010000000",
  26883=>"111111111",
  26884=>"111111111",
  26885=>"111111111",
  26886=>"101111111",
  26887=>"111111111",
  26888=>"101111111",
  26889=>"110000100",
  26890=>"000000101",
  26891=>"111001111",
  26892=>"000000000",
  26893=>"111111000",
  26894=>"001111111",
  26895=>"011111111",
  26896=>"000000000",
  26897=>"011011000",
  26898=>"000000010",
  26899=>"111111111",
  26900=>"000000000",
  26901=>"001000110",
  26902=>"111111111",
  26903=>"001111111",
  26904=>"001000000",
  26905=>"011000000",
  26906=>"111011000",
  26907=>"000000000",
  26908=>"000000000",
  26909=>"111111111",
  26910=>"111111110",
  26911=>"000000110",
  26912=>"110011111",
  26913=>"000000000",
  26914=>"000000000",
  26915=>"111011111",
  26916=>"000000111",
  26917=>"001011111",
  26918=>"000000000",
  26919=>"000000010",
  26920=>"101100100",
  26921=>"000000000",
  26922=>"111000000",
  26923=>"000000100",
  26924=>"000000000",
  26925=>"011011011",
  26926=>"111111111",
  26927=>"000000000",
  26928=>"000100000",
  26929=>"001010000",
  26930=>"111000100",
  26931=>"001111111",
  26932=>"111111111",
  26933=>"011011111",
  26934=>"111111111",
  26935=>"111111111",
  26936=>"000001000",
  26937=>"000000000",
  26938=>"111100000",
  26939=>"011111111",
  26940=>"110110111",
  26941=>"111100000",
  26942=>"110000000",
  26943=>"111111001",
  26944=>"001000100",
  26945=>"100000000",
  26946=>"100000001",
  26947=>"111101111",
  26948=>"111111111",
  26949=>"111111100",
  26950=>"000000000",
  26951=>"000000111",
  26952=>"000000000",
  26953=>"000000000",
  26954=>"000000000",
  26955=>"110001001",
  26956=>"110100100",
  26957=>"111011111",
  26958=>"111100000",
  26959=>"111111111",
  26960=>"001011000",
  26961=>"111111011",
  26962=>"000000000",
  26963=>"111000001",
  26964=>"001000000",
  26965=>"001001001",
  26966=>"000000000",
  26967=>"101101000",
  26968=>"111111100",
  26969=>"111111111",
  26970=>"111111010",
  26971=>"110111011",
  26972=>"111111111",
  26973=>"111100000",
  26974=>"000000001",
  26975=>"110000000",
  26976=>"001011001",
  26977=>"000000000",
  26978=>"000000001",
  26979=>"111111111",
  26980=>"111111111",
  26981=>"000000000",
  26982=>"111111111",
  26983=>"111111111",
  26984=>"001000100",
  26985=>"000000111",
  26986=>"111111000",
  26987=>"011011000",
  26988=>"110111111",
  26989=>"000000000",
  26990=>"000000000",
  26991=>"111111000",
  26992=>"111111111",
  26993=>"011111111",
  26994=>"000111111",
  26995=>"111111111",
  26996=>"110111110",
  26997=>"000011111",
  26998=>"110000000",
  26999=>"001011110",
  27000=>"101101111",
  27001=>"000000011",
  27002=>"000000000",
  27003=>"000110010",
  27004=>"111011000",
  27005=>"111000000",
  27006=>"000001001",
  27007=>"111111111",
  27008=>"110111111",
  27009=>"000000000",
  27010=>"000001011",
  27011=>"111101000",
  27012=>"000000111",
  27013=>"010111010",
  27014=>"000001100",
  27015=>"000000100",
  27016=>"000000000",
  27017=>"111111111",
  27018=>"110100000",
  27019=>"000000000",
  27020=>"111101111",
  27021=>"111111110",
  27022=>"001100110",
  27023=>"010000000",
  27024=>"010000010",
  27025=>"111111111",
  27026=>"000000000",
  27027=>"000000101",
  27028=>"111111111",
  27029=>"000000010",
  27030=>"111010000",
  27031=>"111111111",
  27032=>"000000110",
  27033=>"000000000",
  27034=>"000000010",
  27035=>"101001000",
  27036=>"000000001",
  27037=>"000000000",
  27038=>"000000000",
  27039=>"000000011",
  27040=>"000000010",
  27041=>"111111100",
  27042=>"111001000",
  27043=>"010000010",
  27044=>"011000000",
  27045=>"000000000",
  27046=>"000000001",
  27047=>"000000100",
  27048=>"111111111",
  27049=>"100111111",
  27050=>"110000000",
  27051=>"000000001",
  27052=>"111111110",
  27053=>"111111101",
  27054=>"000000100",
  27055=>"000000000",
  27056=>"111111111",
  27057=>"000101111",
  27058=>"011010010",
  27059=>"001001111",
  27060=>"000101111",
  27061=>"111111111",
  27062=>"111101001",
  27063=>"111111111",
  27064=>"111111111",
  27065=>"111111111",
  27066=>"111011010",
  27067=>"000100000",
  27068=>"000010000",
  27069=>"110110100",
  27070=>"111001001",
  27071=>"110100100",
  27072=>"111111011",
  27073=>"111111111",
  27074=>"111111001",
  27075=>"111111111",
  27076=>"000000001",
  27077=>"111111111",
  27078=>"000000000",
  27079=>"000000100",
  27080=>"000000110",
  27081=>"101111110",
  27082=>"001001011",
  27083=>"000011111",
  27084=>"111111011",
  27085=>"111011111",
  27086=>"111100000",
  27087=>"000010000",
  27088=>"000101101",
  27089=>"000000000",
  27090=>"111110100",
  27091=>"000011111",
  27092=>"111111111",
  27093=>"111111111",
  27094=>"111111011",
  27095=>"111111000",
  27096=>"100100111",
  27097=>"011000000",
  27098=>"010010010",
  27099=>"110110111",
  27100=>"000000000",
  27101=>"111101111",
  27102=>"111111111",
  27103=>"000000011",
  27104=>"001100100",
  27105=>"000100100",
  27106=>"111111111",
  27107=>"001001111",
  27108=>"111110110",
  27109=>"111111111",
  27110=>"000000111",
  27111=>"011011011",
  27112=>"111111111",
  27113=>"111111011",
  27114=>"111111111",
  27115=>"111111111",
  27116=>"111011111",
  27117=>"111111111",
  27118=>"111101111",
  27119=>"110110110",
  27120=>"000000000",
  27121=>"011011111",
  27122=>"011000011",
  27123=>"000000000",
  27124=>"000100111",
  27125=>"111111111",
  27126=>"111111110",
  27127=>"111001100",
  27128=>"011111111",
  27129=>"111011011",
  27130=>"111111111",
  27131=>"011001011",
  27132=>"011110100",
  27133=>"100110100",
  27134=>"111111110",
  27135=>"000000000",
  27136=>"000000110",
  27137=>"011110110",
  27138=>"001001000",
  27139=>"001001001",
  27140=>"110111001",
  27141=>"001001001",
  27142=>"111111010",
  27143=>"001000000",
  27144=>"111111111",
  27145=>"100000000",
  27146=>"000000001",
  27147=>"111111000",
  27148=>"110000111",
  27149=>"111111111",
  27150=>"000000100",
  27151=>"100111111",
  27152=>"100000000",
  27153=>"000100111",
  27154=>"111011000",
  27155=>"000000000",
  27156=>"111110000",
  27157=>"000000000",
  27158=>"011000000",
  27159=>"111011000",
  27160=>"110111001",
  27161=>"100011111",
  27162=>"111111111",
  27163=>"100110111",
  27164=>"111110100",
  27165=>"000100000",
  27166=>"000001001",
  27167=>"111000001",
  27168=>"111111111",
  27169=>"111111000",
  27170=>"100100111",
  27171=>"000001000",
  27172=>"000010111",
  27173=>"111000000",
  27174=>"000010000",
  27175=>"000010000",
  27176=>"111111110",
  27177=>"111111000",
  27178=>"000110000",
  27179=>"111111011",
  27180=>"101100111",
  27181=>"000000001",
  27182=>"001001011",
  27183=>"000000000",
  27184=>"001000000",
  27185=>"000000000",
  27186=>"011111111",
  27187=>"000000100",
  27188=>"100100111",
  27189=>"011011011",
  27190=>"110000000",
  27191=>"111111001",
  27192=>"001001111",
  27193=>"101010011",
  27194=>"100100110",
  27195=>"110111000",
  27196=>"000000000",
  27197=>"011010000",
  27198=>"111111101",
  27199=>"000100111",
  27200=>"000000000",
  27201=>"111101000",
  27202=>"000000001",
  27203=>"000100100",
  27204=>"100000000",
  27205=>"011111111",
  27206=>"001000000",
  27207=>"000000110",
  27208=>"011001000",
  27209=>"111001111",
  27210=>"000000000",
  27211=>"110111111",
  27212=>"111111111",
  27213=>"101001000",
  27214=>"000111110",
  27215=>"111100111",
  27216=>"011111100",
  27217=>"111101000",
  27218=>"000110111",
  27219=>"000011111",
  27220=>"000000001",
  27221=>"000000000",
  27222=>"111111111",
  27223=>"111001001",
  27224=>"110000000",
  27225=>"001101111",
  27226=>"111001101",
  27227=>"100000000",
  27228=>"000100000",
  27229=>"101111101",
  27230=>"000101000",
  27231=>"100000000",
  27232=>"000001101",
  27233=>"111111111",
  27234=>"100100000",
  27235=>"000000010",
  27236=>"111111111",
  27237=>"000001000",
  27238=>"000000101",
  27239=>"000100100",
  27240=>"111111000",
  27241=>"000111000",
  27242=>"011111111",
  27243=>"111110110",
  27244=>"111110100",
  27245=>"100110111",
  27246=>"100000000",
  27247=>"010110000",
  27248=>"000000001",
  27249=>"101000000",
  27250=>"011111111",
  27251=>"000000000",
  27252=>"001001000",
  27253=>"001001000",
  27254=>"111100111",
  27255=>"000000011",
  27256=>"110110011",
  27257=>"111111111",
  27258=>"111111111",
  27259=>"001111000",
  27260=>"001000000",
  27261=>"111111011",
  27262=>"000011111",
  27263=>"000001001",
  27264=>"000000000",
  27265=>"000000000",
  27266=>"000000100",
  27267=>"000010001",
  27268=>"100111111",
  27269=>"100101111",
  27270=>"111111000",
  27271=>"111100000",
  27272=>"000000000",
  27273=>"010000000",
  27274=>"010000111",
  27275=>"011011110",
  27276=>"101001000",
  27277=>"000000111",
  27278=>"000011111",
  27279=>"111111111",
  27280=>"000111111",
  27281=>"001011111",
  27282=>"111111101",
  27283=>"000111110",
  27284=>"000000000",
  27285=>"110111010",
  27286=>"111010000",
  27287=>"111000000",
  27288=>"111111111",
  27289=>"000001111",
  27290=>"100000000",
  27291=>"011111111",
  27292=>"000000000",
  27293=>"111111111",
  27294=>"000000000",
  27295=>"000111010",
  27296=>"111111111",
  27297=>"000000101",
  27298=>"111111111",
  27299=>"000111111",
  27300=>"011011010",
  27301=>"010111111",
  27302=>"000000111",
  27303=>"110110110",
  27304=>"011000000",
  27305=>"000000000",
  27306=>"000000000",
  27307=>"000000111",
  27308=>"101101101",
  27309=>"111011111",
  27310=>"110001000",
  27311=>"001100111",
  27312=>"000000000",
  27313=>"001011111",
  27314=>"010011111",
  27315=>"000100111",
  27316=>"000111111",
  27317=>"100001011",
  27318=>"111111111",
  27319=>"111111100",
  27320=>"111111011",
  27321=>"000000000",
  27322=>"111111101",
  27323=>"011011111",
  27324=>"111111111",
  27325=>"101001111",
  27326=>"000110000",
  27327=>"111111000",
  27328=>"110110000",
  27329=>"111111111",
  27330=>"111111000",
  27331=>"111111111",
  27332=>"000000001",
  27333=>"000000000",
  27334=>"000000000",
  27335=>"111101001",
  27336=>"011111111",
  27337=>"000000000",
  27338=>"000000101",
  27339=>"111111101",
  27340=>"000000000",
  27341=>"111111001",
  27342=>"111111000",
  27343=>"111111100",
  27344=>"111011000",
  27345=>"000111011",
  27346=>"111100000",
  27347=>"111000000",
  27348=>"100000001",
  27349=>"011110110",
  27350=>"000000111",
  27351=>"101110011",
  27352=>"000001001",
  27353=>"100100111",
  27354=>"110110111",
  27355=>"000000000",
  27356=>"111010111",
  27357=>"111111110",
  27358=>"111111111",
  27359=>"000111111",
  27360=>"010111111",
  27361=>"010011000",
  27362=>"111111000",
  27363=>"000000000",
  27364=>"000110000",
  27365=>"011001010",
  27366=>"000001111",
  27367=>"110111000",
  27368=>"001000100",
  27369=>"000001001",
  27370=>"100110110",
  27371=>"111011111",
  27372=>"111110000",
  27373=>"111111111",
  27374=>"000000000",
  27375=>"000000000",
  27376=>"111111111",
  27377=>"111111000",
  27378=>"000000000",
  27379=>"011101000",
  27380=>"111000000",
  27381=>"000001110",
  27382=>"110110100",
  27383=>"111111111",
  27384=>"000100000",
  27385=>"011011011",
  27386=>"010001011",
  27387=>"000011111",
  27388=>"000000001",
  27389=>"111011011",
  27390=>"111001001",
  27391=>"000000000",
  27392=>"111010000",
  27393=>"110110110",
  27394=>"000000010",
  27395=>"110111110",
  27396=>"001111111",
  27397=>"111111111",
  27398=>"111111111",
  27399=>"100110111",
  27400=>"111111111",
  27401=>"101001001",
  27402=>"100110111",
  27403=>"111111111",
  27404=>"100111111",
  27405=>"111101000",
  27406=>"110101100",
  27407=>"111111000",
  27408=>"110100110",
  27409=>"011011111",
  27410=>"000000000",
  27411=>"011000000",
  27412=>"111011001",
  27413=>"111111000",
  27414=>"111111011",
  27415=>"111011000",
  27416=>"110111111",
  27417=>"111011111",
  27418=>"000000000",
  27419=>"000000000",
  27420=>"100000001",
  27421=>"000001111",
  27422=>"110110000",
  27423=>"110011000",
  27424=>"111100100",
  27425=>"100110110",
  27426=>"111111111",
  27427=>"111111000",
  27428=>"000111111",
  27429=>"100000101",
  27430=>"111111101",
  27431=>"101000100",
  27432=>"010111111",
  27433=>"000000000",
  27434=>"001001000",
  27435=>"000001000",
  27436=>"000010111",
  27437=>"111111001",
  27438=>"000000000",
  27439=>"001000001",
  27440=>"101110110",
  27441=>"011001001",
  27442=>"111000000",
  27443=>"011000000",
  27444=>"000000000",
  27445=>"111000111",
  27446=>"111111011",
  27447=>"000000000",
  27448=>"111000000",
  27449=>"000000111",
  27450=>"000000000",
  27451=>"111111000",
  27452=>"111001001",
  27453=>"000000001",
  27454=>"000000000",
  27455=>"000010111",
  27456=>"000000000",
  27457=>"111001111",
  27458=>"111011111",
  27459=>"000100111",
  27460=>"000000101",
  27461=>"111111111",
  27462=>"000000000",
  27463=>"101001101",
  27464=>"010000111",
  27465=>"000111111",
  27466=>"000001100",
  27467=>"000011000",
  27468=>"111111100",
  27469=>"011000110",
  27470=>"000011101",
  27471=>"111011011",
  27472=>"000000000",
  27473=>"011000001",
  27474=>"100111111",
  27475=>"101001000",
  27476=>"000011000",
  27477=>"011111011",
  27478=>"000000011",
  27479=>"000001111",
  27480=>"100101111",
  27481=>"000000000",
  27482=>"000111000",
  27483=>"011011111",
  27484=>"000000000",
  27485=>"110000000",
  27486=>"110111110",
  27487=>"101111100",
  27488=>"001000000",
  27489=>"000000001",
  27490=>"000000111",
  27491=>"111110111",
  27492=>"111011111",
  27493=>"111111101",
  27494=>"111110000",
  27495=>"000000000",
  27496=>"111010001",
  27497=>"000010000",
  27498=>"000011011",
  27499=>"111001000",
  27500=>"000000000",
  27501=>"011000110",
  27502=>"000000000",
  27503=>"000100111",
  27504=>"000000000",
  27505=>"000001000",
  27506=>"111000000",
  27507=>"111111101",
  27508=>"111100000",
  27509=>"111011011",
  27510=>"111001111",
  27511=>"001011000",
  27512=>"100000000",
  27513=>"010110110",
  27514=>"110110110",
  27515=>"110111111",
  27516=>"001001000",
  27517=>"000000111",
  27518=>"100100111",
  27519=>"100111111",
  27520=>"000000000",
  27521=>"000011111",
  27522=>"100110001",
  27523=>"111111110",
  27524=>"011001101",
  27525=>"011000000",
  27526=>"111111111",
  27527=>"000110110",
  27528=>"110111111",
  27529=>"000000001",
  27530=>"000000000",
  27531=>"111111000",
  27532=>"111111111",
  27533=>"111111110",
  27534=>"101001000",
  27535=>"111111000",
  27536=>"000111111",
  27537=>"000000110",
  27538=>"111111000",
  27539=>"010000000",
  27540=>"111111111",
  27541=>"001000000",
  27542=>"000100000",
  27543=>"011001011",
  27544=>"000001111",
  27545=>"011000111",
  27546=>"111111111",
  27547=>"110010000",
  27548=>"111111011",
  27549=>"110000111",
  27550=>"000001001",
  27551=>"000111111",
  27552=>"011111001",
  27553=>"010011111",
  27554=>"111000000",
  27555=>"011000000",
  27556=>"110110000",
  27557=>"000111111",
  27558=>"000001111",
  27559=>"000011111",
  27560=>"000000000",
  27561=>"000011111",
  27562=>"100001001",
  27563=>"111111000",
  27564=>"000000000",
  27565=>"111000000",
  27566=>"111001000",
  27567=>"000111111",
  27568=>"110101111",
  27569=>"111000000",
  27570=>"000000001",
  27571=>"111001000",
  27572=>"000000001",
  27573=>"000011000",
  27574=>"000111101",
  27575=>"111110010",
  27576=>"000000011",
  27577=>"111111000",
  27578=>"000000110",
  27579=>"111000101",
  27580=>"000000111",
  27581=>"110111111",
  27582=>"000111111",
  27583=>"001001001",
  27584=>"000000111",
  27585=>"000000111",
  27586=>"000000000",
  27587=>"000000000",
  27588=>"000000000",
  27589=>"000001101",
  27590=>"110111111",
  27591=>"000000001",
  27592=>"111010111",
  27593=>"111111011",
  27594=>"011011011",
  27595=>"110111001",
  27596=>"000000000",
  27597=>"111111111",
  27598=>"000111111",
  27599=>"000011111",
  27600=>"000000000",
  27601=>"001101111",
  27602=>"000000000",
  27603=>"111111111",
  27604=>"111000000",
  27605=>"000001001",
  27606=>"111111000",
  27607=>"111011000",
  27608=>"010000100",
  27609=>"110000000",
  27610=>"011011000",
  27611=>"111111111",
  27612=>"000000000",
  27613=>"111100000",
  27614=>"011111111",
  27615=>"101000001",
  27616=>"010010111",
  27617=>"001000000",
  27618=>"111000000",
  27619=>"000000000",
  27620=>"000000011",
  27621=>"110100101",
  27622=>"111011111",
  27623=>"110111111",
  27624=>"100111111",
  27625=>"101100111",
  27626=>"000010111",
  27627=>"100100101",
  27628=>"110110000",
  27629=>"011000100",
  27630=>"000000011",
  27631=>"101000000",
  27632=>"000000000",
  27633=>"111111111",
  27634=>"011000011",
  27635=>"000000111",
  27636=>"011001100",
  27637=>"001000101",
  27638=>"111111111",
  27639=>"000000110",
  27640=>"000000000",
  27641=>"110010110",
  27642=>"011111001",
  27643=>"111111000",
  27644=>"000000000",
  27645=>"000000000",
  27646=>"011000000",
  27647=>"110111010",
  27648=>"000001001",
  27649=>"010000111",
  27650=>"011001101",
  27651=>"111101001",
  27652=>"100110110",
  27653=>"011000111",
  27654=>"111111111",
  27655=>"000000000",
  27656=>"000000000",
  27657=>"000000000",
  27658=>"000000000",
  27659=>"010000000",
  27660=>"001111111",
  27661=>"111000000",
  27662=>"101100111",
  27663=>"100111111",
  27664=>"011001000",
  27665=>"000000011",
  27666=>"000100100",
  27667=>"111111111",
  27668=>"111111111",
  27669=>"110110111",
  27670=>"000011111",
  27671=>"000000000",
  27672=>"111111111",
  27673=>"001000100",
  27674=>"011101111",
  27675=>"000100100",
  27676=>"111000000",
  27677=>"111111111",
  27678=>"000100100",
  27679=>"111111111",
  27680=>"001000110",
  27681=>"110100000",
  27682=>"000000000",
  27683=>"000000010",
  27684=>"000000111",
  27685=>"011000000",
  27686=>"111101111",
  27687=>"111110110",
  27688=>"000111111",
  27689=>"111111111",
  27690=>"001000001",
  27691=>"000000000",
  27692=>"111111111",
  27693=>"000101101",
  27694=>"101001000",
  27695=>"100000000",
  27696=>"000001011",
  27697=>"000000000",
  27698=>"111111111",
  27699=>"101100111",
  27700=>"111111011",
  27701=>"111111111",
  27702=>"000000000",
  27703=>"000000000",
  27704=>"011000000",
  27705=>"000110110",
  27706=>"111111111",
  27707=>"000000000",
  27708=>"111111111",
  27709=>"100001000",
  27710=>"111111111",
  27711=>"110110110",
  27712=>"000000000",
  27713=>"000000010",
  27714=>"000000110",
  27715=>"000100000",
  27716=>"000000000",
  27717=>"000000100",
  27718=>"011111111",
  27719=>"111111111",
  27720=>"000001001",
  27721=>"000000000",
  27722=>"000000001",
  27723=>"111111111",
  27724=>"000000000",
  27725=>"001111111",
  27726=>"110011000",
  27727=>"000000000",
  27728=>"110111100",
  27729=>"010000010",
  27730=>"000000000",
  27731=>"011111110",
  27732=>"111111111",
  27733=>"111111000",
  27734=>"101111111",
  27735=>"000000000",
  27736=>"000000000",
  27737=>"111111011",
  27738=>"111111111",
  27739=>"111111111",
  27740=>"011000000",
  27741=>"000000000",
  27742=>"111011011",
  27743=>"111111111",
  27744=>"001000010",
  27745=>"000000001",
  27746=>"111111111",
  27747=>"000010000",
  27748=>"000100000",
  27749=>"001110110",
  27750=>"000000000",
  27751=>"110000000",
  27752=>"000000000",
  27753=>"000000000",
  27754=>"111111011",
  27755=>"011011011",
  27756=>"001001001",
  27757=>"000000000",
  27758=>"111001000",
  27759=>"000000000",
  27760=>"111111111",
  27761=>"001100000",
  27762=>"000100101",
  27763=>"000001000",
  27764=>"111111111",
  27765=>"111111100",
  27766=>"000010000",
  27767=>"000101111",
  27768=>"000000000",
  27769=>"101111111",
  27770=>"111111111",
  27771=>"111001001",
  27772=>"110100100",
  27773=>"000000000",
  27774=>"000000000",
  27775=>"000000000",
  27776=>"111111111",
  27777=>"111111001",
  27778=>"100001001",
  27779=>"110111111",
  27780=>"111111111",
  27781=>"111111111",
  27782=>"111111111",
  27783=>"000000000",
  27784=>"111011000",
  27785=>"111000000",
  27786=>"111111111",
  27787=>"000000000",
  27788=>"000000000",
  27789=>"111111111",
  27790=>"001010111",
  27791=>"000000011",
  27792=>"100000000",
  27793=>"111111111",
  27794=>"101001101",
  27795=>"100111111",
  27796=>"000000000",
  27797=>"000000000",
  27798=>"111111110",
  27799=>"111011111",
  27800=>"001001001",
  27801=>"000000000",
  27802=>"111111111",
  27803=>"000000000",
  27804=>"101101000",
  27805=>"000000101",
  27806=>"101111111",
  27807=>"000000001",
  27808=>"000000000",
  27809=>"111111111",
  27810=>"000110110",
  27811=>"000000011",
  27812=>"000000000",
  27813=>"011111001",
  27814=>"000001001",
  27815=>"001111111",
  27816=>"001000001",
  27817=>"111111110",
  27818=>"000000000",
  27819=>"000000000",
  27820=>"111111000",
  27821=>"100100100",
  27822=>"100100111",
  27823=>"111111101",
  27824=>"111111111",
  27825=>"000111000",
  27826=>"010011010",
  27827=>"000000000",
  27828=>"000000111",
  27829=>"000111111",
  27830=>"100111111",
  27831=>"000000000",
  27832=>"000000110",
  27833=>"111111111",
  27834=>"000000000",
  27835=>"000001111",
  27836=>"000001001",
  27837=>"000001000",
  27838=>"111111111",
  27839=>"001110110",
  27840=>"000000000",
  27841=>"000100100",
  27842=>"000000000",
  27843=>"000000000",
  27844=>"000000000",
  27845=>"011000000",
  27846=>"001101000",
  27847=>"100100101",
  27848=>"111000000",
  27849=>"000111111",
  27850=>"111111111",
  27851=>"110000000",
  27852=>"011111111",
  27853=>"000000000",
  27854=>"011111111",
  27855=>"000000001",
  27856=>"111111111",
  27857=>"110111000",
  27858=>"111111111",
  27859=>"000001111",
  27860=>"000000000",
  27861=>"000000111",
  27862=>"000111111",
  27863=>"010000000",
  27864=>"111111001",
  27865=>"000000000",
  27866=>"011011111",
  27867=>"000000000",
  27868=>"101001001",
  27869=>"111111111",
  27870=>"000000000",
  27871=>"001101101",
  27872=>"000000010",
  27873=>"111011001",
  27874=>"000000010",
  27875=>"001101000",
  27876=>"001111111",
  27877=>"111111111",
  27878=>"000000000",
  27879=>"000000000",
  27880=>"000000000",
  27881=>"111111000",
  27882=>"111111111",
  27883=>"111000101",
  27884=>"111111111",
  27885=>"000000000",
  27886=>"000000111",
  27887=>"110010111",
  27888=>"111111111",
  27889=>"111111111",
  27890=>"111111000",
  27891=>"000100000",
  27892=>"111111111",
  27893=>"100110111",
  27894=>"001000000",
  27895=>"111111111",
  27896=>"111111111",
  27897=>"000000000",
  27898=>"111001001",
  27899=>"000000000",
  27900=>"110100110",
  27901=>"100100111",
  27902=>"000000000",
  27903=>"000000000",
  27904=>"000000000",
  27905=>"101100111",
  27906=>"000001011",
  27907=>"111111111",
  27908=>"000001111",
  27909=>"000100001",
  27910=>"111101111",
  27911=>"111111111",
  27912=>"000000111",
  27913=>"011111111",
  27914=>"111111111",
  27915=>"111111111",
  27916=>"010010000",
  27917=>"011011010",
  27918=>"000000000",
  27919=>"111111110",
  27920=>"111011111",
  27921=>"111111111",
  27922=>"000000011",
  27923=>"111011110",
  27924=>"001000000",
  27925=>"111110110",
  27926=>"001001001",
  27927=>"111111111",
  27928=>"111110111",
  27929=>"000000000",
  27930=>"100101111",
  27931=>"010010111",
  27932=>"111111100",
  27933=>"010000000",
  27934=>"000010000",
  27935=>"000000000",
  27936=>"000000110",
  27937=>"000000000",
  27938=>"111100111",
  27939=>"111111111",
  27940=>"111010001",
  27941=>"000100111",
  27942=>"110110110",
  27943=>"000000000",
  27944=>"111111111",
  27945=>"111110000",
  27946=>"000000100",
  27947=>"100000000",
  27948=>"001011111",
  27949=>"000000000",
  27950=>"111111111",
  27951=>"111111111",
  27952=>"111111100",
  27953=>"111111111",
  27954=>"000000000",
  27955=>"010111000",
  27956=>"011010010",
  27957=>"110111000",
  27958=>"111111111",
  27959=>"000000110",
  27960=>"100111111",
  27961=>"000000000",
  27962=>"000000000",
  27963=>"000011111",
  27964=>"000000000",
  27965=>"111111111",
  27966=>"000000000",
  27967=>"000000000",
  27968=>"000000000",
  27969=>"111111111",
  27970=>"111111111",
  27971=>"111111000",
  27972=>"111100000",
  27973=>"011101101",
  27974=>"000000000",
  27975=>"111111111",
  27976=>"000000111",
  27977=>"000000110",
  27978=>"111000100",
  27979=>"111001111",
  27980=>"001100111",
  27981=>"000111011",
  27982=>"111111111",
  27983=>"000000100",
  27984=>"011011011",
  27985=>"111000001",
  27986=>"011111111",
  27987=>"000000110",
  27988=>"001010000",
  27989=>"111111001",
  27990=>"001001001",
  27991=>"111111111",
  27992=>"111111011",
  27993=>"111111111",
  27994=>"000111000",
  27995=>"011111111",
  27996=>"110111100",
  27997=>"000100100",
  27998=>"011000111",
  27999=>"100000001",
  28000=>"000000000",
  28001=>"000111011",
  28002=>"111111001",
  28003=>"110100000",
  28004=>"000000101",
  28005=>"111111111",
  28006=>"000111111",
  28007=>"000000110",
  28008=>"110100111",
  28009=>"011011111",
  28010=>"001000000",
  28011=>"100100100",
  28012=>"111111001",
  28013=>"111000100",
  28014=>"110111111",
  28015=>"000000000",
  28016=>"000000001",
  28017=>"000000011",
  28018=>"000100111",
  28019=>"010111000",
  28020=>"111111111",
  28021=>"001101110",
  28022=>"000000011",
  28023=>"111100000",
  28024=>"111111111",
  28025=>"100100000",
  28026=>"000000000",
  28027=>"000000111",
  28028=>"111110111",
  28029=>"000000000",
  28030=>"111111111",
  28031=>"111111111",
  28032=>"000100101",
  28033=>"111000000",
  28034=>"000011111",
  28035=>"011000100",
  28036=>"111111111",
  28037=>"010000111",
  28038=>"000000000",
  28039=>"011011111",
  28040=>"001000001",
  28041=>"100000100",
  28042=>"111001001",
  28043=>"111111111",
  28044=>"110110111",
  28045=>"000100110",
  28046=>"110110110",
  28047=>"000110111",
  28048=>"000000000",
  28049=>"111111111",
  28050=>"111111111",
  28051=>"000000001",
  28052=>"111000000",
  28053=>"000000001",
  28054=>"100000000",
  28055=>"100100100",
  28056=>"000001001",
  28057=>"111111101",
  28058=>"111111111",
  28059=>"001000000",
  28060=>"000000001",
  28061=>"000000100",
  28062=>"000000000",
  28063=>"111111111",
  28064=>"000000000",
  28065=>"011000110",
  28066=>"000100000",
  28067=>"100000000",
  28068=>"110110011",
  28069=>"000000000",
  28070=>"000000000",
  28071=>"011110100",
  28072=>"000000000",
  28073=>"000010010",
  28074=>"001000000",
  28075=>"000000000",
  28076=>"000000000",
  28077=>"000000000",
  28078=>"000111111",
  28079=>"111111111",
  28080=>"000100100",
  28081=>"011011000",
  28082=>"111000010",
  28083=>"000000011",
  28084=>"100110110",
  28085=>"111111111",
  28086=>"000000000",
  28087=>"111000100",
  28088=>"011001001",
  28089=>"000000111",
  28090=>"000110111",
  28091=>"100000101",
  28092=>"000000000",
  28093=>"110000000",
  28094=>"001111111",
  28095=>"110100111",
  28096=>"111110011",
  28097=>"000000000",
  28098=>"000000000",
  28099=>"111111111",
  28100=>"111101111",
  28101=>"001001000",
  28102=>"111111111",
  28103=>"000111111",
  28104=>"000000000",
  28105=>"100110111",
  28106=>"101001111",
  28107=>"111111111",
  28108=>"111111011",
  28109=>"000000000",
  28110=>"000000001",
  28111=>"001111111",
  28112=>"000000100",
  28113=>"111111111",
  28114=>"100000000",
  28115=>"111110010",
  28116=>"000111111",
  28117=>"000000100",
  28118=>"111111101",
  28119=>"000001000",
  28120=>"101111101",
  28121=>"011111111",
  28122=>"111111110",
  28123=>"101111111",
  28124=>"000111111",
  28125=>"100100000",
  28126=>"110111111",
  28127=>"111111111",
  28128=>"000000000",
  28129=>"111111011",
  28130=>"011011111",
  28131=>"000000000",
  28132=>"000011111",
  28133=>"000000111",
  28134=>"110111111",
  28135=>"011011111",
  28136=>"111101111",
  28137=>"111111111",
  28138=>"111111100",
  28139=>"000000000",
  28140=>"000000000",
  28141=>"111111111",
  28142=>"100110110",
  28143=>"000000000",
  28144=>"000000000",
  28145=>"111000000",
  28146=>"111111111",
  28147=>"111111110",
  28148=>"111011011",
  28149=>"000000000",
  28150=>"111100100",
  28151=>"100000000",
  28152=>"111111110",
  28153=>"000000000",
  28154=>"000000101",
  28155=>"111111001",
  28156=>"000000000",
  28157=>"111000001",
  28158=>"101111111",
  28159=>"111111111",
  28160=>"110110111",
  28161=>"110111111",
  28162=>"111000111",
  28163=>"111111000",
  28164=>"111111110",
  28165=>"000000000",
  28166=>"000000000",
  28167=>"111111111",
  28168=>"010000011",
  28169=>"000000000",
  28170=>"111111111",
  28171=>"000000000",
  28172=>"100100100",
  28173=>"001111111",
  28174=>"000111001",
  28175=>"000111111",
  28176=>"111100001",
  28177=>"110110110",
  28178=>"111111111",
  28179=>"000000100",
  28180=>"001111101",
  28181=>"001001100",
  28182=>"111111000",
  28183=>"010000000",
  28184=>"000000001",
  28185=>"000000111",
  28186=>"000000000",
  28187=>"100000000",
  28188=>"111111010",
  28189=>"001111110",
  28190=>"011010110",
  28191=>"010110100",
  28192=>"001001000",
  28193=>"011111001",
  28194=>"111110000",
  28195=>"001000000",
  28196=>"110110000",
  28197=>"000000111",
  28198=>"111000000",
  28199=>"011111000",
  28200=>"100010000",
  28201=>"111111111",
  28202=>"111111111",
  28203=>"111111011",
  28204=>"000000001",
  28205=>"000000000",
  28206=>"000000100",
  28207=>"000000110",
  28208=>"100111011",
  28209=>"000000000",
  28210=>"111111000",
  28211=>"111111011",
  28212=>"000010110",
  28213=>"101111111",
  28214=>"110110010",
  28215=>"000011111",
  28216=>"000111011",
  28217=>"111111000",
  28218=>"000111111",
  28219=>"111110000",
  28220=>"000001100",
  28221=>"111111111",
  28222=>"111110010",
  28223=>"110111111",
  28224=>"111111000",
  28225=>"111011001",
  28226=>"000011111",
  28227=>"001101001",
  28228=>"110111000",
  28229=>"000000100",
  28230=>"111011011",
  28231=>"111111111",
  28232=>"000000100",
  28233=>"001000111",
  28234=>"111111000",
  28235=>"100111010",
  28236=>"011111011",
  28237=>"111111001",
  28238=>"000000000",
  28239=>"111111111",
  28240=>"111000000",
  28241=>"111111110",
  28242=>"000000001",
  28243=>"000010110",
  28244=>"000000000",
  28245=>"100100000",
  28246=>"110011001",
  28247=>"000000000",
  28248=>"110111111",
  28249=>"101000111",
  28250=>"111111111",
  28251=>"111101000",
  28252=>"111110111",
  28253=>"101101111",
  28254=>"000000000",
  28255=>"000000001",
  28256=>"111111110",
  28257=>"000000000",
  28258=>"010111111",
  28259=>"000001000",
  28260=>"111111111",
  28261=>"101100000",
  28262=>"111110100",
  28263=>"000010000",
  28264=>"111111111",
  28265=>"100000000",
  28266=>"111111111",
  28267=>"111100000",
  28268=>"110111111",
  28269=>"111111011",
  28270=>"111111111",
  28271=>"011110100",
  28272=>"110110000",
  28273=>"000000000",
  28274=>"010011011",
  28275=>"000000011",
  28276=>"000000000",
  28277=>"000010110",
  28278=>"110110110",
  28279=>"000000001",
  28280=>"000000111",
  28281=>"000011011",
  28282=>"111100100",
  28283=>"111110110",
  28284=>"000000100",
  28285=>"110110100",
  28286=>"000000100",
  28287=>"110111000",
  28288=>"000000101",
  28289=>"000000000",
  28290=>"111111000",
  28291=>"000011111",
  28292=>"111100100",
  28293=>"111100001",
  28294=>"100000000",
  28295=>"001000000",
  28296=>"111111111",
  28297=>"100100000",
  28298=>"000000011",
  28299=>"111101101",
  28300=>"000000000",
  28301=>"000000001",
  28302=>"011001000",
  28303=>"100000000",
  28304=>"000000000",
  28305=>"000000000",
  28306=>"110110110",
  28307=>"001001111",
  28308=>"000000001",
  28309=>"100100111",
  28310=>"000000111",
  28311=>"111001111",
  28312=>"000000000",
  28313=>"111111111",
  28314=>"111111111",
  28315=>"110110110",
  28316=>"000000011",
  28317=>"110110000",
  28318=>"111111111",
  28319=>"110000001",
  28320=>"111111111",
  28321=>"000000111",
  28322=>"110111111",
  28323=>"100111110",
  28324=>"101000000",
  28325=>"000000111",
  28326=>"011011111",
  28327=>"000100101",
  28328=>"001111000",
  28329=>"000000000",
  28330=>"000000000",
  28331=>"111111111",
  28332=>"111111111",
  28333=>"110111001",
  28334=>"000001111",
  28335=>"111110000",
  28336=>"011000100",
  28337=>"000000101",
  28338=>"110110110",
  28339=>"000000000",
  28340=>"000100111",
  28341=>"000000111",
  28342=>"000000111",
  28343=>"111111110",
  28344=>"111111111",
  28345=>"000000000",
  28346=>"111001000",
  28347=>"001100001",
  28348=>"000000000",
  28349=>"001001111",
  28350=>"000000100",
  28351=>"000000000",
  28352=>"000000000",
  28353=>"000001111",
  28354=>"110110111",
  28355=>"011000000",
  28356=>"000000111",
  28357=>"111000000",
  28358=>"000111111",
  28359=>"100110111",
  28360=>"011101111",
  28361=>"000000000",
  28362=>"000000000",
  28363=>"111111000",
  28364=>"110010011",
  28365=>"000000010",
  28366=>"110110100",
  28367=>"101000010",
  28368=>"101111111",
  28369=>"000000100",
  28370=>"000000110",
  28371=>"001000000",
  28372=>"100100111",
  28373=>"111111110",
  28374=>"111101111",
  28375=>"101111111",
  28376=>"000110000",
  28377=>"011111110",
  28378=>"000111111",
  28379=>"000111110",
  28380=>"000101111",
  28381=>"111000100",
  28382=>"000000110",
  28383=>"101101111",
  28384=>"010000000",
  28385=>"000011011",
  28386=>"001000000",
  28387=>"000000000",
  28388=>"111011001",
  28389=>"000100110",
  28390=>"001011001",
  28391=>"000000001",
  28392=>"110110000",
  28393=>"011100100",
  28394=>"111001000",
  28395=>"111111011",
  28396=>"100000000",
  28397=>"111111001",
  28398=>"001001000",
  28399=>"010000000",
  28400=>"000110000",
  28401=>"111111101",
  28402=>"111111000",
  28403=>"110110110",
  28404=>"000000111",
  28405=>"111111111",
  28406=>"001000001",
  28407=>"111110111",
  28408=>"000000000",
  28409=>"011111011",
  28410=>"101100000",
  28411=>"001011111",
  28412=>"000000101",
  28413=>"000011001",
  28414=>"011111000",
  28415=>"111111111",
  28416=>"000000000",
  28417=>"001001001",
  28418=>"111010000",
  28419=>"001000000",
  28420=>"011101100",
  28421=>"100111111",
  28422=>"111111001",
  28423=>"000111111",
  28424=>"111010000",
  28425=>"011011011",
  28426=>"100111111",
  28427=>"010100000",
  28428=>"100100110",
  28429=>"000111111",
  28430=>"000111110",
  28431=>"111111000",
  28432=>"101111001",
  28433=>"000000111",
  28434=>"111111100",
  28435=>"111111010",
  28436=>"001011001",
  28437=>"010010000",
  28438=>"001001011",
  28439=>"001001001",
  28440=>"000000000",
  28441=>"001111110",
  28442=>"010111100",
  28443=>"111111111",
  28444=>"100111110",
  28445=>"000000000",
  28446=>"001000100",
  28447=>"000000111",
  28448=>"111111010",
  28449=>"000110000",
  28450=>"000111111",
  28451=>"110010000",
  28452=>"000110110",
  28453=>"000000000",
  28454=>"000000000",
  28455=>"111111000",
  28456=>"000000000",
  28457=>"010111000",
  28458=>"111010111",
  28459=>"000000100",
  28460=>"100000101",
  28461=>"100000001",
  28462=>"000111000",
  28463=>"000000000",
  28464=>"000100000",
  28465=>"111111111",
  28466=>"001111111",
  28467=>"000000100",
  28468=>"100100000",
  28469=>"000000000",
  28470=>"111111101",
  28471=>"000000000",
  28472=>"000000000",
  28473=>"001101111",
  28474=>"100000000",
  28475=>"101111111",
  28476=>"110110000",
  28477=>"100100000",
  28478=>"111111110",
  28479=>"000000001",
  28480=>"000000000",
  28481=>"000001111",
  28482=>"101100111",
  28483=>"001001000",
  28484=>"110110000",
  28485=>"111101100",
  28486=>"001100111",
  28487=>"000000000",
  28488=>"111001101",
  28489=>"000000001",
  28490=>"011000111",
  28491=>"000110100",
  28492=>"000110110",
  28493=>"100111111",
  28494=>"111111000",
  28495=>"011000001",
  28496=>"101100100",
  28497=>"101101001",
  28498=>"000110000",
  28499=>"011111111",
  28500=>"000000010",
  28501=>"011011001",
  28502=>"000000101",
  28503=>"111111110",
  28504=>"111111111",
  28505=>"000000110",
  28506=>"000000000",
  28507=>"001001011",
  28508=>"000100111",
  28509=>"000000111",
  28510=>"011001000",
  28511=>"001001111",
  28512=>"111111000",
  28513=>"111111110",
  28514=>"110011011",
  28515=>"101001001",
  28516=>"110100100",
  28517=>"000000000",
  28518=>"111111101",
  28519=>"001111011",
  28520=>"001001001",
  28521=>"111111100",
  28522=>"111111011",
  28523=>"000010000",
  28524=>"110111000",
  28525=>"100010111",
  28526=>"000011111",
  28527=>"000111111",
  28528=>"011011111",
  28529=>"000000000",
  28530=>"110111111",
  28531=>"000100111",
  28532=>"000100110",
  28533=>"000000100",
  28534=>"111111011",
  28535=>"001101101",
  28536=>"000000101",
  28537=>"111111111",
  28538=>"111111000",
  28539=>"100101110",
  28540=>"110111111",
  28541=>"110111000",
  28542=>"000010111",
  28543=>"000000100",
  28544=>"000000100",
  28545=>"111111001",
  28546=>"000001111",
  28547=>"111111101",
  28548=>"000000000",
  28549=>"111111001",
  28550=>"011111011",
  28551=>"111000010",
  28552=>"111111111",
  28553=>"001111111",
  28554=>"000000000",
  28555=>"001001000",
  28556=>"100111111",
  28557=>"111111111",
  28558=>"001000001",
  28559=>"001111111",
  28560=>"000000000",
  28561=>"000000000",
  28562=>"110111111",
  28563=>"011001111",
  28564=>"000001110",
  28565=>"010011000",
  28566=>"110011010",
  28567=>"010111000",
  28568=>"000010111",
  28569=>"000000001",
  28570=>"111111111",
  28571=>"111111011",
  28572=>"100110110",
  28573=>"011001000",
  28574=>"011111011",
  28575=>"000000000",
  28576=>"111111111",
  28577=>"000000000",
  28578=>"010110111",
  28579=>"111111101",
  28580=>"000000000",
  28581=>"111001111",
  28582=>"011001011",
  28583=>"000000000",
  28584=>"111100000",
  28585=>"001011111",
  28586=>"000000000",
  28587=>"100100110",
  28588=>"000000000",
  28589=>"100111111",
  28590=>"111111000",
  28591=>"000000011",
  28592=>"000000111",
  28593=>"000000110",
  28594=>"111111111",
  28595=>"100100000",
  28596=>"000000000",
  28597=>"110110010",
  28598=>"000000000",
  28599=>"000010000",
  28600=>"111000001",
  28601=>"111111000",
  28602=>"000000000",
  28603=>"000000101",
  28604=>"100000000",
  28605=>"111000111",
  28606=>"000000000",
  28607=>"001000000",
  28608=>"110010000",
  28609=>"111111111",
  28610=>"000000000",
  28611=>"111011000",
  28612=>"000000011",
  28613=>"000111111",
  28614=>"010110110",
  28615=>"000100111",
  28616=>"101000000",
  28617=>"101101100",
  28618=>"000000000",
  28619=>"111110000",
  28620=>"111011000",
  28621=>"100110000",
  28622=>"111111111",
  28623=>"000000000",
  28624=>"000000110",
  28625=>"110111111",
  28626=>"000000000",
  28627=>"111100100",
  28628=>"111111000",
  28629=>"001000000",
  28630=>"110000000",
  28631=>"000011000",
  28632=>"000000111",
  28633=>"100000110",
  28634=>"000100111",
  28635=>"000000000",
  28636=>"000000111",
  28637=>"000000000",
  28638=>"011100000",
  28639=>"001001001",
  28640=>"000000100",
  28641=>"011011111",
  28642=>"001010000",
  28643=>"000000001",
  28644=>"000000100",
  28645=>"000000000",
  28646=>"111110110",
  28647=>"111000000",
  28648=>"010000000",
  28649=>"000000000",
  28650=>"010110010",
  28651=>"111011011",
  28652=>"000110111",
  28653=>"100110010",
  28654=>"000001111",
  28655=>"000000010",
  28656=>"001000100",
  28657=>"000000000",
  28658=>"000110000",
  28659=>"010110110",
  28660=>"000000000",
  28661=>"000000000",
  28662=>"000000000",
  28663=>"000000100",
  28664=>"010010000",
  28665=>"000000101",
  28666=>"111011000",
  28667=>"100110000",
  28668=>"011000000",
  28669=>"100100110",
  28670=>"000110111",
  28671=>"000100111",
  28672=>"111111111",
  28673=>"001111001",
  28674=>"001000000",
  28675=>"111111110",
  28676=>"111011111",
  28677=>"011001000",
  28678=>"000000000",
  28679=>"111101111",
  28680=>"111111111",
  28681=>"011011011",
  28682=>"111111110",
  28683=>"100000000",
  28684=>"000000000",
  28685=>"000000000",
  28686=>"000000000",
  28687=>"111111111",
  28688=>"110000000",
  28689=>"111011000",
  28690=>"000000000",
  28691=>"111110110",
  28692=>"011001000",
  28693=>"010000000",
  28694=>"100000111",
  28695=>"011001000",
  28696=>"111111001",
  28697=>"001001000",
  28698=>"111111000",
  28699=>"000000000",
  28700=>"111111000",
  28701=>"111111111",
  28702=>"000000010",
  28703=>"111111110",
  28704=>"000111111",
  28705=>"000000000",
  28706=>"000000000",
  28707=>"111111110",
  28708=>"111110001",
  28709=>"111111100",
  28710=>"000000000",
  28711=>"111111111",
  28712=>"111111111",
  28713=>"011011000",
  28714=>"111111111",
  28715=>"111011110",
  28716=>"101000000",
  28717=>"001000000",
  28718=>"000111110",
  28719=>"000000000",
  28720=>"000000100",
  28721=>"111111111",
  28722=>"101101000",
  28723=>"111111111",
  28724=>"111111111",
  28725=>"100100111",
  28726=>"000000000",
  28727=>"011011001",
  28728=>"011011111",
  28729=>"111111000",
  28730=>"101001000",
  28731=>"000000000",
  28732=>"001000111",
  28733=>"111000000",
  28734=>"111111111",
  28735=>"000000000",
  28736=>"100000000",
  28737=>"111001000",
  28738=>"110110100",
  28739=>"100111111",
  28740=>"111111111",
  28741=>"000000000",
  28742=>"000000000",
  28743=>"000100111",
  28744=>"110110000",
  28745=>"000000000",
  28746=>"001000000",
  28747=>"001000000",
  28748=>"111111111",
  28749=>"100111000",
  28750=>"011111111",
  28751=>"101111111",
  28752=>"001000000",
  28753=>"111111001",
  28754=>"000000001",
  28755=>"110111111",
  28756=>"000000000",
  28757=>"000111111",
  28758=>"100100100",
  28759=>"000000000",
  28760=>"100110000",
  28761=>"000000100",
  28762=>"011011000",
  28763=>"010010110",
  28764=>"111111000",
  28765=>"000000000",
  28766=>"100111111",
  28767=>"010110100",
  28768=>"001000000",
  28769=>"110100100",
  28770=>"000000000",
  28771=>"001001111",
  28772=>"000100000",
  28773=>"111111011",
  28774=>"111111000",
  28775=>"000100000",
  28776=>"000100100",
  28777=>"111111111",
  28778=>"100010011",
  28779=>"000000000",
  28780=>"010111111",
  28781=>"000010111",
  28782=>"000000011",
  28783=>"100110111",
  28784=>"001001000",
  28785=>"000000000",
  28786=>"000000111",
  28787=>"000000000",
  28788=>"100000000",
  28789=>"000000110",
  28790=>"111111000",
  28791=>"100111100",
  28792=>"000000000",
  28793=>"100000000",
  28794=>"000000000",
  28795=>"000000000",
  28796=>"000000000",
  28797=>"110000000",
  28798=>"000000000",
  28799=>"111111000",
  28800=>"111111111",
  28801=>"111111111",
  28802=>"000010111",
  28803=>"111111111",
  28804=>"100000000",
  28805=>"010000111",
  28806=>"000000100",
  28807=>"110000000",
  28808=>"111111111",
  28809=>"011000000",
  28810=>"000111111",
  28811=>"111111110",
  28812=>"111111111",
  28813=>"000000000",
  28814=>"001111000",
  28815=>"000100110",
  28816=>"000100000",
  28817=>"000000110",
  28818=>"011001000",
  28819=>"101001001",
  28820=>"000000111",
  28821=>"000000000",
  28822=>"111111111",
  28823=>"000000000",
  28824=>"000000000",
  28825=>"000000000",
  28826=>"111111111",
  28827=>"111111111",
  28828=>"111111111",
  28829=>"000000000",
  28830=>"000000000",
  28831=>"111111111",
  28832=>"000000010",
  28833=>"000110110",
  28834=>"111111000",
  28835=>"000100100",
  28836=>"000000000",
  28837=>"000000000",
  28838=>"111111111",
  28839=>"001000010",
  28840=>"111111111",
  28841=>"000011111",
  28842=>"000000000",
  28843=>"000000000",
  28844=>"011111111",
  28845=>"100100000",
  28846=>"000000100",
  28847=>"010111111",
  28848=>"111100000",
  28849=>"000000000",
  28850=>"111111011",
  28851=>"111111111",
  28852=>"000000000",
  28853=>"000000100",
  28854=>"011000100",
  28855=>"001000000",
  28856=>"111111111",
  28857=>"111001000",
  28858=>"000000000",
  28859=>"111111111",
  28860=>"000000000",
  28861=>"111111011",
  28862=>"000000000",
  28863=>"111111010",
  28864=>"000110110",
  28865=>"001001000",
  28866=>"111011000",
  28867=>"000000111",
  28868=>"100100000",
  28869=>"111111111",
  28870=>"101111011",
  28871=>"000000000",
  28872=>"111111000",
  28873=>"100000000",
  28874=>"101111111",
  28875=>"111111011",
  28876=>"111111111",
  28877=>"001001000",
  28878=>"111111111",
  28879=>"000110111",
  28880=>"000110000",
  28881=>"010000000",
  28882=>"110111111",
  28883=>"000000000",
  28884=>"000000000",
  28885=>"111111011",
  28886=>"000000000",
  28887=>"110111111",
  28888=>"000000100",
  28889=>"111000000",
  28890=>"111111000",
  28891=>"011111111",
  28892=>"110111110",
  28893=>"110110100",
  28894=>"000000000",
  28895=>"001000001",
  28896=>"111111111",
  28897=>"111111111",
  28898=>"010111100",
  28899=>"111111111",
  28900=>"111111111",
  28901=>"100100110",
  28902=>"000001111",
  28903=>"111110010",
  28904=>"000000000",
  28905=>"100100100",
  28906=>"111000100",
  28907=>"000000111",
  28908=>"000000000",
  28909=>"111111111",
  28910=>"011011111",
  28911=>"000000001",
  28912=>"101111111",
  28913=>"100000000",
  28914=>"000000000",
  28915=>"000000001",
  28916=>"111111111",
  28917=>"000000001",
  28918=>"000001000",
  28919=>"000000100",
  28920=>"111111100",
  28921=>"111111111",
  28922=>"111100111",
  28923=>"100100100",
  28924=>"000000000",
  28925=>"000011001",
  28926=>"000000000",
  28927=>"000000000",
  28928=>"111101111",
  28929=>"001101000",
  28930=>"000111111",
  28931=>"100110010",
  28932=>"011001111",
  28933=>"111000000",
  28934=>"000000100",
  28935=>"000000000",
  28936=>"111111111",
  28937=>"111100100",
  28938=>"111101110",
  28939=>"111001011",
  28940=>"000001111",
  28941=>"111110111",
  28942=>"111111111",
  28943=>"100101111",
  28944=>"110100000",
  28945=>"111000000",
  28946=>"111100000",
  28947=>"001000010",
  28948=>"000000000",
  28949=>"000000000",
  28950=>"100100110",
  28951=>"011001111",
  28952=>"011111111",
  28953=>"000010001",
  28954=>"001101000",
  28955=>"111001000",
  28956=>"111111111",
  28957=>"111111001",
  28958=>"111111011",
  28959=>"000000000",
  28960=>"001001000",
  28961=>"011010011",
  28962=>"000000000",
  28963=>"111111111",
  28964=>"000000000",
  28965=>"000001101",
  28966=>"000011111",
  28967=>"000000000",
  28968=>"000000000",
  28969=>"111111111",
  28970=>"111000000",
  28971=>"110100000",
  28972=>"010010110",
  28973=>"110110100",
  28974=>"100100101",
  28975=>"111111111",
  28976=>"101001001",
  28977=>"011000000",
  28978=>"111001000",
  28979=>"000000000",
  28980=>"001000000",
  28981=>"111011000",
  28982=>"010110101",
  28983=>"110110100",
  28984=>"000000000",
  28985=>"110110111",
  28986=>"110111011",
  28987=>"101111111",
  28988=>"001001110",
  28989=>"000000000",
  28990=>"111111111",
  28991=>"001111111",
  28992=>"111110100",
  28993=>"111111111",
  28994=>"000010111",
  28995=>"111110110",
  28996=>"000000100",
  28997=>"011111111",
  28998=>"000000000",
  28999=>"000000000",
  29000=>"000000000",
  29001=>"001111101",
  29002=>"111111111",
  29003=>"011001011",
  29004=>"100100000",
  29005=>"000100101",
  29006=>"110111111",
  29007=>"111111001",
  29008=>"001101001",
  29009=>"000000000",
  29010=>"000000000",
  29011=>"011001111",
  29012=>"000000000",
  29013=>"011011011",
  29014=>"000000110",
  29015=>"100110001",
  29016=>"111111111",
  29017=>"000000001",
  29018=>"000000000",
  29019=>"000000000",
  29020=>"000111001",
  29021=>"000000000",
  29022=>"110111111",
  29023=>"100101000",
  29024=>"010010000",
  29025=>"111100000",
  29026=>"000001000",
  29027=>"111101111",
  29028=>"010010111",
  29029=>"101100101",
  29030=>"111111011",
  29031=>"001001011",
  29032=>"100100000",
  29033=>"000100100",
  29034=>"000000001",
  29035=>"101100000",
  29036=>"001000000",
  29037=>"000000000",
  29038=>"111111111",
  29039=>"111111110",
  29040=>"000000000",
  29041=>"001011011",
  29042=>"000000000",
  29043=>"100000110",
  29044=>"111101111",
  29045=>"000000000",
  29046=>"000000000",
  29047=>"110110111",
  29048=>"000000001",
  29049=>"001111111",
  29050=>"111111011",
  29051=>"100111111",
  29052=>"111111111",
  29053=>"001001001",
  29054=>"000000000",
  29055=>"111111111",
  29056=>"111111001",
  29057=>"101000100",
  29058=>"000000000",
  29059=>"000000000",
  29060=>"000000000",
  29061=>"000000100",
  29062=>"000000000",
  29063=>"010110111",
  29064=>"111111000",
  29065=>"111111111",
  29066=>"000000000",
  29067=>"000000000",
  29068=>"000000111",
  29069=>"110110110",
  29070=>"111100100",
  29071=>"111111111",
  29072=>"000000000",
  29073=>"111111111",
  29074=>"111111111",
  29075=>"110100000",
  29076=>"111111111",
  29077=>"000000000",
  29078=>"001000000",
  29079=>"001011110",
  29080=>"000111111",
  29081=>"111111111",
  29082=>"000000100",
  29083=>"111111111",
  29084=>"111111111",
  29085=>"111111011",
  29086=>"110100100",
  29087=>"000000001",
  29088=>"011111011",
  29089=>"001000010",
  29090=>"000100100",
  29091=>"000000000",
  29092=>"000000110",
  29093=>"110111000",
  29094=>"111110110",
  29095=>"001001111",
  29096=>"011111111",
  29097=>"000000000",
  29098=>"111111111",
  29099=>"000000000",
  29100=>"000000000",
  29101=>"000000000",
  29102=>"000000010",
  29103=>"000000000",
  29104=>"000000100",
  29105=>"000000100",
  29106=>"100100110",
  29107=>"111111111",
  29108=>"111111001",
  29109=>"000000111",
  29110=>"110110000",
  29111=>"011000111",
  29112=>"101000000",
  29113=>"111000000",
  29114=>"000000000",
  29115=>"111111111",
  29116=>"000010110",
  29117=>"000000000",
  29118=>"111010000",
  29119=>"111111100",
  29120=>"000000101",
  29121=>"101101111",
  29122=>"000000000",
  29123=>"000000100",
  29124=>"001001000",
  29125=>"111111111",
  29126=>"100100111",
  29127=>"000000010",
  29128=>"000000111",
  29129=>"000000100",
  29130=>"000000000",
  29131=>"000000000",
  29132=>"000000111",
  29133=>"111111110",
  29134=>"000001000",
  29135=>"001001001",
  29136=>"101101111",
  29137=>"111111000",
  29138=>"111111111",
  29139=>"111111011",
  29140=>"011011000",
  29141=>"000111111",
  29142=>"111111010",
  29143=>"010000000",
  29144=>"111011000",
  29145=>"111000110",
  29146=>"111001001",
  29147=>"111010011",
  29148=>"101100100",
  29149=>"110110111",
  29150=>"111111111",
  29151=>"000000110",
  29152=>"000000000",
  29153=>"111001011",
  29154=>"111111101",
  29155=>"111111000",
  29156=>"100000000",
  29157=>"111111111",
  29158=>"000011111",
  29159=>"000000000",
  29160=>"111111111",
  29161=>"001111111",
  29162=>"001011000",
  29163=>"110110110",
  29164=>"111110100",
  29165=>"010000101",
  29166=>"000000100",
  29167=>"111111111",
  29168=>"111000000",
  29169=>"110111000",
  29170=>"000000000",
  29171=>"101001000",
  29172=>"000011111",
  29173=>"000000000",
  29174=>"111011000",
  29175=>"000000000",
  29176=>"011010110",
  29177=>"001001001",
  29178=>"110111000",
  29179=>"000000000",
  29180=>"000000000",
  29181=>"111111111",
  29182=>"110111111",
  29183=>"000000000",
  29184=>"101000100",
  29185=>"111111111",
  29186=>"111111011",
  29187=>"000000000",
  29188=>"011001111",
  29189=>"111110000",
  29190=>"101101111",
  29191=>"111111111",
  29192=>"000000000",
  29193=>"000011011",
  29194=>"011011111",
  29195=>"111111111",
  29196=>"000000001",
  29197=>"000001111",
  29198=>"110110011",
  29199=>"000000000",
  29200=>"110110000",
  29201=>"000000000",
  29202=>"000011000",
  29203=>"111111111",
  29204=>"100000000",
  29205=>"000000111",
  29206=>"000000000",
  29207=>"111111111",
  29208=>"000000000",
  29209=>"101101111",
  29210=>"000000000",
  29211=>"000110000",
  29212=>"111111111",
  29213=>"000000110",
  29214=>"010111110",
  29215=>"000000111",
  29216=>"001001011",
  29217=>"000000000",
  29218=>"110111111",
  29219=>"101000100",
  29220=>"100000011",
  29221=>"111000000",
  29222=>"000000000",
  29223=>"111111111",
  29224=>"111110010",
  29225=>"101000000",
  29226=>"111101111",
  29227=>"010011111",
  29228=>"011111111",
  29229=>"000100110",
  29230=>"111111111",
  29231=>"111100110",
  29232=>"110111010",
  29233=>"100100101",
  29234=>"111101111",
  29235=>"000000000",
  29236=>"111111111",
  29237=>"000110111",
  29238=>"011011011",
  29239=>"100110111",
  29240=>"111111111",
  29241=>"111111000",
  29242=>"111111111",
  29243=>"010010000",
  29244=>"011000011",
  29245=>"001001000",
  29246=>"111110110",
  29247=>"000000000",
  29248=>"000100110",
  29249=>"000000000",
  29250=>"000010010",
  29251=>"110100110",
  29252=>"001001001",
  29253=>"111101110",
  29254=>"000000000",
  29255=>"000000000",
  29256=>"001000011",
  29257=>"000000111",
  29258=>"111101000",
  29259=>"000000000",
  29260=>"111011111",
  29261=>"000000110",
  29262=>"000001011",
  29263=>"000000000",
  29264=>"000000100",
  29265=>"000000110",
  29266=>"000111111",
  29267=>"010000000",
  29268=>"010111111",
  29269=>"110000000",
  29270=>"111101000",
  29271=>"011000001",
  29272=>"100100011",
  29273=>"111001111",
  29274=>"000010110",
  29275=>"010111011",
  29276=>"010001000",
  29277=>"000010000",
  29278=>"000000000",
  29279=>"000000000",
  29280=>"111000101",
  29281=>"000000000",
  29282=>"111000000",
  29283=>"111111101",
  29284=>"111000000",
  29285=>"000000010",
  29286=>"011000010",
  29287=>"111111111",
  29288=>"110100000",
  29289=>"111111111",
  29290=>"111000000",
  29291=>"111111111",
  29292=>"011101001",
  29293=>"000001111",
  29294=>"111111111",
  29295=>"000000000",
  29296=>"111011010",
  29297=>"000000100",
  29298=>"111111011",
  29299=>"000110110",
  29300=>"001011111",
  29301=>"111110010",
  29302=>"000000111",
  29303=>"000001011",
  29304=>"000010110",
  29305=>"111001000",
  29306=>"000000110",
  29307=>"000100111",
  29308=>"011100100",
  29309=>"000000000",
  29310=>"000000000",
  29311=>"111111111",
  29312=>"111111000",
  29313=>"000000000",
  29314=>"111111111",
  29315=>"000000001",
  29316=>"111111111",
  29317=>"101000000",
  29318=>"010000000",
  29319=>"000000000",
  29320=>"111111000",
  29321=>"000001010",
  29322=>"111001001",
  29323=>"111111111",
  29324=>"111111111",
  29325=>"111111000",
  29326=>"000000000",
  29327=>"011111111",
  29328=>"000000000",
  29329=>"000000001",
  29330=>"000000000",
  29331=>"101000001",
  29332=>"000000000",
  29333=>"000011011",
  29334=>"111111111",
  29335=>"000000000",
  29336=>"000011000",
  29337=>"111111111",
  29338=>"011111110",
  29339=>"001000000",
  29340=>"111110010",
  29341=>"000000000",
  29342=>"011011111",
  29343=>"110111000",
  29344=>"111111111",
  29345=>"000000000",
  29346=>"000000000",
  29347=>"000000000",
  29348=>"000100100",
  29349=>"001111111",
  29350=>"000000000",
  29351=>"000010011",
  29352=>"110000000",
  29353=>"000010000",
  29354=>"000000101",
  29355=>"111111110",
  29356=>"000001101",
  29357=>"010110000",
  29358=>"100100000",
  29359=>"111101000",
  29360=>"111111011",
  29361=>"111111111",
  29362=>"000000000",
  29363=>"111111111",
  29364=>"000000000",
  29365=>"100111111",
  29366=>"000000000",
  29367=>"000010000",
  29368=>"000000010",
  29369=>"000000000",
  29370=>"000000000",
  29371=>"000000100",
  29372=>"111110111",
  29373=>"000101000",
  29374=>"111110111",
  29375=>"000000110",
  29376=>"010000000",
  29377=>"011111110",
  29378=>"000011111",
  29379=>"000000000",
  29380=>"100100000",
  29381=>"011010000",
  29382=>"000000000",
  29383=>"100000000",
  29384=>"000000000",
  29385=>"111111111",
  29386=>"000000000",
  29387=>"111111111",
  29388=>"110110111",
  29389=>"000100100",
  29390=>"111111111",
  29391=>"111111100",
  29392=>"010111111",
  29393=>"100100000",
  29394=>"000010110",
  29395=>"111101111",
  29396=>"111100000",
  29397=>"011001000",
  29398=>"000000000",
  29399=>"111101111",
  29400=>"111111111",
  29401=>"111000000",
  29402=>"110111111",
  29403=>"010010000",
  29404=>"011111011",
  29405=>"110101101",
  29406=>"000000000",
  29407=>"111111000",
  29408=>"000000000",
  29409=>"001001111",
  29410=>"000000000",
  29411=>"111000100",
  29412=>"000000000",
  29413=>"111110110",
  29414=>"111111111",
  29415=>"000000000",
  29416=>"000110111",
  29417=>"000000000",
  29418=>"111111111",
  29419=>"000010110",
  29420=>"000110000",
  29421=>"000000110",
  29422=>"101000100",
  29423=>"001000000",
  29424=>"000000000",
  29425=>"110100110",
  29426=>"111111111",
  29427=>"001000000",
  29428=>"001000101",
  29429=>"001011000",
  29430=>"011111011",
  29431=>"000000000",
  29432=>"101000111",
  29433=>"011011011",
  29434=>"000000000",
  29435=>"000110010",
  29436=>"000000001",
  29437=>"110110010",
  29438=>"001001100",
  29439=>"000000000",
  29440=>"000000000",
  29441=>"000010000",
  29442=>"000000111",
  29443=>"001111000",
  29444=>"111111111",
  29445=>"011011011",
  29446=>"100000000",
  29447=>"111111111",
  29448=>"010011111",
  29449=>"000000100",
  29450=>"100000000",
  29451=>"000001111",
  29452=>"010110110",
  29453=>"000111111",
  29454=>"001000000",
  29455=>"000000101",
  29456=>"111111000",
  29457=>"001000000",
  29458=>"000111111",
  29459=>"111111101",
  29460=>"001111111",
  29461=>"110100000",
  29462=>"011011000",
  29463=>"000001000",
  29464=>"000000000",
  29465=>"111110000",
  29466=>"001001000",
  29467=>"111010000",
  29468=>"000000000",
  29469=>"011111111",
  29470=>"111111111",
  29471=>"000000000",
  29472=>"000000000",
  29473=>"111101100",
  29474=>"111111111",
  29475=>"111111000",
  29476=>"000111111",
  29477=>"001001000",
  29478=>"111110110",
  29479=>"111011111",
  29480=>"000000000",
  29481=>"000000001",
  29482=>"100000000",
  29483=>"111101000",
  29484=>"000011111",
  29485=>"110110110",
  29486=>"111000000",
  29487=>"000000000",
  29488=>"000100000",
  29489=>"000011011",
  29490=>"111111111",
  29491=>"011001000",
  29492=>"010111111",
  29493=>"000000100",
  29494=>"111111111",
  29495=>"100000000",
  29496=>"110000000",
  29497=>"000000000",
  29498=>"111111111",
  29499=>"111000100",
  29500=>"111111110",
  29501=>"000100000",
  29502=>"111111111",
  29503=>"011010011",
  29504=>"100100100",
  29505=>"000000000",
  29506=>"110010000",
  29507=>"000010111",
  29508=>"000000000",
  29509=>"100110111",
  29510=>"000110000",
  29511=>"001001011",
  29512=>"000000001",
  29513=>"000100110",
  29514=>"111000100",
  29515=>"100000000",
  29516=>"011111000",
  29517=>"111000000",
  29518=>"000000000",
  29519=>"101101101",
  29520=>"011011111",
  29521=>"100111100",
  29522=>"001100000",
  29523=>"111111011",
  29524=>"000000000",
  29525=>"010000011",
  29526=>"111111111",
  29527=>"111111011",
  29528=>"010010000",
  29529=>"011011001",
  29530=>"000000000",
  29531=>"000000000",
  29532=>"000000001",
  29533=>"101001111",
  29534=>"000000000",
  29535=>"000000000",
  29536=>"101000000",
  29537=>"000000000",
  29538=>"011111011",
  29539=>"111111111",
  29540=>"100100011",
  29541=>"011011000",
  29542=>"111000000",
  29543=>"000000110",
  29544=>"001001001",
  29545=>"000000011",
  29546=>"111111111",
  29547=>"000000001",
  29548=>"000000100",
  29549=>"000000111",
  29550=>"000000000",
  29551=>"001011001",
  29552=>"001000000",
  29553=>"111111111",
  29554=>"001000011",
  29555=>"000100100",
  29556=>"111001111",
  29557=>"011011011",
  29558=>"100000000",
  29559=>"000000000",
  29560=>"111111111",
  29561=>"000100111",
  29562=>"000010010",
  29563=>"000000000",
  29564=>"000111111",
  29565=>"111111110",
  29566=>"000110110",
  29567=>"000111111",
  29568=>"011001000",
  29569=>"000000000",
  29570=>"011111111",
  29571=>"110111110",
  29572=>"100110111",
  29573=>"000000000",
  29574=>"000011001",
  29575=>"011111111",
  29576=>"000000000",
  29577=>"001000111",
  29578=>"110100100",
  29579=>"000100000",
  29580=>"101111111",
  29581=>"000110010",
  29582=>"000000000",
  29583=>"000111111",
  29584=>"000000000",
  29585=>"010000001",
  29586=>"100000000",
  29587=>"111111111",
  29588=>"000000000",
  29589=>"000000000",
  29590=>"001001100",
  29591=>"110111000",
  29592=>"000100111",
  29593=>"000010010",
  29594=>"000000000",
  29595=>"000100110",
  29596=>"100110011",
  29597=>"111000000",
  29598=>"000000000",
  29599=>"000110110",
  29600=>"000000000",
  29601=>"001000001",
  29602=>"111110110",
  29603=>"100100000",
  29604=>"100100111",
  29605=>"110111010",
  29606=>"000000000",
  29607=>"000111111",
  29608=>"000100111",
  29609=>"000011111",
  29610=>"111101101",
  29611=>"000110000",
  29612=>"000000000",
  29613=>"000000000",
  29614=>"000000000",
  29615=>"000010010",
  29616=>"111111000",
  29617=>"111111111",
  29618=>"111101101",
  29619=>"011111111",
  29620=>"000000110",
  29621=>"000000111",
  29622=>"100011011",
  29623=>"001111100",
  29624=>"111111110",
  29625=>"110111111",
  29626=>"000000000",
  29627=>"000000000",
  29628=>"110000100",
  29629=>"000000000",
  29630=>"100000000",
  29631=>"000010000",
  29632=>"000000000",
  29633=>"110111111",
  29634=>"011111111",
  29635=>"000000000",
  29636=>"000000000",
  29637=>"000000111",
  29638=>"111111110",
  29639=>"000100000",
  29640=>"010000000",
  29641=>"000000011",
  29642=>"101000010",
  29643=>"000000100",
  29644=>"100000000",
  29645=>"011011000",
  29646=>"000000000",
  29647=>"111111000",
  29648=>"000000000",
  29649=>"000000000",
  29650=>"111111111",
  29651=>"111011011",
  29652=>"000110110",
  29653=>"001000000",
  29654=>"011011011",
  29655=>"100101111",
  29656=>"100100100",
  29657=>"111111111",
  29658=>"111111111",
  29659=>"000010011",
  29660=>"111111111",
  29661=>"111111111",
  29662=>"011000000",
  29663=>"111111111",
  29664=>"110111111",
  29665=>"000000000",
  29666=>"000111100",
  29667=>"111111011",
  29668=>"111111111",
  29669=>"000000000",
  29670=>"111100000",
  29671=>"111111110",
  29672=>"111111111",
  29673=>"111111111",
  29674=>"111000001",
  29675=>"111111001",
  29676=>"111111111",
  29677=>"100000000",
  29678=>"111010000",
  29679=>"101100000",
  29680=>"111111111",
  29681=>"000011111",
  29682=>"000001111",
  29683=>"000111111",
  29684=>"100000000",
  29685=>"000000111",
  29686=>"011001000",
  29687=>"100100110",
  29688=>"010000000",
  29689=>"001001001",
  29690=>"010011111",
  29691=>"100100000",
  29692=>"000001000",
  29693=>"100100110",
  29694=>"001001011",
  29695=>"000000111",
  29696=>"000000000",
  29697=>"100000000",
  29698=>"111000111",
  29699=>"111111111",
  29700=>"111111110",
  29701=>"000000001",
  29702=>"000111111",
  29703=>"111000111",
  29704=>"111111111",
  29705=>"111111111",
  29706=>"111111010",
  29707=>"000011011",
  29708=>"000110110",
  29709=>"111110111",
  29710=>"100100111",
  29711=>"000000000",
  29712=>"011000000",
  29713=>"010111111",
  29714=>"000111111",
  29715=>"000000011",
  29716=>"111111100",
  29717=>"111000011",
  29718=>"000000111",
  29719=>"001001000",
  29720=>"000000001",
  29721=>"000000000",
  29722=>"000000000",
  29723=>"000000000",
  29724=>"001000100",
  29725=>"111111111",
  29726=>"101100100",
  29727=>"000000001",
  29728=>"000000010",
  29729=>"001000111",
  29730=>"110111110",
  29731=>"010001000",
  29732=>"110111011",
  29733=>"111000001",
  29734=>"111111111",
  29735=>"111111000",
  29736=>"000000100",
  29737=>"000110111",
  29738=>"000000111",
  29739=>"000000011",
  29740=>"000000111",
  29741=>"110110000",
  29742=>"111111101",
  29743=>"111111111",
  29744=>"111100000",
  29745=>"011111110",
  29746=>"011111000",
  29747=>"110110000",
  29748=>"101111000",
  29749=>"111110000",
  29750=>"000000001",
  29751=>"000000000",
  29752=>"110111110",
  29753=>"000011000",
  29754=>"011111111",
  29755=>"111110101",
  29756=>"100000000",
  29757=>"000000000",
  29758=>"111111100",
  29759=>"111000000",
  29760=>"111011001",
  29761=>"110110000",
  29762=>"111110110",
  29763=>"001111100",
  29764=>"110111110",
  29765=>"111110110",
  29766=>"111111111",
  29767=>"101100101",
  29768=>"000000001",
  29769=>"000000111",
  29770=>"100000000",
  29771=>"111111111",
  29772=>"000000111",
  29773=>"000000111",
  29774=>"111110111",
  29775=>"000111110",
  29776=>"000001000",
  29777=>"000101000",
  29778=>"110111111",
  29779=>"110111111",
  29780=>"001000000",
  29781=>"001000000",
  29782=>"111111111",
  29783=>"000000000",
  29784=>"111111110",
  29785=>"111111111",
  29786=>"111100000",
  29787=>"110110110",
  29788=>"100000000",
  29789=>"111000000",
  29790=>"000000000",
  29791=>"110100000",
  29792=>"111111111",
  29793=>"110110110",
  29794=>"010111111",
  29795=>"000100100",
  29796=>"111110000",
  29797=>"011010111",
  29798=>"011000000",
  29799=>"111110000",
  29800=>"111111111",
  29801=>"110100111",
  29802=>"000000000",
  29803=>"000000000",
  29804=>"111111001",
  29805=>"000111111",
  29806=>"111111111",
  29807=>"000010000",
  29808=>"000000011",
  29809=>"000000001",
  29810=>"111100101",
  29811=>"100101011",
  29812=>"000011111",
  29813=>"000111111",
  29814=>"000000000",
  29815=>"001000111",
  29816=>"111100000",
  29817=>"111111111",
  29818=>"111000000",
  29819=>"000000001",
  29820=>"100101101",
  29821=>"000000000",
  29822=>"111001100",
  29823=>"000000000",
  29824=>"111101000",
  29825=>"111111110",
  29826=>"111101000",
  29827=>"111111000",
  29828=>"100000111",
  29829=>"000000000",
  29830=>"000000000",
  29831=>"000000011",
  29832=>"011000111",
  29833=>"100000000",
  29834=>"111111110",
  29835=>"000000111",
  29836=>"100000101",
  29837=>"000000000",
  29838=>"111111111",
  29839=>"000000111",
  29840=>"111100100",
  29841=>"001000000",
  29842=>"000111000",
  29843=>"111000000",
  29844=>"000000111",
  29845=>"111000000",
  29846=>"001000001",
  29847=>"000000000",
  29848=>"101000101",
  29849=>"111111010",
  29850=>"010111111",
  29851=>"000000000",
  29852=>"000000001",
  29853=>"101001011",
  29854=>"110111111",
  29855=>"111000111",
  29856=>"000010011",
  29857=>"000000000",
  29858=>"000001111",
  29859=>"110000000",
  29860=>"000111111",
  29861=>"000000000",
  29862=>"101000000",
  29863=>"110110100",
  29864=>"000000000",
  29865=>"000000000",
  29866=>"000000000",
  29867=>"001000000",
  29868=>"100100000",
  29869=>"001111111",
  29870=>"000000100",
  29871=>"000101101",
  29872=>"000111111",
  29873=>"100110110",
  29874=>"111111110",
  29875=>"111111000",
  29876=>"000100111",
  29877=>"111111111",
  29878=>"000000000",
  29879=>"100000001",
  29880=>"000000101",
  29881=>"000111111",
  29882=>"111000000",
  29883=>"111011001",
  29884=>"001000000",
  29885=>"111001101",
  29886=>"111111111",
  29887=>"001000000",
  29888=>"010111110",
  29889=>"000000101",
  29890=>"000000111",
  29891=>"101111001",
  29892=>"000000000",
  29893=>"000000000",
  29894=>"000000111",
  29895=>"000001111",
  29896=>"001110010",
  29897=>"111000111",
  29898=>"101100000",
  29899=>"101000000",
  29900=>"000000110",
  29901=>"000000000",
  29902=>"111110000",
  29903=>"111011001",
  29904=>"011111111",
  29905=>"100000000",
  29906=>"111000001",
  29907=>"110000000",
  29908=>"111010000",
  29909=>"000000000",
  29910=>"001000111",
  29911=>"000000000",
  29912=>"000000111",
  29913=>"111101110",
  29914=>"111111111",
  29915=>"011010011",
  29916=>"000000111",
  29917=>"001000001",
  29918=>"000000000",
  29919=>"000111111",
  29920=>"011111111",
  29921=>"000000000",
  29922=>"000010000",
  29923=>"000000000",
  29924=>"110000110",
  29925=>"111111001",
  29926=>"000110110",
  29927=>"001000000",
  29928=>"111111000",
  29929=>"111001000",
  29930=>"111111111",
  29931=>"000100100",
  29932=>"111111111",
  29933=>"000000000",
  29934=>"000100101",
  29935=>"111001000",
  29936=>"111000111",
  29937=>"110000001",
  29938=>"001011001",
  29939=>"101110111",
  29940=>"111111111",
  29941=>"111000000",
  29942=>"000000000",
  29943=>"011111110",
  29944=>"111111111",
  29945=>"011111001",
  29946=>"000000000",
  29947=>"111011111",
  29948=>"000001001",
  29949=>"011001011",
  29950=>"010000000",
  29951=>"001000000",
  29952=>"000000111",
  29953=>"110111100",
  29954=>"111001000",
  29955=>"000000000",
  29956=>"000111111",
  29957=>"000001111",
  29958=>"000000101",
  29959=>"000000101",
  29960=>"111111111",
  29961=>"111111111",
  29962=>"010000000",
  29963=>"000100110",
  29964=>"101001001",
  29965=>"111111101",
  29966=>"000000000",
  29967=>"000000000",
  29968=>"000000000",
  29969=>"000000000",
  29970=>"000000011",
  29971=>"000111111",
  29972=>"000000001",
  29973=>"010111111",
  29974=>"000000100",
  29975=>"111111111",
  29976=>"111111111",
  29977=>"111111111",
  29978=>"000000000",
  29979=>"000110111",
  29980=>"110110110",
  29981=>"111000000",
  29982=>"000000010",
  29983=>"111100111",
  29984=>"111010000",
  29985=>"111111000",
  29986=>"111111001",
  29987=>"000000000",
  29988=>"101000000",
  29989=>"111111111",
  29990=>"000000000",
  29991=>"100001001",
  29992=>"000000000",
  29993=>"010111010",
  29994=>"111111111",
  29995=>"000000001",
  29996=>"111001000",
  29997=>"100000000",
  29998=>"000000000",
  29999=>"000000000",
  30000=>"000111000",
  30001=>"000000000",
  30002=>"000000000",
  30003=>"111001000",
  30004=>"010011000",
  30005=>"111111000",
  30006=>"001001111",
  30007=>"001000000",
  30008=>"000000000",
  30009=>"001000001",
  30010=>"000000101",
  30011=>"111111111",
  30012=>"100000000",
  30013=>"000000000",
  30014=>"000100111",
  30015=>"111111111",
  30016=>"100000000",
  30017=>"000001001",
  30018=>"111111110",
  30019=>"000000000",
  30020=>"111111000",
  30021=>"000110010",
  30022=>"100010111",
  30023=>"000111100",
  30024=>"111100100",
  30025=>"111000111",
  30026=>"110111010",
  30027=>"100100000",
  30028=>"110111111",
  30029=>"000011000",
  30030=>"110001111",
  30031=>"110100000",
  30032=>"101001011",
  30033=>"001000111",
  30034=>"100111111",
  30035=>"000000000",
  30036=>"000110000",
  30037=>"001011001",
  30038=>"111111111",
  30039=>"111100100",
  30040=>"000001011",
  30041=>"000000100",
  30042=>"111111111",
  30043=>"000000001",
  30044=>"000000000",
  30045=>"110110100",
  30046=>"000001111",
  30047=>"000000000",
  30048=>"111111000",
  30049=>"111111111",
  30050=>"100100001",
  30051=>"100101111",
  30052=>"000000110",
  30053=>"000000001",
  30054=>"000100111",
  30055=>"001001011",
  30056=>"111010000",
  30057=>"111111111",
  30058=>"000000000",
  30059=>"111110111",
  30060=>"110111111",
  30061=>"101100101",
  30062=>"011111111",
  30063=>"100101111",
  30064=>"100100111",
  30065=>"000000000",
  30066=>"111111111",
  30067=>"111111001",
  30068=>"000000000",
  30069=>"001101111",
  30070=>"000000000",
  30071=>"111101110",
  30072=>"111111111",
  30073=>"001000000",
  30074=>"101100101",
  30075=>"001000000",
  30076=>"000001000",
  30077=>"111111111",
  30078=>"000110110",
  30079=>"001000101",
  30080=>"001001000",
  30081=>"111000000",
  30082=>"111111011",
  30083=>"000000000",
  30084=>"111000000",
  30085=>"000010011",
  30086=>"100000000",
  30087=>"111100100",
  30088=>"000000000",
  30089=>"111111100",
  30090=>"000000001",
  30091=>"000111111",
  30092=>"111100000",
  30093=>"000100100",
  30094=>"111111010",
  30095=>"111111010",
  30096=>"000000000",
  30097=>"000000000",
  30098=>"000100100",
  30099=>"001000111",
  30100=>"000000011",
  30101=>"010110010",
  30102=>"000000000",
  30103=>"000000100",
  30104=>"000111111",
  30105=>"110111111",
  30106=>"011101101",
  30107=>"111111010",
  30108=>"010001000",
  30109=>"010000001",
  30110=>"111001001",
  30111=>"000000000",
  30112=>"111111111",
  30113=>"111100111",
  30114=>"000000001",
  30115=>"000000000",
  30116=>"000000001",
  30117=>"111111111",
  30118=>"101001110",
  30119=>"111111101",
  30120=>"111000001",
  30121=>"000000001",
  30122=>"000011010",
  30123=>"000000000",
  30124=>"000000111",
  30125=>"110111111",
  30126=>"000000101",
  30127=>"000000000",
  30128=>"000000000",
  30129=>"111110000",
  30130=>"001000101",
  30131=>"000000001",
  30132=>"101000000",
  30133=>"010110110",
  30134=>"111111111",
  30135=>"001000000",
  30136=>"000000000",
  30137=>"000110011",
  30138=>"110100100",
  30139=>"000000111",
  30140=>"001000000",
  30141=>"000000001",
  30142=>"111111111",
  30143=>"101001001",
  30144=>"111111110",
  30145=>"111111111",
  30146=>"111111111",
  30147=>"111000000",
  30148=>"111111111",
  30149=>"001011111",
  30150=>"000000000",
  30151=>"000000101",
  30152=>"000000000",
  30153=>"111111111",
  30154=>"000000101",
  30155=>"000000000",
  30156=>"111111000",
  30157=>"000000011",
  30158=>"111111111",
  30159=>"000000110",
  30160=>"111110000",
  30161=>"110000100",
  30162=>"010000000",
  30163=>"100100000",
  30164=>"111000000",
  30165=>"111111101",
  30166=>"000000000",
  30167=>"011111010",
  30168=>"100000000",
  30169=>"111111111",
  30170=>"111111111",
  30171=>"000000111",
  30172=>"000000000",
  30173=>"000000101",
  30174=>"100000011",
  30175=>"100000000",
  30176=>"000000000",
  30177=>"110111000",
  30178=>"011011011",
  30179=>"000000000",
  30180=>"000000001",
  30181=>"010000111",
  30182=>"000000111",
  30183=>"111001000",
  30184=>"111100000",
  30185=>"000000110",
  30186=>"110000000",
  30187=>"100000101",
  30188=>"000100110",
  30189=>"000001001",
  30190=>"101000001",
  30191=>"000000001",
  30192=>"011001001",
  30193=>"000000000",
  30194=>"000110110",
  30195=>"001000000",
  30196=>"010010010",
  30197=>"011011001",
  30198=>"111000001",
  30199=>"001011111",
  30200=>"001001000",
  30201=>"000000001",
  30202=>"010111110",
  30203=>"011000001",
  30204=>"111011011",
  30205=>"000011111",
  30206=>"111111000",
  30207=>"111001101",
  30208=>"001000111",
  30209=>"000000000",
  30210=>"000000000",
  30211=>"011111111",
  30212=>"000001001",
  30213=>"111110100",
  30214=>"000000000",
  30215=>"111111111",
  30216=>"111011111",
  30217=>"000001001",
  30218=>"111010000",
  30219=>"100000001",
  30220=>"100110100",
  30221=>"110111111",
  30222=>"001001000",
  30223=>"000000000",
  30224=>"010000000",
  30225=>"000000011",
  30226=>"111111110",
  30227=>"010010000",
  30228=>"000000010",
  30229=>"000000111",
  30230=>"000000000",
  30231=>"000000111",
  30232=>"100110110",
  30233=>"000000000",
  30234=>"000100000",
  30235=>"111111000",
  30236=>"000000001",
  30237=>"101101100",
  30238=>"000000000",
  30239=>"111111111",
  30240=>"111101000",
  30241=>"000000000",
  30242=>"000001101",
  30243=>"000000000",
  30244=>"011011111",
  30245=>"000011111",
  30246=>"100000000",
  30247=>"000011011",
  30248=>"000000110",
  30249=>"000000000",
  30250=>"111111111",
  30251=>"100111110",
  30252=>"000000000",
  30253=>"111111110",
  30254=>"000000000",
  30255=>"111001000",
  30256=>"001011111",
  30257=>"000000000",
  30258=>"000100101",
  30259=>"000000100",
  30260=>"111111111",
  30261=>"101100100",
  30262=>"100100000",
  30263=>"000001111",
  30264=>"001101111",
  30265=>"000000100",
  30266=>"001000000",
  30267=>"000000111",
  30268=>"111111111",
  30269=>"100111111",
  30270=>"111101101",
  30271=>"111111111",
  30272=>"011001100",
  30273=>"111110110",
  30274=>"011001011",
  30275=>"000000000",
  30276=>"000011000",
  30277=>"111111111",
  30278=>"000000000",
  30279=>"111111010",
  30280=>"111111111",
  30281=>"011001011",
  30282=>"000000000",
  30283=>"100111111",
  30284=>"001011111",
  30285=>"111011000",
  30286=>"010000000",
  30287=>"000000001",
  30288=>"100110100",
  30289=>"111110011",
  30290=>"011001000",
  30291=>"000000110",
  30292=>"000000000",
  30293=>"000000000",
  30294=>"110111110",
  30295=>"111111111",
  30296=>"000000000",
  30297=>"111101101",
  30298=>"111101000",
  30299=>"110100000",
  30300=>"100010010",
  30301=>"000000000",
  30302=>"000011000",
  30303=>"001000000",
  30304=>"000000000",
  30305=>"110100101",
  30306=>"011100000",
  30307=>"000010110",
  30308=>"000000000",
  30309=>"111111000",
  30310=>"100000000",
  30311=>"111111111",
  30312=>"000000000",
  30313=>"111111111",
  30314=>"110010110",
  30315=>"000000000",
  30316=>"010110001",
  30317=>"011111111",
  30318=>"111111111",
  30319=>"000111100",
  30320=>"111111001",
  30321=>"111111111",
  30322=>"111111111",
  30323=>"010011111",
  30324=>"000100000",
  30325=>"000000000",
  30326=>"000000111",
  30327=>"111101100",
  30328=>"111111111",
  30329=>"001111101",
  30330=>"100100111",
  30331=>"000000001",
  30332=>"110110110",
  30333=>"111111111",
  30334=>"111111111",
  30335=>"000010000",
  30336=>"000110110",
  30337=>"011011111",
  30338=>"000000001",
  30339=>"001011100",
  30340=>"111110000",
  30341=>"001001011",
  30342=>"111111111",
  30343=>"110000000",
  30344=>"000010010",
  30345=>"010010000",
  30346=>"000000000",
  30347=>"000000000",
  30348=>"111111100",
  30349=>"000000000",
  30350=>"000001011",
  30351=>"000000000",
  30352=>"000000111",
  30353=>"000011111",
  30354=>"111110110",
  30355=>"011011010",
  30356=>"100111000",
  30357=>"110100100",
  30358=>"000000000",
  30359=>"111001111",
  30360=>"111011000",
  30361=>"011000000",
  30362=>"000100000",
  30363=>"001000000",
  30364=>"001000000",
  30365=>"100110111",
  30366=>"111111111",
  30367=>"110110110",
  30368=>"111111111",
  30369=>"010011011",
  30370=>"111111111",
  30371=>"011000011",
  30372=>"001001100",
  30373=>"000111111",
  30374=>"000000000",
  30375=>"111101111",
  30376=>"000000000",
  30377=>"011000100",
  30378=>"011001000",
  30379=>"110000011",
  30380=>"101111111",
  30381=>"001000100",
  30382=>"101101100",
  30383=>"000000000",
  30384=>"000000011",
  30385=>"000000000",
  30386=>"011000000",
  30387=>"111111111",
  30388=>"000000000",
  30389=>"000000100",
  30390=>"000000010",
  30391=>"111000010",
  30392=>"111101100",
  30393=>"000000000",
  30394=>"000000111",
  30395=>"100010010",
  30396=>"101101101",
  30397=>"000000000",
  30398=>"000000000",
  30399=>"010000000",
  30400=>"111001000",
  30401=>"100101100",
  30402=>"000000000",
  30403=>"001000000",
  30404=>"000000111",
  30405=>"000111111",
  30406=>"000000000",
  30407=>"000011001",
  30408=>"111111111",
  30409=>"111111111",
  30410=>"111010000",
  30411=>"101111111",
  30412=>"100000000",
  30413=>"000000110",
  30414=>"000000000",
  30415=>"000000110",
  30416=>"000000010",
  30417=>"000000000",
  30418=>"111111110",
  30419=>"111111000",
  30420=>"111100100",
  30421=>"110111111",
  30422=>"000000110",
  30423=>"000000000",
  30424=>"111100100",
  30425=>"000011000",
  30426=>"111010111",
  30427=>"111111001",
  30428=>"110001101",
  30429=>"000000111",
  30430=>"110111111",
  30431=>"111001000",
  30432=>"000000110",
  30433=>"011011000",
  30434=>"011111111",
  30435=>"000000111",
  30436=>"111111001",
  30437=>"000000000",
  30438=>"101000111",
  30439=>"100000111",
  30440=>"001000000",
  30441=>"000000000",
  30442=>"101111111",
  30443=>"100100100",
  30444=>"000000010",
  30445=>"110000000",
  30446=>"000000110",
  30447=>"000000000",
  30448=>"000000000",
  30449=>"000000000",
  30450=>"111111111",
  30451=>"100011111",
  30452=>"111111010",
  30453=>"100000000",
  30454=>"111111111",
  30455=>"000000000",
  30456=>"000000000",
  30457=>"000000000",
  30458=>"000000100",
  30459=>"000000000",
  30460=>"001001001",
  30461=>"001000000",
  30462=>"110000001",
  30463=>"011111111",
  30464=>"110111111",
  30465=>"111101111",
  30466=>"011011111",
  30467=>"100100110",
  30468=>"111111111",
  30469=>"000100000",
  30470=>"111101111",
  30471=>"111111111",
  30472=>"011011111",
  30473=>"010111011",
  30474=>"100100111",
  30475=>"000000000",
  30476=>"111111111",
  30477=>"110000011",
  30478=>"000000000",
  30479=>"000101111",
  30480=>"111111000",
  30481=>"110000110",
  30482=>"000000000",
  30483=>"000001111",
  30484=>"111111110",
  30485=>"000000111",
  30486=>"110100100",
  30487=>"111111000",
  30488=>"000000100",
  30489=>"001000000",
  30490=>"100000000",
  30491=>"000110100",
  30492=>"111111111",
  30493=>"111000000",
  30494=>"110010000",
  30495=>"000000000",
  30496=>"001111111",
  30497=>"000000000",
  30498=>"011101001",
  30499=>"011000000",
  30500=>"111111010",
  30501=>"110000010",
  30502=>"110001101",
  30503=>"001010011",
  30504=>"111011111",
  30505=>"111110110",
  30506=>"000000000",
  30507=>"000101111",
  30508=>"000000111",
  30509=>"000000000",
  30510=>"000000000",
  30511=>"101100000",
  30512=>"111101001",
  30513=>"000000000",
  30514=>"111110000",
  30515=>"111011111",
  30516=>"011000000",
  30517=>"111000001",
  30518=>"001000100",
  30519=>"111100100",
  30520=>"111111111",
  30521=>"111111111",
  30522=>"111111111",
  30523=>"010011011",
  30524=>"100101111",
  30525=>"100000000",
  30526=>"001000000",
  30527=>"000110111",
  30528=>"111000000",
  30529=>"000000000",
  30530=>"111001100",
  30531=>"101101101",
  30532=>"110100100",
  30533=>"000000000",
  30534=>"001101101",
  30535=>"101000000",
  30536=>"111010011",
  30537=>"000010000",
  30538=>"111111000",
  30539=>"111101111",
  30540=>"000000000",
  30541=>"001000000",
  30542=>"000000100",
  30543=>"101101001",
  30544=>"111101111",
  30545=>"001000000",
  30546=>"100000100",
  30547=>"110100100",
  30548=>"111111011",
  30549=>"011011011",
  30550=>"000000000",
  30551=>"111110110",
  30552=>"001011011",
  30553=>"000000000",
  30554=>"111011000",
  30555=>"100011000",
  30556=>"000000000",
  30557=>"110111100",
  30558=>"000111001",
  30559=>"011000000",
  30560=>"011011111",
  30561=>"111001000",
  30562=>"000000100",
  30563=>"001001011",
  30564=>"111111111",
  30565=>"111111111",
  30566=>"010000000",
  30567=>"001001000",
  30568=>"100100101",
  30569=>"011011001",
  30570=>"000000000",
  30571=>"010011010",
  30572=>"010110000",
  30573=>"100011110",
  30574=>"000000000",
  30575=>"000000011",
  30576=>"111111111",
  30577=>"010011011",
  30578=>"100110000",
  30579=>"011011011",
  30580=>"011011000",
  30581=>"100110110",
  30582=>"100111111",
  30583=>"000000000",
  30584=>"000000000",
  30585=>"000110111",
  30586=>"111111000",
  30587=>"101100101",
  30588=>"001001000",
  30589=>"111111100",
  30590=>"111111111",
  30591=>"001001000",
  30592=>"100110100",
  30593=>"011001001",
  30594=>"111001000",
  30595=>"111111111",
  30596=>"000000011",
  30597=>"011000000",
  30598=>"000000101",
  30599=>"111011000",
  30600=>"000000000",
  30601=>"000001011",
  30602=>"011111111",
  30603=>"000000000",
  30604=>"110110111",
  30605=>"110110110",
  30606=>"111111111",
  30607=>"000000000",
  30608=>"011011011",
  30609=>"110000000",
  30610=>"011011011",
  30611=>"111111111",
  30612=>"111011000",
  30613=>"010010010",
  30614=>"000111100",
  30615=>"111111000",
  30616=>"001000111",
  30617=>"000011001",
  30618=>"000000000",
  30619=>"000011011",
  30620=>"000000101",
  30621=>"000000000",
  30622=>"000000001",
  30623=>"000000000",
  30624=>"111111111",
  30625=>"111110110",
  30626=>"100001111",
  30627=>"011011001",
  30628=>"111111100",
  30629=>"000000001",
  30630=>"111111111",
  30631=>"011011001",
  30632=>"100000000",
  30633=>"111111011",
  30634=>"110111111",
  30635=>"000000100",
  30636=>"000000110",
  30637=>"110000100",
  30638=>"000000101",
  30639=>"111110011",
  30640=>"000010111",
  30641=>"111111011",
  30642=>"111011110",
  30643=>"000000000",
  30644=>"011111111",
  30645=>"000000000",
  30646=>"100111000",
  30647=>"111111111",
  30648=>"111111001",
  30649=>"000000000",
  30650=>"111011111",
  30651=>"001101001",
  30652=>"011011111",
  30653=>"000000000",
  30654=>"000110111",
  30655=>"101100100",
  30656=>"101000000",
  30657=>"111111000",
  30658=>"101001000",
  30659=>"101001000",
  30660=>"100000000",
  30661=>"101111111",
  30662=>"111011000",
  30663=>"111111110",
  30664=>"110111011",
  30665=>"100000000",
  30666=>"110010000",
  30667=>"000010000",
  30668=>"100000000",
  30669=>"100010000",
  30670=>"111000000",
  30671=>"000010000",
  30672=>"011011110",
  30673=>"111111111",
  30674=>"111111101",
  30675=>"111111111",
  30676=>"100000000",
  30677=>"101111111",
  30678=>"100110001",
  30679=>"110000010",
  30680=>"000000100",
  30681=>"010111111",
  30682=>"000010000",
  30683=>"000000000",
  30684=>"111110000",
  30685=>"111111111",
  30686=>"111100000",
  30687=>"111111111",
  30688=>"111110110",
  30689=>"011011111",
  30690=>"110111011",
  30691=>"111001101",
  30692=>"000000000",
  30693=>"111111111",
  30694=>"000001101",
  30695=>"000010010",
  30696=>"000000111",
  30697=>"000000111",
  30698=>"000000101",
  30699=>"111111111",
  30700=>"101111000",
  30701=>"100110111",
  30702=>"000000101",
  30703=>"110111111",
  30704=>"001011011",
  30705=>"000000000",
  30706=>"111111111",
  30707=>"000100101",
  30708=>"001011011",
  30709=>"010111000",
  30710=>"100000000",
  30711=>"111111101",
  30712=>"011001000",
  30713=>"100000000",
  30714=>"111111111",
  30715=>"111000011",
  30716=>"000000110",
  30717=>"111110100",
  30718=>"100100100",
  30719=>"000000000",
  30720=>"101101101",
  30721=>"011000100",
  30722=>"101000000",
  30723=>"000000010",
  30724=>"111001011",
  30725=>"111111111",
  30726=>"000000000",
  30727=>"111111111",
  30728=>"000111111",
  30729=>"001000000",
  30730=>"010100111",
  30731=>"111111011",
  30732=>"000000000",
  30733=>"000000000",
  30734=>"110111111",
  30735=>"111111011",
  30736=>"000110111",
  30737=>"110000000",
  30738=>"001111111",
  30739=>"000000000",
  30740=>"000000000",
  30741=>"111100111",
  30742=>"000001000",
  30743=>"000111111",
  30744=>"111111111",
  30745=>"111111100",
  30746=>"111100000",
  30747=>"000000111",
  30748=>"100000000",
  30749=>"000001111",
  30750=>"000110110",
  30751=>"000000001",
  30752=>"000001000",
  30753=>"000111111",
  30754=>"111111110",
  30755=>"111101111",
  30756=>"111111111",
  30757=>"111111111",
  30758=>"001000000",
  30759=>"111111110",
  30760=>"000000000",
  30761=>"111110000",
  30762=>"100100110",
  30763=>"100000111",
  30764=>"110111111",
  30765=>"000111111",
  30766=>"001000100",
  30767=>"111000000",
  30768=>"111111000",
  30769=>"000000000",
  30770=>"111111000",
  30771=>"111111111",
  30772=>"000000000",
  30773=>"110001000",
  30774=>"000000000",
  30775=>"000001001",
  30776=>"111111000",
  30777=>"000111111",
  30778=>"101000000",
  30779=>"000100111",
  30780=>"000001001",
  30781=>"000111111",
  30782=>"110001011",
  30783=>"110110111",
  30784=>"000000000",
  30785=>"000001000",
  30786=>"000001111",
  30787=>"000000000",
  30788=>"100001000",
  30789=>"000000000",
  30790=>"111010110",
  30791=>"111111111",
  30792=>"000001001",
  30793=>"000000000",
  30794=>"000111111",
  30795=>"101101111",
  30796=>"000111111",
  30797=>"100000000",
  30798=>"000100110",
  30799=>"101000000",
  30800=>"111111000",
  30801=>"000000000",
  30802=>"111111110",
  30803=>"000000110",
  30804=>"000110011",
  30805=>"000111011",
  30806=>"000000001",
  30807=>"000000000",
  30808=>"111111110",
  30809=>"111000000",
  30810=>"000011111",
  30811=>"111001011",
  30812=>"111111111",
  30813=>"111111000",
  30814=>"000000111",
  30815=>"110111111",
  30816=>"000000000",
  30817=>"000111111",
  30818=>"000000000",
  30819=>"111011111",
  30820=>"001000110",
  30821=>"111110111",
  30822=>"000001000",
  30823=>"010000000",
  30824=>"111111000",
  30825=>"110000000",
  30826=>"000000111",
  30827=>"001000001",
  30828=>"101100000",
  30829=>"111111111",
  30830=>"001000000",
  30831=>"001000000",
  30832=>"111011111",
  30833=>"011011000",
  30834=>"000000000",
  30835=>"011011111",
  30836=>"000111111",
  30837=>"000000000",
  30838=>"110111111",
  30839=>"111111000",
  30840=>"111101000",
  30841=>"000000000",
  30842=>"100100000",
  30843=>"111111111",
  30844=>"100111101",
  30845=>"001101101",
  30846=>"000000111",
  30847=>"000000000",
  30848=>"111101111",
  30849=>"111111111",
  30850=>"011111111",
  30851=>"111111111",
  30852=>"111111100",
  30853=>"111111111",
  30854=>"111001001",
  30855=>"010110011",
  30856=>"000000000",
  30857=>"001001000",
  30858=>"100000000",
  30859=>"011001001",
  30860=>"001011111",
  30861=>"001000000",
  30862=>"111111000",
  30863=>"011011000",
  30864=>"000111111",
  30865=>"000111110",
  30866=>"000000000",
  30867=>"000011111",
  30868=>"000000000",
  30869=>"100101101",
  30870=>"000000000",
  30871=>"111111111",
  30872=>"001011111",
  30873=>"000000000",
  30874=>"011011111",
  30875=>"000000011",
  30876=>"001001111",
  30877=>"100000100",
  30878=>"001111111",
  30879=>"001001111",
  30880=>"000010010",
  30881=>"000011011",
  30882=>"111110001",
  30883=>"101001000",
  30884=>"100000001",
  30885=>"111111001",
  30886=>"000111111",
  30887=>"001001001",
  30888=>"000000000",
  30889=>"011000000",
  30890=>"111111001",
  30891=>"000111111",
  30892=>"000000100",
  30893=>"100101001",
  30894=>"101010000",
  30895=>"000000111",
  30896=>"000000111",
  30897=>"111111101",
  30898=>"110111111",
  30899=>"111111111",
  30900=>"001001101",
  30901=>"111111111",
  30902=>"000000111",
  30903=>"111111010",
  30904=>"110100111",
  30905=>"111101101",
  30906=>"111001000",
  30907=>"111100000",
  30908=>"111000000",
  30909=>"001111001",
  30910=>"101000001",
  30911=>"110110111",
  30912=>"000010000",
  30913=>"110000000",
  30914=>"000001001",
  30915=>"111111111",
  30916=>"000000111",
  30917=>"000110000",
  30918=>"111101000",
  30919=>"110111000",
  30920=>"000111111",
  30921=>"111000000",
  30922=>"000101000",
  30923=>"111000000",
  30924=>"000000000",
  30925=>"000110110",
  30926=>"111111000",
  30927=>"100000000",
  30928=>"000111111",
  30929=>"111000000",
  30930=>"000111111",
  30931=>"000000000",
  30932=>"100001000",
  30933=>"100111111",
  30934=>"000000001",
  30935=>"101101000",
  30936=>"100111111",
  30937=>"011001001",
  30938=>"000000000",
  30939=>"000100110",
  30940=>"111000000",
  30941=>"001000001",
  30942=>"011011000",
  30943=>"000111111",
  30944=>"111000000",
  30945=>"000011000",
  30946=>"111111001",
  30947=>"000000111",
  30948=>"111100000",
  30949=>"000000100",
  30950=>"100000001",
  30951=>"111000000",
  30952=>"000000111",
  30953=>"111111100",
  30954=>"000000111",
  30955=>"111000000",
  30956=>"001100000",
  30957=>"011000000",
  30958=>"000001001",
  30959=>"111101111",
  30960=>"100101100",
  30961=>"001111111",
  30962=>"111011001",
  30963=>"101111111",
  30964=>"100110000",
  30965=>"011111111",
  30966=>"001111111",
  30967=>"111111111",
  30968=>"111001000",
  30969=>"000110000",
  30970=>"000000000",
  30971=>"000001011",
  30972=>"001000001",
  30973=>"111011111",
  30974=>"000111110",
  30975=>"111111111",
  30976=>"000101111",
  30977=>"001001000",
  30978=>"111111000",
  30979=>"111111110",
  30980=>"100000000",
  30981=>"100111111",
  30982=>"111101111",
  30983=>"000001100",
  30984=>"111111111",
  30985=>"000000000",
  30986=>"111000000",
  30987=>"110000100",
  30988=>"111101101",
  30989=>"000111111",
  30990=>"011111000",
  30991=>"000101000",
  30992=>"111111001",
  30993=>"111011000",
  30994=>"000000000",
  30995=>"100111111",
  30996=>"111111111",
  30997=>"111010000",
  30998=>"111111111",
  30999=>"000000000",
  31000=>"000000000",
  31001=>"111111001",
  31002=>"000000000",
  31003=>"001000111",
  31004=>"011111111",
  31005=>"011000000",
  31006=>"111111111",
  31007=>"010000000",
  31008=>"100101001",
  31009=>"011111111",
  31010=>"011110111",
  31011=>"110100111",
  31012=>"001000000",
  31013=>"111111111",
  31014=>"100111111",
  31015=>"001000000",
  31016=>"000000001",
  31017=>"000001111",
  31018=>"110111111",
  31019=>"100101101",
  31020=>"111111000",
  31021=>"001111100",
  31022=>"110111111",
  31023=>"000000000",
  31024=>"000001001",
  31025=>"111111111",
  31026=>"000111111",
  31027=>"000000000",
  31028=>"110101111",
  31029=>"100111110",
  31030=>"000000000",
  31031=>"111000101",
  31032=>"001111000",
  31033=>"111111000",
  31034=>"000110110",
  31035=>"111011000",
  31036=>"111110000",
  31037=>"001001111",
  31038=>"000000110",
  31039=>"111110001",
  31040=>"111111001",
  31041=>"111000000",
  31042=>"000001001",
  31043=>"000111111",
  31044=>"000100111",
  31045=>"100100000",
  31046=>"000000000",
  31047=>"111000001",
  31048=>"000000010",
  31049=>"111111111",
  31050=>"000010111",
  31051=>"000111001",
  31052=>"110111111",
  31053=>"001000000",
  31054=>"000001111",
  31055=>"110000000",
  31056=>"000100000",
  31057=>"100001111",
  31058=>"011011111",
  31059=>"110000000",
  31060=>"000000000",
  31061=>"011111010",
  31062=>"111001001",
  31063=>"000000111",
  31064=>"010111111",
  31065=>"111101111",
  31066=>"111100110",
  31067=>"111111111",
  31068=>"000000000",
  31069=>"111111011",
  31070=>"111110110",
  31071=>"111111001",
  31072=>"111000000",
  31073=>"000000000",
  31074=>"011111111",
  31075=>"111101000",
  31076=>"000000001",
  31077=>"000000000",
  31078=>"000000000",
  31079=>"000111111",
  31080=>"000110110",
  31081=>"110110111",
  31082=>"111000000",
  31083=>"101111001",
  31084=>"000100111",
  31085=>"111111111",
  31086=>"100100111",
  31087=>"000000110",
  31088=>"000000000",
  31089=>"000111000",
  31090=>"000000010",
  31091=>"111111111",
  31092=>"000100100",
  31093=>"000000000",
  31094=>"000110111",
  31095=>"000000000",
  31096=>"111111111",
  31097=>"111111100",
  31098=>"111111111",
  31099=>"000000000",
  31100=>"101111111",
  31101=>"111100000",
  31102=>"000000000",
  31103=>"001000101",
  31104=>"111111111",
  31105=>"001000000",
  31106=>"100100000",
  31107=>"001101111",
  31108=>"111111000",
  31109=>"000111110",
  31110=>"100110110",
  31111=>"111000000",
  31112=>"100110111",
  31113=>"100111001",
  31114=>"100101111",
  31115=>"111111111",
  31116=>"111110111",
  31117=>"000110111",
  31118=>"001010000",
  31119=>"000000110",
  31120=>"000000000",
  31121=>"000000111",
  31122=>"111110100",
  31123=>"111011000",
  31124=>"111111110",
  31125=>"000000000",
  31126=>"100000111",
  31127=>"101111111",
  31128=>"111001111",
  31129=>"000100111",
  31130=>"110000001",
  31131=>"111111000",
  31132=>"000000000",
  31133=>"110110100",
  31134=>"000000001",
  31135=>"000000000",
  31136=>"001011010",
  31137=>"111111111",
  31138=>"000000000",
  31139=>"000000001",
  31140=>"111011111",
  31141=>"110111111",
  31142=>"110110110",
  31143=>"000110111",
  31144=>"001111111",
  31145=>"000010111",
  31146=>"111111000",
  31147=>"000100000",
  31148=>"000000000",
  31149=>"101111111",
  31150=>"000000111",
  31151=>"110000000",
  31152=>"111111111",
  31153=>"111100100",
  31154=>"101101111",
  31155=>"000000000",
  31156=>"000000000",
  31157=>"000000000",
  31158=>"111011000",
  31159=>"011000000",
  31160=>"101111111",
  31161=>"111111111",
  31162=>"111001000",
  31163=>"111000000",
  31164=>"001000000",
  31165=>"001000000",
  31166=>"111111000",
  31167=>"101001111",
  31168=>"111111111",
  31169=>"000101111",
  31170=>"000000000",
  31171=>"000000000",
  31172=>"011111111",
  31173=>"110110101",
  31174=>"000110000",
  31175=>"000111111",
  31176=>"000000000",
  31177=>"110111111",
  31178=>"000000001",
  31179=>"000000000",
  31180=>"111111111",
  31181=>"100000000",
  31182=>"000000001",
  31183=>"111100100",
  31184=>"001000000",
  31185=>"111001001",
  31186=>"110011011",
  31187=>"110100001",
  31188=>"111110000",
  31189=>"001000000",
  31190=>"000110110",
  31191=>"010001001",
  31192=>"000000110",
  31193=>"000101111",
  31194=>"000000110",
  31195=>"001001011",
  31196=>"111111111",
  31197=>"100100100",
  31198=>"111000100",
  31199=>"111101000",
  31200=>"000000000",
  31201=>"101111111",
  31202=>"000000001",
  31203=>"111000110",
  31204=>"111111111",
  31205=>"111111111",
  31206=>"011111100",
  31207=>"111111111",
  31208=>"111111111",
  31209=>"111111111",
  31210=>"000000000",
  31211=>"110000000",
  31212=>"000000100",
  31213=>"011111100",
  31214=>"111101000",
  31215=>"111000000",
  31216=>"111001000",
  31217=>"111000000",
  31218=>"110011011",
  31219=>"011011011",
  31220=>"110111111",
  31221=>"000000000",
  31222=>"110111001",
  31223=>"111101001",
  31224=>"000000111",
  31225=>"100111011",
  31226=>"100111111",
  31227=>"000111000",
  31228=>"000111111",
  31229=>"111111000",
  31230=>"111001001",
  31231=>"111111110",
  31232=>"111111111",
  31233=>"001000001",
  31234=>"001000000",
  31235=>"001001000",
  31236=>"000000101",
  31237=>"011011111",
  31238=>"001000100",
  31239=>"000000000",
  31240=>"111010000",
  31241=>"011000000",
  31242=>"110110001",
  31243=>"111001001",
  31244=>"000001000",
  31245=>"111100100",
  31246=>"100111111",
  31247=>"000000000",
  31248=>"111011011",
  31249=>"000111111",
  31250=>"111111110",
  31251=>"111111111",
  31252=>"011100111",
  31253=>"111000000",
  31254=>"111010010",
  31255=>"000111111",
  31256=>"000001100",
  31257=>"111000000",
  31258=>"000000010",
  31259=>"000001111",
  31260=>"111110100",
  31261=>"000110111",
  31262=>"011111111",
  31263=>"000000000",
  31264=>"000000000",
  31265=>"000111111",
  31266=>"111001000",
  31267=>"000000101",
  31268=>"111111111",
  31269=>"000000000",
  31270=>"111010000",
  31271=>"110011000",
  31272=>"001111111",
  31273=>"000000110",
  31274=>"000111111",
  31275=>"000000000",
  31276=>"011000001",
  31277=>"011001001",
  31278=>"111000000",
  31279=>"001000001",
  31280=>"000000000",
  31281=>"000011000",
  31282=>"000000000",
  31283=>"000000000",
  31284=>"000110111",
  31285=>"000001011",
  31286=>"001001001",
  31287=>"011100000",
  31288=>"110100001",
  31289=>"111110000",
  31290=>"000000111",
  31291=>"011011000",
  31292=>"000000000",
  31293=>"011111110",
  31294=>"110111000",
  31295=>"001011111",
  31296=>"100100000",
  31297=>"110110000",
  31298=>"000000111",
  31299=>"000000000",
  31300=>"011011011",
  31301=>"100100000",
  31302=>"000011111",
  31303=>"110100000",
  31304=>"110011011",
  31305=>"111111111",
  31306=>"111111111",
  31307=>"000000000",
  31308=>"111110000",
  31309=>"111110000",
  31310=>"001101101",
  31311=>"001001101",
  31312=>"111100111",
  31313=>"000000111",
  31314=>"011111111",
  31315=>"101111100",
  31316=>"111111111",
  31317=>"011100111",
  31318=>"101000000",
  31319=>"000010010",
  31320=>"101111110",
  31321=>"100000000",
  31322=>"111111111",
  31323=>"111011011",
  31324=>"000000100",
  31325=>"000111011",
  31326=>"001001111",
  31327=>"111100100",
  31328=>"111000000",
  31329=>"000111111",
  31330=>"111111111",
  31331=>"000000000",
  31332=>"000111111",
  31333=>"000000110",
  31334=>"010011111",
  31335=>"000111111",
  31336=>"000110000",
  31337=>"110001000",
  31338=>"111111000",
  31339=>"111111111",
  31340=>"001111111",
  31341=>"011011111",
  31342=>"111110000",
  31343=>"111000000",
  31344=>"111111001",
  31345=>"000110111",
  31346=>"111111001",
  31347=>"111100000",
  31348=>"111110100",
  31349=>"111111000",
  31350=>"000000000",
  31351=>"000000000",
  31352=>"000000000",
  31353=>"111111011",
  31354=>"000000000",
  31355=>"000000000",
  31356=>"110001000",
  31357=>"010111011",
  31358=>"000000000",
  31359=>"111111111",
  31360=>"001001111",
  31361=>"111111111",
  31362=>"111111111",
  31363=>"110111001",
  31364=>"111101000",
  31365=>"111001111",
  31366=>"001111000",
  31367=>"111101000",
  31368=>"011001111",
  31369=>"000000001",
  31370=>"000000000",
  31371=>"100110000",
  31372=>"000000011",
  31373=>"001010010",
  31374=>"101000000",
  31375=>"101000110",
  31376=>"000000100",
  31377=>"111111000",
  31378=>"001001011",
  31379=>"000110111",
  31380=>"110000000",
  31381=>"111001000",
  31382=>"110000000",
  31383=>"000010110",
  31384=>"000001001",
  31385=>"111011000",
  31386=>"000000111",
  31387=>"111111000",
  31388=>"111100101",
  31389=>"011001100",
  31390=>"000000000",
  31391=>"000000000",
  31392=>"111101100",
  31393=>"001001111",
  31394=>"001000111",
  31395=>"000000000",
  31396=>"000001000",
  31397=>"000100111",
  31398=>"000111111",
  31399=>"100100111",
  31400=>"000000000",
  31401=>"000000000",
  31402=>"000000000",
  31403=>"000000000",
  31404=>"111011011",
  31405=>"011011001",
  31406=>"001000000",
  31407=>"000000000",
  31408=>"000000111",
  31409=>"011011011",
  31410=>"010111111",
  31411=>"000000100",
  31412=>"010000001",
  31413=>"111111001",
  31414=>"111111101",
  31415=>"110111111",
  31416=>"111111011",
  31417=>"000111000",
  31418=>"000000001",
  31419=>"100110000",
  31420=>"111001111",
  31421=>"111111110",
  31422=>"111111111",
  31423=>"111000000",
  31424=>"001011011",
  31425=>"000000010",
  31426=>"111111111",
  31427=>"101001000",
  31428=>"000000111",
  31429=>"001000011",
  31430=>"000100100",
  31431=>"001101110",
  31432=>"110000000",
  31433=>"000001111",
  31434=>"101111111",
  31435=>"000000000",
  31436=>"001110111",
  31437=>"100111011",
  31438=>"111100000",
  31439=>"100111111",
  31440=>"111111000",
  31441=>"011000000",
  31442=>"000000101",
  31443=>"011000000",
  31444=>"000000101",
  31445=>"000000000",
  31446=>"111011011",
  31447=>"000111111",
  31448=>"101101000",
  31449=>"000111111",
  31450=>"000000000",
  31451=>"111100000",
  31452=>"111111011",
  31453=>"010010000",
  31454=>"000000010",
  31455=>"001101100",
  31456=>"000000100",
  31457=>"111111011",
  31458=>"110000111",
  31459=>"111000000",
  31460=>"100100101",
  31461=>"111111100",
  31462=>"000011001",
  31463=>"111110110",
  31464=>"000101101",
  31465=>"110100110",
  31466=>"111101111",
  31467=>"000000000",
  31468=>"000000000",
  31469=>"111110111",
  31470=>"000000001",
  31471=>"111000100",
  31472=>"111111110",
  31473=>"000110101",
  31474=>"000000000",
  31475=>"101101010",
  31476=>"000111111",
  31477=>"011011001",
  31478=>"111101101",
  31479=>"011010111",
  31480=>"111000000",
  31481=>"111111111",
  31482=>"001000000",
  31483=>"000000111",
  31484=>"000000110",
  31485=>"001111111",
  31486=>"011111111",
  31487=>"000000100",
  31488=>"000000000",
  31489=>"000011110",
  31490=>"110111111",
  31491=>"000000000",
  31492=>"111111110",
  31493=>"001111111",
  31494=>"000000000",
  31495=>"000111111",
  31496=>"101000000",
  31497=>"111111011",
  31498=>"111011111",
  31499=>"000000000",
  31500=>"011011011",
  31501=>"001000011",
  31502=>"000000000",
  31503=>"001001000",
  31504=>"111000000",
  31505=>"100000000",
  31506=>"000000111",
  31507=>"000001000",
  31508=>"011111111",
  31509=>"000000001",
  31510=>"011011001",
  31511=>"000000000",
  31512=>"000010110",
  31513=>"111111110",
  31514=>"000000000",
  31515=>"111111111",
  31516=>"001110100",
  31517=>"110110010",
  31518=>"000111111",
  31519=>"100000000",
  31520=>"111101000",
  31521=>"000000000",
  31522=>"000000000",
  31523=>"111111001",
  31524=>"000000000",
  31525=>"010010111",
  31526=>"111111101",
  31527=>"111011000",
  31528=>"100111110",
  31529=>"000000111",
  31530=>"111111111",
  31531=>"110111011",
  31532=>"000000111",
  31533=>"000011010",
  31534=>"111111111",
  31535=>"000000111",
  31536=>"111111010",
  31537=>"000000111",
  31538=>"011000001",
  31539=>"000000000",
  31540=>"000000000",
  31541=>"100111000",
  31542=>"000110110",
  31543=>"000111111",
  31544=>"110000011",
  31545=>"110000011",
  31546=>"111111000",
  31547=>"110000000",
  31548=>"000000000",
  31549=>"111111001",
  31550=>"110111100",
  31551=>"111010000",
  31552=>"100100100",
  31553=>"000100000",
  31554=>"000111000",
  31555=>"000000001",
  31556=>"000000110",
  31557=>"000000000",
  31558=>"111111111",
  31559=>"101111111",
  31560=>"000000010",
  31561=>"111000000",
  31562=>"001111111",
  31563=>"010111111",
  31564=>"011000000",
  31565=>"100110111",
  31566=>"111001000",
  31567=>"000000000",
  31568=>"111111110",
  31569=>"111101101",
  31570=>"111110000",
  31571=>"000000001",
  31572=>"000000000",
  31573=>"110100000",
  31574=>"111100000",
  31575=>"110000011",
  31576=>"001000000",
  31577=>"101100111",
  31578=>"111111000",
  31579=>"111111111",
  31580=>"111010000",
  31581=>"111110100",
  31582=>"001111111",
  31583=>"101000000",
  31584=>"101111111",
  31585=>"001001111",
  31586=>"100111111",
  31587=>"011001111",
  31588=>"100111111",
  31589=>"000000111",
  31590=>"000000101",
  31591=>"000111111",
  31592=>"011111111",
  31593=>"010000000",
  31594=>"000111111",
  31595=>"111101111",
  31596=>"100000000",
  31597=>"001001000",
  31598=>"000001111",
  31599=>"111111000",
  31600=>"001000000",
  31601=>"111011000",
  31602=>"000000000",
  31603=>"111100000",
  31604=>"111001000",
  31605=>"000000111",
  31606=>"000000000",
  31607=>"111110000",
  31608=>"001000001",
  31609=>"111111000",
  31610=>"000101111",
  31611=>"001000100",
  31612=>"111111110",
  31613=>"000000111",
  31614=>"011001100",
  31615=>"000000111",
  31616=>"000111110",
  31617=>"101000000",
  31618=>"001001001",
  31619=>"110000000",
  31620=>"000000001",
  31621=>"000011010",
  31622=>"111111111",
  31623=>"111000000",
  31624=>"001001111",
  31625=>"110111100",
  31626=>"111000000",
  31627=>"010111111",
  31628=>"111111111",
  31629=>"001001001",
  31630=>"111111111",
  31631=>"000001011",
  31632=>"000001000",
  31633=>"111111001",
  31634=>"111011110",
  31635=>"000000000",
  31636=>"000011111",
  31637=>"000010000",
  31638=>"111111011",
  31639=>"001001000",
  31640=>"111101000",
  31641=>"111011001",
  31642=>"111111111",
  31643=>"111110110",
  31644=>"101111001",
  31645=>"001111001",
  31646=>"000000101",
  31647=>"000000111",
  31648=>"111111111",
  31649=>"110110100",
  31650=>"100110010",
  31651=>"001000001",
  31652=>"000000000",
  31653=>"111110000",
  31654=>"100100100",
  31655=>"001111111",
  31656=>"000010011",
  31657=>"000011111",
  31658=>"000000000",
  31659=>"001101001",
  31660=>"111111111",
  31661=>"111001000",
  31662=>"000101000",
  31663=>"001000000",
  31664=>"111111111",
  31665=>"010001000",
  31666=>"001111111",
  31667=>"011000000",
  31668=>"111100000",
  31669=>"000000111",
  31670=>"100100111",
  31671=>"100000000",
  31672=>"110000000",
  31673=>"111111001",
  31674=>"000000000",
  31675=>"101000000",
  31676=>"111111110",
  31677=>"110101111",
  31678=>"000110111",
  31679=>"111111111",
  31680=>"111001001",
  31681=>"001000000",
  31682=>"011001000",
  31683=>"000110010",
  31684=>"111111001",
  31685=>"100011001",
  31686=>"111101000",
  31687=>"111111111",
  31688=>"000111111",
  31689=>"100100011",
  31690=>"000000000",
  31691=>"000000110",
  31692=>"100111001",
  31693=>"111111111",
  31694=>"001000001",
  31695=>"111000000",
  31696=>"010000000",
  31697=>"001111111",
  31698=>"110111111",
  31699=>"000101100",
  31700=>"110000111",
  31701=>"000000000",
  31702=>"011111111",
  31703=>"000110111",
  31704=>"100001001",
  31705=>"111000001",
  31706=>"111100000",
  31707=>"110001001",
  31708=>"000111111",
  31709=>"001111111",
  31710=>"000010000",
  31711=>"000000000",
  31712=>"111011000",
  31713=>"000010000",
  31714=>"001000111",
  31715=>"001000000",
  31716=>"111111000",
  31717=>"100110000",
  31718=>"010000010",
  31719=>"011000111",
  31720=>"101101100",
  31721=>"111111000",
  31722=>"110000000",
  31723=>"001011011",
  31724=>"000111111",
  31725=>"110111110",
  31726=>"000100100",
  31727=>"000111111",
  31728=>"001111000",
  31729=>"000000000",
  31730=>"101111110",
  31731=>"000110111",
  31732=>"001011011",
  31733=>"001001111",
  31734=>"000110111",
  31735=>"011011011",
  31736=>"100111111",
  31737=>"011111101",
  31738=>"010010011",
  31739=>"111111111",
  31740=>"111111111",
  31741=>"011111111",
  31742=>"111011000",
  31743=>"000001000",
  31744=>"111111111",
  31745=>"010010010",
  31746=>"000000111",
  31747=>"000000000",
  31748=>"111111111",
  31749=>"010000000",
  31750=>"000000111",
  31751=>"100000111",
  31752=>"000000000",
  31753=>"000000111",
  31754=>"000000000",
  31755=>"111111100",
  31756=>"100100110",
  31757=>"111100001",
  31758=>"111011111",
  31759=>"000000111",
  31760=>"000000000",
  31761=>"000000000",
  31762=>"111111111",
  31763=>"000000000",
  31764=>"010010000",
  31765=>"000000111",
  31766=>"000000000",
  31767=>"000000000",
  31768=>"111111111",
  31769=>"000000000",
  31770=>"000100000",
  31771=>"110111111",
  31772=>"111110100",
  31773=>"111111111",
  31774=>"000000000",
  31775=>"001000000",
  31776=>"110110111",
  31777=>"001001111",
  31778=>"110110110",
  31779=>"100100100",
  31780=>"110000000",
  31781=>"000000000",
  31782=>"111111111",
  31783=>"111111010",
  31784=>"001001111",
  31785=>"111000000",
  31786=>"110111111",
  31787=>"000110111",
  31788=>"110010000",
  31789=>"000000100",
  31790=>"111111111",
  31791=>"100101111",
  31792=>"000011111",
  31793=>"111101100",
  31794=>"011111011",
  31795=>"111000011",
  31796=>"000000000",
  31797=>"011000000",
  31798=>"000001000",
  31799=>"111111111",
  31800=>"101101101",
  31801=>"000000000",
  31802=>"010001110",
  31803=>"111111111",
  31804=>"000000111",
  31805=>"111111100",
  31806=>"111111111",
  31807=>"000000000",
  31808=>"111111000",
  31809=>"011101100",
  31810=>"000000000",
  31811=>"010010010",
  31812=>"111111111",
  31813=>"110100100",
  31814=>"111111011",
  31815=>"111111111",
  31816=>"000000000",
  31817=>"001101111",
  31818=>"000000000",
  31819=>"000000000",
  31820=>"000000000",
  31821=>"000000000",
  31822=>"000000100",
  31823=>"000000000",
  31824=>"111111000",
  31825=>"001000000",
  31826=>"111110000",
  31827=>"111100100",
  31828=>"000111011",
  31829=>"001111111",
  31830=>"011011000",
  31831=>"000000101",
  31832=>"100111111",
  31833=>"111001101",
  31834=>"111110100",
  31835=>"000011001",
  31836=>"111111111",
  31837=>"011111011",
  31838=>"011000000",
  31839=>"111111011",
  31840=>"111100100",
  31841=>"111101000",
  31842=>"000000000",
  31843=>"001001111",
  31844=>"111101111",
  31845=>"111111111",
  31846=>"111110111",
  31847=>"000010111",
  31848=>"111111111",
  31849=>"100000000",
  31850=>"011011000",
  31851=>"111100000",
  31852=>"111111111",
  31853=>"000000000",
  31854=>"000000000",
  31855=>"111111111",
  31856=>"101000000",
  31857=>"011011111",
  31858=>"100110111",
  31859=>"111111111",
  31860=>"000000000",
  31861=>"111100000",
  31862=>"000110111",
  31863=>"111111110",
  31864=>"111111111",
  31865=>"000000000",
  31866=>"111100101",
  31867=>"111111011",
  31868=>"111000000",
  31869=>"011011000",
  31870=>"001001001",
  31871=>"111000000",
  31872=>"000000000",
  31873=>"111111000",
  31874=>"111111000",
  31875=>"111111011",
  31876=>"000000000",
  31877=>"110001001",
  31878=>"111111111",
  31879=>"111111111",
  31880=>"000000001",
  31881=>"101111111",
  31882=>"000000000",
  31883=>"111111111",
  31884=>"010010110",
  31885=>"000000000",
  31886=>"000111001",
  31887=>"111111000",
  31888=>"000000000",
  31889=>"110000000",
  31890=>"111111111",
  31891=>"110110111",
  31892=>"000000000",
  31893=>"000100100",
  31894=>"101000000",
  31895=>"000001111",
  31896=>"101101010",
  31897=>"111111111",
  31898=>"000000011",
  31899=>"111100111",
  31900=>"100110100",
  31901=>"000000111",
  31902=>"000000000",
  31903=>"000000000",
  31904=>"000001111",
  31905=>"111110100",
  31906=>"111111111",
  31907=>"001011000",
  31908=>"000000001",
  31909=>"000000000",
  31910=>"111111111",
  31911=>"100000100",
  31912=>"110110000",
  31913=>"000000000",
  31914=>"000000000",
  31915=>"011000000",
  31916=>"110010111",
  31917=>"011111010",
  31918=>"110111111",
  31919=>"111000000",
  31920=>"100110100",
  31921=>"011000000",
  31922=>"110111111",
  31923=>"100100100",
  31924=>"000010111",
  31925=>"111111111",
  31926=>"111111111",
  31927=>"111111000",
  31928=>"000000110",
  31929=>"111000000",
  31930=>"111011000",
  31931=>"000111000",
  31932=>"001101000",
  31933=>"010000111",
  31934=>"000000000",
  31935=>"000111111",
  31936=>"111101101",
  31937=>"000000000",
  31938=>"100101101",
  31939=>"000000000",
  31940=>"100110000",
  31941=>"111111000",
  31942=>"011111111",
  31943=>"111111111",
  31944=>"111111000",
  31945=>"111100110",
  31946=>"111111001",
  31947=>"000000110",
  31948=>"000000000",
  31949=>"111100111",
  31950=>"000000100",
  31951=>"000000000",
  31952=>"000000000",
  31953=>"111111110",
  31954=>"111111111",
  31955=>"111111100",
  31956=>"111110111",
  31957=>"111111110",
  31958=>"111111111",
  31959=>"100000000",
  31960=>"100000000",
  31961=>"111111110",
  31962=>"100101110",
  31963=>"000000000",
  31964=>"111111001",
  31965=>"111111111",
  31966=>"000000000",
  31967=>"110110111",
  31968=>"111000110",
  31969=>"101001111",
  31970=>"000000000",
  31971=>"000000000",
  31972=>"110110000",
  31973=>"000000100",
  31974=>"111111111",
  31975=>"111001000",
  31976=>"111111111",
  31977=>"111111111",
  31978=>"111100100",
  31979=>"111111111",
  31980=>"111111011",
  31981=>"000000000",
  31982=>"000000000",
  31983=>"000000111",
  31984=>"011110000",
  31985=>"100111111",
  31986=>"111111111",
  31987=>"011111000",
  31988=>"111111111",
  31989=>"111111111",
  31990=>"001111111",
  31991=>"111000000",
  31992=>"000000000",
  31993=>"000001001",
  31994=>"111111000",
  31995=>"110100100",
  31996=>"111001011",
  31997=>"000000001",
  31998=>"000000000",
  31999=>"000010000",
  32000=>"000100110",
  32001=>"111111011",
  32002=>"000000000",
  32003=>"000000000",
  32004=>"000000000",
  32005=>"110110111",
  32006=>"111011000",
  32007=>"000000001",
  32008=>"111111000",
  32009=>"000000000",
  32010=>"000110000",
  32011=>"111001000",
  32012=>"111101001",
  32013=>"111111111",
  32014=>"000111111",
  32015=>"111111110",
  32016=>"000011011",
  32017=>"000000000",
  32018=>"101100000",
  32019=>"111111111",
  32020=>"000010000",
  32021=>"000000000",
  32022=>"000000000",
  32023=>"111111000",
  32024=>"111010000",
  32025=>"000000000",
  32026=>"100100100",
  32027=>"111111101",
  32028=>"100100000",
  32029=>"000000000",
  32030=>"010111100",
  32031=>"111111001",
  32032=>"111110000",
  32033=>"111111111",
  32034=>"000010000",
  32035=>"111000000",
  32036=>"000100110",
  32037=>"110110100",
  32038=>"000111111",
  32039=>"001001011",
  32040=>"111111111",
  32041=>"111110000",
  32042=>"100000100",
  32043=>"110111111",
  32044=>"111111111",
  32045=>"011000000",
  32046=>"000010111",
  32047=>"000000000",
  32048=>"111111111",
  32049=>"011111001",
  32050=>"111111111",
  32051=>"010000000",
  32052=>"111001000",
  32053=>"111011001",
  32054=>"000100000",
  32055=>"000100000",
  32056=>"000000000",
  32057=>"110100000",
  32058=>"111111111",
  32059=>"000000000",
  32060=>"010010011",
  32061=>"110110000",
  32062=>"000001001",
  32063=>"000000001",
  32064=>"000000000",
  32065=>"110111000",
  32066=>"111111111",
  32067=>"000000000",
  32068=>"000000000",
  32069=>"000000001",
  32070=>"100000000",
  32071=>"000000001",
  32072=>"000001000",
  32073=>"100100000",
  32074=>"010000011",
  32075=>"011111001",
  32076=>"100010000",
  32077=>"000000111",
  32078=>"111111001",
  32079=>"111000000",
  32080=>"111011000",
  32081=>"001000000",
  32082=>"000000000",
  32083=>"111111111",
  32084=>"000000000",
  32085=>"001000000",
  32086=>"000001001",
  32087=>"000000000",
  32088=>"000000000",
  32089=>"111111111",
  32090=>"000010111",
  32091=>"000000000",
  32092=>"000000001",
  32093=>"101000000",
  32094=>"111000000",
  32095=>"000000110",
  32096=>"111111111",
  32097=>"000111111",
  32098=>"000010000",
  32099=>"111100000",
  32100=>"111111111",
  32101=>"111111011",
  32102=>"000000000",
  32103=>"000001101",
  32104=>"010011010",
  32105=>"000000010",
  32106=>"111111111",
  32107=>"001111111",
  32108=>"000000000",
  32109=>"000000000",
  32110=>"001000000",
  32111=>"111111111",
  32112=>"111111111",
  32113=>"000000000",
  32114=>"110010001",
  32115=>"111111111",
  32116=>"000000000",
  32117=>"000000000",
  32118=>"111011001",
  32119=>"110111000",
  32120=>"111000101",
  32121=>"110110000",
  32122=>"111111111",
  32123=>"000000000",
  32124=>"111111111",
  32125=>"000000000",
  32126=>"001100101",
  32127=>"000000000",
  32128=>"001001000",
  32129=>"111000001",
  32130=>"011001000",
  32131=>"001000000",
  32132=>"000100111",
  32133=>"001000000",
  32134=>"111101101",
  32135=>"011001011",
  32136=>"000000111",
  32137=>"000000000",
  32138=>"111101000",
  32139=>"111100000",
  32140=>"111111111",
  32141=>"011011011",
  32142=>"110100111",
  32143=>"111111111",
  32144=>"111111111",
  32145=>"000000000",
  32146=>"111111111",
  32147=>"100110110",
  32148=>"111111111",
  32149=>"111111001",
  32150=>"111111111",
  32151=>"111111110",
  32152=>"000000001",
  32153=>"111001001",
  32154=>"101100100",
  32155=>"111111111",
  32156=>"111111111",
  32157=>"111111110",
  32158=>"000011011",
  32159=>"000000000",
  32160=>"100100000",
  32161=>"000000000",
  32162=>"111001000",
  32163=>"110000000",
  32164=>"111111110",
  32165=>"011111111",
  32166=>"111111111",
  32167=>"111111111",
  32168=>"000000000",
  32169=>"000000000",
  32170=>"011111101",
  32171=>"111111111",
  32172=>"111111111",
  32173=>"000001000",
  32174=>"000000000",
  32175=>"111101010",
  32176=>"011001001",
  32177=>"000000000",
  32178=>"011111111",
  32179=>"000000000",
  32180=>"111000000",
  32181=>"011000101",
  32182=>"111111111",
  32183=>"110111010",
  32184=>"000000111",
  32185=>"000000000",
  32186=>"000000000",
  32187=>"011010000",
  32188=>"100100111",
  32189=>"010000100",
  32190=>"010000000",
  32191=>"111110010",
  32192=>"111000000",
  32193=>"111111111",
  32194=>"000111111",
  32195=>"000110010",
  32196=>"111110111",
  32197=>"000000000",
  32198=>"110110000",
  32199=>"110100100",
  32200=>"000100111",
  32201=>"101111111",
  32202=>"111111111",
  32203=>"010110110",
  32204=>"100000110",
  32205=>"111111111",
  32206=>"110110000",
  32207=>"111111111",
  32208=>"100000000",
  32209=>"111011001",
  32210=>"000000000",
  32211=>"100000000",
  32212=>"111111111",
  32213=>"110100100",
  32214=>"111111101",
  32215=>"000000010",
  32216=>"000000000",
  32217=>"000000001",
  32218=>"000000000",
  32219=>"111111111",
  32220=>"000000001",
  32221=>"000010001",
  32222=>"000000111",
  32223=>"000100100",
  32224=>"000100111",
  32225=>"000000000",
  32226=>"011011001",
  32227=>"111111111",
  32228=>"110011001",
  32229=>"100100001",
  32230=>"001001011",
  32231=>"000010010",
  32232=>"000000000",
  32233=>"000111010",
  32234=>"000000000",
  32235=>"000000001",
  32236=>"010110011",
  32237=>"111110111",
  32238=>"000111111",
  32239=>"000000000",
  32240=>"111000011",
  32241=>"000110100",
  32242=>"111111111",
  32243=>"111111110",
  32244=>"111111111",
  32245=>"101101111",
  32246=>"111111111",
  32247=>"000000110",
  32248=>"000000000",
  32249=>"000011001",
  32250=>"111111111",
  32251=>"000000000",
  32252=>"110000000",
  32253=>"000000100",
  32254=>"000011011",
  32255=>"111011111",
  32256=>"000000100",
  32257=>"100111111",
  32258=>"000000010",
  32259=>"111111111",
  32260=>"111111111",
  32261=>"000000001",
  32262=>"100100100",
  32263=>"000000000",
  32264=>"000000000",
  32265=>"000111111",
  32266=>"100000100",
  32267=>"000110110",
  32268=>"100101111",
  32269=>"000001011",
  32270=>"111011111",
  32271=>"000000000",
  32272=>"000000001",
  32273=>"000000111",
  32274=>"100100110",
  32275=>"000000000",
  32276=>"111111101",
  32277=>"000000001",
  32278=>"000000000",
  32279=>"111111000",
  32280=>"000000111",
  32281=>"100111111",
  32282=>"111111000",
  32283=>"011001000",
  32284=>"000000111",
  32285=>"001000000",
  32286=>"110110110",
  32287=>"111111011",
  32288=>"110110111",
  32289=>"111111111",
  32290=>"011011010",
  32291=>"111111111",
  32292=>"111111111",
  32293=>"111110111",
  32294=>"010010110",
  32295=>"111000000",
  32296=>"011011011",
  32297=>"111000000",
  32298=>"111111111",
  32299=>"000000000",
  32300=>"000000001",
  32301=>"001111111",
  32302=>"000000000",
  32303=>"111111000",
  32304=>"010110110",
  32305=>"110100100",
  32306=>"111111111",
  32307=>"000000110",
  32308=>"101111111",
  32309=>"000000000",
  32310=>"110001000",
  32311=>"010000100",
  32312=>"111000000",
  32313=>"111111000",
  32314=>"001001111",
  32315=>"000000001",
  32316=>"000000111",
  32317=>"001111111",
  32318=>"111000000",
  32319=>"001001001",
  32320=>"011011111",
  32321=>"000110111",
  32322=>"000000000",
  32323=>"001000111",
  32324=>"111111111",
  32325=>"111111110",
  32326=>"111111101",
  32327=>"000000000",
  32328=>"111111111",
  32329=>"000000000",
  32330=>"001011100",
  32331=>"000110111",
  32332=>"111111111",
  32333=>"110010110",
  32334=>"000000110",
  32335=>"111111111",
  32336=>"111111111",
  32337=>"011011111",
  32338=>"010111111",
  32339=>"011111001",
  32340=>"000000000",
  32341=>"001000000",
  32342=>"011010000",
  32343=>"111111111",
  32344=>"000000111",
  32345=>"001001001",
  32346=>"111111000",
  32347=>"110110110",
  32348=>"110000000",
  32349=>"110110100",
  32350=>"000001011",
  32351=>"101101101",
  32352=>"000000000",
  32353=>"000000000",
  32354=>"111000000",
  32355=>"110100111",
  32356=>"000100001",
  32357=>"110110000",
  32358=>"000010000",
  32359=>"000000000",
  32360=>"000101111",
  32361=>"001111111",
  32362=>"011000110",
  32363=>"000000000",
  32364=>"001000000",
  32365=>"111111000",
  32366=>"000000000",
  32367=>"111110010",
  32368=>"001111111",
  32369=>"011110111",
  32370=>"011111111",
  32371=>"110000111",
  32372=>"011000000",
  32373=>"110110000",
  32374=>"001001111",
  32375=>"000000000",
  32376=>"000000000",
  32377=>"000000000",
  32378=>"100000000",
  32379=>"000000000",
  32380=>"000110100",
  32381=>"000000000",
  32382=>"110000000",
  32383=>"111111111",
  32384=>"111111010",
  32385=>"000000000",
  32386=>"011011111",
  32387=>"011110100",
  32388=>"111010000",
  32389=>"000001001",
  32390=>"001100111",
  32391=>"011001001",
  32392=>"100111111",
  32393=>"000000000",
  32394=>"110111111",
  32395=>"100000000",
  32396=>"101000001",
  32397=>"000010111",
  32398=>"000000011",
  32399=>"101101101",
  32400=>"100100101",
  32401=>"000000000",
  32402=>"000101000",
  32403=>"000000000",
  32404=>"000000000",
  32405=>"011111111",
  32406=>"000000111",
  32407=>"000000010",
  32408=>"000000111",
  32409=>"001101111",
  32410=>"111111110",
  32411=>"011001111",
  32412=>"000001000",
  32413=>"000100111",
  32414=>"000001000",
  32415=>"111111011",
  32416=>"111001101",
  32417=>"100000111",
  32418=>"000000000",
  32419=>"000000000",
  32420=>"100000000",
  32421=>"101000000",
  32422=>"001111000",
  32423=>"000100001",
  32424=>"000000100",
  32425=>"000111111",
  32426=>"100100100",
  32427=>"111111101",
  32428=>"001000101",
  32429=>"011011000",
  32430=>"000110111",
  32431=>"111111111",
  32432=>"011111010",
  32433=>"110110001",
  32434=>"011011011",
  32435=>"111111111",
  32436=>"010111111",
  32437=>"001000100",
  32438=>"111111000",
  32439=>"000100111",
  32440=>"111111001",
  32441=>"000000000",
  32442=>"110100100",
  32443=>"000000011",
  32444=>"111000000",
  32445=>"110111001",
  32446=>"111011001",
  32447=>"100000101",
  32448=>"010000000",
  32449=>"000111100",
  32450=>"000000000",
  32451=>"101011110",
  32452=>"011111111",
  32453=>"000011111",
  32454=>"000000000",
  32455=>"010110100",
  32456=>"000001111",
  32457=>"101101111",
  32458=>"000000111",
  32459=>"111111110",
  32460=>"101101001",
  32461=>"111111001",
  32462=>"000000111",
  32463=>"000000000",
  32464=>"001111111",
  32465=>"000011111",
  32466=>"000000111",
  32467=>"110100100",
  32468=>"110000000",
  32469=>"000000000",
  32470=>"000000000",
  32471=>"011000000",
  32472=>"111111111",
  32473=>"001000111",
  32474=>"000000011",
  32475=>"110000000",
  32476=>"011111111",
  32477=>"111111110",
  32478=>"001001011",
  32479=>"000000000",
  32480=>"000000000",
  32481=>"000010000",
  32482=>"111011001",
  32483=>"111110110",
  32484=>"100010000",
  32485=>"111011011",
  32486=>"111111011",
  32487=>"000000000",
  32488=>"000000000",
  32489=>"111000000",
  32490=>"000111111",
  32491=>"111111001",
  32492=>"000000001",
  32493=>"101000111",
  32494=>"100100100",
  32495=>"000111111",
  32496=>"001000000",
  32497=>"111111000",
  32498=>"110100111",
  32499=>"001000000",
  32500=>"001000111",
  32501=>"000111111",
  32502=>"000011111",
  32503=>"000000111",
  32504=>"111111011",
  32505=>"000000000",
  32506=>"000000000",
  32507=>"000000010",
  32508=>"011011000",
  32509=>"101100111",
  32510=>"011000000",
  32511=>"111011011",
  32512=>"110110110",
  32513=>"100100000",
  32514=>"111111111",
  32515=>"000000100",
  32516=>"110100110",
  32517=>"000000000",
  32518=>"000000000",
  32519=>"011111110",
  32520=>"001000000",
  32521=>"000111111",
  32522=>"111111011",
  32523=>"000100111",
  32524=>"101001111",
  32525=>"000010110",
  32526=>"111010110",
  32527=>"000011111",
  32528=>"111111110",
  32529=>"000000111",
  32530=>"001000000",
  32531=>"100111111",
  32532=>"110111111",
  32533=>"011000000",
  32534=>"001100100",
  32535=>"101001111",
  32536=>"001111111",
  32537=>"100110000",
  32538=>"110010000",
  32539=>"001000110",
  32540=>"001000000",
  32541=>"000001111",
  32542=>"100111111",
  32543=>"101001101",
  32544=>"000000000",
  32545=>"110111010",
  32546=>"001100110",
  32547=>"001001101",
  32548=>"110110110",
  32549=>"110100111",
  32550=>"000111111",
  32551=>"000000111",
  32552=>"111111100",
  32553=>"100101111",
  32554=>"000001011",
  32555=>"000001111",
  32556=>"111111111",
  32557=>"000000000",
  32558=>"111000111",
  32559=>"101101111",
  32560=>"110111111",
  32561=>"000110010",
  32562=>"011001111",
  32563=>"000110110",
  32564=>"110000000",
  32565=>"011111111",
  32566=>"111001101",
  32567=>"000000011",
  32568=>"011011001",
  32569=>"001001000",
  32570=>"111110000",
  32571=>"110111111",
  32572=>"111111000",
  32573=>"000111001",
  32574=>"111111111",
  32575=>"111111001",
  32576=>"000000000",
  32577=>"111011000",
  32578=>"000000111",
  32579=>"001001000",
  32580=>"000000111",
  32581=>"111111111",
  32582=>"111111110",
  32583=>"000000000",
  32584=>"111110000",
  32585=>"101101111",
  32586=>"000001101",
  32587=>"001001011",
  32588=>"000110110",
  32589=>"111111111",
  32590=>"001001001",
  32591=>"111101101",
  32592=>"011111001",
  32593=>"000000000",
  32594=>"000000010",
  32595=>"000000000",
  32596=>"111000111",
  32597=>"000011001",
  32598=>"000000111",
  32599=>"100111101",
  32600=>"000000111",
  32601=>"111111111",
  32602=>"110111111",
  32603=>"111111111",
  32604=>"000100111",
  32605=>"100100111",
  32606=>"000001111",
  32607=>"000001000",
  32608=>"000000110",
  32609=>"100000111",
  32610=>"111111110",
  32611=>"000000000",
  32612=>"000000000",
  32613=>"000001001",
  32614=>"111111000",
  32615=>"000000111",
  32616=>"000000000",
  32617=>"110111111",
  32618=>"000000000",
  32619=>"000000000",
  32620=>"000000000",
  32621=>"100000000",
  32622=>"111100110",
  32623=>"000000000",
  32624=>"111111111",
  32625=>"010010000",
  32626=>"000001111",
  32627=>"011001001",
  32628=>"010110110",
  32629=>"111011111",
  32630=>"111111111",
  32631=>"111111001",
  32632=>"100100000",
  32633=>"111111111",
  32634=>"111011000",
  32635=>"011000000",
  32636=>"000000110",
  32637=>"011011100",
  32638=>"111100100",
  32639=>"000111111",
  32640=>"000111111",
  32641=>"011011101",
  32642=>"110101000",
  32643=>"000000111",
  32644=>"111111000",
  32645=>"000100000",
  32646=>"100100111",
  32647=>"100000111",
  32648=>"100100000",
  32649=>"011011000",
  32650=>"000000001",
  32651=>"000011001",
  32652=>"111111101",
  32653=>"111111111",
  32654=>"011011011",
  32655=>"000000000",
  32656=>"110110000",
  32657=>"000100000",
  32658=>"111111100",
  32659=>"111111000",
  32660=>"000000000",
  32661=>"010010000",
  32662=>"111111111",
  32663=>"000000110",
  32664=>"000000000",
  32665=>"000000000",
  32666=>"000000000",
  32667=>"111111111",
  32668=>"000000000",
  32669=>"111111011",
  32670=>"000010000",
  32671=>"111111001",
  32672=>"101100100",
  32673=>"111111011",
  32674=>"000000111",
  32675=>"111111111",
  32676=>"011111111",
  32677=>"000001111",
  32678=>"111111001",
  32679=>"000000000",
  32680=>"000001000",
  32681=>"001000000",
  32682=>"000110111",
  32683=>"000000010",
  32684=>"111111100",
  32685=>"111000000",
  32686=>"110111000",
  32687=>"111111111",
  32688=>"000000000",
  32689=>"111111111",
  32690=>"000100111",
  32691=>"111111110",
  32692=>"101001001",
  32693=>"000000110",
  32694=>"000011111",
  32695=>"111111111",
  32696=>"000000100",
  32697=>"011111111",
  32698=>"000000011",
  32699=>"000000101",
  32700=>"011001001",
  32701=>"000101111",
  32702=>"000000001",
  32703=>"001101000",
  32704=>"000110111",
  32705=>"000001001",
  32706=>"000000000",
  32707=>"111111111",
  32708=>"111111111",
  32709=>"111000000",
  32710=>"111110000",
  32711=>"111111011",
  32712=>"000000100",
  32713=>"000000000",
  32714=>"000000110",
  32715=>"101001111",
  32716=>"011011000",
  32717=>"111111011",
  32718=>"011001000",
  32719=>"010111111",
  32720=>"100111111",
  32721=>"111111111",
  32722=>"101111110",
  32723=>"000000001",
  32724=>"001000000",
  32725=>"110110111",
  32726=>"111111010",
  32727=>"111111111",
  32728=>"000010110",
  32729=>"100000110",
  32730=>"000000001",
  32731=>"000000000",
  32732=>"011111111",
  32733=>"101111111",
  32734=>"111111000",
  32735=>"100100000",
  32736=>"001101111",
  32737=>"000000000",
  32738=>"111111000",
  32739=>"011111111",
  32740=>"000000000",
  32741=>"111111001",
  32742=>"000000001",
  32743=>"111111101",
  32744=>"001000111",
  32745=>"111110100",
  32746=>"000000000",
  32747=>"000000000",
  32748=>"000001001",
  32749=>"111111011",
  32750=>"111100000",
  32751=>"000001111",
  32752=>"111111111",
  32753=>"000010000",
  32754=>"000101111",
  32755=>"000001001",
  32756=>"000000100",
  32757=>"111110111",
  32758=>"111111111",
  32759=>"000000011",
  32760=>"011000000",
  32761=>"111101001",
  32762=>"000100000",
  32763=>"001001000",
  32764=>"000000000",
  32765=>"000000000",
  32766=>"111000000",
  32767=>"000000111",
  32768=>"101111111",
  32769=>"001010000",
  32770=>"000000000",
  32771=>"000111111",
  32772=>"100010000",
  32773=>"000000001",
  32774=>"000000000",
  32775=>"111101100",
  32776=>"000000000",
  32777=>"110111011",
  32778=>"000000100",
  32779=>"111111111",
  32780=>"110110110",
  32781=>"111000000",
  32782=>"000001111",
  32783=>"000000001",
  32784=>"000000000",
  32785=>"000100000",
  32786=>"000101101",
  32787=>"111111110",
  32788=>"111000011",
  32789=>"110000001",
  32790=>"111111100",
  32791=>"001001001",
  32792=>"110000000",
  32793=>"101100111",
  32794=>"011110111",
  32795=>"000000000",
  32796=>"111111011",
  32797=>"000111111",
  32798=>"000000011",
  32799=>"100000000",
  32800=>"111000100",
  32801=>"000100111",
  32802=>"000100000",
  32803=>"000000000",
  32804=>"000000111",
  32805=>"111111111",
  32806=>"001001001",
  32807=>"111000001",
  32808=>"000100101",
  32809=>"000000000",
  32810=>"000000000",
  32811=>"000000000",
  32812=>"110111111",
  32813=>"110110110",
  32814=>"000000000",
  32815=>"111001000",
  32816=>"111111111",
  32817=>"111111111",
  32818=>"001001001",
  32819=>"001011111",
  32820=>"111000000",
  32821=>"001000000",
  32822=>"000001001",
  32823=>"000111110",
  32824=>"111111111",
  32825=>"110000001",
  32826=>"111111000",
  32827=>"111111111",
  32828=>"011011101",
  32829=>"000000000",
  32830=>"100100000",
  32831=>"101101001",
  32832=>"110111011",
  32833=>"110010000",
  32834=>"010010111",
  32835=>"100001001",
  32836=>"001000000",
  32837=>"111111111",
  32838=>"111111000",
  32839=>"000000000",
  32840=>"011011011",
  32841=>"010010000",
  32842=>"000001001",
  32843=>"100100110",
  32844=>"111111111",
  32845=>"111111000",
  32846=>"000010011",
  32847=>"111111111",
  32848=>"111111000",
  32849=>"000000010",
  32850=>"001000000",
  32851=>"111111101",
  32852=>"001000101",
  32853=>"100000000",
  32854=>"111011011",
  32855=>"011111110",
  32856=>"001001001",
  32857=>"000000000",
  32858=>"001001000",
  32859=>"110110110",
  32860=>"001000000",
  32861=>"000000000",
  32862=>"000000000",
  32863=>"111111111",
  32864=>"001001000",
  32865=>"011011000",
  32866=>"010000000",
  32867=>"111000111",
  32868=>"110110110",
  32869=>"001010000",
  32870=>"000001001",
  32871=>"000000111",
  32872=>"111000000",
  32873=>"111111111",
  32874=>"010011110",
  32875=>"000000000",
  32876=>"000000000",
  32877=>"000000000",
  32878=>"000000001",
  32879=>"000001001",
  32880=>"010001011",
  32881=>"000011111",
  32882=>"000100100",
  32883=>"000000101",
  32884=>"011011000",
  32885=>"001011111",
  32886=>"010000000",
  32887=>"011111111",
  32888=>"000000011",
  32889=>"111101000",
  32890=>"000000000",
  32891=>"011001000",
  32892=>"001111111",
  32893=>"101101111",
  32894=>"000000000",
  32895=>"111111001",
  32896=>"101101101",
  32897=>"111000000",
  32898=>"111011001",
  32899=>"001011000",
  32900=>"000000000",
  32901=>"000000000",
  32902=>"111111111",
  32903=>"111010000",
  32904=>"000000010",
  32905=>"000001001",
  32906=>"111111111",
  32907=>"111111000",
  32908=>"000000000",
  32909=>"111100000",
  32910=>"111111011",
  32911=>"111110010",
  32912=>"100000000",
  32913=>"001000100",
  32914=>"000000001",
  32915=>"001110110",
  32916=>"110110100",
  32917=>"111000011",
  32918=>"111111111",
  32919=>"111111111",
  32920=>"000000000",
  32921=>"000000000",
  32922=>"000001111",
  32923=>"000000000",
  32924=>"001001000",
  32925=>"010000001",
  32926=>"001000000",
  32927=>"111111111",
  32928=>"000000101",
  32929=>"101100000",
  32930=>"111000100",
  32931=>"111111011",
  32932=>"000000011",
  32933=>"111111111",
  32934=>"111000000",
  32935=>"000100111",
  32936=>"111110110",
  32937=>"111001001",
  32938=>"000000000",
  32939=>"110000000",
  32940=>"101111111",
  32941=>"111000000",
  32942=>"111111111",
  32943=>"111111001",
  32944=>"010111001",
  32945=>"100111111",
  32946=>"001010000",
  32947=>"000000000",
  32948=>"011001011",
  32949=>"111111000",
  32950=>"101000001",
  32951=>"000000000",
  32952=>"110111111",
  32953=>"111111111",
  32954=>"001000101",
  32955=>"000110011",
  32956=>"110111001",
  32957=>"000000000",
  32958=>"000000000",
  32959=>"111111000",
  32960=>"000000000",
  32961=>"000000011",
  32962=>"010010010",
  32963=>"111111100",
  32964=>"111111100",
  32965=>"000000000",
  32966=>"000111111",
  32967=>"000000011",
  32968=>"111111111",
  32969=>"111001011",
  32970=>"000000000",
  32971=>"111100110",
  32972=>"000000111",
  32973=>"000110111",
  32974=>"000110111",
  32975=>"000000000",
  32976=>"111010000",
  32977=>"000000011",
  32978=>"001111111",
  32979=>"000000000",
  32980=>"111100000",
  32981=>"010111111",
  32982=>"000000100",
  32983=>"011001001",
  32984=>"000000111",
  32985=>"100111101",
  32986=>"000000000",
  32987=>"111111010",
  32988=>"111001001",
  32989=>"001001001",
  32990=>"000000100",
  32991=>"110010000",
  32992=>"000110110",
  32993=>"000000000",
  32994=>"111111111",
  32995=>"111111010",
  32996=>"011011011",
  32997=>"111110111",
  32998=>"000000001",
  32999=>"111110110",
  33000=>"111111010",
  33001=>"111111111",
  33002=>"101001111",
  33003=>"110111011",
  33004=>"111000000",
  33005=>"110100000",
  33006=>"111110111",
  33007=>"111111111",
  33008=>"101001000",
  33009=>"111111111",
  33010=>"000010011",
  33011=>"000000011",
  33012=>"111111111",
  33013=>"111110110",
  33014=>"001000111",
  33015=>"110110000",
  33016=>"111111111",
  33017=>"111110000",
  33018=>"000001000",
  33019=>"110110000",
  33020=>"000000100",
  33021=>"000110110",
  33022=>"001000000",
  33023=>"000000000",
  33024=>"001111010",
  33025=>"000010111",
  33026=>"000000000",
  33027=>"111111010",
  33028=>"001001000",
  33029=>"111111011",
  33030=>"011111111",
  33031=>"101111011",
  33032=>"001001000",
  33033=>"000000000",
  33034=>"000000111",
  33035=>"000000000",
  33036=>"000000000",
  33037=>"111000000",
  33038=>"001001111",
  33039=>"000110110",
  33040=>"000111001",
  33041=>"101101111",
  33042=>"001001001",
  33043=>"000000000",
  33044=>"000000000",
  33045=>"111111111",
  33046=>"001000000",
  33047=>"000101000",
  33048=>"000000000",
  33049=>"000000111",
  33050=>"100111011",
  33051=>"110111111",
  33052=>"001001010",
  33053=>"000000000",
  33054=>"000000000",
  33055=>"000000001",
  33056=>"111111111",
  33057=>"001011111",
  33058=>"110110111",
  33059=>"111111111",
  33060=>"111101001",
  33061=>"000000000",
  33062=>"111111011",
  33063=>"111111111",
  33064=>"000000000",
  33065=>"001001111",
  33066=>"000000000",
  33067=>"111111111",
  33068=>"111111111",
  33069=>"100100000",
  33070=>"111011000",
  33071=>"111111111",
  33072=>"000111111",
  33073=>"000000000",
  33074=>"000000001",
  33075=>"000000110",
  33076=>"000000110",
  33077=>"111000000",
  33078=>"110111110",
  33079=>"111100100",
  33080=>"000010000",
  33081=>"000000000",
  33082=>"000000000",
  33083=>"100110000",
  33084=>"111111111",
  33085=>"001111100",
  33086=>"111111111",
  33087=>"111111000",
  33088=>"001001000",
  33089=>"001000100",
  33090=>"010111010",
  33091=>"000000000",
  33092=>"000001000",
  33093=>"000011111",
  33094=>"000000000",
  33095=>"000010110",
  33096=>"000000101",
  33097=>"011000000",
  33098=>"100101101",
  33099=>"001101101",
  33100=>"111111111",
  33101=>"010000000",
  33102=>"110110000",
  33103=>"111100111",
  33104=>"101011011",
  33105=>"010011000",
  33106=>"000000110",
  33107=>"111000011",
  33108=>"110000000",
  33109=>"011011111",
  33110=>"110110000",
  33111=>"111111111",
  33112=>"111111111",
  33113=>"111111111",
  33114=>"111111001",
  33115=>"111111111",
  33116=>"111000000",
  33117=>"111111111",
  33118=>"001010000",
  33119=>"110110000",
  33120=>"111111111",
  33121=>"111001001",
  33122=>"001000100",
  33123=>"101111011",
  33124=>"000000000",
  33125=>"011001001",
  33126=>"011011001",
  33127=>"110110110",
  33128=>"001000000",
  33129=>"000000010",
  33130=>"111111001",
  33131=>"000011111",
  33132=>"000000000",
  33133=>"011111011",
  33134=>"001000000",
  33135=>"111111101",
  33136=>"111111111",
  33137=>"111001000",
  33138=>"111111011",
  33139=>"100100100",
  33140=>"000000000",
  33141=>"011011000",
  33142=>"111000001",
  33143=>"111110100",
  33144=>"000000001",
  33145=>"110111111",
  33146=>"111111011",
  33147=>"110100110",
  33148=>"111100111",
  33149=>"111111111",
  33150=>"011111010",
  33151=>"001111111",
  33152=>"010010011",
  33153=>"110110000",
  33154=>"111111111",
  33155=>"110001000",
  33156=>"111111111",
  33157=>"000110000",
  33158=>"011000001",
  33159=>"001101111",
  33160=>"110111111",
  33161=>"111100100",
  33162=>"000000011",
  33163=>"000110110",
  33164=>"111111111",
  33165=>"000110111",
  33166=>"110110110",
  33167=>"000000000",
  33168=>"000000000",
  33169=>"001001000",
  33170=>"100101001",
  33171=>"111111111",
  33172=>"000000011",
  33173=>"000010110",
  33174=>"000000000",
  33175=>"000000010",
  33176=>"000000100",
  33177=>"000000000",
  33178=>"101111111",
  33179=>"111000000",
  33180=>"111111111",
  33181=>"000000000",
  33182=>"111111100",
  33183=>"111111111",
  33184=>"001000111",
  33185=>"011011001",
  33186=>"000100100",
  33187=>"111111010",
  33188=>"100111000",
  33189=>"010010110",
  33190=>"111101111",
  33191=>"110111001",
  33192=>"011000000",
  33193=>"000010010",
  33194=>"000000000",
  33195=>"111111111",
  33196=>"100101001",
  33197=>"000000000",
  33198=>"111011111",
  33199=>"000110011",
  33200=>"000000000",
  33201=>"000000111",
  33202=>"000000000",
  33203=>"111111110",
  33204=>"111001001",
  33205=>"000000000",
  33206=>"010000010",
  33207=>"100000000",
  33208=>"000010010",
  33209=>"000000000",
  33210=>"001000000",
  33211=>"111111111",
  33212=>"110100110",
  33213=>"001000000",
  33214=>"000000000",
  33215=>"010010010",
  33216=>"100100000",
  33217=>"111100111",
  33218=>"111000000",
  33219=>"111111000",
  33220=>"000110111",
  33221=>"001001111",
  33222=>"110000000",
  33223=>"111110100",
  33224=>"000000000",
  33225=>"000011011",
  33226=>"100000111",
  33227=>"111111011",
  33228=>"000111111",
  33229=>"000000000",
  33230=>"100000000",
  33231=>"000000000",
  33232=>"000000100",
  33233=>"111111111",
  33234=>"000110111",
  33235=>"111000000",
  33236=>"110110110",
  33237=>"111111000",
  33238=>"000000000",
  33239=>"000011011",
  33240=>"000001001",
  33241=>"111011000",
  33242=>"000000001",
  33243=>"000000000",
  33244=>"101000000",
  33245=>"111111011",
  33246=>"001000111",
  33247=>"001010111",
  33248=>"000001101",
  33249=>"111111111",
  33250=>"000001000",
  33251=>"111111001",
  33252=>"001000000",
  33253=>"001101111",
  33254=>"111111100",
  33255=>"011001001",
  33256=>"110001001",
  33257=>"001001001",
  33258=>"010000000",
  33259=>"000000111",
  33260=>"000000000",
  33261=>"100100100",
  33262=>"000100111",
  33263=>"000000000",
  33264=>"111100110",
  33265=>"000111111",
  33266=>"000000000",
  33267=>"000000010",
  33268=>"100000000",
  33269=>"000000001",
  33270=>"111111111",
  33271=>"111110100",
  33272=>"000000010",
  33273=>"000000000",
  33274=>"000000000",
  33275=>"000000001",
  33276=>"111111111",
  33277=>"110001011",
  33278=>"000100001",
  33279=>"000000100",
  33280=>"000000000",
  33281=>"000110110",
  33282=>"111100111",
  33283=>"000100000",
  33284=>"000000001",
  33285=>"111000000",
  33286=>"011111011",
  33287=>"111111111",
  33288=>"111111111",
  33289=>"000001000",
  33290=>"111011001",
  33291=>"000000000",
  33292=>"111111111",
  33293=>"000000100",
  33294=>"111110111",
  33295=>"000000111",
  33296=>"100111011",
  33297=>"011000011",
  33298=>"000000111",
  33299=>"111010000",
  33300=>"000000000",
  33301=>"000001111",
  33302=>"000000111",
  33303=>"000101100",
  33304=>"111101000",
  33305=>"100000000",
  33306=>"001111111",
  33307=>"000000100",
  33308=>"000101111",
  33309=>"001001101",
  33310=>"110110100",
  33311=>"111111111",
  33312=>"011111111",
  33313=>"111110110",
  33314=>"101000000",
  33315=>"100001101",
  33316=>"111111010",
  33317=>"001000000",
  33318=>"001000000",
  33319=>"000000111",
  33320=>"000000000",
  33321=>"111111111",
  33322=>"111000000",
  33323=>"001001111",
  33324=>"000001111",
  33325=>"000000110",
  33326=>"110000000",
  33327=>"000000111",
  33328=>"111111111",
  33329=>"000000000",
  33330=>"110000000",
  33331=>"111111010",
  33332=>"010110010",
  33333=>"100110110",
  33334=>"000000000",
  33335=>"111111111",
  33336=>"011001111",
  33337=>"001001001",
  33338=>"001000000",
  33339=>"000000000",
  33340=>"111101111",
  33341=>"010000111",
  33342=>"000000111",
  33343=>"111000000",
  33344=>"110111110",
  33345=>"011000111",
  33346=>"111100110",
  33347=>"000000000",
  33348=>"000000100",
  33349=>"000000000",
  33350=>"001000000",
  33351=>"000000000",
  33352=>"001000000",
  33353=>"111000111",
  33354=>"000000111",
  33355=>"111111111",
  33356=>"111000000",
  33357=>"000000000",
  33358=>"111000111",
  33359=>"110100101",
  33360=>"000111111",
  33361=>"000000000",
  33362=>"111000000",
  33363=>"111111111",
  33364=>"111111110",
  33365=>"111011000",
  33366=>"111111111",
  33367=>"001001000",
  33368=>"000000000",
  33369=>"111000111",
  33370=>"101000000",
  33371=>"111000001",
  33372=>"000000000",
  33373=>"111011111",
  33374=>"011000001",
  33375=>"110111000",
  33376=>"000000111",
  33377=>"000111111",
  33378=>"000100000",
  33379=>"000000111",
  33380=>"111101000",
  33381=>"111111111",
  33382=>"000000001",
  33383=>"011000001",
  33384=>"111111110",
  33385=>"011001011",
  33386=>"000000111",
  33387=>"111000000",
  33388=>"101111111",
  33389=>"000000000",
  33390=>"000000000",
  33391=>"011011011",
  33392=>"111000001",
  33393=>"000000000",
  33394=>"010110010",
  33395=>"111111100",
  33396=>"111101111",
  33397=>"000000111",
  33398=>"000000000",
  33399=>"111110100",
  33400=>"000011111",
  33401=>"011001000",
  33402=>"111111000",
  33403=>"000000000",
  33404=>"000110111",
  33405=>"000110111",
  33406=>"111111011",
  33407=>"000011011",
  33408=>"111111111",
  33409=>"000000000",
  33410=>"000000111",
  33411=>"111111000",
  33412=>"000000000",
  33413=>"000001111",
  33414=>"111111110",
  33415=>"111100000",
  33416=>"111111111",
  33417=>"111111101",
  33418=>"000000000",
  33419=>"010000011",
  33420=>"110000000",
  33421=>"111111110",
  33422=>"111000000",
  33423=>"000000000",
  33424=>"100110111",
  33425=>"111110000",
  33426=>"100101101",
  33427=>"100100000",
  33428=>"011000000",
  33429=>"010110000",
  33430=>"000000111",
  33431=>"101000001",
  33432=>"101001111",
  33433=>"111111000",
  33434=>"111011000",
  33435=>"011000000",
  33436=>"111111111",
  33437=>"111111100",
  33438=>"000000111",
  33439=>"111111111",
  33440=>"011110000",
  33441=>"111111000",
  33442=>"111111111",
  33443=>"011011010",
  33444=>"111111000",
  33445=>"110110100",
  33446=>"111111111",
  33447=>"000001111",
  33448=>"111011111",
  33449=>"100101111",
  33450=>"111111000",
  33451=>"000100100",
  33452=>"110000101",
  33453=>"100100111",
  33454=>"111111000",
  33455=>"000000011",
  33456=>"111111011",
  33457=>"000100111",
  33458=>"111111011",
  33459=>"111111111",
  33460=>"011000110",
  33461=>"000011011",
  33462=>"000000000",
  33463=>"101000000",
  33464=>"000110110",
  33465=>"111111111",
  33466=>"111100101",
  33467=>"011001011",
  33468=>"001001000",
  33469=>"111111010",
  33470=>"011111110",
  33471=>"111111011",
  33472=>"111111111",
  33473=>"111111111",
  33474=>"111000000",
  33475=>"111000010",
  33476=>"111001111",
  33477=>"000000001",
  33478=>"110101111",
  33479=>"000000000",
  33480=>"000111111",
  33481=>"111101111",
  33482=>"000000000",
  33483=>"000111111",
  33484=>"111111100",
  33485=>"000110100",
  33486=>"110111111",
  33487=>"111110111",
  33488=>"111111100",
  33489=>"011000000",
  33490=>"000000000",
  33491=>"111011011",
  33492=>"101100111",
  33493=>"111111111",
  33494=>"000000000",
  33495=>"111011000",
  33496=>"110111001",
  33497=>"111001001",
  33498=>"111011001",
  33499=>"111111111",
  33500=>"111110110",
  33501=>"111011110",
  33502=>"111000000",
  33503=>"011011011",
  33504=>"000000000",
  33505=>"000001111",
  33506=>"010111111",
  33507=>"000000011",
  33508=>"000110111",
  33509=>"000000000",
  33510=>"000001011",
  33511=>"000000000",
  33512=>"111111100",
  33513=>"000000000",
  33514=>"000001111",
  33515=>"010100000",
  33516=>"000010100",
  33517=>"111111000",
  33518=>"101100111",
  33519=>"111111111",
  33520=>"100111111",
  33521=>"001001001",
  33522=>"000001011",
  33523=>"111111111",
  33524=>"111111111",
  33525=>"101101000",
  33526=>"110111000",
  33527=>"111011000",
  33528=>"111111000",
  33529=>"000111111",
  33530=>"001001111",
  33531=>"001000000",
  33532=>"110110110",
  33533=>"111111000",
  33534=>"101000000",
  33535=>"111111111",
  33536=>"000000001",
  33537=>"000000011",
  33538=>"111111011",
  33539=>"000000010",
  33540=>"111111111",
  33541=>"011111111",
  33542=>"000111100",
  33543=>"111010000",
  33544=>"001000000",
  33545=>"010000000",
  33546=>"101100000",
  33547=>"111111111",
  33548=>"011001011",
  33549=>"000000000",
  33550=>"111111111",
  33551=>"111000000",
  33552=>"111111001",
  33553=>"011111111",
  33554=>"011110110",
  33555=>"000000001",
  33556=>"011011000",
  33557=>"000010001",
  33558=>"100110101",
  33559=>"111000000",
  33560=>"011100000",
  33561=>"111111001",
  33562=>"000000000",
  33563=>"001000000",
  33564=>"111110000",
  33565=>"110000000",
  33566=>"010000000",
  33567=>"000011111",
  33568=>"101000000",
  33569=>"111111000",
  33570=>"001100000",
  33571=>"000110111",
  33572=>"001001111",
  33573=>"000000111",
  33574=>"011111110",
  33575=>"011001001",
  33576=>"101100100",
  33577=>"000000001",
  33578=>"011111011",
  33579=>"001000000",
  33580=>"010010011",
  33581=>"111101000",
  33582=>"111111000",
  33583=>"111000111",
  33584=>"000000000",
  33585=>"110000000",
  33586=>"111111111",
  33587=>"111100011",
  33588=>"010110000",
  33589=>"011000000",
  33590=>"000111111",
  33591=>"000000001",
  33592=>"000000000",
  33593=>"011000000",
  33594=>"111000000",
  33595=>"111111111",
  33596=>"000001001",
  33597=>"111101111",
  33598=>"111111111",
  33599=>"111011111",
  33600=>"101100111",
  33601=>"011001000",
  33602=>"111111000",
  33603=>"000000000",
  33604=>"111111111",
  33605=>"001000000",
  33606=>"000000001",
  33607=>"001001011",
  33608=>"111000000",
  33609=>"111011001",
  33610=>"111000101",
  33611=>"000000100",
  33612=>"111011000",
  33613=>"000000001",
  33614=>"111111111",
  33615=>"000000100",
  33616=>"001001001",
  33617=>"001111001",
  33618=>"111111111",
  33619=>"000000000",
  33620=>"100000000",
  33621=>"011111001",
  33622=>"000000011",
  33623=>"100100101",
  33624=>"001101100",
  33625=>"101000000",
  33626=>"000000100",
  33627=>"111111100",
  33628=>"111111011",
  33629=>"000000000",
  33630=>"111001101",
  33631=>"000011010",
  33632=>"000000000",
  33633=>"000101100",
  33634=>"111111111",
  33635=>"111001001",
  33636=>"000110110",
  33637=>"111110000",
  33638=>"000011111",
  33639=>"111011011",
  33640=>"101011111",
  33641=>"011111111",
  33642=>"111000000",
  33643=>"010000101",
  33644=>"111111000",
  33645=>"111111111",
  33646=>"111111111",
  33647=>"111001001",
  33648=>"001000000",
  33649=>"010011111",
  33650=>"110110111",
  33651=>"100110100",
  33652=>"110010010",
  33653=>"001100100",
  33654=>"111101111",
  33655=>"001111111",
  33656=>"100000000",
  33657=>"000000000",
  33658=>"111111000",
  33659=>"111111000",
  33660=>"111000101",
  33661=>"000111000",
  33662=>"000000000",
  33663=>"001111111",
  33664=>"011111111",
  33665=>"111111111",
  33666=>"100100100",
  33667=>"111101000",
  33668=>"100111111",
  33669=>"011110111",
  33670=>"111000110",
  33671=>"111111101",
  33672=>"111111100",
  33673=>"011011111",
  33674=>"011011000",
  33675=>"000001111",
  33676=>"111000000",
  33677=>"111111111",
  33678=>"111100000",
  33679=>"100110110",
  33680=>"011111111",
  33681=>"000111111",
  33682=>"001011011",
  33683=>"111110110",
  33684=>"111000000",
  33685=>"000011000",
  33686=>"111111000",
  33687=>"111111111",
  33688=>"111111111",
  33689=>"111111111",
  33690=>"000000001",
  33691=>"111111011",
  33692=>"111111111",
  33693=>"111111111",
  33694=>"000000000",
  33695=>"010111111",
  33696=>"000000111",
  33697=>"111111101",
  33698=>"111010000",
  33699=>"101000101",
  33700=>"111111111",
  33701=>"111000000",
  33702=>"000000000",
  33703=>"000000001",
  33704=>"001011000",
  33705=>"000000110",
  33706=>"111111111",
  33707=>"000010000",
  33708=>"111111111",
  33709=>"011111111",
  33710=>"101000111",
  33711=>"000100111",
  33712=>"000000111",
  33713=>"111001000",
  33714=>"010010010",
  33715=>"001000000",
  33716=>"011000000",
  33717=>"000000000",
  33718=>"000000000",
  33719=>"111011001",
  33720=>"111111111",
  33721=>"111111111",
  33722=>"000000000",
  33723=>"001011111",
  33724=>"000000000",
  33725=>"000000000",
  33726=>"111111111",
  33727=>"001001000",
  33728=>"111111111",
  33729=>"000000000",
  33730=>"111111111",
  33731=>"000111111",
  33732=>"011111000",
  33733=>"000000111",
  33734=>"000000000",
  33735=>"111010010",
  33736=>"111111111",
  33737=>"000000001",
  33738=>"110110111",
  33739=>"000000000",
  33740=>"000000111",
  33741=>"000100111",
  33742=>"000000000",
  33743=>"000000001",
  33744=>"110000100",
  33745=>"011000000",
  33746=>"111111011",
  33747=>"101100111",
  33748=>"000000000",
  33749=>"000000111",
  33750=>"011011111",
  33751=>"011010000",
  33752=>"111111100",
  33753=>"111111110",
  33754=>"111011111",
  33755=>"111111111",
  33756=>"110111001",
  33757=>"000000000",
  33758=>"111111110",
  33759=>"110000111",
  33760=>"011001111",
  33761=>"100000000",
  33762=>"000001111",
  33763=>"111110100",
  33764=>"111111111",
  33765=>"000000111",
  33766=>"000000100",
  33767=>"111011000",
  33768=>"000000000",
  33769=>"001001011",
  33770=>"000001001",
  33771=>"111111100",
  33772=>"100000000",
  33773=>"000001111",
  33774=>"111000000",
  33775=>"000000000",
  33776=>"010110111",
  33777=>"011111111",
  33778=>"111111000",
  33779=>"011011111",
  33780=>"110111111",
  33781=>"001000111",
  33782=>"111111000",
  33783=>"000111110",
  33784=>"011011001",
  33785=>"011001100",
  33786=>"110111000",
  33787=>"001011000",
  33788=>"000100100",
  33789=>"111001101",
  33790=>"111111111",
  33791=>"000000000",
  33792=>"011000000",
  33793=>"100000011",
  33794=>"101000000",
  33795=>"000110111",
  33796=>"000111001",
  33797=>"001011111",
  33798=>"111111110",
  33799=>"000000000",
  33800=>"111111000",
  33801=>"111000111",
  33802=>"000111101",
  33803=>"000000000",
  33804=>"000000111",
  33805=>"111111111",
  33806=>"100111111",
  33807=>"110010000",
  33808=>"000000000",
  33809=>"000000110",
  33810=>"111110000",
  33811=>"000000000",
  33812=>"111000001",
  33813=>"000000100",
  33814=>"111000000",
  33815=>"111011011",
  33816=>"111111110",
  33817=>"011111110",
  33818=>"111111111",
  33819=>"111111111",
  33820=>"000000101",
  33821=>"000000001",
  33822=>"010000000",
  33823=>"011111010",
  33824=>"100110110",
  33825=>"110110110",
  33826=>"111111100",
  33827=>"101011101",
  33828=>"001001001",
  33829=>"001000111",
  33830=>"110111111",
  33831=>"000000000",
  33832=>"001111111",
  33833=>"111111111",
  33834=>"100100111",
  33835=>"000111111",
  33836=>"000011111",
  33837=>"111011001",
  33838=>"100000001",
  33839=>"111011000",
  33840=>"000000000",
  33841=>"110111000",
  33842=>"110111111",
  33843=>"000000111",
  33844=>"000001000",
  33845=>"001000000",
  33846=>"000000111",
  33847=>"101100100",
  33848=>"001111111",
  33849=>"010111001",
  33850=>"111111111",
  33851=>"000111111",
  33852=>"001000000",
  33853=>"011111111",
  33854=>"110111100",
  33855=>"000000000",
  33856=>"000011111",
  33857=>"000000111",
  33858=>"111111100",
  33859=>"000000011",
  33860=>"011001000",
  33861=>"000100000",
  33862=>"111000010",
  33863=>"111111000",
  33864=>"000000001",
  33865=>"111111111",
  33866=>"111000000",
  33867=>"111111101",
  33868=>"100110110",
  33869=>"000010110",
  33870=>"111111110",
  33871=>"111111111",
  33872=>"101111001",
  33873=>"001111111",
  33874=>"000000111",
  33875=>"000000000",
  33876=>"000000010",
  33877=>"000000000",
  33878=>"100100011",
  33879=>"100111000",
  33880=>"111111010",
  33881=>"111101111",
  33882=>"111000000",
  33883=>"011011001",
  33884=>"000100111",
  33885=>"000000000",
  33886=>"011000001",
  33887=>"111011111",
  33888=>"011111010",
  33889=>"001001001",
  33890=>"000000011",
  33891=>"111111111",
  33892=>"110110000",
  33893=>"000000010",
  33894=>"001000001",
  33895=>"110110000",
  33896=>"111000001",
  33897=>"111001111",
  33898=>"111110111",
  33899=>"100110000",
  33900=>"011111011",
  33901=>"111111111",
  33902=>"000001111",
  33903=>"000000000",
  33904=>"010111111",
  33905=>"000000000",
  33906=>"000111111",
  33907=>"111001000",
  33908=>"000000000",
  33909=>"110111111",
  33910=>"111111000",
  33911=>"110111011",
  33912=>"001101111",
  33913=>"001000010",
  33914=>"000000000",
  33915=>"011001001",
  33916=>"000000000",
  33917=>"100100000",
  33918=>"000011010",
  33919=>"000000001",
  33920=>"111011000",
  33921=>"000000000",
  33922=>"000000011",
  33923=>"111110010",
  33924=>"001011111",
  33925=>"111101000",
  33926=>"000000100",
  33927=>"000111111",
  33928=>"111111010",
  33929=>"001001000",
  33930=>"111111111",
  33931=>"000100000",
  33932=>"001000000",
  33933=>"000000000",
  33934=>"110010000",
  33935=>"000000000",
  33936=>"000000000",
  33937=>"000000000",
  33938=>"011111011",
  33939=>"101000000",
  33940=>"000110111",
  33941=>"000000100",
  33942=>"111001000",
  33943=>"101001001",
  33944=>"001001111",
  33945=>"101101101",
  33946=>"111111111",
  33947=>"111111001",
  33948=>"111111110",
  33949=>"101000001",
  33950=>"000100011",
  33951=>"111111111",
  33952=>"101101101",
  33953=>"001000000",
  33954=>"111111111",
  33955=>"000110110",
  33956=>"001111110",
  33957=>"001001100",
  33958=>"101001101",
  33959=>"000100000",
  33960=>"010000000",
  33961=>"001001101",
  33962=>"000000000",
  33963=>"001001111",
  33964=>"001001000",
  33965=>"110111111",
  33966=>"000000101",
  33967=>"001000101",
  33968=>"000111111",
  33969=>"110111011",
  33970=>"111111110",
  33971=>"101101101",
  33972=>"111101001",
  33973=>"000010010",
  33974=>"000000000",
  33975=>"001100110",
  33976=>"000111111",
  33977=>"011111111",
  33978=>"101000000",
  33979=>"111111011",
  33980=>"000000000",
  33981=>"111111010",
  33982=>"111000000",
  33983=>"000000000",
  33984=>"010111010",
  33985=>"111111011",
  33986=>"000000010",
  33987=>"000000000",
  33988=>"111111111",
  33989=>"000000000",
  33990=>"110000000",
  33991=>"001000000",
  33992=>"000000000",
  33993=>"000100100",
  33994=>"001000001",
  33995=>"111011011",
  33996=>"001011011",
  33997=>"101111111",
  33998=>"000001111",
  33999=>"000011001",
  34000=>"100101110",
  34001=>"001000111",
  34002=>"000000001",
  34003=>"001011000",
  34004=>"001000000",
  34005=>"111000000",
  34006=>"111001001",
  34007=>"000000000",
  34008=>"011011000",
  34009=>"011111001",
  34010=>"011110000",
  34011=>"111000000",
  34012=>"110111111",
  34013=>"000000011",
  34014=>"111111111",
  34015=>"010110010",
  34016=>"111001101",
  34017=>"000011111",
  34018=>"000111111",
  34019=>"111111111",
  34020=>"000000000",
  34021=>"100110110",
  34022=>"001000111",
  34023=>"001000000",
  34024=>"000000111",
  34025=>"000000000",
  34026=>"000000000",
  34027=>"111000000",
  34028=>"000000111",
  34029=>"111111100",
  34030=>"101000000",
  34031=>"101100111",
  34032=>"111011000",
  34033=>"111111111",
  34034=>"111111111",
  34035=>"001000110",
  34036=>"111111111",
  34037=>"111100110",
  34038=>"000010110",
  34039=>"001000000",
  34040=>"111111111",
  34041=>"000000100",
  34042=>"000000010",
  34043=>"000111111",
  34044=>"011001011",
  34045=>"001011011",
  34046=>"111000000",
  34047=>"011111110",
  34048=>"001000101",
  34049=>"111111111",
  34050=>"000000011",
  34051=>"111111001",
  34052=>"111111111",
  34053=>"011111111",
  34054=>"000000000",
  34055=>"010111010",
  34056=>"111111111",
  34057=>"111000000",
  34058=>"001000100",
  34059=>"101101111",
  34060=>"110110110",
  34061=>"111111111",
  34062=>"110111010",
  34063=>"111001011",
  34064=>"000000000",
  34065=>"001111111",
  34066=>"000001111",
  34067=>"011011111",
  34068=>"000101100",
  34069=>"000111111",
  34070=>"001001000",
  34071=>"110110110",
  34072=>"001011011",
  34073=>"011011000",
  34074=>"000000000",
  34075=>"000000000",
  34076=>"001000000",
  34077=>"111110000",
  34078=>"001000000",
  34079=>"011111111",
  34080=>"111111100",
  34081=>"000000000",
  34082=>"100111111",
  34083=>"101110111",
  34084=>"100111111",
  34085=>"000000000",
  34086=>"100000000",
  34087=>"001111000",
  34088=>"100100100",
  34089=>"101000000",
  34090=>"010111010",
  34091=>"000000000",
  34092=>"000111110",
  34093=>"010110000",
  34094=>"000001000",
  34095=>"000000000",
  34096=>"000000111",
  34097=>"110111001",
  34098=>"100000000",
  34099=>"011000000",
  34100=>"000111111",
  34101=>"000001011",
  34102=>"001010100",
  34103=>"000000000",
  34104=>"111010010",
  34105=>"111001000",
  34106=>"000000000",
  34107=>"110011111",
  34108=>"000001000",
  34109=>"000000110",
  34110=>"111111100",
  34111=>"101000001",
  34112=>"000000110",
  34113=>"000001101",
  34114=>"000000101",
  34115=>"001001000",
  34116=>"111111110",
  34117=>"111111000",
  34118=>"000111111",
  34119=>"000001101",
  34120=>"000000010",
  34121=>"111101111",
  34122=>"000000101",
  34123=>"111000000",
  34124=>"111100000",
  34125=>"111000000",
  34126=>"000100001",
  34127=>"001011011",
  34128=>"000010110",
  34129=>"001000111",
  34130=>"100110111",
  34131=>"000000111",
  34132=>"000000000",
  34133=>"011000000",
  34134=>"000000000",
  34135=>"000000001",
  34136=>"111111110",
  34137=>"000000000",
  34138=>"110010000",
  34139=>"111000000",
  34140=>"000000001",
  34141=>"000000000",
  34142=>"001000000",
  34143=>"110110000",
  34144=>"000000000",
  34145=>"000000000",
  34146=>"001000000",
  34147=>"001001001",
  34148=>"110111111",
  34149=>"111111001",
  34150=>"111000111",
  34151=>"000000001",
  34152=>"111110100",
  34153=>"000110111",
  34154=>"011001111",
  34155=>"000000000",
  34156=>"111110110",
  34157=>"000001111",
  34158=>"111110000",
  34159=>"101001011",
  34160=>"101000001",
  34161=>"111110100",
  34162=>"000000000",
  34163=>"010010000",
  34164=>"110110010",
  34165=>"001111111",
  34166=>"000000000",
  34167=>"011001111",
  34168=>"111111001",
  34169=>"010001001",
  34170=>"111100101",
  34171=>"111101100",
  34172=>"101101111",
  34173=>"000000001",
  34174=>"000001011",
  34175=>"111011001",
  34176=>"011010000",
  34177=>"101000000",
  34178=>"000000011",
  34179=>"111111111",
  34180=>"000000111",
  34181=>"111111111",
  34182=>"111000000",
  34183=>"101000101",
  34184=>"000000000",
  34185=>"000010011",
  34186=>"001001001",
  34187=>"011111111",
  34188=>"000100111",
  34189=>"100111111",
  34190=>"011111010",
  34191=>"010000000",
  34192=>"000000000",
  34193=>"111101111",
  34194=>"111111101",
  34195=>"000100100",
  34196=>"000000000",
  34197=>"010010000",
  34198=>"000101001",
  34199=>"111110100",
  34200=>"001101111",
  34201=>"111110110",
  34202=>"111111010",
  34203=>"110110000",
  34204=>"111111111",
  34205=>"000001111",
  34206=>"101101000",
  34207=>"111111000",
  34208=>"111001000",
  34209=>"100100000",
  34210=>"000011000",
  34211=>"111101111",
  34212=>"111111111",
  34213=>"101001000",
  34214=>"101101101",
  34215=>"111111111",
  34216=>"101001001",
  34217=>"000000011",
  34218=>"000111111",
  34219=>"001000000",
  34220=>"000000111",
  34221=>"111111111",
  34222=>"101000111",
  34223=>"000000000",
  34224=>"000000111",
  34225=>"010111000",
  34226=>"000000000",
  34227=>"010011010",
  34228=>"000000100",
  34229=>"010010000",
  34230=>"001111111",
  34231=>"101101000",
  34232=>"001000000",
  34233=>"000000111",
  34234=>"110110111",
  34235=>"000000111",
  34236=>"000111111",
  34237=>"001011000",
  34238=>"111001011",
  34239=>"000101111",
  34240=>"011011001",
  34241=>"000000000",
  34242=>"011000010",
  34243=>"000000000",
  34244=>"111111010",
  34245=>"000100100",
  34246=>"010000000",
  34247=>"000001000",
  34248=>"011110110",
  34249=>"000000111",
  34250=>"111111011",
  34251=>"111111111",
  34252=>"000000000",
  34253=>"000000111",
  34254=>"101000000",
  34255=>"001000001",
  34256=>"101000000",
  34257=>"100011000",
  34258=>"011011101",
  34259=>"000010000",
  34260=>"000000000",
  34261=>"100000000",
  34262=>"011001000",
  34263=>"000110110",
  34264=>"101101101",
  34265=>"111111100",
  34266=>"000111111",
  34267=>"111110000",
  34268=>"001100110",
  34269=>"111000000",
  34270=>"011000001",
  34271=>"100100000",
  34272=>"000000000",
  34273=>"111111000",
  34274=>"000000000",
  34275=>"111111001",
  34276=>"000000010",
  34277=>"001000001",
  34278=>"000001111",
  34279=>"011000000",
  34280=>"100111111",
  34281=>"111111111",
  34282=>"000000110",
  34283=>"001001101",
  34284=>"000001111",
  34285=>"111001000",
  34286=>"000001001",
  34287=>"000000110",
  34288=>"000000000",
  34289=>"110111111",
  34290=>"000000000",
  34291=>"100101101",
  34292=>"111111011",
  34293=>"000000000",
  34294=>"000000010",
  34295=>"011001001",
  34296=>"111111000",
  34297=>"000010010",
  34298=>"111101000",
  34299=>"000000000",
  34300=>"001000000",
  34301=>"101000000",
  34302=>"111011000",
  34303=>"101000000",
  34304=>"000000000",
  34305=>"111111111",
  34306=>"011011111",
  34307=>"001011001",
  34308=>"111010011",
  34309=>"011001111",
  34310=>"010000000",
  34311=>"111111111",
  34312=>"001000100",
  34313=>"000111111",
  34314=>"111101001",
  34315=>"000110111",
  34316=>"000100110",
  34317=>"000000000",
  34318=>"000110111",
  34319=>"000000111",
  34320=>"111111011",
  34321=>"000111111",
  34322=>"000000000",
  34323=>"111111001",
  34324=>"000101111",
  34325=>"001001111",
  34326=>"001000001",
  34327=>"111111101",
  34328=>"000000000",
  34329=>"100111111",
  34330=>"001011010",
  34331=>"001000010",
  34332=>"000000000",
  34333=>"101111101",
  34334=>"111111111",
  34335=>"001000010",
  34336=>"010110110",
  34337=>"001101001",
  34338=>"000000001",
  34339=>"011111101",
  34340=>"110111110",
  34341=>"111110000",
  34342=>"001001100",
  34343=>"011001001",
  34344=>"001000100",
  34345=>"000000000",
  34346=>"000100101",
  34347=>"000000101",
  34348=>"101001000",
  34349=>"111111010",
  34350=>"000000000",
  34351=>"111111011",
  34352=>"000000001",
  34353=>"000111111",
  34354=>"110100000",
  34355=>"111111010",
  34356=>"111111001",
  34357=>"000001011",
  34358=>"000000000",
  34359=>"111111011",
  34360=>"101111011",
  34361=>"000000101",
  34362=>"000110110",
  34363=>"101111111",
  34364=>"000000001",
  34365=>"111000000",
  34366=>"011001111",
  34367=>"001001111",
  34368=>"000000000",
  34369=>"001111111",
  34370=>"101111100",
  34371=>"011001111",
  34372=>"110110110",
  34373=>"011111111",
  34374=>"000000111",
  34375=>"100101111",
  34376=>"111111111",
  34377=>"000000000",
  34378=>"000000100",
  34379=>"000000101",
  34380=>"000000000",
  34381=>"111010000",
  34382=>"111011011",
  34383=>"110100110",
  34384=>"000000000",
  34385=>"110110111",
  34386=>"100110000",
  34387=>"110110000",
  34388=>"000111110",
  34389=>"000001111",
  34390=>"000000101",
  34391=>"001000000",
  34392=>"001111010",
  34393=>"000000001",
  34394=>"000100000",
  34395=>"001001111",
  34396=>"100000000",
  34397=>"001000110",
  34398=>"000001001",
  34399=>"000000000",
  34400=>"000011000",
  34401=>"001111111",
  34402=>"000000000",
  34403=>"000111111",
  34404=>"001001001",
  34405=>"000000111",
  34406=>"011001000",
  34407=>"000001000",
  34408=>"000111111",
  34409=>"100000001",
  34410=>"100111000",
  34411=>"000010110",
  34412=>"000000001",
  34413=>"110111111",
  34414=>"000001001",
  34415=>"000111111",
  34416=>"110100000",
  34417=>"000101111",
  34418=>"001001111",
  34419=>"010000111",
  34420=>"001000111",
  34421=>"110111110",
  34422=>"000000000",
  34423=>"001001111",
  34424=>"000000000",
  34425=>"000000000",
  34426=>"111111111",
  34427=>"111000000",
  34428=>"111111111",
  34429=>"000010000",
  34430=>"100101111",
  34431=>"010111000",
  34432=>"111101101",
  34433=>"011000000",
  34434=>"111111111",
  34435=>"000100011",
  34436=>"000000000",
  34437=>"000000111",
  34438=>"001001001",
  34439=>"111001111",
  34440=>"000000011",
  34441=>"000000001",
  34442=>"000000001",
  34443=>"110110000",
  34444=>"000101001",
  34445=>"001001101",
  34446=>"001001100",
  34447=>"110111100",
  34448=>"111101100",
  34449=>"100110110",
  34450=>"100100000",
  34451=>"111111111",
  34452=>"000000000",
  34453=>"111111111",
  34454=>"101000101",
  34455=>"000000111",
  34456=>"001000000",
  34457=>"000100111",
  34458=>"011000000",
  34459=>"000000000",
  34460=>"001000000",
  34461=>"000000101",
  34462=>"010000111",
  34463=>"000110111",
  34464=>"111111111",
  34465=>"011111111",
  34466=>"111111111",
  34467=>"111111010",
  34468=>"111011111",
  34469=>"111111111",
  34470=>"000000000",
  34471=>"001111111",
  34472=>"000001011",
  34473=>"001000111",
  34474=>"000000000",
  34475=>"111111011",
  34476=>"111110000",
  34477=>"000110111",
  34478=>"111111111",
  34479=>"011111111",
  34480=>"111110000",
  34481=>"000001000",
  34482=>"111111000",
  34483=>"000000000",
  34484=>"000000011",
  34485=>"001001001",
  34486=>"000001111",
  34487=>"000000000",
  34488=>"001111111",
  34489=>"111111101",
  34490=>"111001000",
  34491=>"011011011",
  34492=>"000000000",
  34493=>"111111111",
  34494=>"111111100",
  34495=>"000000001",
  34496=>"111000000",
  34497=>"000001000",
  34498=>"011000000",
  34499=>"111111101",
  34500=>"111101111",
  34501=>"001000000",
  34502=>"000001010",
  34503=>"010100000",
  34504=>"000000000",
  34505=>"000000000",
  34506=>"110100110",
  34507=>"101000100",
  34508=>"000000110",
  34509=>"000000101",
  34510=>"111110111",
  34511=>"000000110",
  34512=>"111011000",
  34513=>"000000100",
  34514=>"000000000",
  34515=>"100000000",
  34516=>"001000000",
  34517=>"111111000",
  34518=>"000111001",
  34519=>"111111010",
  34520=>"000101111",
  34521=>"111110000",
  34522=>"011111111",
  34523=>"100111101",
  34524=>"111111000",
  34525=>"001000111",
  34526=>"000001000",
  34527=>"111111000",
  34528=>"000001011",
  34529=>"000000110",
  34530=>"111100000",
  34531=>"010000101",
  34532=>"000001011",
  34533=>"000000000",
  34534=>"111111000",
  34535=>"101111111",
  34536=>"000111111",
  34537=>"111111000",
  34538=>"110111110",
  34539=>"001000111",
  34540=>"111111111",
  34541=>"000000000",
  34542=>"100100111",
  34543=>"000100111",
  34544=>"111011001",
  34545=>"001011100",
  34546=>"000011011",
  34547=>"010000000",
  34548=>"000000011",
  34549=>"000010011",
  34550=>"000000011",
  34551=>"000010010",
  34552=>"000111111",
  34553=>"000000000",
  34554=>"000110111",
  34555=>"111111011",
  34556=>"001100111",
  34557=>"011111000",
  34558=>"101001001",
  34559=>"100101010",
  34560=>"000000000",
  34561=>"001001001",
  34562=>"000000000",
  34563=>"111000000",
  34564=>"111111000",
  34565=>"001000000",
  34566=>"000100100",
  34567=>"000000101",
  34568=>"111100000",
  34569=>"111110000",
  34570=>"001000111",
  34571=>"111111010",
  34572=>"001000001",
  34573=>"011001000",
  34574=>"000111111",
  34575=>"001000000",
  34576=>"000011011",
  34577=>"001000111",
  34578=>"001001101",
  34579=>"100111111",
  34580=>"111011011",
  34581=>"000100110",
  34582=>"110111000",
  34583=>"000001001",
  34584=>"011010000",
  34585=>"000110001",
  34586=>"001001111",
  34587=>"111110000",
  34588=>"001001000",
  34589=>"001101111",
  34590=>"000000000",
  34591=>"000000111",
  34592=>"111011000",
  34593=>"000000000",
  34594=>"010000000",
  34595=>"001000111",
  34596=>"111110100",
  34597=>"000101111",
  34598=>"111111111",
  34599=>"000000011",
  34600=>"000000110",
  34601=>"000000000",
  34602=>"011011011",
  34603=>"000000111",
  34604=>"000000000",
  34605=>"011011011",
  34606=>"000000110",
  34607=>"000000010",
  34608=>"111111111",
  34609=>"111111000",
  34610=>"001000001",
  34611=>"001000000",
  34612=>"000000000",
  34613=>"001000000",
  34614=>"000000000",
  34615=>"111011101",
  34616=>"011011000",
  34617=>"011010111",
  34618=>"000000001",
  34619=>"101101110",
  34620=>"100110001",
  34621=>"011111111",
  34622=>"101001111",
  34623=>"011000000",
  34624=>"000001111",
  34625=>"000000110",
  34626=>"111001101",
  34627=>"001001111",
  34628=>"001001111",
  34629=>"001001111",
  34630=>"010001001",
  34631=>"100110111",
  34632=>"000000001",
  34633=>"000000100",
  34634=>"000000000",
  34635=>"100100000",
  34636=>"011011000",
  34637=>"011111111",
  34638=>"000000000",
  34639=>"000100100",
  34640=>"111100110",
  34641=>"111111011",
  34642=>"111111000",
  34643=>"000000111",
  34644=>"010110100",
  34645=>"001011011",
  34646=>"111111010",
  34647=>"000000001",
  34648=>"001011011",
  34649=>"101000001",
  34650=>"001001111",
  34651=>"000000100",
  34652=>"000000000",
  34653=>"000000111",
  34654=>"000000000",
  34655=>"001001111",
  34656=>"011111111",
  34657=>"100001011",
  34658=>"101101100",
  34659=>"001000001",
  34660=>"101001000",
  34661=>"111010000",
  34662=>"000000111",
  34663=>"110110110",
  34664=>"001011000",
  34665=>"000000000",
  34666=>"110100110",
  34667=>"000110110",
  34668=>"110110000",
  34669=>"111111101",
  34670=>"000100110",
  34671=>"001111111",
  34672=>"111111110",
  34673=>"111101111",
  34674=>"011000001",
  34675=>"001111110",
  34676=>"000000000",
  34677=>"001101000",
  34678=>"110110111",
  34679=>"110000100",
  34680=>"000000000",
  34681=>"111101111",
  34682=>"001000011",
  34683=>"000000000",
  34684=>"100100111",
  34685=>"001000001",
  34686=>"000011111",
  34687=>"111111111",
  34688=>"011111111",
  34689=>"000000111",
  34690=>"111111111",
  34691=>"111001101",
  34692=>"101111111",
  34693=>"000001111",
  34694=>"010001010",
  34695=>"111111111",
  34696=>"000000010",
  34697=>"111000001",
  34698=>"100000000",
  34699=>"000110111",
  34700=>"000000000",
  34701=>"000000000",
  34702=>"001101111",
  34703=>"000000111",
  34704=>"000000000",
  34705=>"000111111",
  34706=>"001001001",
  34707=>"111111111",
  34708=>"000000000",
  34709=>"000000000",
  34710=>"110110110",
  34711=>"111111011",
  34712=>"001001111",
  34713=>"000000100",
  34714=>"111000000",
  34715=>"111110111",
  34716=>"010111011",
  34717=>"100110111",
  34718=>"101000000",
  34719=>"111111111",
  34720=>"000000000",
  34721=>"111110011",
  34722=>"111000001",
  34723=>"001111111",
  34724=>"111111110",
  34725=>"110111111",
  34726=>"001001111",
  34727=>"100000001",
  34728=>"100000000",
  34729=>"000000111",
  34730=>"000111111",
  34731=>"110110110",
  34732=>"000000111",
  34733=>"000000111",
  34734=>"000000000",
  34735=>"110110110",
  34736=>"000000000",
  34737=>"101001111",
  34738=>"110110110",
  34739=>"000000101",
  34740=>"111111111",
  34741=>"111110101",
  34742=>"000000001",
  34743=>"110110100",
  34744=>"111111111",
  34745=>"111111110",
  34746=>"111111101",
  34747=>"000000111",
  34748=>"111101000",
  34749=>"000001111",
  34750=>"011011011",
  34751=>"000101101",
  34752=>"000000101",
  34753=>"100111111",
  34754=>"000000000",
  34755=>"010111100",
  34756=>"000000000",
  34757=>"000000000",
  34758=>"000001101",
  34759=>"111111101",
  34760=>"001001000",
  34761=>"000000010",
  34762=>"000000111",
  34763=>"111111111",
  34764=>"111111011",
  34765=>"001011001",
  34766=>"000000000",
  34767=>"010000000",
  34768=>"100110000",
  34769=>"110110001",
  34770=>"000111111",
  34771=>"111111111",
  34772=>"000100100",
  34773=>"000110110",
  34774=>"011011111",
  34775=>"001101001",
  34776=>"000000000",
  34777=>"111000000",
  34778=>"111101110",
  34779=>"111110101",
  34780=>"111101111",
  34781=>"011001001",
  34782=>"111111001",
  34783=>"111000000",
  34784=>"111000000",
  34785=>"110111111",
  34786=>"110110100",
  34787=>"110111111",
  34788=>"111111111",
  34789=>"011010000",
  34790=>"110110110",
  34791=>"000000111",
  34792=>"011010111",
  34793=>"001001100",
  34794=>"011011000",
  34795=>"110110100",
  34796=>"000100101",
  34797=>"001000110",
  34798=>"011111111",
  34799=>"000011111",
  34800=>"000100000",
  34801=>"000000000",
  34802=>"101100000",
  34803=>"100100000",
  34804=>"000000000",
  34805=>"000000011",
  34806=>"111111101",
  34807=>"001000000",
  34808=>"011111111",
  34809=>"011000000",
  34810=>"000000000",
  34811=>"000000001",
  34812=>"000111011",
  34813=>"001000100",
  34814=>"001000100",
  34815=>"111001001",
  34816=>"111111111",
  34817=>"000110110",
  34818=>"101111111",
  34819=>"001000000",
  34820=>"110000000",
  34821=>"011011001",
  34822=>"010000000",
  34823=>"111001111",
  34824=>"011010111",
  34825=>"000000001",
  34826=>"000110110",
  34827=>"110110110",
  34828=>"100000000",
  34829=>"111111001",
  34830=>"000000000",
  34831=>"000011101",
  34832=>"000000111",
  34833=>"011011111",
  34834=>"011010111",
  34835=>"101000000",
  34836=>"000000001",
  34837=>"100000100",
  34838=>"101001000",
  34839=>"110000000",
  34840=>"111111111",
  34841=>"000000001",
  34842=>"010011000",
  34843=>"111111111",
  34844=>"000011111",
  34845=>"000000000",
  34846=>"101101101",
  34847=>"100000000",
  34848=>"111110100",
  34849=>"001111000",
  34850=>"000000110",
  34851=>"011111111",
  34852=>"000000000",
  34853=>"100001001",
  34854=>"111110000",
  34855=>"000010010",
  34856=>"111111110",
  34857=>"000000000",
  34858=>"111011111",
  34859=>"000000100",
  34860=>"001111111",
  34861=>"100110000",
  34862=>"000001000",
  34863=>"000100000",
  34864=>"110100100",
  34865=>"011111011",
  34866=>"110100100",
  34867=>"000000000",
  34868=>"111111101",
  34869=>"010011011",
  34870=>"010111100",
  34871=>"011111000",
  34872=>"111000110",
  34873=>"000000000",
  34874=>"000000000",
  34875=>"111000000",
  34876=>"101111111",
  34877=>"111110110",
  34878=>"010110110",
  34879=>"000000000",
  34880=>"110111111",
  34881=>"000000111",
  34882=>"010000000",
  34883=>"000000000",
  34884=>"000000000",
  34885=>"001000000",
  34886=>"110011001",
  34887=>"100100110",
  34888=>"010000011",
  34889=>"000000111",
  34890=>"111111111",
  34891=>"111111111",
  34892=>"000000011",
  34893=>"111100111",
  34894=>"101000000",
  34895=>"110100000",
  34896=>"111111110",
  34897=>"000001011",
  34898=>"000010000",
  34899=>"010000000",
  34900=>"000000000",
  34901=>"110000000",
  34902=>"010110111",
  34903=>"011001000",
  34904=>"111111111",
  34905=>"111111000",
  34906=>"000111111",
  34907=>"010000100",
  34908=>"001000000",
  34909=>"000000110",
  34910=>"000000110",
  34911=>"000110000",
  34912=>"111001000",
  34913=>"000111001",
  34914=>"001001101",
  34915=>"100000111",
  34916=>"111111000",
  34917=>"001000000",
  34918=>"110110010",
  34919=>"000000000",
  34920=>"111111111",
  34921=>"100000000",
  34922=>"111111001",
  34923=>"000001001",
  34924=>"111011011",
  34925=>"111111111",
  34926=>"001001111",
  34927=>"000000000",
  34928=>"000000000",
  34929=>"101101111",
  34930=>"000011001",
  34931=>"111100111",
  34932=>"001000000",
  34933=>"000000000",
  34934=>"000000000",
  34935=>"011001111",
  34936=>"011111111",
  34937=>"111111111",
  34938=>"000000111",
  34939=>"000100110",
  34940=>"111011010",
  34941=>"011111101",
  34942=>"011111111",
  34943=>"000101111",
  34944=>"000000000",
  34945=>"000000000",
  34946=>"000111111",
  34947=>"111110111",
  34948=>"111111000",
  34949=>"000000100",
  34950=>"101111001",
  34951=>"000000110",
  34952=>"000000000",
  34953=>"000100100",
  34954=>"001001001",
  34955=>"111111111",
  34956=>"001000000",
  34957=>"000000000",
  34958=>"001001001",
  34959=>"000000000",
  34960=>"000000000",
  34961=>"111111111",
  34962=>"000000010",
  34963=>"000110000",
  34964=>"111111110",
  34965=>"111110111",
  34966=>"000000000",
  34967=>"000000000",
  34968=>"000000000",
  34969=>"000000000",
  34970=>"000000000",
  34971=>"000000000",
  34972=>"000000000",
  34973=>"111111111",
  34974=>"111111111",
  34975=>"000000100",
  34976=>"111111111",
  34977=>"111111000",
  34978=>"000000000",
  34979=>"000000000",
  34980=>"111000101",
  34981=>"111000000",
  34982=>"111111110",
  34983=>"110100000",
  34984=>"110011110",
  34985=>"000000000",
  34986=>"100000000",
  34987=>"111111011",
  34988=>"000000000",
  34989=>"100100110",
  34990=>"110110100",
  34991=>"000011111",
  34992=>"001000000",
  34993=>"001000110",
  34994=>"111111111",
  34995=>"111010010",
  34996=>"000101111",
  34997=>"000010000",
  34998=>"111111000",
  34999=>"111111110",
  35000=>"111110111",
  35001=>"010000111",
  35002=>"000001101",
  35003=>"010000000",
  35004=>"000000000",
  35005=>"000100111",
  35006=>"111111011",
  35007=>"000000000",
  35008=>"000000000",
  35009=>"000000100",
  35010=>"010000000",
  35011=>"000000000",
  35012=>"000000000",
  35013=>"000100111",
  35014=>"111011000",
  35015=>"000100110",
  35016=>"111111111",
  35017=>"111000000",
  35018=>"111111111",
  35019=>"111111111",
  35020=>"111110000",
  35021=>"000000000",
  35022=>"111111011",
  35023=>"000000000",
  35024=>"001011011",
  35025=>"000000001",
  35026=>"000000000",
  35027=>"000000000",
  35028=>"100110000",
  35029=>"111101001",
  35030=>"000000000",
  35031=>"101001000",
  35032=>"010011111",
  35033=>"101000000",
  35034=>"111111110",
  35035=>"111101111",
  35036=>"100000000",
  35037=>"101111001",
  35038=>"110010111",
  35039=>"101000000",
  35040=>"111111111",
  35041=>"111111011",
  35042=>"000000000",
  35043=>"000000111",
  35044=>"000000000",
  35045=>"000000000",
  35046=>"111111111",
  35047=>"111001001",
  35048=>"000110110",
  35049=>"100000000",
  35050=>"110110111",
  35051=>"000000000",
  35052=>"000000111",
  35053=>"110010010",
  35054=>"111111110",
  35055=>"111111111",
  35056=>"000000100",
  35057=>"001000000",
  35058=>"001000000",
  35059=>"110111101",
  35060=>"000000111",
  35061=>"111111111",
  35062=>"001000000",
  35063=>"111011111",
  35064=>"110111111",
  35065=>"000000000",
  35066=>"000000111",
  35067=>"111111111",
  35068=>"100111111",
  35069=>"110000111",
  35070=>"110110000",
  35071=>"000001000",
  35072=>"000000000",
  35073=>"111101111",
  35074=>"100110100",
  35075=>"000100111",
  35076=>"000000111",
  35077=>"101110110",
  35078=>"111111111",
  35079=>"000001101",
  35080=>"111111111",
  35081=>"001100100",
  35082=>"000000000",
  35083=>"111111111",
  35084=>"111011011",
  35085=>"000011011",
  35086=>"110100100",
  35087=>"000000011",
  35088=>"011111110",
  35089=>"000001111",
  35090=>"001001011",
  35091=>"000001001",
  35092=>"110110000",
  35093=>"011011011",
  35094=>"110110110",
  35095=>"111111111",
  35096=>"111111111",
  35097=>"011000000",
  35098=>"101111111",
  35099=>"111110010",
  35100=>"111111111",
  35101=>"000000011",
  35102=>"011011000",
  35103=>"111111111",
  35104=>"110010000",
  35105=>"111110000",
  35106=>"000000001",
  35107=>"000000111",
  35108=>"111000010",
  35109=>"011111111",
  35110=>"000000000",
  35111=>"101101001",
  35112=>"000000000",
  35113=>"000000011",
  35114=>"111111110",
  35115=>"111111010",
  35116=>"001011111",
  35117=>"001001001",
  35118=>"100001001",
  35119=>"011000000",
  35120=>"011001111",
  35121=>"011001111",
  35122=>"011000000",
  35123=>"111111011",
  35124=>"111000000",
  35125=>"111111111",
  35126=>"111001100",
  35127=>"111110100",
  35128=>"000010000",
  35129=>"001111111",
  35130=>"111111111",
  35131=>"000000011",
  35132=>"001001111",
  35133=>"000111111",
  35134=>"010000000",
  35135=>"111111111",
  35136=>"000000000",
  35137=>"110111111",
  35138=>"111100111",
  35139=>"000011111",
  35140=>"111111111",
  35141=>"110100000",
  35142=>"000000000",
  35143=>"000000001",
  35144=>"111111111",
  35145=>"000000000",
  35146=>"000111111",
  35147=>"100000000",
  35148=>"000000100",
  35149=>"000000111",
  35150=>"000000000",
  35151=>"000000111",
  35152=>"111011001",
  35153=>"000000000",
  35154=>"000000000",
  35155=>"000000000",
  35156=>"111111111",
  35157=>"000000000",
  35158=>"111111000",
  35159=>"000000000",
  35160=>"111111111",
  35161=>"111111111",
  35162=>"100111110",
  35163=>"000110100",
  35164=>"100001000",
  35165=>"000000000",
  35166=>"000000000",
  35167=>"111100100",
  35168=>"101101111",
  35169=>"000011011",
  35170=>"001000000",
  35171=>"111111101",
  35172=>"001001000",
  35173=>"111111111",
  35174=>"101000110",
  35175=>"011111101",
  35176=>"000000000",
  35177=>"000111111",
  35178=>"110000000",
  35179=>"100111111",
  35180=>"000000000",
  35181=>"111010000",
  35182=>"000000000",
  35183=>"000000000",
  35184=>"111111111",
  35185=>"111111010",
  35186=>"101101001",
  35187=>"000011011",
  35188=>"000000111",
  35189=>"111100100",
  35190=>"111111111",
  35191=>"110111111",
  35192=>"000000000",
  35193=>"111111111",
  35194=>"111111111",
  35195=>"111111111",
  35196=>"010000010",
  35197=>"000000100",
  35198=>"000000000",
  35199=>"000000001",
  35200=>"110110100",
  35201=>"111011111",
  35202=>"100000001",
  35203=>"111111111",
  35204=>"100000000",
  35205=>"111111011",
  35206=>"000100100",
  35207=>"111110110",
  35208=>"111100000",
  35209=>"000000100",
  35210=>"111101001",
  35211=>"001011001",
  35212=>"100100000",
  35213=>"001001001",
  35214=>"111111111",
  35215=>"010111000",
  35216=>"111000000",
  35217=>"000000000",
  35218=>"000000000",
  35219=>"111100111",
  35220=>"111000000",
  35221=>"000000110",
  35222=>"110000001",
  35223=>"110110000",
  35224=>"110110110",
  35225=>"001110110",
  35226=>"111011111",
  35227=>"010000100",
  35228=>"000000000",
  35229=>"111111111",
  35230=>"000000000",
  35231=>"000000000",
  35232=>"110010111",
  35233=>"100100110",
  35234=>"111111111",
  35235=>"000000000",
  35236=>"001001001",
  35237=>"111111011",
  35238=>"000000111",
  35239=>"000000011",
  35240=>"000000000",
  35241=>"111001111",
  35242=>"000000000",
  35243=>"000000000",
  35244=>"000000000",
  35245=>"111000000",
  35246=>"110110000",
  35247=>"111111111",
  35248=>"111111110",
  35249=>"000000000",
  35250=>"111111111",
  35251=>"111000111",
  35252=>"000000000",
  35253=>"010000000",
  35254=>"101101101",
  35255=>"100111010",
  35256=>"001000110",
  35257=>"000000000",
  35258=>"100100110",
  35259=>"110111011",
  35260=>"100010110",
  35261=>"111111000",
  35262=>"100100000",
  35263=>"110110111",
  35264=>"100110111",
  35265=>"000011011",
  35266=>"111111111",
  35267=>"011010010",
  35268=>"111111111",
  35269=>"110000000",
  35270=>"000000000",
  35271=>"111111000",
  35272=>"000000111",
  35273=>"000011011",
  35274=>"111001100",
  35275=>"111111101",
  35276=>"111111111",
  35277=>"000000001",
  35278=>"111100110",
  35279=>"111000000",
  35280=>"001111111",
  35281=>"000000000",
  35282=>"001010000",
  35283=>"000000111",
  35284=>"110000000",
  35285=>"100000111",
  35286=>"111111111",
  35287=>"000000010",
  35288=>"000000110",
  35289=>"111011011",
  35290=>"111010011",
  35291=>"000000000",
  35292=>"011111111",
  35293=>"000000000",
  35294=>"010000011",
  35295=>"110110111",
  35296=>"111011111",
  35297=>"111111111",
  35298=>"000000000",
  35299=>"111111000",
  35300=>"111111111",
  35301=>"111111111",
  35302=>"111111111",
  35303=>"111111111",
  35304=>"111111001",
  35305=>"111000001",
  35306=>"111111110",
  35307=>"111100000",
  35308=>"000111111",
  35309=>"011111001",
  35310=>"001011011",
  35311=>"001000000",
  35312=>"111111111",
  35313=>"000111111",
  35314=>"001001111",
  35315=>"000000000",
  35316=>"100111111",
  35317=>"000000000",
  35318=>"111111000",
  35319=>"001011000",
  35320=>"000000000",
  35321=>"010011011",
  35322=>"110110000",
  35323=>"000111111",
  35324=>"111111111",
  35325=>"110110110",
  35326=>"101100110",
  35327=>"111111111",
  35328=>"000000000",
  35329=>"111110111",
  35330=>"000000000",
  35331=>"101000100",
  35332=>"000111111",
  35333=>"000000001",
  35334=>"000000010",
  35335=>"001001111",
  35336=>"111111000",
  35337=>"100000110",
  35338=>"111111011",
  35339=>"000100111",
  35340=>"100110110",
  35341=>"010111111",
  35342=>"110111011",
  35343=>"000000100",
  35344=>"101111000",
  35345=>"000000000",
  35346=>"111100000",
  35347=>"000000000",
  35348=>"110000101",
  35349=>"000000001",
  35350=>"111111000",
  35351=>"010111011",
  35352=>"000110110",
  35353=>"001001000",
  35354=>"111111001",
  35355=>"111001000",
  35356=>"001011111",
  35357=>"001101000",
  35358=>"111110110",
  35359=>"001000111",
  35360=>"000111111",
  35361=>"000000000",
  35362=>"111111010",
  35363=>"110110111",
  35364=>"111111111",
  35365=>"000000000",
  35366=>"111110000",
  35367=>"111111000",
  35368=>"100000100",
  35369=>"100100100",
  35370=>"000000000",
  35371=>"111100000",
  35372=>"000000000",
  35373=>"111111000",
  35374=>"111111111",
  35375=>"000111111",
  35376=>"000100110",
  35377=>"000000100",
  35378=>"000000000",
  35379=>"000011111",
  35380=>"111111111",
  35381=>"100000000",
  35382=>"111111111",
  35383=>"000110111",
  35384=>"000000000",
  35385=>"100111001",
  35386=>"000000000",
  35387=>"000000000",
  35388=>"000000100",
  35389=>"100000011",
  35390=>"100100001",
  35391=>"000000000",
  35392=>"111111111",
  35393=>"000001000",
  35394=>"111111111",
  35395=>"100000001",
  35396=>"100110110",
  35397=>"100100100",
  35398=>"010110111",
  35399=>"111010000",
  35400=>"000000001",
  35401=>"111111010",
  35402=>"000000000",
  35403=>"011000101",
  35404=>"000000100",
  35405=>"001000000",
  35406=>"111000000",
  35407=>"111111111",
  35408=>"111111000",
  35409=>"101000001",
  35410=>"000000011",
  35411=>"111111001",
  35412=>"111111111",
  35413=>"000000100",
  35414=>"000111110",
  35415=>"001000000",
  35416=>"100110010",
  35417=>"101000000",
  35418=>"111111111",
  35419=>"111001000",
  35420=>"111100000",
  35421=>"001000100",
  35422=>"000010000",
  35423=>"111111111",
  35424=>"001000001",
  35425=>"000111111",
  35426=>"110111000",
  35427=>"100000000",
  35428=>"000000000",
  35429=>"000000001",
  35430=>"000000111",
  35431=>"111111110",
  35432=>"111111000",
  35433=>"111111000",
  35434=>"111011111",
  35435=>"000000001",
  35436=>"110110000",
  35437=>"000000100",
  35438=>"000000000",
  35439=>"010000000",
  35440=>"000000000",
  35441=>"000110011",
  35442=>"111111111",
  35443=>"110110001",
  35444=>"011111111",
  35445=>"110110000",
  35446=>"101101001",
  35447=>"000110000",
  35448=>"111110110",
  35449=>"000010100",
  35450=>"000110000",
  35451=>"000000000",
  35452=>"111110111",
  35453=>"000000101",
  35454=>"110111000",
  35455=>"000000001",
  35456=>"000000000",
  35457=>"110110100",
  35458=>"111111111",
  35459=>"001000000",
  35460=>"111111011",
  35461=>"111111001",
  35462=>"110111111",
  35463=>"100000000",
  35464=>"000000001",
  35465=>"000110100",
  35466=>"110000000",
  35467=>"000000000",
  35468=>"110011011",
  35469=>"111111110",
  35470=>"110110111",
  35471=>"000110110",
  35472=>"000000000",
  35473=>"011000000",
  35474=>"000100101",
  35475=>"000000111",
  35476=>"001100110",
  35477=>"111110000",
  35478=>"010000000",
  35479=>"111101111",
  35480=>"000000001",
  35481=>"111111111",
  35482=>"111111111",
  35483=>"111000000",
  35484=>"110000001",
  35485=>"111110000",
  35486=>"000111111",
  35487=>"000000000",
  35488=>"011001111",
  35489=>"101111011",
  35490=>"000011111",
  35491=>"111111110",
  35492=>"000000100",
  35493=>"100000000",
  35494=>"100101111",
  35495=>"111011111",
  35496=>"111111111",
  35497=>"000000000",
  35498=>"001000000",
  35499=>"000000000",
  35500=>"110111111",
  35501=>"101101111",
  35502=>"110111011",
  35503=>"111111001",
  35504=>"010000000",
  35505=>"111111110",
  35506=>"111111011",
  35507=>"111111000",
  35508=>"110111110",
  35509=>"111000111",
  35510=>"000000000",
  35511=>"000000000",
  35512=>"110110000",
  35513=>"110111111",
  35514=>"001000001",
  35515=>"111111111",
  35516=>"100000000",
  35517=>"000000000",
  35518=>"111111111",
  35519=>"000000000",
  35520=>"010000000",
  35521=>"000000111",
  35522=>"000000111",
  35523=>"111000000",
  35524=>"000000000",
  35525=>"111111111",
  35526=>"010110111",
  35527=>"111111111",
  35528=>"000000000",
  35529=>"000000111",
  35530=>"001100100",
  35531=>"000000000",
  35532=>"010000111",
  35533=>"001011111",
  35534=>"000100101",
  35535=>"000000110",
  35536=>"100000000",
  35537=>"000000000",
  35538=>"111000000",
  35539=>"111111100",
  35540=>"000000100",
  35541=>"000000000",
  35542=>"000000001",
  35543=>"111111011",
  35544=>"000000001",
  35545=>"000000000",
  35546=>"111111111",
  35547=>"011110111",
  35548=>"000100010",
  35549=>"000011011",
  35550=>"111000000",
  35551=>"010010111",
  35552=>"111111001",
  35553=>"000000000",
  35554=>"000000000",
  35555=>"000000001",
  35556=>"000000100",
  35557=>"111000100",
  35558=>"111110110",
  35559=>"100001000",
  35560=>"111111000",
  35561=>"111111111",
  35562=>"111110110",
  35563=>"000000000",
  35564=>"101000000",
  35565=>"000000000",
  35566=>"000000000",
  35567=>"000010111",
  35568=>"010111111",
  35569=>"111111110",
  35570=>"111111111",
  35571=>"111111111",
  35572=>"000111111",
  35573=>"011111111",
  35574=>"110000000",
  35575=>"111111111",
  35576=>"111111110",
  35577=>"111110111",
  35578=>"000100111",
  35579=>"111111111",
  35580=>"111011111",
  35581=>"000001000",
  35582=>"101000000",
  35583=>"110000000",
  35584=>"000000000",
  35585=>"000011111",
  35586=>"000000111",
  35587=>"111111010",
  35588=>"000111111",
  35589=>"000000111",
  35590=>"000000000",
  35591=>"000001011",
  35592=>"111111011",
  35593=>"000000000",
  35594=>"100000111",
  35595=>"000001100",
  35596=>"101000000",
  35597=>"000000000",
  35598=>"000011011",
  35599=>"111111111",
  35600=>"111111111",
  35601=>"000000000",
  35602=>"111001000",
  35603=>"001000000",
  35604=>"000001111",
  35605=>"011111111",
  35606=>"110110110",
  35607=>"111111000",
  35608=>"111111111",
  35609=>"000000000",
  35610=>"111000000",
  35611=>"000000000",
  35612=>"000000000",
  35613=>"010001111",
  35614=>"000000000",
  35615=>"000000000",
  35616=>"000000000",
  35617=>"100001001",
  35618=>"000000000",
  35619=>"110100110",
  35620=>"100110111",
  35621=>"110100111",
  35622=>"001111010",
  35623=>"001001011",
  35624=>"011001000",
  35625=>"111000000",
  35626=>"111001001",
  35627=>"111111111",
  35628=>"111111111",
  35629=>"001011011",
  35630=>"111000111",
  35631=>"111111100",
  35632=>"000000000",
  35633=>"111001101",
  35634=>"111111111",
  35635=>"010010000",
  35636=>"000000111",
  35637=>"111111000",
  35638=>"011001011",
  35639=>"000000001",
  35640=>"111001001",
  35641=>"100000111",
  35642=>"111111111",
  35643=>"111111001",
  35644=>"111110100",
  35645=>"111111000",
  35646=>"110111010",
  35647=>"110110111",
  35648=>"000001001",
  35649=>"000100111",
  35650=>"111011011",
  35651=>"001011000",
  35652=>"100101111",
  35653=>"111011000",
  35654=>"000000110",
  35655=>"111111000",
  35656=>"000000101",
  35657=>"000111111",
  35658=>"111000111",
  35659=>"100001111",
  35660=>"001000000",
  35661=>"000000000",
  35662=>"000000000",
  35663=>"100010000",
  35664=>"111111111",
  35665=>"000000110",
  35666=>"110100111",
  35667=>"001111111",
  35668=>"000000100",
  35669=>"011011001",
  35670=>"001111111",
  35671=>"000100100",
  35672=>"111010100",
  35673=>"111111111",
  35674=>"111110000",
  35675=>"110110111",
  35676=>"100000001",
  35677=>"000000000",
  35678=>"111101001",
  35679=>"000000000",
  35680=>"111010000",
  35681=>"001000111",
  35682=>"110111011",
  35683=>"000111111",
  35684=>"000000011",
  35685=>"000000000",
  35686=>"111101000",
  35687=>"111111110",
  35688=>"000000111",
  35689=>"000000111",
  35690=>"001000001",
  35691=>"001000000",
  35692=>"000000000",
  35693=>"001010111",
  35694=>"000000000",
  35695=>"011000011",
  35696=>"110110111",
  35697=>"000000000",
  35698=>"111111110",
  35699=>"001001011",
  35700=>"001000000",
  35701=>"000110000",
  35702=>"001000000",
  35703=>"111011000",
  35704=>"000000111",
  35705=>"111000111",
  35706=>"110111111",
  35707=>"000110100",
  35708=>"011111111",
  35709=>"000000000",
  35710=>"100110000",
  35711=>"000000000",
  35712=>"111110110",
  35713=>"111110110",
  35714=>"001000000",
  35715=>"000000000",
  35716=>"100111111",
  35717=>"111111110",
  35718=>"001001111",
  35719=>"000000000",
  35720=>"001011111",
  35721=>"111111111",
  35722=>"000000101",
  35723=>"000010111",
  35724=>"111101111",
  35725=>"100011011",
  35726=>"110000000",
  35727=>"000000111",
  35728=>"000000000",
  35729=>"110011011",
  35730=>"110000001",
  35731=>"111111010",
  35732=>"011011111",
  35733=>"010111010",
  35734=>"100000000",
  35735=>"000000000",
  35736=>"111111111",
  35737=>"000000111",
  35738=>"110111111",
  35739=>"000000000",
  35740=>"101111111",
  35741=>"111000111",
  35742=>"001101101",
  35743=>"111011001",
  35744=>"111000100",
  35745=>"111000000",
  35746=>"000000110",
  35747=>"000000101",
  35748=>"110111111",
  35749=>"111111001",
  35750=>"001001111",
  35751=>"111000110",
  35752=>"111111111",
  35753=>"000000100",
  35754=>"111111111",
  35755=>"101000000",
  35756=>"000100111",
  35757=>"000011110",
  35758=>"000000111",
  35759=>"000000000",
  35760=>"000100000",
  35761=>"001001101",
  35762=>"111111110",
  35763=>"000000000",
  35764=>"000100101",
  35765=>"111111111",
  35766=>"000110110",
  35767=>"111111111",
  35768=>"000000111",
  35769=>"100101111",
  35770=>"010110111",
  35771=>"011111111",
  35772=>"101111011",
  35773=>"100111111",
  35774=>"111100000",
  35775=>"100111110",
  35776=>"110110000",
  35777=>"000000011",
  35778=>"111111111",
  35779=>"000000111",
  35780=>"110110111",
  35781=>"000000000",
  35782=>"100100111",
  35783=>"111001001",
  35784=>"011010111",
  35785=>"111010111",
  35786=>"111110111",
  35787=>"000100111",
  35788=>"110110000",
  35789=>"000000000",
  35790=>"000000011",
  35791=>"000000000",
  35792=>"000011011",
  35793=>"111111111",
  35794=>"000010110",
  35795=>"111001111",
  35796=>"111111110",
  35797=>"111010000",
  35798=>"000000001",
  35799=>"111111011",
  35800=>"100000100",
  35801=>"000000000",
  35802=>"111111111",
  35803=>"000000000",
  35804=>"111111111",
  35805=>"111001001",
  35806=>"111000111",
  35807=>"001001000",
  35808=>"111111111",
  35809=>"000000000",
  35810=>"000101111",
  35811=>"100000010",
  35812=>"000110111",
  35813=>"100000000",
  35814=>"111000000",
  35815=>"000000000",
  35816=>"010011111",
  35817=>"000111110",
  35818=>"000011111",
  35819=>"000000000",
  35820=>"010000000",
  35821=>"000001001",
  35822=>"000000101",
  35823=>"000000110",
  35824=>"000100100",
  35825=>"110110110",
  35826=>"111101111",
  35827=>"000000010",
  35828=>"111101011",
  35829=>"001000111",
  35830=>"100111100",
  35831=>"000101110",
  35832=>"000011000",
  35833=>"000101111",
  35834=>"110000000",
  35835=>"000110111",
  35836=>"011011110",
  35837=>"111110111",
  35838=>"000000111",
  35839=>"000000111",
  35840=>"001011111",
  35841=>"111000110",
  35842=>"101000000",
  35843=>"001000111",
  35844=>"110110000",
  35845=>"011011111",
  35846=>"001001011",
  35847=>"111111111",
  35848=>"001001000",
  35849=>"111011001",
  35850=>"000000000",
  35851=>"111111111",
  35852=>"011011011",
  35853=>"100000000",
  35854=>"111111111",
  35855=>"000011011",
  35856=>"010000000",
  35857=>"111111111",
  35858=>"000000111",
  35859=>"000000000",
  35860=>"100000000",
  35861=>"000000000",
  35862=>"111111001",
  35863=>"111111001",
  35864=>"111111111",
  35865=>"111110111",
  35866=>"000000100",
  35867=>"111111001",
  35868=>"010000000",
  35869=>"111111111",
  35870=>"010011001",
  35871=>"000000000",
  35872=>"110111000",
  35873=>"001001001",
  35874=>"111111111",
  35875=>"111101000",
  35876=>"011001111",
  35877=>"111111110",
  35878=>"000011111",
  35879=>"110110111",
  35880=>"111001010",
  35881=>"111111001",
  35882=>"011011000",
  35883=>"110000100",
  35884=>"100000000",
  35885=>"111001111",
  35886=>"000000000",
  35887=>"111000000",
  35888=>"001001011",
  35889=>"001000011",
  35890=>"000011011",
  35891=>"000011110",
  35892=>"000110111",
  35893=>"111000001",
  35894=>"000011011",
  35895=>"001001001",
  35896=>"111111000",
  35897=>"011000000",
  35898=>"000000000",
  35899=>"000000001",
  35900=>"101101111",
  35901=>"010011111",
  35902=>"011011111",
  35903=>"111111111",
  35904=>"000000101",
  35905=>"000000000",
  35906=>"001011001",
  35907=>"000110000",
  35908=>"110110110",
  35909=>"011000000",
  35910=>"000000000",
  35911=>"000000000",
  35912=>"000001011",
  35913=>"000000000",
  35914=>"111111111",
  35915=>"000000000",
  35916=>"000000000",
  35917=>"010111111",
  35918=>"000000011",
  35919=>"000001111",
  35920=>"000011000",
  35921=>"000000000",
  35922=>"100000000",
  35923=>"010000111",
  35924=>"000000101",
  35925=>"000000000",
  35926=>"000000000",
  35927=>"110000000",
  35928=>"000000000",
  35929=>"111101101",
  35930=>"000000110",
  35931=>"000001111",
  35932=>"110111111",
  35933=>"111111111",
  35934=>"000110110",
  35935=>"100100100",
  35936=>"000000000",
  35937=>"000000000",
  35938=>"111000000",
  35939=>"000000000",
  35940=>"111000000",
  35941=>"000000000",
  35942=>"111111111",
  35943=>"000000000",
  35944=>"000000000",
  35945=>"010010000",
  35946=>"111111111",
  35947=>"000000000",
  35948=>"001111000",
  35949=>"111111111",
  35950=>"111011000",
  35951=>"111111110",
  35952=>"000000000",
  35953=>"110010000",
  35954=>"000000111",
  35955=>"111100100",
  35956=>"111111111",
  35957=>"000001111",
  35958=>"001100100",
  35959=>"000000000",
  35960=>"000000000",
  35961=>"000000000",
  35962=>"110111101",
  35963=>"110111010",
  35964=>"000001110",
  35965=>"000000000",
  35966=>"000000000",
  35967=>"000000000",
  35968=>"000000000",
  35969=>"110000001",
  35970=>"000000001",
  35971=>"000000100",
  35972=>"000000000",
  35973=>"111101101",
  35974=>"111111000",
  35975=>"110111000",
  35976=>"000000000",
  35977=>"101001001",
  35978=>"000000000",
  35979=>"000000000",
  35980=>"000000001",
  35981=>"001001111",
  35982=>"111001001",
  35983=>"010000000",
  35984=>"110110111",
  35985=>"000000101",
  35986=>"000000011",
  35987=>"001111111",
  35988=>"000000000",
  35989=>"000000111",
  35990=>"001000001",
  35991=>"111111111",
  35992=>"001111111",
  35993=>"000000000",
  35994=>"111111111",
  35995=>"000000000",
  35996=>"101111110",
  35997=>"110110000",
  35998=>"010111111",
  35999=>"000001111",
  36000=>"000000111",
  36001=>"111001000",
  36002=>"111111111",
  36003=>"000000000",
  36004=>"110000011",
  36005=>"000011101",
  36006=>"011111011",
  36007=>"001011111",
  36008=>"111111111",
  36009=>"000000000",
  36010=>"111111111",
  36011=>"111000011",
  36012=>"110110000",
  36013=>"100100100",
  36014=>"100111111",
  36015=>"001001001",
  36016=>"001001000",
  36017=>"001001100",
  36018=>"010010011",
  36019=>"111110000",
  36020=>"111011000",
  36021=>"000000011",
  36022=>"000000111",
  36023=>"111111111",
  36024=>"000011010",
  36025=>"000111111",
  36026=>"111000000",
  36027=>"111111011",
  36028=>"000000000",
  36029=>"111111011",
  36030=>"111111111",
  36031=>"001000000",
  36032=>"111111101",
  36033=>"011000000",
  36034=>"000000000",
  36035=>"111111111",
  36036=>"000000000",
  36037=>"000000000",
  36038=>"000011001",
  36039=>"111111111",
  36040=>"111101111",
  36041=>"000000000",
  36042=>"000000111",
  36043=>"110010100",
  36044=>"000000100",
  36045=>"110110100",
  36046=>"101110111",
  36047=>"111110000",
  36048=>"111111001",
  36049=>"000001000",
  36050=>"000000000",
  36051=>"000100000",
  36052=>"111111110",
  36053=>"111111011",
  36054=>"111111000",
  36055=>"011111010",
  36056=>"111111111",
  36057=>"000000000",
  36058=>"000000000",
  36059=>"011111111",
  36060=>"011000100",
  36061=>"000000100",
  36062=>"111111111",
  36063=>"000001101",
  36064=>"001111111",
  36065=>"111100101",
  36066=>"101000100",
  36067=>"000101110",
  36068=>"110111111",
  36069=>"110100000",
  36070=>"000000111",
  36071=>"110111001",
  36072=>"111101000",
  36073=>"111011111",
  36074=>"111111111",
  36075=>"110110000",
  36076=>"000000000",
  36077=>"111111111",
  36078=>"111010000",
  36079=>"000101000",
  36080=>"000001000",
  36081=>"000001000",
  36082=>"111100100",
  36083=>"111111111",
  36084=>"111111101",
  36085=>"011001111",
  36086=>"100100100",
  36087=>"111111001",
  36088=>"101101101",
  36089=>"000000000",
  36090=>"001001111",
  36091=>"000000111",
  36092=>"011001001",
  36093=>"000000000",
  36094=>"111110110",
  36095=>"111111101",
  36096=>"111111101",
  36097=>"011111011",
  36098=>"111111110",
  36099=>"011011011",
  36100=>"000111100",
  36101=>"001010010",
  36102=>"000000011",
  36103=>"000000011",
  36104=>"000000000",
  36105=>"001111100",
  36106=>"001001101",
  36107=>"011111111",
  36108=>"111111111",
  36109=>"000000001",
  36110=>"000000000",
  36111=>"000000000",
  36112=>"000000001",
  36113=>"111111111",
  36114=>"000000000",
  36115=>"000000001",
  36116=>"001001000",
  36117=>"111001000",
  36118=>"000000000",
  36119=>"000011011",
  36120=>"111111110",
  36121=>"111100110",
  36122=>"001001000",
  36123=>"000000101",
  36124=>"000000000",
  36125=>"111100110",
  36126=>"011001000",
  36127=>"100110110",
  36128=>"001000111",
  36129=>"100111110",
  36130=>"000000110",
  36131=>"010000000",
  36132=>"100100100",
  36133=>"001011000",
  36134=>"111111111",
  36135=>"110111111",
  36136=>"111111111",
  36137=>"011000000",
  36138=>"000001000",
  36139=>"000011111",
  36140=>"001001100",
  36141=>"010011000",
  36142=>"000000000",
  36143=>"101101001",
  36144=>"001001001",
  36145=>"111111111",
  36146=>"011001100",
  36147=>"111111111",
  36148=>"000000111",
  36149=>"111111111",
  36150=>"101101101",
  36151=>"111101000",
  36152=>"001000001",
  36153=>"111010111",
  36154=>"111111111",
  36155=>"000000100",
  36156=>"111111111",
  36157=>"111101111",
  36158=>"110110011",
  36159=>"011011001",
  36160=>"111000000",
  36161=>"111111111",
  36162=>"001000111",
  36163=>"000100000",
  36164=>"111111101",
  36165=>"000101101",
  36166=>"110100110",
  36167=>"001001111",
  36168=>"000000011",
  36169=>"111000000",
  36170=>"000110110",
  36171=>"111110100",
  36172=>"000001111",
  36173=>"101000111",
  36174=>"000000111",
  36175=>"000000100",
  36176=>"000001001",
  36177=>"011000011",
  36178=>"100100100",
  36179=>"111111000",
  36180=>"110111111",
  36181=>"111000000",
  36182=>"001001000",
  36183=>"111111000",
  36184=>"000000000",
  36185=>"101111000",
  36186=>"001111111",
  36187=>"100111110",
  36188=>"000000010",
  36189=>"000000010",
  36190=>"000000111",
  36191=>"111111011",
  36192=>"000111011",
  36193=>"111111111",
  36194=>"001101100",
  36195=>"101001001",
  36196=>"111011110",
  36197=>"111011111",
  36198=>"001000111",
  36199=>"011011001",
  36200=>"000000001",
  36201=>"000000000",
  36202=>"011000000",
  36203=>"000001001",
  36204=>"000011111",
  36205=>"010000011",
  36206=>"000010111",
  36207=>"001001001",
  36208=>"000000000",
  36209=>"001111011",
  36210=>"101000000",
  36211=>"111111111",
  36212=>"111111111",
  36213=>"111111001",
  36214=>"000000000",
  36215=>"001001000",
  36216=>"111100010",
  36217=>"110100100",
  36218=>"000000000",
  36219=>"111111111",
  36220=>"100000000",
  36221=>"110000000",
  36222=>"111111111",
  36223=>"100000000",
  36224=>"000001001",
  36225=>"111101001",
  36226=>"111111010",
  36227=>"000000000",
  36228=>"011110000",
  36229=>"111011111",
  36230=>"000000000",
  36231=>"000000000",
  36232=>"000000000",
  36233=>"110000000",
  36234=>"101101001",
  36235=>"111111011",
  36236=>"111100111",
  36237=>"000000110",
  36238=>"001001111",
  36239=>"111011000",
  36240=>"000000000",
  36241=>"111111111",
  36242=>"111111111",
  36243=>"000001011",
  36244=>"011000000",
  36245=>"000000000",
  36246=>"110000111",
  36247=>"110100101",
  36248=>"000101001",
  36249=>"001001111",
  36250=>"111111110",
  36251=>"000000000",
  36252=>"001101000",
  36253=>"110010000",
  36254=>"111111111",
  36255=>"000000000",
  36256=>"100100100",
  36257=>"000101101",
  36258=>"010000000",
  36259=>"111111111",
  36260=>"011001000",
  36261=>"000100110",
  36262=>"111111111",
  36263=>"000111111",
  36264=>"000000000",
  36265=>"000010011",
  36266=>"111001100",
  36267=>"111111111",
  36268=>"000000000",
  36269=>"000000001",
  36270=>"000000000",
  36271=>"010010000",
  36272=>"000000000",
  36273=>"001000000",
  36274=>"000000100",
  36275=>"000111111",
  36276=>"111111111",
  36277=>"000011000",
  36278=>"111111011",
  36279=>"001000000",
  36280=>"011000000",
  36281=>"000000000",
  36282=>"111111100",
  36283=>"000001000",
  36284=>"000011111",
  36285=>"111111001",
  36286=>"001100011",
  36287=>"110000010",
  36288=>"111111111",
  36289=>"000111010",
  36290=>"111111111",
  36291=>"000000001",
  36292=>"000010100",
  36293=>"111100100",
  36294=>"111111101",
  36295=>"011111111",
  36296=>"000001000",
  36297=>"000000000",
  36298=>"000000000",
  36299=>"111111111",
  36300=>"000000000",
  36301=>"111111001",
  36302=>"001111111",
  36303=>"000000101",
  36304=>"000110111",
  36305=>"111111011",
  36306=>"111111111",
  36307=>"000110000",
  36308=>"000111111",
  36309=>"111111111",
  36310=>"000000111",
  36311=>"000000100",
  36312=>"011011000",
  36313=>"000111110",
  36314=>"111111000",
  36315=>"101101100",
  36316=>"000001000",
  36317=>"000011000",
  36318=>"111000000",
  36319=>"110110000",
  36320=>"100111111",
  36321=>"000011111",
  36322=>"111111111",
  36323=>"010000011",
  36324=>"000000000",
  36325=>"100000010",
  36326=>"111100100",
  36327=>"111101100",
  36328=>"011011010",
  36329=>"111111111",
  36330=>"111111111",
  36331=>"000000001",
  36332=>"101111010",
  36333=>"001001011",
  36334=>"111111111",
  36335=>"011011111",
  36336=>"111111111",
  36337=>"100000000",
  36338=>"001000010",
  36339=>"000000010",
  36340=>"000101111",
  36341=>"001000101",
  36342=>"000000101",
  36343=>"101101101",
  36344=>"001001111",
  36345=>"001000000",
  36346=>"000000111",
  36347=>"100110111",
  36348=>"000000100",
  36349=>"001001001",
  36350=>"111111111",
  36351=>"000000000",
  36352=>"111110111",
  36353=>"111111001",
  36354=>"111010000",
  36355=>"110111111",
  36356=>"111111001",
  36357=>"000000000",
  36358=>"111101001",
  36359=>"010111111",
  36360=>"001000001",
  36361=>"110111111",
  36362=>"111111111",
  36363=>"101001000",
  36364=>"111000000",
  36365=>"011111111",
  36366=>"100000001",
  36367=>"100100000",
  36368=>"110100000",
  36369=>"111111010",
  36370=>"000001011",
  36371=>"111111011",
  36372=>"000000100",
  36373=>"111101111",
  36374=>"011000011",
  36375=>"000100100",
  36376=>"111111111",
  36377=>"110110101",
  36378=>"111111111",
  36379=>"111111000",
  36380=>"001000000",
  36381=>"110101100",
  36382=>"000100110",
  36383=>"111111111",
  36384=>"001100111",
  36385=>"111111000",
  36386=>"000000000",
  36387=>"001001001",
  36388=>"111110100",
  36389=>"111111111",
  36390=>"100000000",
  36391=>"000000000",
  36392=>"111111111",
  36393=>"111111111",
  36394=>"001001001",
  36395=>"111100000",
  36396=>"100100000",
  36397=>"000000000",
  36398=>"000000000",
  36399=>"111111001",
  36400=>"111111011",
  36401=>"100100001",
  36402=>"001001000",
  36403=>"100111111",
  36404=>"110010000",
  36405=>"111111110",
  36406=>"101000000",
  36407=>"111111111",
  36408=>"000100100",
  36409=>"000011111",
  36410=>"100000111",
  36411=>"011111111",
  36412=>"000000000",
  36413=>"000010111",
  36414=>"111111111",
  36415=>"001000000",
  36416=>"000000101",
  36417=>"111111110",
  36418=>"111111000",
  36419=>"000001001",
  36420=>"000010010",
  36421=>"001001111",
  36422=>"000000000",
  36423=>"111000000",
  36424=>"011001001",
  36425=>"111111111",
  36426=>"001011111",
  36427=>"001001111",
  36428=>"000000011",
  36429=>"100111111",
  36430=>"110000000",
  36431=>"000000000",
  36432=>"000000000",
  36433=>"000000110",
  36434=>"111111111",
  36435=>"111110110",
  36436=>"000000000",
  36437=>"110000000",
  36438=>"111011001",
  36439=>"001011111",
  36440=>"110111111",
  36441=>"101111000",
  36442=>"000000110",
  36443=>"111111111",
  36444=>"010110111",
  36445=>"000000001",
  36446=>"111111111",
  36447=>"000011011",
  36448=>"010110000",
  36449=>"001001101",
  36450=>"011001001",
  36451=>"100110111",
  36452=>"110110011",
  36453=>"100000101",
  36454=>"111001000",
  36455=>"001111111",
  36456=>"111000000",
  36457=>"000100100",
  36458=>"111111000",
  36459=>"011001001",
  36460=>"110111110",
  36461=>"000000111",
  36462=>"000000000",
  36463=>"000000000",
  36464=>"000000000",
  36465=>"001011011",
  36466=>"010010110",
  36467=>"111000000",
  36468=>"110110111",
  36469=>"000100000",
  36470=>"000111111",
  36471=>"000000000",
  36472=>"010000100",
  36473=>"000000000",
  36474=>"000000000",
  36475=>"000000000",
  36476=>"100110110",
  36477=>"111101111",
  36478=>"000000000",
  36479=>"000000000",
  36480=>"100100000",
  36481=>"111111111",
  36482=>"001100000",
  36483=>"001000001",
  36484=>"000000001",
  36485=>"011000100",
  36486=>"000000001",
  36487=>"000000101",
  36488=>"000000000",
  36489=>"010110111",
  36490=>"000110111",
  36491=>"000111111",
  36492=>"011101111",
  36493=>"011001001",
  36494=>"000000010",
  36495=>"101011001",
  36496=>"000001001",
  36497=>"010111000",
  36498=>"000000000",
  36499=>"000001001",
  36500=>"111111011",
  36501=>"001100111",
  36502=>"010110111",
  36503=>"001000001",
  36504=>"110000000",
  36505=>"111111011",
  36506=>"111111111",
  36507=>"010001001",
  36508=>"111111111",
  36509=>"000110100",
  36510=>"111011011",
  36511=>"100100111",
  36512=>"000000000",
  36513=>"110110000",
  36514=>"000000100",
  36515=>"000000111",
  36516=>"001011011",
  36517=>"100101101",
  36518=>"100100000",
  36519=>"110011000",
  36520=>"001111111",
  36521=>"000000000",
  36522=>"011001101",
  36523=>"100011111",
  36524=>"100100100",
  36525=>"000100000",
  36526=>"011011011",
  36527=>"111011110",
  36528=>"111111110",
  36529=>"011010000",
  36530=>"000111000",
  36531=>"000000000",
  36532=>"000000001",
  36533=>"110110110",
  36534=>"111111111",
  36535=>"001000001",
  36536=>"110000100",
  36537=>"000000000",
  36538=>"100010000",
  36539=>"110111110",
  36540=>"001001011",
  36541=>"010111111",
  36542=>"110111000",
  36543=>"100101111",
  36544=>"010011100",
  36545=>"000100100",
  36546=>"000000000",
  36547=>"001000000",
  36548=>"111111111",
  36549=>"011111111",
  36550=>"111000000",
  36551=>"100000111",
  36552=>"000010010",
  36553=>"001000111",
  36554=>"011001001",
  36555=>"111111011",
  36556=>"111111111",
  36557=>"100000000",
  36558=>"111111100",
  36559=>"000000000",
  36560=>"011111111",
  36561=>"111000000",
  36562=>"100100100",
  36563=>"000001111",
  36564=>"000000000",
  36565=>"001001011",
  36566=>"000110110",
  36567=>"100001111",
  36568=>"000000100",
  36569=>"111110110",
  36570=>"111111111",
  36571=>"100100000",
  36572=>"110100101",
  36573=>"000001111",
  36574=>"000101111",
  36575=>"000000000",
  36576=>"111011010",
  36577=>"111111111",
  36578=>"010110000",
  36579=>"010110111",
  36580=>"001000011",
  36581=>"111111111",
  36582=>"100000000",
  36583=>"111111111",
  36584=>"000000000",
  36585=>"001001111",
  36586=>"111001001",
  36587=>"111111101",
  36588=>"000000000",
  36589=>"000000000",
  36590=>"000100110",
  36591=>"010010000",
  36592=>"111101000",
  36593=>"001000000",
  36594=>"001011111",
  36595=>"101111001",
  36596=>"110100011",
  36597=>"000100100",
  36598=>"111000001",
  36599=>"011111111",
  36600=>"000000001",
  36601=>"001001000",
  36602=>"100000000",
  36603=>"111111100",
  36604=>"011001011",
  36605=>"001001011",
  36606=>"000111111",
  36607=>"100100000",
  36608=>"111111111",
  36609=>"000000000",
  36610=>"111111111",
  36611=>"000111111",
  36612=>"000000100",
  36613=>"000000000",
  36614=>"000000000",
  36615=>"111011011",
  36616=>"111111111",
  36617=>"000000000",
  36618=>"001001111",
  36619=>"000000111",
  36620=>"110110110",
  36621=>"100111101",
  36622=>"011011111",
  36623=>"000000000",
  36624=>"000000000",
  36625=>"000001111",
  36626=>"000000100",
  36627=>"000011000",
  36628=>"001001111",
  36629=>"001111001",
  36630=>"000110100",
  36631=>"100000000",
  36632=>"000110110",
  36633=>"011000000",
  36634=>"100000101",
  36635=>"000110110",
  36636=>"111111111",
  36637=>"000000000",
  36638=>"010000000",
  36639=>"110111111",
  36640=>"000010011",
  36641=>"001000000",
  36642=>"111011011",
  36643=>"000001111",
  36644=>"100100100",
  36645=>"111101111",
  36646=>"001000101",
  36647=>"000000000",
  36648=>"111110111",
  36649=>"111001001",
  36650=>"010011000",
  36651=>"000000000",
  36652=>"001011000",
  36653=>"000001011",
  36654=>"110000000",
  36655=>"100000000",
  36656=>"000000000",
  36657=>"111111111",
  36658=>"000000000",
  36659=>"000000000",
  36660=>"010000000",
  36661=>"000010010",
  36662=>"000111111",
  36663=>"111100100",
  36664=>"010010000",
  36665=>"111111111",
  36666=>"000000000",
  36667=>"000111111",
  36668=>"000000001",
  36669=>"111111000",
  36670=>"000011111",
  36671=>"100100000",
  36672=>"000110111",
  36673=>"100110110",
  36674=>"111111111",
  36675=>"000000000",
  36676=>"000000000",
  36677=>"111011000",
  36678=>"000000000",
  36679=>"000100000",
  36680=>"100110000",
  36681=>"000100000",
  36682=>"101000000",
  36683=>"000000001",
  36684=>"000010000",
  36685=>"111111011",
  36686=>"111001011",
  36687=>"101111011",
  36688=>"001001011",
  36689=>"000010110",
  36690=>"001000000",
  36691=>"111111111",
  36692=>"111111111",
  36693=>"011011011",
  36694=>"000000000",
  36695=>"000110110",
  36696=>"000000001",
  36697=>"111111111",
  36698=>"001101001",
  36699=>"111100001",
  36700=>"000000001",
  36701=>"100100110",
  36702=>"111011000",
  36703=>"001001001",
  36704=>"011111111",
  36705=>"000000000",
  36706=>"011011001",
  36707=>"111111111",
  36708=>"100111111",
  36709=>"000000000",
  36710=>"000000000",
  36711=>"100111111",
  36712=>"000000100",
  36713=>"111111110",
  36714=>"000000000",
  36715=>"001001100",
  36716=>"110110100",
  36717=>"000011001",
  36718=>"001111111",
  36719=>"000111111",
  36720=>"000000000",
  36721=>"110110000",
  36722=>"001001011",
  36723=>"111101100",
  36724=>"111111101",
  36725=>"100000000",
  36726=>"000000000",
  36727=>"110110011",
  36728=>"000011000",
  36729=>"000000000",
  36730=>"000001111",
  36731=>"000000000",
  36732=>"111010000",
  36733=>"111111000",
  36734=>"000000000",
  36735=>"001000111",
  36736=>"111111111",
  36737=>"000001010",
  36738=>"001100000",
  36739=>"110110100",
  36740=>"001000100",
  36741=>"110110110",
  36742=>"101111110",
  36743=>"110110110",
  36744=>"000001000",
  36745=>"111111111",
  36746=>"111011000",
  36747=>"110110110",
  36748=>"000111111",
  36749=>"101000000",
  36750=>"000000000",
  36751=>"100111111",
  36752=>"000000000",
  36753=>"000000000",
  36754=>"000000000",
  36755=>"100110110",
  36756=>"000000000",
  36757=>"110110110",
  36758=>"001001111",
  36759=>"011010000",
  36760=>"111011001",
  36761=>"000000110",
  36762=>"000000100",
  36763=>"000111111",
  36764=>"001001000",
  36765=>"111000000",
  36766=>"100000000",
  36767=>"111111000",
  36768=>"000110010",
  36769=>"000011011",
  36770=>"101000000",
  36771=>"000000011",
  36772=>"100000011",
  36773=>"010111000",
  36774=>"001000000",
  36775=>"000100101",
  36776=>"111011111",
  36777=>"111010100",
  36778=>"001001111",
  36779=>"100111111",
  36780=>"001000100",
  36781=>"111111111",
  36782=>"100000000",
  36783=>"000111111",
  36784=>"111111111",
  36785=>"100101111",
  36786=>"000000000",
  36787=>"000100001",
  36788=>"100100000",
  36789=>"000110111",
  36790=>"000000000",
  36791=>"000111111",
  36792=>"000111111",
  36793=>"001000000",
  36794=>"111111100",
  36795=>"111111111",
  36796=>"111111011",
  36797=>"101001001",
  36798=>"000000000",
  36799=>"000010000",
  36800=>"001000001",
  36801=>"101100000",
  36802=>"010111010",
  36803=>"000111111",
  36804=>"111111111",
  36805=>"000000010",
  36806=>"111101000",
  36807=>"111111111",
  36808=>"000100100",
  36809=>"111111011",
  36810=>"000010111",
  36811=>"100000000",
  36812=>"000111110",
  36813=>"000000000",
  36814=>"111111111",
  36815=>"010011000",
  36816=>"000110100",
  36817=>"111110100",
  36818=>"000100111",
  36819=>"111111111",
  36820=>"101000000",
  36821=>"001000000",
  36822=>"111111000",
  36823=>"110000000",
  36824=>"001011001",
  36825=>"000000000",
  36826=>"111111011",
  36827=>"101001001",
  36828=>"001001001",
  36829=>"100000000",
  36830=>"110111111",
  36831=>"000000000",
  36832=>"100000000",
  36833=>"100111111",
  36834=>"011001001",
  36835=>"111111111",
  36836=>"111111111",
  36837=>"100100000",
  36838=>"111111100",
  36839=>"000000111",
  36840=>"111111100",
  36841=>"111001000",
  36842=>"111111111",
  36843=>"110110100",
  36844=>"101100111",
  36845=>"110110000",
  36846=>"000001000",
  36847=>"000000000",
  36848=>"000000000",
  36849=>"111111111",
  36850=>"111000111",
  36851=>"010000000",
  36852=>"001000110",
  36853=>"110111111",
  36854=>"001111111",
  36855=>"000000000",
  36856=>"001001001",
  36857=>"100110010",
  36858=>"011111111",
  36859=>"000000000",
  36860=>"111111111",
  36861=>"001111111",
  36862=>"110111111",
  36863=>"001000000",
  36864=>"111111111",
  36865=>"000000000",
  36866=>"000111111",
  36867=>"100111111",
  36868=>"110111011",
  36869=>"000000000",
  36870=>"001000000",
  36871=>"111111111",
  36872=>"000000000",
  36873=>"001000001",
  36874=>"110101001",
  36875=>"001111111",
  36876=>"000000100",
  36877=>"111011001",
  36878=>"001111111",
  36879=>"111000000",
  36880=>"011011011",
  36881=>"111101000",
  36882=>"100000000",
  36883=>"011011011",
  36884=>"000000000",
  36885=>"110111001",
  36886=>"000000000",
  36887=>"111001000",
  36888=>"100001001",
  36889=>"101001011",
  36890=>"111001001",
  36891=>"111001000",
  36892=>"011011011",
  36893=>"111111111",
  36894=>"001000101",
  36895=>"000010111",
  36896=>"111111000",
  36897=>"000000000",
  36898=>"000111011",
  36899=>"111011110",
  36900=>"111111111",
  36901=>"001001000",
  36902=>"110100000",
  36903=>"000011111",
  36904=>"000100000",
  36905=>"000000000",
  36906=>"111101001",
  36907=>"100100000",
  36908=>"111111011",
  36909=>"010111111",
  36910=>"000010111",
  36911=>"110111111",
  36912=>"100100101",
  36913=>"111011001",
  36914=>"011111001",
  36915=>"000000000",
  36916=>"000010111",
  36917=>"011100000",
  36918=>"111111111",
  36919=>"001101101",
  36920=>"011111111",
  36921=>"000000000",
  36922=>"000000000",
  36923=>"000000110",
  36924=>"000111111",
  36925=>"110100000",
  36926=>"100000000",
  36927=>"000000101",
  36928=>"100010011",
  36929=>"011010111",
  36930=>"010000001",
  36931=>"000001111",
  36932=>"000000000",
  36933=>"011011110",
  36934=>"111000000",
  36935=>"000000000",
  36936=>"000000000",
  36937=>"000000000",
  36938=>"111111011",
  36939=>"110000111",
  36940=>"000000000",
  36941=>"111111010",
  36942=>"111111111",
  36943=>"110110111",
  36944=>"000110111",
  36945=>"000000000",
  36946=>"110000000",
  36947=>"000000000",
  36948=>"000001011",
  36949=>"000000011",
  36950=>"110110000",
  36951=>"110011010",
  36952=>"000000001",
  36953=>"000000111",
  36954=>"111011111",
  36955=>"000000000",
  36956=>"001000000",
  36957=>"000000000",
  36958=>"001111111",
  36959=>"010110111",
  36960=>"111111111",
  36961=>"101101001",
  36962=>"000000000",
  36963=>"111110000",
  36964=>"010000110",
  36965=>"111110111",
  36966=>"000000000",
  36967=>"000000000",
  36968=>"000010011",
  36969=>"100110000",
  36970=>"111111111",
  36971=>"111111111",
  36972=>"111110111",
  36973=>"111011111",
  36974=>"111111111",
  36975=>"111010000",
  36976=>"000010111",
  36977=>"000011111",
  36978=>"000001111",
  36979=>"111110000",
  36980=>"111001101",
  36981=>"000100110",
  36982=>"111111111",
  36983=>"000000100",
  36984=>"101111111",
  36985=>"000111011",
  36986=>"111000000",
  36987=>"011001001",
  36988=>"010111110",
  36989=>"000000000",
  36990=>"000000000",
  36991=>"111111111",
  36992=>"011010111",
  36993=>"111111111",
  36994=>"110000111",
  36995=>"000000000",
  36996=>"111111111",
  36997=>"000000111",
  36998=>"111111111",
  36999=>"000000001",
  37000=>"000000011",
  37001=>"000000111",
  37002=>"000000100",
  37003=>"000000000",
  37004=>"000000000",
  37005=>"000000100",
  37006=>"101001011",
  37007=>"000000100",
  37008=>"000000000",
  37009=>"000000100",
  37010=>"110010010",
  37011=>"111111100",
  37012=>"111001000",
  37013=>"000110101",
  37014=>"110111000",
  37015=>"000000000",
  37016=>"111111111",
  37017=>"000000011",
  37018=>"111111011",
  37019=>"111111111",
  37020=>"000001101",
  37021=>"111111011",
  37022=>"000101111",
  37023=>"111111111",
  37024=>"100100110",
  37025=>"000110111",
  37026=>"100111011",
  37027=>"100111001",
  37028=>"111000000",
  37029=>"001001001",
  37030=>"111111111",
  37031=>"100110100",
  37032=>"001000000",
  37033=>"100000010",
  37034=>"111001000",
  37035=>"000110111",
  37036=>"101111010",
  37037=>"000001001",
  37038=>"111000000",
  37039=>"000000000",
  37040=>"100111111",
  37041=>"000100100",
  37042=>"110111111",
  37043=>"011000111",
  37044=>"111111011",
  37045=>"110000000",
  37046=>"000000011",
  37047=>"000000000",
  37048=>"100000001",
  37049=>"000000000",
  37050=>"101000100",
  37051=>"000000111",
  37052=>"100100000",
  37053=>"010000111",
  37054=>"111111111",
  37055=>"110000100",
  37056=>"000110110",
  37057=>"111111111",
  37058=>"111011011",
  37059=>"000000000",
  37060=>"000000011",
  37061=>"000000110",
  37062=>"111110100",
  37063=>"111111111",
  37064=>"000110111",
  37065=>"111111111",
  37066=>"111111000",
  37067=>"111111000",
  37068=>"111111111",
  37069=>"111111111",
  37070=>"111111000",
  37071=>"111000000",
  37072=>"111011000",
  37073=>"000000000",
  37074=>"001000000",
  37075=>"000000001",
  37076=>"000001000",
  37077=>"101111111",
  37078=>"000000000",
  37079=>"011111001",
  37080=>"111111111",
  37081=>"000111000",
  37082=>"110110000",
  37083=>"101000000",
  37084=>"111111011",
  37085=>"011111111",
  37086=>"000000111",
  37087=>"000000000",
  37088=>"000000001",
  37089=>"110000110",
  37090=>"110111111",
  37091=>"000111111",
  37092=>"111110100",
  37093=>"000000001",
  37094=>"000111100",
  37095=>"000000000",
  37096=>"111100000",
  37097=>"000000000",
  37098=>"101101101",
  37099=>"100100100",
  37100=>"000010010",
  37101=>"000000000",
  37102=>"111101111",
  37103=>"111011000",
  37104=>"100101001",
  37105=>"000000000",
  37106=>"000111111",
  37107=>"000000000",
  37108=>"011000000",
  37109=>"000000000",
  37110=>"111111111",
  37111=>"111111111",
  37112=>"111000000",
  37113=>"111111001",
  37114=>"010111111",
  37115=>"010011001",
  37116=>"100110011",
  37117=>"110100101",
  37118=>"101001000",
  37119=>"100000000",
  37120=>"000000100",
  37121=>"100101111",
  37122=>"111111011",
  37123=>"000011111",
  37124=>"111101101",
  37125=>"010101100",
  37126=>"000000000",
  37127=>"110111001",
  37128=>"110111000",
  37129=>"111110110",
  37130=>"000011111",
  37131=>"000111111",
  37132=>"100100100",
  37133=>"000001111",
  37134=>"111111011",
  37135=>"010000111",
  37136=>"000000100",
  37137=>"000001001",
  37138=>"000011111",
  37139=>"111111111",
  37140=>"000000000",
  37141=>"111111111",
  37142=>"100100000",
  37143=>"000000111",
  37144=>"000110110",
  37145=>"000011111",
  37146=>"000000111",
  37147=>"110100000",
  37148=>"110110111",
  37149=>"000010001",
  37150=>"111101111",
  37151=>"111010000",
  37152=>"001000100",
  37153=>"111000000",
  37154=>"000110111",
  37155=>"100000000",
  37156=>"110010000",
  37157=>"111100100",
  37158=>"111011001",
  37159=>"110110111",
  37160=>"111111111",
  37161=>"111111111",
  37162=>"010010010",
  37163=>"011011001",
  37164=>"111111111",
  37165=>"100110000",
  37166=>"011001000",
  37167=>"000000111",
  37168=>"001000011",
  37169=>"001100110",
  37170=>"111001100",
  37171=>"011000100",
  37172=>"110000000",
  37173=>"000011111",
  37174=>"000111101",
  37175=>"110000000",
  37176=>"110010000",
  37177=>"111111111",
  37178=>"111111111",
  37179=>"110000000",
  37180=>"111110111",
  37181=>"010111000",
  37182=>"000111111",
  37183=>"001111111",
  37184=>"001001000",
  37185=>"000111111",
  37186=>"000000000",
  37187=>"111111111",
  37188=>"000001111",
  37189=>"100101101",
  37190=>"101011111",
  37191=>"100100100",
  37192=>"000000000",
  37193=>"001000000",
  37194=>"000000000",
  37195=>"000100100",
  37196=>"000000000",
  37197=>"011111011",
  37198=>"000101001",
  37199=>"000001000",
  37200=>"101111011",
  37201=>"000111000",
  37202=>"000000001",
  37203=>"111111111",
  37204=>"111111111",
  37205=>"001001001",
  37206=>"111111100",
  37207=>"111111110",
  37208=>"010010111",
  37209=>"111111111",
  37210=>"000000000",
  37211=>"111011000",
  37212=>"000000001",
  37213=>"111110111",
  37214=>"100111000",
  37215=>"000000100",
  37216=>"111011011",
  37217=>"000000000",
  37218=>"000011011",
  37219=>"011000000",
  37220=>"000100100",
  37221=>"111111111",
  37222=>"000000000",
  37223=>"000001001",
  37224=>"100101000",
  37225=>"000000000",
  37226=>"000100000",
  37227=>"111111111",
  37228=>"000110010",
  37229=>"000000110",
  37230=>"001000000",
  37231=>"001000000",
  37232=>"100111111",
  37233=>"111111111",
  37234=>"000001001",
  37235=>"000000110",
  37236=>"111111111",
  37237=>"111001000",
  37238=>"111111111",
  37239=>"000000000",
  37240=>"110000111",
  37241=>"000111111",
  37242=>"000000000",
  37243=>"111111100",
  37244=>"011011111",
  37245=>"100111111",
  37246=>"000100000",
  37247=>"111000000",
  37248=>"000000000",
  37249=>"100111111",
  37250=>"000000001",
  37251=>"000011111",
  37252=>"000000000",
  37253=>"000010111",
  37254=>"111111011",
  37255=>"000011111",
  37256=>"100101000",
  37257=>"110010000",
  37258=>"000001011",
  37259=>"110011111",
  37260=>"111111101",
  37261=>"000000000",
  37262=>"000000000",
  37263=>"011000000",
  37264=>"111111111",
  37265=>"001001111",
  37266=>"000110110",
  37267=>"001001011",
  37268=>"000000111",
  37269=>"000000000",
  37270=>"111111001",
  37271=>"001000000",
  37272=>"111001000",
  37273=>"111111111",
  37274=>"000011111",
  37275=>"000000000",
  37276=>"100100110",
  37277=>"000010010",
  37278=>"100100110",
  37279=>"011000000",
  37280=>"011000000",
  37281=>"111111100",
  37282=>"000111111",
  37283=>"000001001",
  37284=>"100111111",
  37285=>"000111011",
  37286=>"011000000",
  37287=>"000000000",
  37288=>"000000000",
  37289=>"000111111",
  37290=>"101111111",
  37291=>"000111010",
  37292=>"000000000",
  37293=>"100111111",
  37294=>"000001000",
  37295=>"000000000",
  37296=>"111011011",
  37297=>"100000000",
  37298=>"000100000",
  37299=>"000110000",
  37300=>"111111111",
  37301=>"111111100",
  37302=>"100110101",
  37303=>"111111001",
  37304=>"010010001",
  37305=>"111000000",
  37306=>"100110000",
  37307=>"100101111",
  37308=>"010000000",
  37309=>"111100101",
  37310=>"000011011",
  37311=>"000100111",
  37312=>"000110110",
  37313=>"000100000",
  37314=>"111011011",
  37315=>"011000000",
  37316=>"111111111",
  37317=>"111111111",
  37318=>"111111111",
  37319=>"000111000",
  37320=>"101100101",
  37321=>"111100111",
  37322=>"000000111",
  37323=>"000000000",
  37324=>"011011000",
  37325=>"111011111",
  37326=>"000011111",
  37327=>"111111111",
  37328=>"001001000",
  37329=>"001001001",
  37330=>"111111000",
  37331=>"111111111",
  37332=>"000111111",
  37333=>"111111111",
  37334=>"000000001",
  37335=>"011000000",
  37336=>"000100100",
  37337=>"000010010",
  37338=>"010111111",
  37339=>"000000110",
  37340=>"011011111",
  37341=>"110111011",
  37342=>"111001000",
  37343=>"111111111",
  37344=>"110111110",
  37345=>"000000111",
  37346=>"000000000",
  37347=>"000111101",
  37348=>"000111111",
  37349=>"100000000",
  37350=>"010010000",
  37351=>"000000000",
  37352=>"000010000",
  37353=>"100100011",
  37354=>"111111111",
  37355=>"001101101",
  37356=>"000011000",
  37357=>"000000100",
  37358=>"000000010",
  37359=>"110101101",
  37360=>"111111101",
  37361=>"111000000",
  37362=>"111111111",
  37363=>"000000111",
  37364=>"000100100",
  37365=>"011111111",
  37366=>"101100100",
  37367=>"011000001",
  37368=>"000000000",
  37369=>"000000100",
  37370=>"111111000",
  37371=>"100100000",
  37372=>"010000001",
  37373=>"100100110",
  37374=>"000000000",
  37375=>"111000100",
  37376=>"111100000",
  37377=>"111111000",
  37378=>"001111111",
  37379=>"000111110",
  37380=>"111111111",
  37381=>"010100000",
  37382=>"001001001",
  37383=>"111111111",
  37384=>"001000000",
  37385=>"000000101",
  37386=>"000000000",
  37387=>"110111111",
  37388=>"110111101",
  37389=>"100100111",
  37390=>"111111001",
  37391=>"000000000",
  37392=>"000110111",
  37393=>"001111101",
  37394=>"000000000",
  37395=>"110000010",
  37396=>"111111011",
  37397=>"111111111",
  37398=>"000111110",
  37399=>"111111000",
  37400=>"111111111",
  37401=>"111111011",
  37402=>"101100111",
  37403=>"111111001",
  37404=>"001000101",
  37405=>"111000001",
  37406=>"001001001",
  37407=>"011011001",
  37408=>"110111001",
  37409=>"110110000",
  37410=>"110111010",
  37411=>"000111101",
  37412=>"000110101",
  37413=>"000000100",
  37414=>"000000000",
  37415=>"000000100",
  37416=>"001001001",
  37417=>"000000110",
  37418=>"000000001",
  37419=>"111111010",
  37420=>"100000000",
  37421=>"111111010",
  37422=>"000000000",
  37423=>"000000000",
  37424=>"010111111",
  37425=>"110111001",
  37426=>"000111111",
  37427=>"000100011",
  37428=>"100111100",
  37429=>"101000011",
  37430=>"111011000",
  37431=>"110111111",
  37432=>"110111111",
  37433=>"111001111",
  37434=>"011011111",
  37435=>"111100000",
  37436=>"000000000",
  37437=>"001000000",
  37438=>"000111101",
  37439=>"000000000",
  37440=>"001000100",
  37441=>"001111111",
  37442=>"000000111",
  37443=>"000001111",
  37444=>"111110000",
  37445=>"001000010",
  37446=>"000011001",
  37447=>"111111100",
  37448=>"100100100",
  37449=>"000000001",
  37450=>"011010111",
  37451=>"101100111",
  37452=>"110111110",
  37453=>"000010011",
  37454=>"001010000",
  37455=>"000000000",
  37456=>"000000000",
  37457=>"000100100",
  37458=>"000000000",
  37459=>"011000000",
  37460=>"011011011",
  37461=>"000111111",
  37462=>"111000101",
  37463=>"000000000",
  37464=>"000000000",
  37465=>"101000101",
  37466=>"000000010",
  37467=>"100000001",
  37468=>"111000000",
  37469=>"000111111",
  37470=>"011011111",
  37471=>"011011111",
  37472=>"000101000",
  37473=>"110111100",
  37474=>"000000000",
  37475=>"111111110",
  37476=>"110110110",
  37477=>"001000001",
  37478=>"011111111",
  37479=>"100101111",
  37480=>"111000000",
  37481=>"111111101",
  37482=>"000000011",
  37483=>"110111111",
  37484=>"000111110",
  37485=>"001000111",
  37486=>"000000101",
  37487=>"100110111",
  37488=>"011000000",
  37489=>"101101111",
  37490=>"111110100",
  37491=>"111000001",
  37492=>"000000000",
  37493=>"001000000",
  37494=>"111101111",
  37495=>"000000010",
  37496=>"000000000",
  37497=>"111111010",
  37498=>"000000000",
  37499=>"000000000",
  37500=>"110110110",
  37501=>"111111011",
  37502=>"000000000",
  37503=>"111111010",
  37504=>"000000111",
  37505=>"110110111",
  37506=>"111111110",
  37507=>"000000000",
  37508=>"110110100",
  37509=>"000000111",
  37510=>"000000100",
  37511=>"000000000",
  37512=>"000110111",
  37513=>"110100000",
  37514=>"000000000",
  37515=>"001000111",
  37516=>"000000000",
  37517=>"001000000",
  37518=>"001111111",
  37519=>"000010000",
  37520=>"000000101",
  37521=>"111000100",
  37522=>"111111111",
  37523=>"111111000",
  37524=>"011111111",
  37525=>"111011000",
  37526=>"111111101",
  37527=>"001001111",
  37528=>"001000101",
  37529=>"000000000",
  37530=>"111111111",
  37531=>"010111111",
  37532=>"001001011",
  37533=>"011001000",
  37534=>"111111111",
  37535=>"000100111",
  37536=>"111111111",
  37537=>"111111000",
  37538=>"000000111",
  37539=>"011000000",
  37540=>"011001001",
  37541=>"111111111",
  37542=>"000111111",
  37543=>"110110110",
  37544=>"001000000",
  37545=>"001001001",
  37546=>"111111111",
  37547=>"011000000",
  37548=>"110101111",
  37549=>"110111111",
  37550=>"111000000",
  37551=>"000000000",
  37552=>"000000000",
  37553=>"111111111",
  37554=>"110111011",
  37555=>"111011011",
  37556=>"011011011",
  37557=>"000001011",
  37558=>"000000001",
  37559=>"000000000",
  37560=>"001000111",
  37561=>"000000000",
  37562=>"000000000",
  37563=>"010000000",
  37564=>"001000000",
  37565=>"000111011",
  37566=>"111110111",
  37567=>"111111000",
  37568=>"111111111",
  37569=>"001001101",
  37570=>"110100000",
  37571=>"000000000",
  37572=>"000000000",
  37573=>"000000000",
  37574=>"001000000",
  37575=>"110110110",
  37576=>"000000000",
  37577=>"110111010",
  37578=>"000000000",
  37579=>"011000111",
  37580=>"100000000",
  37581=>"000100100",
  37582=>"000000111",
  37583=>"011000000",
  37584=>"111111011",
  37585=>"100100110",
  37586=>"111111000",
  37587=>"010000000",
  37588=>"100000011",
  37589=>"110111010",
  37590=>"000000110",
  37591=>"000001101",
  37592=>"000111110",
  37593=>"001001001",
  37594=>"111000111",
  37595=>"111111001",
  37596=>"111001000",
  37597=>"000000001",
  37598=>"000000100",
  37599=>"011011001",
  37600=>"000000000",
  37601=>"000000111",
  37602=>"000111111",
  37603=>"000000001",
  37604=>"011111111",
  37605=>"000000111",
  37606=>"000100111",
  37607=>"001111111",
  37608=>"111011011",
  37609=>"111110111",
  37610=>"001011011",
  37611=>"111101111",
  37612=>"000000000",
  37613=>"001000100",
  37614=>"000000000",
  37615=>"000000000",
  37616=>"000000000",
  37617=>"011000000",
  37618=>"111100000",
  37619=>"111001000",
  37620=>"000000000",
  37621=>"100110110",
  37622=>"111111011",
  37623=>"110100100",
  37624=>"000000111",
  37625=>"010011011",
  37626=>"001000001",
  37627=>"110111111",
  37628=>"110111111",
  37629=>"000000000",
  37630=>"000110110",
  37631=>"110000100",
  37632=>"000000000",
  37633=>"111111111",
  37634=>"001000111",
  37635=>"111111000",
  37636=>"000000000",
  37637=>"000000000",
  37638=>"000110111",
  37639=>"000001001",
  37640=>"000000000",
  37641=>"000000000",
  37642=>"000000100",
  37643=>"111111001",
  37644=>"000001111",
  37645=>"000000010",
  37646=>"000000000",
  37647=>"111100110",
  37648=>"110000000",
  37649=>"000000011",
  37650=>"001001001",
  37651=>"010111111",
  37652=>"111000000",
  37653=>"011000000",
  37654=>"111011011",
  37655=>"011111000",
  37656=>"001011111",
  37657=>"011000001",
  37658=>"000000000",
  37659=>"011111011",
  37660=>"111000000",
  37661=>"111111111",
  37662=>"000000000",
  37663=>"011001000",
  37664=>"111011000",
  37665=>"100111111",
  37666=>"000000000",
  37667=>"111100001",
  37668=>"000000000",
  37669=>"111011001",
  37670=>"000000000",
  37671=>"111110000",
  37672=>"000000110",
  37673=>"010011011",
  37674=>"111111010",
  37675=>"000000000",
  37676=>"100111111",
  37677=>"000000000",
  37678=>"000000001",
  37679=>"000000000",
  37680=>"000100110",
  37681=>"000000000",
  37682=>"111111000",
  37683=>"000000000",
  37684=>"000000000",
  37685=>"110011111",
  37686=>"111100100",
  37687=>"111111001",
  37688=>"000000000",
  37689=>"111100101",
  37690=>"111011000",
  37691=>"111111000",
  37692=>"000000000",
  37693=>"000110110",
  37694=>"001111111",
  37695=>"000000000",
  37696=>"001000101",
  37697=>"110111000",
  37698=>"001000000",
  37699=>"001111001",
  37700=>"000000100",
  37701=>"111111111",
  37702=>"111111111",
  37703=>"110000110",
  37704=>"000000100",
  37705=>"000001001",
  37706=>"000000000",
  37707=>"011000100",
  37708=>"111011000",
  37709=>"000000100",
  37710=>"000000100",
  37711=>"110111111",
  37712=>"000000100",
  37713=>"011001101",
  37714=>"010000110",
  37715=>"110111010",
  37716=>"000001001",
  37717=>"011011011",
  37718=>"000000000",
  37719=>"000000000",
  37720=>"000000000",
  37721=>"111111111",
  37722=>"111111000",
  37723=>"110111010",
  37724=>"000000000",
  37725=>"000000000",
  37726=>"001001000",
  37727=>"111111111",
  37728=>"111111111",
  37729=>"111111100",
  37730=>"110100100",
  37731=>"000000101",
  37732=>"000000100",
  37733=>"000011000",
  37734=>"000101111",
  37735=>"010111111",
  37736=>"010000000",
  37737=>"100000101",
  37738=>"000100111",
  37739=>"111000000",
  37740=>"001011110",
  37741=>"111110010",
  37742=>"000000000",
  37743=>"000000000",
  37744=>"000000111",
  37745=>"000110000",
  37746=>"110111100",
  37747=>"111111011",
  37748=>"111111011",
  37749=>"111111111",
  37750=>"000000000",
  37751=>"000000001",
  37752=>"111111111",
  37753=>"111111111",
  37754=>"010111011",
  37755=>"111000110",
  37756=>"000000011",
  37757=>"000000010",
  37758=>"110000000",
  37759=>"000000000",
  37760=>"000000000",
  37761=>"110111011",
  37762=>"110011011",
  37763=>"000000010",
  37764=>"111101000",
  37765=>"000001011",
  37766=>"101000001",
  37767=>"000000000",
  37768=>"011000011",
  37769=>"000000100",
  37770=>"111111111",
  37771=>"000000000",
  37772=>"000000111",
  37773=>"000000000",
  37774=>"000100000",
  37775=>"000000100",
  37776=>"010111111",
  37777=>"000000001",
  37778=>"100100000",
  37779=>"100000100",
  37780=>"110110000",
  37781=>"000000000",
  37782=>"000011111",
  37783=>"111111001",
  37784=>"000111110",
  37785=>"011001011",
  37786=>"001000001",
  37787=>"111111000",
  37788=>"000000101",
  37789=>"000110110",
  37790=>"111111011",
  37791=>"000000100",
  37792=>"000000011",
  37793=>"000000100",
  37794=>"001111100",
  37795=>"000000000",
  37796=>"000000111",
  37797=>"111111111",
  37798=>"011111010",
  37799=>"111110110",
  37800=>"000100110",
  37801=>"101000000",
  37802=>"111111111",
  37803=>"011001000",
  37804=>"000000000",
  37805=>"101111111",
  37806=>"100000111",
  37807=>"000000000",
  37808=>"001000000",
  37809=>"000000111",
  37810=>"100110000",
  37811=>"010000000",
  37812=>"110110100",
  37813=>"111111111",
  37814=>"110111111",
  37815=>"000000000",
  37816=>"000000000",
  37817=>"110110110",
  37818=>"100000000",
  37819=>"000111111",
  37820=>"000001000",
  37821=>"101000000",
  37822=>"111110000",
  37823=>"010000100",
  37824=>"000000000",
  37825=>"000000111",
  37826=>"000001000",
  37827=>"111111011",
  37828=>"111000001",
  37829=>"000000100",
  37830=>"100110111",
  37831=>"000100100",
  37832=>"001001000",
  37833=>"001011111",
  37834=>"000000000",
  37835=>"110110110",
  37836=>"001000000",
  37837=>"110110100",
  37838=>"100110000",
  37839=>"111111110",
  37840=>"111011000",
  37841=>"000000100",
  37842=>"100100100",
  37843=>"111101100",
  37844=>"111100000",
  37845=>"011000000",
  37846=>"011111111",
  37847=>"000000110",
  37848=>"000000000",
  37849=>"011001111",
  37850=>"000000100",
  37851=>"011000000",
  37852=>"110111111",
  37853=>"000000000",
  37854=>"101000101",
  37855=>"111110100",
  37856=>"110000100",
  37857=>"000000100",
  37858=>"000100111",
  37859=>"000000100",
  37860=>"111111111",
  37861=>"000111111",
  37862=>"000000110",
  37863=>"000000111",
  37864=>"100100000",
  37865=>"000101111",
  37866=>"110000100",
  37867=>"110111010",
  37868=>"111111101",
  37869=>"111111100",
  37870=>"000000000",
  37871=>"011011000",
  37872=>"100000000",
  37873=>"010111111",
  37874=>"111101000",
  37875=>"111111000",
  37876=>"111000110",
  37877=>"000000000",
  37878=>"111111000",
  37879=>"000111111",
  37880=>"001101111",
  37881=>"010011001",
  37882=>"000000000",
  37883=>"000000000",
  37884=>"111111111",
  37885=>"111111100",
  37886=>"000000000",
  37887=>"000000111",
  37888=>"111111001",
  37889=>"000000000",
  37890=>"000000000",
  37891=>"011001111",
  37892=>"100000011",
  37893=>"011101101",
  37894=>"001111111",
  37895=>"000000000",
  37896=>"001001111",
  37897=>"000000001",
  37898=>"111111111",
  37899=>"111100101",
  37900=>"110110110",
  37901=>"100100000",
  37902=>"101001111",
  37903=>"001111111",
  37904=>"000110111",
  37905=>"111111011",
  37906=>"000000000",
  37907=>"110111011",
  37908=>"101100100",
  37909=>"000111111",
  37910=>"000111111",
  37911=>"011111011",
  37912=>"000000100",
  37913=>"111011111",
  37914=>"000111111",
  37915=>"011000100",
  37916=>"001001111",
  37917=>"000000110",
  37918=>"001001101",
  37919=>"000000000",
  37920=>"111111111",
  37921=>"111111111",
  37922=>"111111110",
  37923=>"110110010",
  37924=>"000000000",
  37925=>"111001001",
  37926=>"000000000",
  37927=>"000100101",
  37928=>"111110010",
  37929=>"000110000",
  37930=>"001000000",
  37931=>"000000001",
  37932=>"000000101",
  37933=>"110111010",
  37934=>"001001011",
  37935=>"111111000",
  37936=>"111001001",
  37937=>"111111111",
  37938=>"111111100",
  37939=>"000000000",
  37940=>"110010000",
  37941=>"001001000",
  37942=>"000000000",
  37943=>"000000000",
  37944=>"111111111",
  37945=>"000000000",
  37946=>"000111111",
  37947=>"111100110",
  37948=>"000000000",
  37949=>"010100000",
  37950=>"001011111",
  37951=>"000000111",
  37952=>"011000011",
  37953=>"110000001",
  37954=>"111111111",
  37955=>"110000100",
  37956=>"001000000",
  37957=>"001011011",
  37958=>"000000000",
  37959=>"000000000",
  37960=>"001100000",
  37961=>"111111111",
  37962=>"001101111",
  37963=>"111100100",
  37964=>"101001111",
  37965=>"000000000",
  37966=>"011010110",
  37967=>"001001000",
  37968=>"000000000",
  37969=>"000000000",
  37970=>"011011111",
  37971=>"000000000",
  37972=>"001011001",
  37973=>"000000000",
  37974=>"111110111",
  37975=>"110110110",
  37976=>"111111110",
  37977=>"101100111",
  37978=>"000000111",
  37979=>"110000110",
  37980=>"000111111",
  37981=>"000000000",
  37982=>"111110110",
  37983=>"011001001",
  37984=>"011111010",
  37985=>"011000000",
  37986=>"000000100",
  37987=>"111111111",
  37988=>"111111011",
  37989=>"001001111",
  37990=>"000000111",
  37991=>"110110110",
  37992=>"111111010",
  37993=>"001001111",
  37994=>"000001110",
  37995=>"100111011",
  37996=>"111111110",
  37997=>"111111111",
  37998=>"000000000",
  37999=>"111100000",
  38000=>"111101101",
  38001=>"000000000",
  38002=>"000100100",
  38003=>"101111011",
  38004=>"000000100",
  38005=>"111111111",
  38006=>"000000000",
  38007=>"001101000",
  38008=>"001000101",
  38009=>"111111000",
  38010=>"000000000",
  38011=>"111111001",
  38012=>"100101000",
  38013=>"100110110",
  38014=>"000000000",
  38015=>"111111111",
  38016=>"000000001",
  38017=>"110010011",
  38018=>"111000000",
  38019=>"110010001",
  38020=>"000000001",
  38021=>"111000000",
  38022=>"000000100",
  38023=>"000000000",
  38024=>"111111111",
  38025=>"111111111",
  38026=>"000001011",
  38027=>"000111111",
  38028=>"000000000",
  38029=>"000010010",
  38030=>"000101110",
  38031=>"111111110",
  38032=>"000000000",
  38033=>"000000111",
  38034=>"111011001",
  38035=>"111011011",
  38036=>"011011001",
  38037=>"000000101",
  38038=>"000111111",
  38039=>"100000000",
  38040=>"101001101",
  38041=>"111111111",
  38042=>"110111110",
  38043=>"111111111",
  38044=>"001000000",
  38045=>"101000101",
  38046=>"111101111",
  38047=>"000000000",
  38048=>"010000110",
  38049=>"011111111",
  38050=>"000110111",
  38051=>"000000000",
  38052=>"000110110",
  38053=>"000001101",
  38054=>"111111101",
  38055=>"100100100",
  38056=>"000000100",
  38057=>"101000001",
  38058=>"000000000",
  38059=>"111111111",
  38060=>"000110101",
  38061=>"111111011",
  38062=>"000000000",
  38063=>"000000000",
  38064=>"000110111",
  38065=>"011111111",
  38066=>"011011010",
  38067=>"000000000",
  38068=>"111100011",
  38069=>"110000000",
  38070=>"111111111",
  38071=>"001001011",
  38072=>"000000000",
  38073=>"110111111",
  38074=>"001000000",
  38075=>"111111111",
  38076=>"000000000",
  38077=>"001001111",
  38078=>"001000000",
  38079=>"000011001",
  38080=>"111111111",
  38081=>"001111001",
  38082=>"010110010",
  38083=>"000000000",
  38084=>"000000000",
  38085=>"000000000",
  38086=>"100000000",
  38087=>"111100111",
  38088=>"000100111",
  38089=>"000000111",
  38090=>"101000000",
  38091=>"111111011",
  38092=>"110110110",
  38093=>"000111111",
  38094=>"100110100",
  38095=>"100111111",
  38096=>"110111101",
  38097=>"111001000",
  38098=>"000100111",
  38099=>"000000000",
  38100=>"110100000",
  38101=>"100000111",
  38102=>"100111111",
  38103=>"001000000",
  38104=>"011011011",
  38105=>"110110110",
  38106=>"000000000",
  38107=>"000000111",
  38108=>"000000111",
  38109=>"000000100",
  38110=>"000000011",
  38111=>"000100000",
  38112=>"010000000",
  38113=>"000000000",
  38114=>"111111111",
  38115=>"111111111",
  38116=>"000001101",
  38117=>"111111111",
  38118=>"111111110",
  38119=>"000000001",
  38120=>"000000001",
  38121=>"001001000",
  38122=>"000000000",
  38123=>"111000100",
  38124=>"000000101",
  38125=>"001011000",
  38126=>"110111111",
  38127=>"000000001",
  38128=>"101000000",
  38129=>"001011111",
  38130=>"111110110",
  38131=>"000000000",
  38132=>"000011001",
  38133=>"110110100",
  38134=>"011011101",
  38135=>"010010010",
  38136=>"001111111",
  38137=>"101111111",
  38138=>"000010000",
  38139=>"100001001",
  38140=>"011011011",
  38141=>"011011111",
  38142=>"000000000",
  38143=>"010110110",
  38144=>"000000000",
  38145=>"101001000",
  38146=>"001011000",
  38147=>"000000010",
  38148=>"110111110",
  38149=>"000111111",
  38150=>"000000100",
  38151=>"111111110",
  38152=>"000000000",
  38153=>"100100000",
  38154=>"000000000",
  38155=>"111111111",
  38156=>"000000000",
  38157=>"110111101",
  38158=>"000000001",
  38159=>"010010000",
  38160=>"000000000",
  38161=>"011000111",
  38162=>"000000110",
  38163=>"111110111",
  38164=>"100100111",
  38165=>"110000000",
  38166=>"111111111",
  38167=>"000000000",
  38168=>"110111011",
  38169=>"111111000",
  38170=>"000000100",
  38171=>"010010000",
  38172=>"111110110",
  38173=>"010110111",
  38174=>"000000000",
  38175=>"000000100",
  38176=>"111111000",
  38177=>"110000000",
  38178=>"010000000",
  38179=>"000000100",
  38180=>"101001001",
  38181=>"000000000",
  38182=>"110110110",
  38183=>"001001011",
  38184=>"000000000",
  38185=>"000000000",
  38186=>"010110000",
  38187=>"000000000",
  38188=>"000000000",
  38189=>"010111110",
  38190=>"111111000",
  38191=>"111101001",
  38192=>"000111001",
  38193=>"000001011",
  38194=>"101000001",
  38195=>"111111010",
  38196=>"000010000",
  38197=>"111110000",
  38198=>"011001000",
  38199=>"001111000",
  38200=>"110010010",
  38201=>"111001100",
  38202=>"000000000",
  38203=>"111111111",
  38204=>"111111111",
  38205=>"100110111",
  38206=>"100111111",
  38207=>"001001100",
  38208=>"111000000",
  38209=>"000001001",
  38210=>"111111110",
  38211=>"000000000",
  38212=>"111111110",
  38213=>"000000000",
  38214=>"111111111",
  38215=>"001111111",
  38216=>"000000010",
  38217=>"000000000",
  38218=>"111111100",
  38219=>"000100100",
  38220=>"111000000",
  38221=>"110011000",
  38222=>"111100000",
  38223=>"000011111",
  38224=>"001000000",
  38225=>"000000010",
  38226=>"111111110",
  38227=>"000001111",
  38228=>"010010000",
  38229=>"001001001",
  38230=>"001001111",
  38231=>"000000000",
  38232=>"101111100",
  38233=>"001011001",
  38234=>"110100000",
  38235=>"001010000",
  38236=>"111111001",
  38237=>"000110000",
  38238=>"010011111",
  38239=>"000000010",
  38240=>"011001000",
  38241=>"100000001",
  38242=>"000000000",
  38243=>"000000000",
  38244=>"000000000",
  38245=>"000000000",
  38246=>"000000000",
  38247=>"000000111",
  38248=>"001000111",
  38249=>"011011111",
  38250=>"000101111",
  38251=>"111010011",
  38252=>"110111111",
  38253=>"000000111",
  38254=>"111100101",
  38255=>"001001001",
  38256=>"111111111",
  38257=>"011011011",
  38258=>"000011101",
  38259=>"111111010",
  38260=>"110110111",
  38261=>"001001101",
  38262=>"011110000",
  38263=>"100110010",
  38264=>"000000000",
  38265=>"100000100",
  38266=>"000000001",
  38267=>"011111111",
  38268=>"000011001",
  38269=>"101100101",
  38270=>"100000100",
  38271=>"111111111",
  38272=>"111111111",
  38273=>"111111111",
  38274=>"110111110",
  38275=>"000000000",
  38276=>"001111111",
  38277=>"000000000",
  38278=>"011001000",
  38279=>"001000000",
  38280=>"001000000",
  38281=>"111111111",
  38282=>"011001001",
  38283=>"010110111",
  38284=>"000011111",
  38285=>"111001001",
  38286=>"000000000",
  38287=>"000000000",
  38288=>"101001000",
  38289=>"000000100",
  38290=>"111111111",
  38291=>"110111111",
  38292=>"111011011",
  38293=>"000010000",
  38294=>"101000101",
  38295=>"100001001",
  38296=>"010000110",
  38297=>"111011001",
  38298=>"111111111",
  38299=>"110010000",
  38300=>"001000100",
  38301=>"111111100",
  38302=>"100100100",
  38303=>"111111111",
  38304=>"000011001",
  38305=>"100000000",
  38306=>"110110000",
  38307=>"000000000",
  38308=>"110110110",
  38309=>"001011011",
  38310=>"101100111",
  38311=>"000000000",
  38312=>"111000000",
  38313=>"100110110",
  38314=>"110011111",
  38315=>"111010000",
  38316=>"111000000",
  38317=>"110000101",
  38318=>"001011111",
  38319=>"011111111",
  38320=>"100110111",
  38321=>"111111111",
  38322=>"000000000",
  38323=>"110110110",
  38324=>"010000000",
  38325=>"010110110",
  38326=>"000000011",
  38327=>"110111111",
  38328=>"110110100",
  38329=>"110000000",
  38330=>"111111001",
  38331=>"111111111",
  38332=>"000110110",
  38333=>"100111111",
  38334=>"011011000",
  38335=>"001000101",
  38336=>"100011011",
  38337=>"001001001",
  38338=>"000111011",
  38339=>"000000000",
  38340=>"110111110",
  38341=>"111011010",
  38342=>"000000010",
  38343=>"100100110",
  38344=>"000000010",
  38345=>"000010000",
  38346=>"101111001",
  38347=>"110111111",
  38348=>"010000000",
  38349=>"000000111",
  38350=>"111110001",
  38351=>"111111110",
  38352=>"111111000",
  38353=>"000000001",
  38354=>"000000000",
  38355=>"000011111",
  38356=>"100010111",
  38357=>"000000100",
  38358=>"000001011",
  38359=>"011111011",
  38360=>"100100101",
  38361=>"000000001",
  38362=>"111000101",
  38363=>"111001000",
  38364=>"011111110",
  38365=>"010000000",
  38366=>"111111111",
  38367=>"100100100",
  38368=>"111111000",
  38369=>"111111111",
  38370=>"111100111",
  38371=>"111001001",
  38372=>"111000000",
  38373=>"011111111",
  38374=>"111111111",
  38375=>"110011010",
  38376=>"000000001",
  38377=>"111110110",
  38378=>"000000000",
  38379=>"000101111",
  38380=>"101101101",
  38381=>"100110000",
  38382=>"010111000",
  38383=>"000010010",
  38384=>"000001000",
  38385=>"001000000",
  38386=>"001000000",
  38387=>"000000000",
  38388=>"111111111",
  38389=>"111111111",
  38390=>"001011001",
  38391=>"000000000",
  38392=>"110000000",
  38393=>"000100000",
  38394=>"001000001",
  38395=>"000000000",
  38396=>"111111111",
  38397=>"000000000",
  38398=>"111001001",
  38399=>"101001111",
  38400=>"101111011",
  38401=>"000000000",
  38402=>"011111100",
  38403=>"011011000",
  38404=>"111100111",
  38405=>"000000001",
  38406=>"111111111",
  38407=>"000001001",
  38408=>"000000000",
  38409=>"111111111",
  38410=>"000000000",
  38411=>"001000010",
  38412=>"000000000",
  38413=>"011111110",
  38414=>"110111111",
  38415=>"111111111",
  38416=>"110000000",
  38417=>"111111111",
  38418=>"111101001",
  38419=>"101100000",
  38420=>"100100000",
  38421=>"011001000",
  38422=>"000000000",
  38423=>"100000000",
  38424=>"010000111",
  38425=>"001001011",
  38426=>"111110000",
  38427=>"111111000",
  38428=>"111111100",
  38429=>"111000000",
  38430=>"100110000",
  38431=>"000000100",
  38432=>"111111000",
  38433=>"111110000",
  38434=>"001000000",
  38435=>"000000000",
  38436=>"100011000",
  38437=>"111111111",
  38438=>"111111111",
  38439=>"100101111",
  38440=>"000000000",
  38441=>"000000000",
  38442=>"100000000",
  38443=>"110111000",
  38444=>"010000000",
  38445=>"000001010",
  38446=>"111111111",
  38447=>"111111101",
  38448=>"000110010",
  38449=>"111000000",
  38450=>"000000101",
  38451=>"111001101",
  38452=>"000111000",
  38453=>"000000000",
  38454=>"001101011",
  38455=>"000100100",
  38456=>"111111111",
  38457=>"000000000",
  38458=>"000000110",
  38459=>"000000000",
  38460=>"111111111",
  38461=>"000000000",
  38462=>"111111111",
  38463=>"111000000",
  38464=>"000000000",
  38465=>"110111111",
  38466=>"111101000",
  38467=>"000000000",
  38468=>"111000000",
  38469=>"111111001",
  38470=>"111000000",
  38471=>"000000000",
  38472=>"011001001",
  38473=>"111000000",
  38474=>"111111111",
  38475=>"001111011",
  38476=>"011011110",
  38477=>"110000000",
  38478=>"000000011",
  38479=>"000000011",
  38480=>"111111100",
  38481=>"111111111",
  38482=>"100110000",
  38483=>"000000000",
  38484=>"111000001",
  38485=>"111111111",
  38486=>"000010011",
  38487=>"000000100",
  38488=>"100111011",
  38489=>"000000000",
  38490=>"100000000",
  38491=>"110110000",
  38492=>"111111110",
  38493=>"111111111",
  38494=>"111111111",
  38495=>"011111100",
  38496=>"000001011",
  38497=>"111001000",
  38498=>"000000001",
  38499=>"110110110",
  38500=>"110010110",
  38501=>"110100000",
  38502=>"111111111",
  38503=>"111111001",
  38504=>"110000000",
  38505=>"000000000",
  38506=>"100110110",
  38507=>"000010010",
  38508=>"111111101",
  38509=>"111111111",
  38510=>"111111111",
  38511=>"000000000",
  38512=>"111000000",
  38513=>"100101000",
  38514=>"000111111",
  38515=>"011111100",
  38516=>"111111111",
  38517=>"000011011",
  38518=>"110111111",
  38519=>"111111000",
  38520=>"111111111",
  38521=>"111000100",
  38522=>"111111111",
  38523=>"111111111",
  38524=>"000010000",
  38525=>"000000111",
  38526=>"000000001",
  38527=>"001011011",
  38528=>"110110110",
  38529=>"111110000",
  38530=>"000000000",
  38531=>"111111111",
  38532=>"111111111",
  38533=>"110000100",
  38534=>"100101000",
  38535=>"111111111",
  38536=>"001011001",
  38537=>"001000000",
  38538=>"000000000",
  38539=>"111111111",
  38540=>"010111100",
  38541=>"001111111",
  38542=>"110110100",
  38543=>"100100010",
  38544=>"000000000",
  38545=>"111111111",
  38546=>"111111111",
  38547=>"111111001",
  38548=>"111111110",
  38549=>"001011011",
  38550=>"111111011",
  38551=>"110110000",
  38552=>"000000101",
  38553=>"111000001",
  38554=>"111110111",
  38555=>"111111111",
  38556=>"111110110",
  38557=>"101001001",
  38558=>"101110110",
  38559=>"000000000",
  38560=>"100000111",
  38561=>"111111000",
  38562=>"111000000",
  38563=>"111111111",
  38564=>"000000000",
  38565=>"101001000",
  38566=>"000000000",
  38567=>"011011011",
  38568=>"110111011",
  38569=>"000000000",
  38570=>"110100000",
  38571=>"011011111",
  38572=>"111000000",
  38573=>"111111111",
  38574=>"111111111",
  38575=>"111111111",
  38576=>"000100111",
  38577=>"111100110",
  38578=>"011001000",
  38579=>"000000000",
  38580=>"000001001",
  38581=>"000000000",
  38582=>"000000000",
  38583=>"000000000",
  38584=>"010100100",
  38585=>"111011000",
  38586=>"000000111",
  38587=>"000010001",
  38588=>"000000111",
  38589=>"100111001",
  38590=>"111111111",
  38591=>"011101100",
  38592=>"111111111",
  38593=>"111111111",
  38594=>"001111111",
  38595=>"010111111",
  38596=>"110111011",
  38597=>"111111000",
  38598=>"110110110",
  38599=>"111111110",
  38600=>"111100100",
  38601=>"000110110",
  38602=>"011000001",
  38603=>"001001000",
  38604=>"111111011",
  38605=>"111111111",
  38606=>"001001011",
  38607=>"111111111",
  38608=>"111011011",
  38609=>"010000000",
  38610=>"111001001",
  38611=>"001000000",
  38612=>"111000000",
  38613=>"111100000",
  38614=>"000000111",
  38615=>"001001000",
  38616=>"000000000",
  38617=>"000011111",
  38618=>"000000111",
  38619=>"111111110",
  38620=>"111100100",
  38621=>"111111011",
  38622=>"011011111",
  38623=>"001110110",
  38624=>"010110010",
  38625=>"000111111",
  38626=>"111111110",
  38627=>"101001001",
  38628=>"111100000",
  38629=>"111111111",
  38630=>"111111111",
  38631=>"111111011",
  38632=>"111001011",
  38633=>"001001111",
  38634=>"111111011",
  38635=>"111000000",
  38636=>"000000000",
  38637=>"111111111",
  38638=>"000111001",
  38639=>"000001000",
  38640=>"000000000",
  38641=>"111011000",
  38642=>"111111111",
  38643=>"000100100",
  38644=>"000110000",
  38645=>"010010000",
  38646=>"100000011",
  38647=>"000000001",
  38648=>"111111110",
  38649=>"001000100",
  38650=>"000000000",
  38651=>"010000000",
  38652=>"011011011",
  38653=>"000110110",
  38654=>"000000000",
  38655=>"111111001",
  38656=>"000000000",
  38657=>"000011011",
  38658=>"111111100",
  38659=>"110000000",
  38660=>"100110110",
  38661=>"000000000",
  38662=>"000000000",
  38663=>"000000000",
  38664=>"000000000",
  38665=>"110111110",
  38666=>"001001001",
  38667=>"000011111",
  38668=>"000000110",
  38669=>"111111110",
  38670=>"111010000",
  38671=>"000111111",
  38672=>"000010111",
  38673=>"000001111",
  38674=>"111000000",
  38675=>"000000001",
  38676=>"000011001",
  38677=>"110111111",
  38678=>"110100110",
  38679=>"110100101",
  38680=>"111111111",
  38681=>"000000000",
  38682=>"111010000",
  38683=>"111111010",
  38684=>"000011011",
  38685=>"000000000",
  38686=>"001111111",
  38687=>"001000001",
  38688=>"100101111",
  38689=>"000000011",
  38690=>"000000111",
  38691=>"111111000",
  38692=>"000000000",
  38693=>"000000000",
  38694=>"000000000",
  38695=>"000010000",
  38696=>"111011010",
  38697=>"111111111",
  38698=>"111111000",
  38699=>"000111111",
  38700=>"100111011",
  38701=>"111111111",
  38702=>"000000000",
  38703=>"000000000",
  38704=>"000000001",
  38705=>"001010000",
  38706=>"000000000",
  38707=>"000111111",
  38708=>"000000111",
  38709=>"000111111",
  38710=>"000000000",
  38711=>"111110000",
  38712=>"111111000",
  38713=>"100100100",
  38714=>"111111111",
  38715=>"110110101",
  38716=>"000000011",
  38717=>"111000001",
  38718=>"000000000",
  38719=>"110110000",
  38720=>"111111111",
  38721=>"110110100",
  38722=>"111111100",
  38723=>"110100111",
  38724=>"000000111",
  38725=>"110011011",
  38726=>"011111100",
  38727=>"000000000",
  38728=>"000000000",
  38729=>"100110000",
  38730=>"110000110",
  38731=>"010011110",
  38732=>"000000111",
  38733=>"000100111",
  38734=>"000010000",
  38735=>"011111111",
  38736=>"100101100",
  38737=>"000100011",
  38738=>"000100101",
  38739=>"000000110",
  38740=>"000000001",
  38741=>"011001001",
  38742=>"111111111",
  38743=>"000000000",
  38744=>"111111001",
  38745=>"000000000",
  38746=>"110100000",
  38747=>"111000001",
  38748=>"111101111",
  38749=>"111111111",
  38750=>"111111011",
  38751=>"110111111",
  38752=>"110000000",
  38753=>"111111111",
  38754=>"000000110",
  38755=>"000000100",
  38756=>"001011111",
  38757=>"001011111",
  38758=>"010011000",
  38759=>"111110110",
  38760=>"001000000",
  38761=>"111110010",
  38762=>"000000110",
  38763=>"011111111",
  38764=>"001001000",
  38765=>"100111111",
  38766=>"000000000",
  38767=>"010010000",
  38768=>"000000000",
  38769=>"100000000",
  38770=>"000000000",
  38771=>"001001011",
  38772=>"000000101",
  38773=>"000000110",
  38774=>"000000111",
  38775=>"000100000",
  38776=>"011111000",
  38777=>"000000011",
  38778=>"001111111",
  38779=>"000000111",
  38780=>"000000110",
  38781=>"000000001",
  38782=>"001011001",
  38783=>"111111110",
  38784=>"000000000",
  38785=>"110110111",
  38786=>"111000000",
  38787=>"111111100",
  38788=>"000100000",
  38789=>"111011000",
  38790=>"111111010",
  38791=>"111000000",
  38792=>"111111110",
  38793=>"000110000",
  38794=>"001001111",
  38795=>"000000110",
  38796=>"111111111",
  38797=>"011011000",
  38798=>"000001011",
  38799=>"000110110",
  38800=>"111111111",
  38801=>"111001011",
  38802=>"010011111",
  38803=>"000000000",
  38804=>"111111111",
  38805=>"000000000",
  38806=>"011010000",
  38807=>"000000001",
  38808=>"011000000",
  38809=>"100100110",
  38810=>"101111111",
  38811=>"000000000",
  38812=>"000000000",
  38813=>"111111011",
  38814=>"110000010",
  38815=>"000000001",
  38816=>"100100101",
  38817=>"111111111",
  38818=>"100010001",
  38819=>"000000000",
  38820=>"000000110",
  38821=>"111111001",
  38822=>"000000000",
  38823=>"110110110",
  38824=>"000010000",
  38825=>"000000000",
  38826=>"111111011",
  38827=>"001111111",
  38828=>"000000000",
  38829=>"001001111",
  38830=>"111110010",
  38831=>"000000000",
  38832=>"100100000",
  38833=>"111111111",
  38834=>"101111111",
  38835=>"000111111",
  38836=>"000010110",
  38837=>"000000000",
  38838=>"010010000",
  38839=>"111011011",
  38840=>"111011001",
  38841=>"111111011",
  38842=>"111100010",
  38843=>"001000000",
  38844=>"000000000",
  38845=>"110100000",
  38846=>"000000011",
  38847=>"010010010",
  38848=>"001111111",
  38849=>"110000111",
  38850=>"000000000",
  38851=>"110100000",
  38852=>"000100110",
  38853=>"110100100",
  38854=>"110010000",
  38855=>"010000000",
  38856=>"000000001",
  38857=>"000000110",
  38858=>"100100100",
  38859=>"000000000",
  38860=>"111101111",
  38861=>"010000000",
  38862=>"111110110",
  38863=>"011111111",
  38864=>"011111111",
  38865=>"000000100",
  38866=>"011111111",
  38867=>"111111111",
  38868=>"011001111",
  38869=>"111111111",
  38870=>"011111111",
  38871=>"100000100",
  38872=>"000001001",
  38873=>"111100011",
  38874=>"000000000",
  38875=>"110100000",
  38876=>"001011111",
  38877=>"000000000",
  38878=>"000000000",
  38879=>"001011001",
  38880=>"000000000",
  38881=>"111111110",
  38882=>"000000110",
  38883=>"111101111",
  38884=>"111111111",
  38885=>"111111111",
  38886=>"010110110",
  38887=>"000000110",
  38888=>"111111101",
  38889=>"111110111",
  38890=>"000100111",
  38891=>"000000000",
  38892=>"111100000",
  38893=>"101111011",
  38894=>"000000100",
  38895=>"111111000",
  38896=>"000000000",
  38897=>"100111111",
  38898=>"111111001",
  38899=>"000000001",
  38900=>"000000000",
  38901=>"001111111",
  38902=>"000000000",
  38903=>"001001111",
  38904=>"000000110",
  38905=>"100100110",
  38906=>"111011001",
  38907=>"110110111",
  38908=>"000111111",
  38909=>"111110110",
  38910=>"111011011",
  38911=>"000000001",
  38912=>"111011011",
  38913=>"000000111",
  38914=>"000000000",
  38915=>"000000111",
  38916=>"111100100",
  38917=>"111001000",
  38918=>"001000000",
  38919=>"111111111",
  38920=>"000000000",
  38921=>"111010000",
  38922=>"110111001",
  38923=>"101111110",
  38924=>"100110010",
  38925=>"000000001",
  38926=>"111111000",
  38927=>"000000111",
  38928=>"111000111",
  38929=>"010110111",
  38930=>"000000000",
  38931=>"111100111",
  38932=>"110000110",
  38933=>"000000000",
  38934=>"001101111",
  38935=>"000111111",
  38936=>"001111111",
  38937=>"000000100",
  38938=>"001000000",
  38939=>"001011100",
  38940=>"100000000",
  38941=>"000001000",
  38942=>"111111111",
  38943=>"111111110",
  38944=>"111000110",
  38945=>"000000011",
  38946=>"110111000",
  38947=>"111101001",
  38948=>"000100111",
  38949=>"111111000",
  38950=>"000100000",
  38951=>"000000111",
  38952=>"110111111",
  38953=>"000100111",
  38954=>"111111000",
  38955=>"111111011",
  38956=>"000000000",
  38957=>"000000000",
  38958=>"101001001",
  38959=>"011000000",
  38960=>"111001111",
  38961=>"000000000",
  38962=>"001001011",
  38963=>"000000101",
  38964=>"111111001",
  38965=>"111011011",
  38966=>"111111000",
  38967=>"001000000",
  38968=>"000000111",
  38969=>"111111111",
  38970=>"010010110",
  38971=>"000000000",
  38972=>"111001001",
  38973=>"101111111",
  38974=>"001001111",
  38975=>"000000000",
  38976=>"000000010",
  38977=>"111111001",
  38978=>"111000111",
  38979=>"000111111",
  38980=>"111001000",
  38981=>"110111110",
  38982=>"000110110",
  38983=>"011000000",
  38984=>"111111100",
  38985=>"111111110",
  38986=>"111111011",
  38987=>"001001000",
  38988=>"001001000",
  38989=>"001000100",
  38990=>"000110100",
  38991=>"111111001",
  38992=>"000000100",
  38993=>"111111111",
  38994=>"111111000",
  38995=>"001001001",
  38996=>"001000000",
  38997=>"101110100",
  38998=>"111111001",
  38999=>"001001001",
  39000=>"001100110",
  39001=>"111001111",
  39002=>"010010011",
  39003=>"000000000",
  39004=>"100111111",
  39005=>"001000111",
  39006=>"000001000",
  39007=>"011011000",
  39008=>"000100111",
  39009=>"000110000",
  39010=>"000011010",
  39011=>"110011000",
  39012=>"110111110",
  39013=>"001001011",
  39014=>"011001000",
  39015=>"000000000",
  39016=>"110000000",
  39017=>"111001111",
  39018=>"111111110",
  39019=>"000000000",
  39020=>"001001111",
  39021=>"010111111",
  39022=>"101101111",
  39023=>"001000000",
  39024=>"100111100",
  39025=>"000000000",
  39026=>"111111000",
  39027=>"000010110",
  39028=>"111111010",
  39029=>"111111111",
  39030=>"000011111",
  39031=>"111111111",
  39032=>"000000000",
  39033=>"000000100",
  39034=>"001000000",
  39035=>"000111111",
  39036=>"000100000",
  39037=>"001001111",
  39038=>"000000000",
  39039=>"000000000",
  39040=>"000000000",
  39041=>"111111100",
  39042=>"000111110",
  39043=>"001111110",
  39044=>"000001111",
  39045=>"111001000",
  39046=>"111111000",
  39047=>"111011011",
  39048=>"110001011",
  39049=>"110111111",
  39050=>"110110111",
  39051=>"111111111",
  39052=>"111111110",
  39053=>"001111111",
  39054=>"011011111",
  39055=>"000100000",
  39056=>"111111111",
  39057=>"111111111",
  39058=>"000000001",
  39059=>"000101111",
  39060=>"111111111",
  39061=>"111111111",
  39062=>"111000000",
  39063=>"000000100",
  39064=>"000000000",
  39065=>"111111010",
  39066=>"000000000",
  39067=>"110100100",
  39068=>"010011111",
  39069=>"000000011",
  39070=>"111111101",
  39071=>"100100100",
  39072=>"001111000",
  39073=>"111000000",
  39074=>"011000000",
  39075=>"111111110",
  39076=>"001001001",
  39077=>"000011111",
  39078=>"011000100",
  39079=>"100110110",
  39080=>"111111111",
  39081=>"000000111",
  39082=>"111000011",
  39083=>"111111111",
  39084=>"111111000",
  39085=>"000100111",
  39086=>"001000001",
  39087=>"000010111",
  39088=>"110111111",
  39089=>"000000000",
  39090=>"111111111",
  39091=>"000000000",
  39092=>"000000000",
  39093=>"000000100",
  39094=>"000001111",
  39095=>"010110000",
  39096=>"111111000",
  39097=>"111111101",
  39098=>"000000000",
  39099=>"001000000",
  39100=>"000000000",
  39101=>"110111000",
  39102=>"011011011",
  39103=>"001000000",
  39104=>"001000100",
  39105=>"111111111",
  39106=>"111111111",
  39107=>"000000110",
  39108=>"011111111",
  39109=>"001011011",
  39110=>"000000000",
  39111=>"101110111",
  39112=>"001000111",
  39113=>"111001101",
  39114=>"101111000",
  39115=>"000000000",
  39116=>"000111110",
  39117=>"000000000",
  39118=>"111111000",
  39119=>"000000000",
  39120=>"111010000",
  39121=>"111100100",
  39122=>"011111111",
  39123=>"000100000",
  39124=>"000000000",
  39125=>"110111001",
  39126=>"000000000",
  39127=>"000000000",
  39128=>"100110100",
  39129=>"000000100",
  39130=>"011111111",
  39131=>"000000000",
  39132=>"011011001",
  39133=>"001011111",
  39134=>"111111111",
  39135=>"111111110",
  39136=>"000110000",
  39137=>"000000000",
  39138=>"000011000",
  39139=>"000000000",
  39140=>"000110111",
  39141=>"000001011",
  39142=>"111110111",
  39143=>"110111000",
  39144=>"000000111",
  39145=>"111111110",
  39146=>"101000101",
  39147=>"000000001",
  39148=>"000111111",
  39149=>"000111111",
  39150=>"011000110",
  39151=>"000000000",
  39152=>"000110000",
  39153=>"111000000",
  39154=>"000001111",
  39155=>"111101000",
  39156=>"011001111",
  39157=>"100110000",
  39158=>"010111110",
  39159=>"000000001",
  39160=>"000000000",
  39161=>"000000111",
  39162=>"110111000",
  39163=>"111011001",
  39164=>"001001001",
  39165=>"001111000",
  39166=>"001111000",
  39167=>"000000000",
  39168=>"000110111",
  39169=>"111100111",
  39170=>"111001111",
  39171=>"000110000",
  39172=>"001000111",
  39173=>"100110000",
  39174=>"111111100",
  39175=>"111111011",
  39176=>"000000111",
  39177=>"110111111",
  39178=>"010000111",
  39179=>"001000000",
  39180=>"001001011",
  39181=>"001011011",
  39182=>"111111000",
  39183=>"000001000",
  39184=>"001101001",
  39185=>"110111111",
  39186=>"111011111",
  39187=>"000000000",
  39188=>"000000000",
  39189=>"000100000",
  39190=>"001001001",
  39191=>"011100100",
  39192=>"111111001",
  39193=>"011011011",
  39194=>"111111111",
  39195=>"000111001",
  39196=>"110110000",
  39197=>"110000000",
  39198=>"001000100",
  39199=>"111100101",
  39200=>"000001111",
  39201=>"001000000",
  39202=>"111011011",
  39203=>"111111111",
  39204=>"000100100",
  39205=>"000100000",
  39206=>"001000000",
  39207=>"000111011",
  39208=>"000000000",
  39209=>"000000000",
  39210=>"100000000",
  39211=>"111001101",
  39212=>"110110111",
  39213=>"001111011",
  39214=>"111110110",
  39215=>"100111000",
  39216=>"000111111",
  39217=>"111111000",
  39218=>"000011001",
  39219=>"111111111",
  39220=>"100000000",
  39221=>"000000011",
  39222=>"011000000",
  39223=>"000111111",
  39224=>"000000100",
  39225=>"111001111",
  39226=>"001000111",
  39227=>"101000000",
  39228=>"001111111",
  39229=>"001100100",
  39230=>"000100111",
  39231=>"000000000",
  39232=>"111111000",
  39233=>"101101111",
  39234=>"000000111",
  39235=>"111001000",
  39236=>"011010000",
  39237=>"000110110",
  39238=>"000001111",
  39239=>"000000000",
  39240=>"110111110",
  39241=>"000010000",
  39242=>"110110000",
  39243=>"000101101",
  39244=>"111100110",
  39245=>"111111111",
  39246=>"000001101",
  39247=>"000001001",
  39248=>"111111111",
  39249=>"001101100",
  39250=>"000000111",
  39251=>"111111111",
  39252=>"000000000",
  39253=>"011011111",
  39254=>"000000101",
  39255=>"100111111",
  39256=>"000111000",
  39257=>"000000010",
  39258=>"101101111",
  39259=>"000000001",
  39260=>"000000010",
  39261=>"111111111",
  39262=>"000000001",
  39263=>"110111000",
  39264=>"011011011",
  39265=>"001101111",
  39266=>"100111111",
  39267=>"001101111",
  39268=>"011011001",
  39269=>"000000001",
  39270=>"110010011",
  39271=>"101001000",
  39272=>"100100000",
  39273=>"111111111",
  39274=>"111111111",
  39275=>"110000000",
  39276=>"111001000",
  39277=>"000100000",
  39278=>"110111110",
  39279=>"111000100",
  39280=>"000000000",
  39281=>"111110111",
  39282=>"111111111",
  39283=>"111110100",
  39284=>"010000000",
  39285=>"111001110",
  39286=>"001111111",
  39287=>"110100000",
  39288=>"001000100",
  39289=>"011111111",
  39290=>"001001001",
  39291=>"111111111",
  39292=>"000000111",
  39293=>"111111111",
  39294=>"001000000",
  39295=>"000000000",
  39296=>"110111000",
  39297=>"011000000",
  39298=>"001001000",
  39299=>"111000111",
  39300=>"001111111",
  39301=>"100000111",
  39302=>"111100000",
  39303=>"110111111",
  39304=>"000000000",
  39305=>"100111111",
  39306=>"000100100",
  39307=>"000010000",
  39308=>"111000000",
  39309=>"111111111",
  39310=>"110111011",
  39311=>"000000000",
  39312=>"000000100",
  39313=>"111011001",
  39314=>"000100000",
  39315=>"001111111",
  39316=>"000000111",
  39317=>"000010000",
  39318=>"001000000",
  39319=>"000101001",
  39320=>"000111111",
  39321=>"111111010",
  39322=>"000000111",
  39323=>"000000000",
  39324=>"000000111",
  39325=>"001111111",
  39326=>"111101001",
  39327=>"111111111",
  39328=>"011000000",
  39329=>"110100000",
  39330=>"111000000",
  39331=>"111110000",
  39332=>"111111111",
  39333=>"000011001",
  39334=>"001000001",
  39335=>"111000000",
  39336=>"000000000",
  39337=>"001000000",
  39338=>"000000000",
  39339=>"101001101",
  39340=>"010110110",
  39341=>"000111110",
  39342=>"100100000",
  39343=>"111111111",
  39344=>"000100110",
  39345=>"111111111",
  39346=>"111111101",
  39347=>"000000000",
  39348=>"101101101",
  39349=>"000000000",
  39350=>"001000100",
  39351=>"001000111",
  39352=>"000001001",
  39353=>"001000001",
  39354=>"010110010",
  39355=>"001000000",
  39356=>"000000000",
  39357=>"110111111",
  39358=>"101001000",
  39359=>"100100101",
  39360=>"000000000",
  39361=>"111101111",
  39362=>"000000000",
  39363=>"000000000",
  39364=>"111111001",
  39365=>"100011011",
  39366=>"000000111",
  39367=>"111111000",
  39368=>"000000001",
  39369=>"000000000",
  39370=>"000000010",
  39371=>"000000111",
  39372=>"111110111",
  39373=>"110111001",
  39374=>"000110100",
  39375=>"000000000",
  39376=>"111111100",
  39377=>"111111111",
  39378=>"101000000",
  39379=>"111111111",
  39380=>"111111101",
  39381=>"000000000",
  39382=>"000000101",
  39383=>"011111110",
  39384=>"000000000",
  39385=>"000000000",
  39386=>"111111111",
  39387=>"111110111",
  39388=>"001000000",
  39389=>"001001000",
  39390=>"011011111",
  39391=>"100111111",
  39392=>"000001111",
  39393=>"111111111",
  39394=>"000000000",
  39395=>"010000100",
  39396=>"111001001",
  39397=>"110000000",
  39398=>"000000000",
  39399=>"110000000",
  39400=>"111111111",
  39401=>"111111001",
  39402=>"111110101",
  39403=>"000000100",
  39404=>"000000000",
  39405=>"000000100",
  39406=>"111111111",
  39407=>"011010001",
  39408=>"101000000",
  39409=>"111111000",
  39410=>"000001001",
  39411=>"000000100",
  39412=>"011000000",
  39413=>"000111110",
  39414=>"000100110",
  39415=>"000000000",
  39416=>"000000000",
  39417=>"000001000",
  39418=>"111000000",
  39419=>"000110111",
  39420=>"000000000",
  39421=>"111000001",
  39422=>"000101000",
  39423=>"000000000",
  39424=>"000000011",
  39425=>"111111110",
  39426=>"111111010",
  39427=>"111001111",
  39428=>"110110000",
  39429=>"000100000",
  39430=>"110110100",
  39431=>"011001001",
  39432=>"000001000",
  39433=>"000001001",
  39434=>"011001001",
  39435=>"111111111",
  39436=>"011001001",
  39437=>"110110111",
  39438=>"100000100",
  39439=>"111001111",
  39440=>"111111011",
  39441=>"111111111",
  39442=>"000100000",
  39443=>"111011011",
  39444=>"100111111",
  39445=>"111111111",
  39446=>"110110111",
  39447=>"100100101",
  39448=>"010010000",
  39449=>"111001011",
  39450=>"011000000",
  39451=>"111011111",
  39452=>"000101011",
  39453=>"000000100",
  39454=>"000100111",
  39455=>"000010011",
  39456=>"000001101",
  39457=>"000000000",
  39458=>"001111011",
  39459=>"110110010",
  39460=>"011011011",
  39461=>"000101111",
  39462=>"100100000",
  39463=>"000110111",
  39464=>"110010000",
  39465=>"111111111",
  39466=>"111111111",
  39467=>"111110000",
  39468=>"000111010",
  39469=>"111111110",
  39470=>"111110111",
  39471=>"111111111",
  39472=>"011011111",
  39473=>"000000001",
  39474=>"010100000",
  39475=>"111111111",
  39476=>"001011011",
  39477=>"010000000",
  39478=>"111001000",
  39479=>"101111001",
  39480=>"010111011",
  39481=>"111111011",
  39482=>"100000000",
  39483=>"000000000",
  39484=>"111111111",
  39485=>"110100101",
  39486=>"111111111",
  39487=>"111111111",
  39488=>"011000000",
  39489=>"011001001",
  39490=>"110100011",
  39491=>"100100111",
  39492=>"010001001",
  39493=>"111111111",
  39494=>"111110000",
  39495=>"111111011",
  39496=>"000000010",
  39497=>"000000111",
  39498=>"111111011",
  39499=>"101100000",
  39500=>"000001111",
  39501=>"110111001",
  39502=>"111100100",
  39503=>"000010000",
  39504=>"100110011",
  39505=>"001011010",
  39506=>"111001000",
  39507=>"000000000",
  39508=>"111111110",
  39509=>"100100111",
  39510=>"101000011",
  39511=>"000000000",
  39512=>"000000010",
  39513=>"111111111",
  39514=>"100000000",
  39515=>"100101011",
  39516=>"110111111",
  39517=>"111011000",
  39518=>"100110111",
  39519=>"000000100",
  39520=>"010000111",
  39521=>"001000001",
  39522=>"000000000",
  39523=>"000000001",
  39524=>"011000000",
  39525=>"011011011",
  39526=>"101111111",
  39527=>"111111110",
  39528=>"000000111",
  39529=>"000011000",
  39530=>"111111111",
  39531=>"100100110",
  39532=>"000000111",
  39533=>"010000000",
  39534=>"111111111",
  39535=>"111000100",
  39536=>"001001000",
  39537=>"011011000",
  39538=>"000000001",
  39539=>"110111001",
  39540=>"111111111",
  39541=>"100100001",
  39542=>"001111111",
  39543=>"111111111",
  39544=>"000000011",
  39545=>"111001001",
  39546=>"110110000",
  39547=>"111100000",
  39548=>"111011111",
  39549=>"111011000",
  39550=>"111111011",
  39551=>"110111111",
  39552=>"000000000",
  39553=>"101111000",
  39554=>"111001000",
  39555=>"101101111",
  39556=>"111000011",
  39557=>"000000001",
  39558=>"010010010",
  39559=>"010000110",
  39560=>"000110010",
  39561=>"000000000",
  39562=>"100101101",
  39563=>"000000001",
  39564=>"011111011",
  39565=>"111111110",
  39566=>"011010111",
  39567=>"111111001",
  39568=>"000001001",
  39569=>"111111111",
  39570=>"000000110",
  39571=>"110111111",
  39572=>"001001111",
  39573=>"111111001",
  39574=>"000000110",
  39575=>"000000000",
  39576=>"111010011",
  39577=>"110010010",
  39578=>"111111110",
  39579=>"000000110",
  39580=>"111111111",
  39581=>"111111011",
  39582=>"111111111",
  39583=>"110100000",
  39584=>"111100111",
  39585=>"011111111",
  39586=>"111111111",
  39587=>"000000000",
  39588=>"110111000",
  39589=>"100100110",
  39590=>"001000000",
  39591=>"101101101",
  39592=>"100000000",
  39593=>"001000010",
  39594=>"000111010",
  39595=>"011111111",
  39596=>"110110011",
  39597=>"001001001",
  39598=>"000000010",
  39599=>"001011011",
  39600=>"111111111",
  39601=>"100100100",
  39602=>"101001001",
  39603=>"111111111",
  39604=>"111001000",
  39605=>"110110001",
  39606=>"000000000",
  39607=>"110111011",
  39608=>"000101111",
  39609=>"010110110",
  39610=>"110110110",
  39611=>"011111111",
  39612=>"000010011",
  39613=>"110100001",
  39614=>"010000000",
  39615=>"111111001",
  39616=>"111111111",
  39617=>"111000000",
  39618=>"000000000",
  39619=>"000110000",
  39620=>"011110001",
  39621=>"000011111",
  39622=>"110100000",
  39623=>"000000011",
  39624=>"000010000",
  39625=>"000001011",
  39626=>"111111010",
  39627=>"000100111",
  39628=>"111000000",
  39629=>"001111110",
  39630=>"000000000",
  39631=>"000000001",
  39632=>"111100100",
  39633=>"111111111",
  39634=>"001000000",
  39635=>"000000000",
  39636=>"111001100",
  39637=>"001111101",
  39638=>"011010010",
  39639=>"111111011",
  39640=>"000000000",
  39641=>"011000011",
  39642=>"000100101",
  39643=>"000000011",
  39644=>"000000001",
  39645=>"100000000",
  39646=>"111011001",
  39647=>"110100001",
  39648=>"001000000",
  39649=>"001101111",
  39650=>"111011010",
  39651=>"111100101",
  39652=>"000000000",
  39653=>"000001001",
  39654=>"000000000",
  39655=>"110110010",
  39656=>"111001111",
  39657=>"111111111",
  39658=>"111011111",
  39659=>"111111111",
  39660=>"111111111",
  39661=>"000000111",
  39662=>"111111111",
  39663=>"000000000",
  39664=>"011010111",
  39665=>"110000111",
  39666=>"000111010",
  39667=>"000000011",
  39668=>"010110111",
  39669=>"011011111",
  39670=>"101101111",
  39671=>"010000000",
  39672=>"111111111",
  39673=>"111001011",
  39674=>"111101111",
  39675=>"011111111",
  39676=>"000010110",
  39677=>"001000000",
  39678=>"110000010",
  39679=>"011010010",
  39680=>"101000000",
  39681=>"101100100",
  39682=>"011000000",
  39683=>"111000000",
  39684=>"000001111",
  39685=>"001000100",
  39686=>"000000000",
  39687=>"001011111",
  39688=>"110100011",
  39689=>"010000000",
  39690=>"111011111",
  39691=>"000000010",
  39692=>"011111010",
  39693=>"001001001",
  39694=>"000000111",
  39695=>"011000000",
  39696=>"011011011",
  39697=>"111001001",
  39698=>"000000111",
  39699=>"000000000",
  39700=>"000000111",
  39701=>"000011111",
  39702=>"101001111",
  39703=>"110000000",
  39704=>"011001101",
  39705=>"110000011",
  39706=>"100101000",
  39707=>"011111001",
  39708=>"000011011",
  39709=>"110011001",
  39710=>"000011111",
  39711=>"011001001",
  39712=>"001001101",
  39713=>"111111110",
  39714=>"111111111",
  39715=>"011011000",
  39716=>"111110110",
  39717=>"111111111",
  39718=>"111101100",
  39719=>"111111111",
  39720=>"111111111",
  39721=>"000001111",
  39722=>"001111111",
  39723=>"000000011",
  39724=>"100000000",
  39725=>"010010110",
  39726=>"000000111",
  39727=>"110010010",
  39728=>"000111111",
  39729=>"110010010",
  39730=>"001001001",
  39731=>"011111111",
  39732=>"001001000",
  39733=>"111011010",
  39734=>"111110000",
  39735=>"101001000",
  39736=>"010000000",
  39737=>"110000000",
  39738=>"000000110",
  39739=>"110000000",
  39740=>"110110111",
  39741=>"111111111",
  39742=>"110110110",
  39743=>"000000000",
  39744=>"111011011",
  39745=>"000000110",
  39746=>"101001011",
  39747=>"000110111",
  39748=>"100001000",
  39749=>"111111111",
  39750=>"010110110",
  39751=>"000000000",
  39752=>"110111101",
  39753=>"000111111",
  39754=>"111011011",
  39755=>"010011011",
  39756=>"110110000",
  39757=>"110111101",
  39758=>"101101101",
  39759=>"100010000",
  39760=>"011010000",
  39761=>"110011011",
  39762=>"001001111",
  39763=>"111110000",
  39764=>"000001000",
  39765=>"001000110",
  39766=>"101000000",
  39767=>"000000000",
  39768=>"000001001",
  39769=>"000000000",
  39770=>"100000100",
  39771=>"110100111",
  39772=>"010111111",
  39773=>"111111111",
  39774=>"111011001",
  39775=>"100000001",
  39776=>"111001011",
  39777=>"111111111",
  39778=>"110000001",
  39779=>"000000000",
  39780=>"000111111",
  39781=>"101111111",
  39782=>"001100110",
  39783=>"000000011",
  39784=>"001001111",
  39785=>"111011010",
  39786=>"001011000",
  39787=>"101001101",
  39788=>"110110111",
  39789=>"010110110",
  39790=>"000010000",
  39791=>"111001001",
  39792=>"111100111",
  39793=>"111111111",
  39794=>"000000000",
  39795=>"101000000",
  39796=>"110101000",
  39797=>"111111011",
  39798=>"111111011",
  39799=>"101001001",
  39800=>"111111111",
  39801=>"001001101",
  39802=>"100100111",
  39803=>"111001000",
  39804=>"000000111",
  39805=>"000000000",
  39806=>"111111011",
  39807=>"010001000",
  39808=>"101100000",
  39809=>"000000001",
  39810=>"111111111",
  39811=>"111101000",
  39812=>"000110000",
  39813=>"000010010",
  39814=>"111100111",
  39815=>"011010000",
  39816=>"000011111",
  39817=>"111011000",
  39818=>"000011010",
  39819=>"011011000",
  39820=>"000000000",
  39821=>"101001101",
  39822=>"111111001",
  39823=>"000000001",
  39824=>"011111011",
  39825=>"000110000",
  39826=>"111010011",
  39827=>"111001001",
  39828=>"111111110",
  39829=>"101111111",
  39830=>"111000000",
  39831=>"000000000",
  39832=>"000000000",
  39833=>"010000001",
  39834=>"110000000",
  39835=>"100000001",
  39836=>"000000100",
  39837=>"000011111",
  39838=>"110110110",
  39839=>"111111111",
  39840=>"110010000",
  39841=>"001101111",
  39842=>"001000000",
  39843=>"111111000",
  39844=>"100000000",
  39845=>"000000110",
  39846=>"000010111",
  39847=>"111111100",
  39848=>"000011001",
  39849=>"111111111",
  39850=>"111111111",
  39851=>"110001000",
  39852=>"000000000",
  39853=>"001001111",
  39854=>"000010000",
  39855=>"111101001",
  39856=>"111101111",
  39857=>"001111000",
  39858=>"011001111",
  39859=>"100100100",
  39860=>"111111111",
  39861=>"011111111",
  39862=>"100011111",
  39863=>"000000000",
  39864=>"111111111",
  39865=>"001101100",
  39866=>"110110000",
  39867=>"011011111",
  39868=>"010000000",
  39869=>"110010011",
  39870=>"001000000",
  39871=>"100101101",
  39872=>"111111001",
  39873=>"011011000",
  39874=>"111000000",
  39875=>"000000000",
  39876=>"101010010",
  39877=>"111011000",
  39878=>"000000010",
  39879=>"011000000",
  39880=>"110001001",
  39881=>"110011111",
  39882=>"111000000",
  39883=>"001111111",
  39884=>"000000000",
  39885=>"000001011",
  39886=>"011001111",
  39887=>"100100110",
  39888=>"001000000",
  39889=>"001011001",
  39890=>"000000000",
  39891=>"100100000",
  39892=>"000000000",
  39893=>"111001111",
  39894=>"100111111",
  39895=>"101101111",
  39896=>"101001011",
  39897=>"111101011",
  39898=>"010110110",
  39899=>"010010110",
  39900=>"011111111",
  39901=>"100111111",
  39902=>"100110111",
  39903=>"110110110",
  39904=>"000001001",
  39905=>"000000000",
  39906=>"010100110",
  39907=>"111110011",
  39908=>"111110110",
  39909=>"111101100",
  39910=>"000001011",
  39911=>"111111100",
  39912=>"000000001",
  39913=>"000000000",
  39914=>"011111111",
  39915=>"110100000",
  39916=>"010111111",
  39917=>"100100001",
  39918=>"001001111",
  39919=>"011000000",
  39920=>"000010111",
  39921=>"000101111",
  39922=>"111000000",
  39923=>"000000000",
  39924=>"100000000",
  39925=>"100110110",
  39926=>"000000000",
  39927=>"000001111",
  39928=>"011000000",
  39929=>"011010010",
  39930=>"111011111",
  39931=>"011001111",
  39932=>"001010010",
  39933=>"011001111",
  39934=>"001001101",
  39935=>"001000000",
  39936=>"110000010",
  39937=>"111000000",
  39938=>"100100000",
  39939=>"111000000",
  39940=>"011000111",
  39941=>"000111001",
  39942=>"100110100",
  39943=>"111111111",
  39944=>"111111111",
  39945=>"111111111",
  39946=>"000000000",
  39947=>"111111111",
  39948=>"101100000",
  39949=>"101001000",
  39950=>"001011001",
  39951=>"111100001",
  39952=>"110000001",
  39953=>"111111000",
  39954=>"000000000",
  39955=>"000100100",
  39956=>"111110110",
  39957=>"000000111",
  39958=>"000000110",
  39959=>"111100001",
  39960=>"000000001",
  39961=>"001001000",
  39962=>"011000000",
  39963=>"111000000",
  39964=>"000011111",
  39965=>"001000011",
  39966=>"111111011",
  39967=>"000000000",
  39968=>"000010000",
  39969=>"000001111",
  39970=>"110111111",
  39971=>"111111111",
  39972=>"000000000",
  39973=>"101100111",
  39974=>"000001111",
  39975=>"000100101",
  39976=>"001001111",
  39977=>"000000000",
  39978=>"011011001",
  39979=>"111001001",
  39980=>"111111101",
  39981=>"000000000",
  39982=>"000000111",
  39983=>"111111000",
  39984=>"111111111",
  39985=>"000000110",
  39986=>"000110110",
  39987=>"111111111",
  39988=>"000011011",
  39989=>"110111111",
  39990=>"111110000",
  39991=>"001111110",
  39992=>"111110000",
  39993=>"111011001",
  39994=>"000000000",
  39995=>"100110111",
  39996=>"111000000",
  39997=>"000000000",
  39998=>"100100001",
  39999=>"000000111",
  40000=>"111111000",
  40001=>"001001111",
  40002=>"011011000",
  40003=>"001101000",
  40004=>"000000000",
  40005=>"100100110",
  40006=>"101101000",
  40007=>"110111111",
  40008=>"001011110",
  40009=>"101000101",
  40010=>"111111111",
  40011=>"010011111",
  40012=>"111000010",
  40013=>"111111000",
  40014=>"000000001",
  40015=>"000000000",
  40016=>"000000111",
  40017=>"000000000",
  40018=>"000000000",
  40019=>"110111010",
  40020=>"001000000",
  40021=>"100000000",
  40022=>"001000101",
  40023=>"000000000",
  40024=>"111001001",
  40025=>"110000001",
  40026=>"000001110",
  40027=>"110100000",
  40028=>"001000000",
  40029=>"000111111",
  40030=>"011011111",
  40031=>"000110100",
  40032=>"000000000",
  40033=>"111000000",
  40034=>"001101001",
  40035=>"111000000",
  40036=>"000000000",
  40037=>"000000111",
  40038=>"001000000",
  40039=>"100000111",
  40040=>"011111111",
  40041=>"000111111",
  40042=>"000000111",
  40043=>"000000000",
  40044=>"000100110",
  40045=>"110000100",
  40046=>"111111000",
  40047=>"111111110",
  40048=>"111111111",
  40049=>"111111000",
  40050=>"111101111",
  40051=>"110110000",
  40052=>"111111111",
  40053=>"000000001",
  40054=>"000000000",
  40055=>"000100100",
  40056=>"111000000",
  40057=>"001000000",
  40058=>"000000000",
  40059=>"111000000",
  40060=>"010111110",
  40061=>"000000000",
  40062=>"000000000",
  40063=>"000100100",
  40064=>"000000100",
  40065=>"111100000",
  40066=>"010010111",
  40067=>"001000111",
  40068=>"111111111",
  40069=>"000000101",
  40070=>"000100111",
  40071=>"100000000",
  40072=>"000000011",
  40073=>"000000001",
  40074=>"000000111",
  40075=>"100111111",
  40076=>"111000011",
  40077=>"111111010",
  40078=>"111111111",
  40079=>"111100000",
  40080=>"001111000",
  40081=>"111000000",
  40082=>"111111000",
  40083=>"001011111",
  40084=>"000000000",
  40085=>"000000000",
  40086=>"101111100",
  40087=>"111000000",
  40088=>"111111101",
  40089=>"111110100",
  40090=>"000111111",
  40091=>"011011011",
  40092=>"000111111",
  40093=>"111000001",
  40094=>"000000000",
  40095=>"000000011",
  40096=>"100000000",
  40097=>"000000000",
  40098=>"000000000",
  40099=>"011111111",
  40100=>"001000000",
  40101=>"101011011",
  40102=>"110110110",
  40103=>"011001001",
  40104=>"111011000",
  40105=>"101000000",
  40106=>"111111000",
  40107=>"111111111",
  40108=>"000000000",
  40109=>"110010000",
  40110=>"111000000",
  40111=>"000101101",
  40112=>"000100001",
  40113=>"010110111",
  40114=>"101111111",
  40115=>"011000000",
  40116=>"111001000",
  40117=>"111100111",
  40118=>"000000111",
  40119=>"001000000",
  40120=>"111111111",
  40121=>"001000000",
  40122=>"000000010",
  40123=>"111001111",
  40124=>"111111000",
  40125=>"111111111",
  40126=>"111111101",
  40127=>"000000111",
  40128=>"011111000",
  40129=>"000001111",
  40130=>"011011001",
  40131=>"000000000",
  40132=>"000000001",
  40133=>"000000000",
  40134=>"000000010",
  40135=>"111111000",
  40136=>"110000011",
  40137=>"001111111",
  40138=>"000001101",
  40139=>"001111000",
  40140=>"110111111",
  40141=>"000000000",
  40142=>"100000110",
  40143=>"110110000",
  40144=>"000111111",
  40145=>"100000001",
  40146=>"111111111",
  40147=>"000000111",
  40148=>"111001000",
  40149=>"011111111",
  40150=>"110110000",
  40151=>"111110000",
  40152=>"100000000",
  40153=>"111001101",
  40154=>"000000111",
  40155=>"111110100",
  40156=>"000000001",
  40157=>"001101101",
  40158=>"111111111",
  40159=>"000000000",
  40160=>"001000000",
  40161=>"111110110",
  40162=>"110111011",
  40163=>"000001000",
  40164=>"000000001",
  40165=>"100100101",
  40166=>"000000001",
  40167=>"011000001",
  40168=>"011111111",
  40169=>"111101011",
  40170=>"110111111",
  40171=>"110000111",
  40172=>"111111000",
  40173=>"111000101",
  40174=>"111111101",
  40175=>"111001000",
  40176=>"000000001",
  40177=>"001101111",
  40178=>"111111111",
  40179=>"001000111",
  40180=>"111111000",
  40181=>"000001000",
  40182=>"111111001",
  40183=>"111011000",
  40184=>"000111110",
  40185=>"111110110",
  40186=>"000000000",
  40187=>"000000000",
  40188=>"001000000",
  40189=>"110010010",
  40190=>"000000111",
  40191=>"101000000",
  40192=>"000000001",
  40193=>"011001001",
  40194=>"010000000",
  40195=>"111111000",
  40196=>"100000000",
  40197=>"111110111",
  40198=>"111111000",
  40199=>"001101110",
  40200=>"110100111",
  40201=>"111100000",
  40202=>"001001001",
  40203=>"110111001",
  40204=>"000100100",
  40205=>"000111111",
  40206=>"000000110",
  40207=>"110111110",
  40208=>"110111000",
  40209=>"000000000",
  40210=>"000000000",
  40211=>"000111111",
  40212=>"111111000",
  40213=>"111011100",
  40214=>"000111001",
  40215=>"000000110",
  40216=>"000000111",
  40217=>"110111111",
  40218=>"000000111",
  40219=>"000000000",
  40220=>"011011111",
  40221=>"101000100",
  40222=>"111111011",
  40223=>"111111101",
  40224=>"100011000",
  40225=>"111111001",
  40226=>"101111000",
  40227=>"000000000",
  40228=>"111001001",
  40229=>"001000000",
  40230=>"000000000",
  40231=>"101000100",
  40232=>"000000000",
  40233=>"100000101",
  40234=>"111100101",
  40235=>"100100000",
  40236=>"101111111",
  40237=>"011111110",
  40238=>"000111101",
  40239=>"000000000",
  40240=>"011011000",
  40241=>"111110111",
  40242=>"111111111",
  40243=>"111111111",
  40244=>"111100110",
  40245=>"001111111",
  40246=>"110000000",
  40247=>"100000001",
  40248=>"111111000",
  40249=>"101001000",
  40250=>"111000100",
  40251=>"000000000",
  40252=>"111111111",
  40253=>"000000110",
  40254=>"000001111",
  40255=>"111111111",
  40256=>"111111011",
  40257=>"111110110",
  40258=>"000100000",
  40259=>"000000111",
  40260=>"000000000",
  40261=>"111000000",
  40262=>"111001001",
  40263=>"000000111",
  40264=>"111111111",
  40265=>"111000000",
  40266=>"110010000",
  40267=>"011111011",
  40268=>"000000001",
  40269=>"000000000",
  40270=>"110111111",
  40271=>"000111111",
  40272=>"001011011",
  40273=>"000000000",
  40274=>"111111111",
  40275=>"110100000",
  40276=>"000000111",
  40277=>"001101111",
  40278=>"011111111",
  40279=>"100100111",
  40280=>"111111111",
  40281=>"100111111",
  40282=>"110110111",
  40283=>"000000000",
  40284=>"111111001",
  40285=>"000000000",
  40286=>"001000000",
  40287=>"000000000",
  40288=>"101100000",
  40289=>"110111110",
  40290=>"111111111",
  40291=>"001000000",
  40292=>"000000000",
  40293=>"011011000",
  40294=>"000101101",
  40295=>"010111111",
  40296=>"000010001",
  40297=>"011100101",
  40298=>"000000000",
  40299=>"000000100",
  40300=>"111101111",
  40301=>"011001000",
  40302=>"001111111",
  40303=>"011011010",
  40304=>"000000000",
  40305=>"000011000",
  40306=>"001110111",
  40307=>"000000000",
  40308=>"001001000",
  40309=>"111111000",
  40310=>"111011001",
  40311=>"111111111",
  40312=>"000000111",
  40313=>"111000000",
  40314=>"000101111",
  40315=>"010000001",
  40316=>"001001001",
  40317=>"001111111",
  40318=>"000000000",
  40319=>"000000000",
  40320=>"110111111",
  40321=>"100101101",
  40322=>"111111111",
  40323=>"111111111",
  40324=>"111111111",
  40325=>"110100110",
  40326=>"000000000",
  40327=>"001000111",
  40328=>"100000000",
  40329=>"111111101",
  40330=>"001011001",
  40331=>"000101111",
  40332=>"000111111",
  40333=>"111011011",
  40334=>"000001000",
  40335=>"000000000",
  40336=>"110111111",
  40337=>"000000000",
  40338=>"000000001",
  40339=>"110110110",
  40340=>"111000110",
  40341=>"000011000",
  40342=>"011111000",
  40343=>"111111101",
  40344=>"011011000",
  40345=>"000110000",
  40346=>"001000111",
  40347=>"111111111",
  40348=>"000000000",
  40349=>"000000111",
  40350=>"000000111",
  40351=>"000001000",
  40352=>"000000000",
  40353=>"111111011",
  40354=>"010000101",
  40355=>"000000000",
  40356=>"111111111",
  40357=>"000000000",
  40358=>"000000000",
  40359=>"011111111",
  40360=>"111000111",
  40361=>"111111110",
  40362=>"110100100",
  40363=>"000000000",
  40364=>"000000000",
  40365=>"011000000",
  40366=>"100111111",
  40367=>"011111111",
  40368=>"111111000",
  40369=>"000100000",
  40370=>"111111011",
  40371=>"110000000",
  40372=>"001101111",
  40373=>"111111111",
  40374=>"111101000",
  40375=>"010111111",
  40376=>"111001000",
  40377=>"000001111",
  40378=>"100000000",
  40379=>"111000111",
  40380=>"111110000",
  40381=>"111000111",
  40382=>"000000000",
  40383=>"011011011",
  40384=>"011100100",
  40385=>"111001001",
  40386=>"111111000",
  40387=>"000101011",
  40388=>"011001111",
  40389=>"000000100",
  40390=>"000010010",
  40391=>"000010110",
  40392=>"111111111",
  40393=>"000110111",
  40394=>"000000000",
  40395=>"110111000",
  40396=>"111000000",
  40397=>"111110000",
  40398=>"111000000",
  40399=>"111111010",
  40400=>"000000011",
  40401=>"110100100",
  40402=>"111011111",
  40403=>"111111000",
  40404=>"110110011",
  40405=>"000000000",
  40406=>"100111111",
  40407=>"011000111",
  40408=>"000001111",
  40409=>"000000000",
  40410=>"111111111",
  40411=>"001000101",
  40412=>"000001001",
  40413=>"000000111",
  40414=>"111101000",
  40415=>"010011001",
  40416=>"111111100",
  40417=>"111000000",
  40418=>"000100111",
  40419=>"000000111",
  40420=>"011000001",
  40421=>"100100111",
  40422=>"111000000",
  40423=>"000101111",
  40424=>"110100001",
  40425=>"100000000",
  40426=>"001001011",
  40427=>"000111011",
  40428=>"111101111",
  40429=>"111111001",
  40430=>"111000000",
  40431=>"001000000",
  40432=>"000000100",
  40433=>"111111111",
  40434=>"000000000",
  40435=>"000000000",
  40436=>"000000111",
  40437=>"111000000",
  40438=>"111111111",
  40439=>"011111111",
  40440=>"111111000",
  40441=>"100100100",
  40442=>"001001000",
  40443=>"110110000",
  40444=>"111111000",
  40445=>"111000111",
  40446=>"111011000",
  40447=>"111000000",
  40448=>"110110110",
  40449=>"000000100",
  40450=>"011111111",
  40451=>"000000111",
  40452=>"100000000",
  40453=>"111111111",
  40454=>"101100111",
  40455=>"111111111",
  40456=>"111000000",
  40457=>"110111000",
  40458=>"000000111",
  40459=>"000000011",
  40460=>"100100000",
  40461=>"111001000",
  40462=>"011111111",
  40463=>"000000011",
  40464=>"111000111",
  40465=>"010000000",
  40466=>"011011000",
  40467=>"111111111",
  40468=>"100100111",
  40469=>"111111100",
  40470=>"000000000",
  40471=>"001111001",
  40472=>"010000111",
  40473=>"011000100",
  40474=>"000000000",
  40475=>"001110100",
  40476=>"111100000",
  40477=>"111111000",
  40478=>"001100110",
  40479=>"001101101",
  40480=>"000000000",
  40481=>"111000000",
  40482=>"000000000",
  40483=>"111111111",
  40484=>"111110000",
  40485=>"111111111",
  40486=>"111111111",
  40487=>"111011111",
  40488=>"010100100",
  40489=>"000000000",
  40490=>"000110111",
  40491=>"000001001",
  40492=>"111111000",
  40493=>"111111111",
  40494=>"000011001",
  40495=>"111111111",
  40496=>"000100111",
  40497=>"001111111",
  40498=>"110000100",
  40499=>"011111111",
  40500=>"000011000",
  40501=>"010011000",
  40502=>"000000011",
  40503=>"000000001",
  40504=>"111111000",
  40505=>"000000000",
  40506=>"000000000",
  40507=>"000000000",
  40508=>"111111111",
  40509=>"000110110",
  40510=>"101000001",
  40511=>"100110111",
  40512=>"010111000",
  40513=>"100110110",
  40514=>"000000000",
  40515=>"011111100",
  40516=>"000000000",
  40517=>"000001111",
  40518=>"110111000",
  40519=>"000100100",
  40520=>"010011010",
  40521=>"000000111",
  40522=>"111111111",
  40523=>"110111111",
  40524=>"011110110",
  40525=>"000000000",
  40526=>"000000110",
  40527=>"011111000",
  40528=>"000000000",
  40529=>"111100110",
  40530=>"110110000",
  40531=>"000011111",
  40532=>"000000000",
  40533=>"000000000",
  40534=>"010000000",
  40535=>"111111111",
  40536=>"000000000",
  40537=>"000000000",
  40538=>"111100000",
  40539=>"001001001",
  40540=>"000001111",
  40541=>"111010000",
  40542=>"111010010",
  40543=>"110000000",
  40544=>"000000100",
  40545=>"000010011",
  40546=>"000000000",
  40547=>"000000000",
  40548=>"000010011",
  40549=>"111000000",
  40550=>"000100111",
  40551=>"010111011",
  40552=>"000111111",
  40553=>"011000101",
  40554=>"000011111",
  40555=>"111111110",
  40556=>"000000000",
  40557=>"000000100",
  40558=>"000000000",
  40559=>"000011111",
  40560=>"111100000",
  40561=>"000111111",
  40562=>"000000111",
  40563=>"000110100",
  40564=>"100000110",
  40565=>"010001000",
  40566=>"111111000",
  40567=>"010011011",
  40568=>"110111000",
  40569=>"111011011",
  40570=>"111001000",
  40571=>"000000011",
  40572=>"110110101",
  40573=>"000110110",
  40574=>"111110000",
  40575=>"000011111",
  40576=>"000000000",
  40577=>"111011100",
  40578=>"111111001",
  40579=>"000111011",
  40580=>"000000111",
  40581=>"100000000",
  40582=>"100110110",
  40583=>"011000000",
  40584=>"111000000",
  40585=>"000000101",
  40586=>"000000000",
  40587=>"111111111",
  40588=>"000101111",
  40589=>"000011111",
  40590=>"111010111",
  40591=>"111110111",
  40592=>"111111000",
  40593=>"011111001",
  40594=>"111000000",
  40595=>"111111000",
  40596=>"111110000",
  40597=>"000000000",
  40598=>"000000000",
  40599=>"000000111",
  40600=>"101101101",
  40601=>"111000000",
  40602=>"111111000",
  40603=>"111111011",
  40604=>"000000111",
  40605=>"110011010",
  40606=>"111111101",
  40607=>"101111111",
  40608=>"000000000",
  40609=>"110101000",
  40610=>"001001011",
  40611=>"111111111",
  40612=>"111000000",
  40613=>"111110000",
  40614=>"111111110",
  40615=>"011000000",
  40616=>"000100111",
  40617=>"011001011",
  40618=>"111111100",
  40619=>"110111111",
  40620=>"111111100",
  40621=>"011000000",
  40622=>"000000000",
  40623=>"111011110",
  40624=>"110000011",
  40625=>"001010011",
  40626=>"111111111",
  40627=>"000000010",
  40628=>"111000000",
  40629=>"000000000",
  40630=>"111000010",
  40631=>"101111111",
  40632=>"111001000",
  40633=>"111111000",
  40634=>"111001111",
  40635=>"111111100",
  40636=>"111010110",
  40637=>"100100101",
  40638=>"111110111",
  40639=>"110010000",
  40640=>"111111000",
  40641=>"100000000",
  40642=>"111000000",
  40643=>"010010010",
  40644=>"000000000",
  40645=>"001000001",
  40646=>"000000000",
  40647=>"000000000",
  40648=>"000100100",
  40649=>"000110111",
  40650=>"100000000",
  40651=>"100110111",
  40652=>"000001001",
  40653=>"000111111",
  40654=>"000100111",
  40655=>"001111111",
  40656=>"001000111",
  40657=>"000111111",
  40658=>"000011111",
  40659=>"111100100",
  40660=>"000000000",
  40661=>"111000100",
  40662=>"100111111",
  40663=>"000000100",
  40664=>"111110000",
  40665=>"000000100",
  40666=>"000000000",
  40667=>"111111010",
  40668=>"111011101",
  40669=>"000000000",
  40670=>"000111111",
  40671=>"000000000",
  40672=>"101000000",
  40673=>"001111011",
  40674=>"111110000",
  40675=>"000111111",
  40676=>"111111001",
  40677=>"100000110",
  40678=>"000111111",
  40679=>"111111110",
  40680=>"111111111",
  40681=>"110111111",
  40682=>"011000000",
  40683=>"111000110",
  40684=>"011000100",
  40685=>"111111111",
  40686=>"101100111",
  40687=>"000000000",
  40688=>"000000011",
  40689=>"111110111",
  40690=>"111111000",
  40691=>"000000000",
  40692=>"000000110",
  40693=>"001001000",
  40694=>"010011110",
  40695=>"111111110",
  40696=>"101001011",
  40697=>"011111111",
  40698=>"001000000",
  40699=>"001101111",
  40700=>"000000000",
  40701=>"000000000",
  40702=>"011110111",
  40703=>"100110100",
  40704=>"111111110",
  40705=>"001000001",
  40706=>"111011011",
  40707=>"011010000",
  40708=>"111111000",
  40709=>"101101111",
  40710=>"000000000",
  40711=>"000110111",
  40712=>"001000000",
  40713=>"000000000",
  40714=>"001000000",
  40715=>"000000000",
  40716=>"101111111",
  40717=>"000000000",
  40718=>"111000000",
  40719=>"111111000",
  40720=>"000000011",
  40721=>"000000000",
  40722=>"000000000",
  40723=>"000110111",
  40724=>"110111111",
  40725=>"010110000",
  40726=>"000000000",
  40727=>"111111111",
  40728=>"000011110",
  40729=>"000000011",
  40730=>"011011011",
  40731=>"001111111",
  40732=>"000000000",
  40733=>"000000111",
  40734=>"111111101",
  40735=>"000000000",
  40736=>"001011001",
  40737=>"100111111",
  40738=>"011111111",
  40739=>"111011111",
  40740=>"111111011",
  40741=>"111101111",
  40742=>"100100000",
  40743=>"000000011",
  40744=>"101100000",
  40745=>"111111111",
  40746=>"111000000",
  40747=>"110100101",
  40748=>"000001001",
  40749=>"110110010",
  40750=>"000000111",
  40751=>"000000001",
  40752=>"011010000",
  40753=>"000000000",
  40754=>"000111111",
  40755=>"000000111",
  40756=>"000000000",
  40757=>"001000001",
  40758=>"111000000",
  40759=>"111111101",
  40760=>"111100000",
  40761=>"111000000",
  40762=>"000000111",
  40763=>"010000000",
  40764=>"100000000",
  40765=>"111111111",
  40766=>"111011000",
  40767=>"011000111",
  40768=>"111000000",
  40769=>"111110000",
  40770=>"000000000",
  40771=>"110111111",
  40772=>"000001001",
  40773=>"000000000",
  40774=>"001000001",
  40775=>"000001111",
  40776=>"001000000",
  40777=>"000111111",
  40778=>"100100011",
  40779=>"001111111",
  40780=>"000000000",
  40781=>"111111111",
  40782=>"000000000",
  40783=>"000111111",
  40784=>"111000100",
  40785=>"111111100",
  40786=>"100000010",
  40787=>"110111111",
  40788=>"000010000",
  40789=>"001011011",
  40790=>"000000000",
  40791=>"011111111",
  40792=>"111111111",
  40793=>"111000000",
  40794=>"000001000",
  40795=>"111000100",
  40796=>"110111110",
  40797=>"001000000",
  40798=>"110011111",
  40799=>"101101111",
  40800=>"000000111",
  40801=>"011111010",
  40802=>"000000001",
  40803=>"111111111",
  40804=>"000110100",
  40805=>"000000000",
  40806=>"111000011",
  40807=>"111111110",
  40808=>"110110111",
  40809=>"100000000",
  40810=>"000110010",
  40811=>"110010110",
  40812=>"001111011",
  40813=>"100110111",
  40814=>"111000000",
  40815=>"000110000",
  40816=>"101111110",
  40817=>"111101100",
  40818=>"000000000",
  40819=>"000110010",
  40820=>"111100000",
  40821=>"000000000",
  40822=>"111000000",
  40823=>"000000000",
  40824=>"111000000",
  40825=>"111111111",
  40826=>"010111111",
  40827=>"000010000",
  40828=>"111001000",
  40829=>"111111111",
  40830=>"001000000",
  40831=>"100100000",
  40832=>"000000000",
  40833=>"110111111",
  40834=>"001001111",
  40835=>"000010011",
  40836=>"000000111",
  40837=>"000000000",
  40838=>"110000000",
  40839=>"000100101",
  40840=>"000000010",
  40841=>"111011000",
  40842=>"111111111",
  40843=>"111100111",
  40844=>"111001111",
  40845=>"011011011",
  40846=>"000111110",
  40847=>"111111111",
  40848=>"111111111",
  40849=>"111111111",
  40850=>"011111111",
  40851=>"001000000",
  40852=>"001100111",
  40853=>"000000000",
  40854=>"111000100",
  40855=>"010010010",
  40856=>"000000000",
  40857=>"000111000",
  40858=>"000000100",
  40859=>"111011010",
  40860=>"000011111",
  40861=>"000000000",
  40862=>"000000000",
  40863=>"000000010",
  40864=>"000000100",
  40865=>"110110101",
  40866=>"011111111",
  40867=>"000000000",
  40868=>"001000101",
  40869=>"000100111",
  40870=>"100101111",
  40871=>"010110111",
  40872=>"111111111",
  40873=>"111011011",
  40874=>"000000101",
  40875=>"011000000",
  40876=>"000000000",
  40877=>"001000000",
  40878=>"111111000",
  40879=>"110110000",
  40880=>"111111110",
  40881=>"000000000",
  40882=>"111000001",
  40883=>"000111111",
  40884=>"000110111",
  40885=>"101101111",
  40886=>"111111111",
  40887=>"000000011",
  40888=>"010011001",
  40889=>"111111110",
  40890=>"001011011",
  40891=>"111111011",
  40892=>"000000111",
  40893=>"000000101",
  40894=>"100100000",
  40895=>"011001001",
  40896=>"001100000",
  40897=>"111111000",
  40898=>"000000111",
  40899=>"000000111",
  40900=>"111110111",
  40901=>"011000100",
  40902=>"111111110",
  40903=>"100000100",
  40904=>"111100100",
  40905=>"001011111",
  40906=>"000001000",
  40907=>"000110000",
  40908=>"111100000",
  40909=>"000110000",
  40910=>"001000111",
  40911=>"010001000",
  40912=>"000111111",
  40913=>"001101000",
  40914=>"111111110",
  40915=>"000000011",
  40916=>"000000011",
  40917=>"001000100",
  40918=>"011111100",
  40919=>"000001011",
  40920=>"000111011",
  40921=>"011000000",
  40922=>"000111111",
  40923=>"101000000",
  40924=>"000111011",
  40925=>"011000110",
  40926=>"000000000",
  40927=>"001001011",
  40928=>"110000000",
  40929=>"000000000",
  40930=>"000000011",
  40931=>"000000001",
  40932=>"100000000",
  40933=>"101000000",
  40934=>"011000111",
  40935=>"000000001",
  40936=>"001011011",
  40937=>"000000001",
  40938=>"000000000",
  40939=>"000000000",
  40940=>"000000001",
  40941=>"010000001",
  40942=>"100100111",
  40943=>"001001111",
  40944=>"100000000",
  40945=>"111111111",
  40946=>"001000000",
  40947=>"000111011",
  40948=>"010010000",
  40949=>"011011111",
  40950=>"000111011",
  40951=>"111111011",
  40952=>"111111000",
  40953=>"110111000",
  40954=>"100000000",
  40955=>"010111110",
  40956=>"111001000",
  40957=>"101101000",
  40958=>"111111010",
  40959=>"111000111",
  40960=>"000000001",
  40961=>"001000000",
  40962=>"111111001",
  40963=>"000100111",
  40964=>"001111011",
  40965=>"000001111",
  40966=>"111000000",
  40967=>"011011011",
  40968=>"111011000",
  40969=>"111100100",
  40970=>"000111111",
  40971=>"000000000",
  40972=>"000111001",
  40973=>"111011010",
  40974=>"000110110",
  40975=>"111000000",
  40976=>"111111111",
  40977=>"000011111",
  40978=>"001111111",
  40979=>"111010111",
  40980=>"000000000",
  40981=>"111011011",
  40982=>"000000000",
  40983=>"111110011",
  40984=>"110000000",
  40985=>"100000000",
  40986=>"111000000",
  40987=>"111110110",
  40988=>"000000000",
  40989=>"111111111",
  40990=>"000001000",
  40991=>"000000000",
  40992=>"111111101",
  40993=>"000111111",
  40994=>"000111111",
  40995=>"000010010",
  40996=>"000100100",
  40997=>"000000010",
  40998=>"101101100",
  40999=>"000100111",
  41000=>"100100100",
  41001=>"000000000",
  41002=>"111111000",
  41003=>"000001110",
  41004=>"101111111",
  41005=>"111111111",
  41006=>"111111111",
  41007=>"000000000",
  41008=>"111111111",
  41009=>"000000000",
  41010=>"100110100",
  41011=>"111111111",
  41012=>"000000000",
  41013=>"111001000",
  41014=>"001100100",
  41015=>"101100001",
  41016=>"000000000",
  41017=>"010111111",
  41018=>"110001111",
  41019=>"011011111",
  41020=>"111111111",
  41021=>"001011100",
  41022=>"111011011",
  41023=>"100000101",
  41024=>"111111001",
  41025=>"111111000",
  41026=>"000111111",
  41027=>"111111111",
  41028=>"111111000",
  41029=>"001000000",
  41030=>"111000111",
  41031=>"111111111",
  41032=>"111111010",
  41033=>"000000100",
  41034=>"111111110",
  41035=>"100101001",
  41036=>"001010000",
  41037=>"111111000",
  41038=>"001101100",
  41039=>"111111111",
  41040=>"000010111",
  41041=>"010011111",
  41042=>"001000101",
  41043=>"000000100",
  41044=>"000000000",
  41045=>"000110111",
  41046=>"001000000",
  41047=>"111111011",
  41048=>"110110000",
  41049=>"111000000",
  41050=>"011010111",
  41051=>"111011001",
  41052=>"000000000",
  41053=>"111111000",
  41054=>"111101001",
  41055=>"111111000",
  41056=>"000000000",
  41057=>"001011111",
  41058=>"001101001",
  41059=>"010010111",
  41060=>"000000011",
  41061=>"010010001",
  41062=>"011000000",
  41063=>"000000001",
  41064=>"011011000",
  41065=>"111111010",
  41066=>"000000111",
  41067=>"000000000",
  41068=>"001000000",
  41069=>"100000000",
  41070=>"001000000",
  41071=>"000101000",
  41072=>"110110110",
  41073=>"111000000",
  41074=>"110110110",
  41075=>"111111000",
  41076=>"000000000",
  41077=>"101011111",
  41078=>"000111111",
  41079=>"000000000",
  41080=>"111001000",
  41081=>"000000000",
  41082=>"001011010",
  41083=>"111000000",
  41084=>"111011011",
  41085=>"111100001",
  41086=>"100000000",
  41087=>"000000000",
  41088=>"000100101",
  41089=>"110010111",
  41090=>"110000010",
  41091=>"001001000",
  41092=>"110011000",
  41093=>"101011011",
  41094=>"000000110",
  41095=>"100110111",
  41096=>"111111111",
  41097=>"001000000",
  41098=>"110111111",
  41099=>"000000000",
  41100=>"101111111",
  41101=>"001001000",
  41102=>"111111111",
  41103=>"110111111",
  41104=>"000000000",
  41105=>"000011010",
  41106=>"000000000",
  41107=>"010111110",
  41108=>"001001001",
  41109=>"000111111",
  41110=>"010101111",
  41111=>"111000000",
  41112=>"101000001",
  41113=>"111111111",
  41114=>"111001111",
  41115=>"111101001",
  41116=>"111100000",
  41117=>"110100000",
  41118=>"111110000",
  41119=>"110000111",
  41120=>"111000000",
  41121=>"001011000",
  41122=>"000111111",
  41123=>"000000100",
  41124=>"011001001",
  41125=>"000000110",
  41126=>"000010111",
  41127=>"111110010",
  41128=>"000000111",
  41129=>"000000000",
  41130=>"111111100",
  41131=>"000100110",
  41132=>"011000011",
  41133=>"100110010",
  41134=>"000000000",
  41135=>"000000000",
  41136=>"010000000",
  41137=>"100011000",
  41138=>"010111111",
  41139=>"010000000",
  41140=>"111100100",
  41141=>"000000000",
  41142=>"000000001",
  41143=>"111000000",
  41144=>"000100100",
  41145=>"111111111",
  41146=>"001001001",
  41147=>"111111111",
  41148=>"000000000",
  41149=>"101111111",
  41150=>"111000000",
  41151=>"000100111",
  41152=>"111111111",
  41153=>"001011001",
  41154=>"111111111",
  41155=>"111011000",
  41156=>"001100110",
  41157=>"000001111",
  41158=>"111000000",
  41159=>"000111000",
  41160=>"000000011",
  41161=>"000001000",
  41162=>"111111111",
  41163=>"000100111",
  41164=>"111111001",
  41165=>"110101111",
  41166=>"000000100",
  41167=>"111111000",
  41168=>"000000001",
  41169=>"001000000",
  41170=>"000001000",
  41171=>"001000001",
  41172=>"111111111",
  41173=>"100111111",
  41174=>"001111011",
  41175=>"111110010",
  41176=>"000110111",
  41177=>"111111111",
  41178=>"111111000",
  41179=>"000001101",
  41180=>"001000000",
  41181=>"000111100",
  41182=>"111111111",
  41183=>"000000000",
  41184=>"010000000",
  41185=>"000000011",
  41186=>"011011000",
  41187=>"101000101",
  41188=>"101011111",
  41189=>"110100100",
  41190=>"011111111",
  41191=>"000000000",
  41192=>"000000001",
  41193=>"111000000",
  41194=>"111011000",
  41195=>"100001000",
  41196=>"111100111",
  41197=>"000011111",
  41198=>"111000000",
  41199=>"000111111",
  41200=>"110110110",
  41201=>"111110000",
  41202=>"111110000",
  41203=>"001001011",
  41204=>"111111011",
  41205=>"111110111",
  41206=>"110110110",
  41207=>"111000110",
  41208=>"001111111",
  41209=>"011111010",
  41210=>"000000000",
  41211=>"111111011",
  41212=>"111111110",
  41213=>"111011001",
  41214=>"001001001",
  41215=>"111111110",
  41216=>"111001111",
  41217=>"011000000",
  41218=>"000010101",
  41219=>"000000001",
  41220=>"011011000",
  41221=>"001001001",
  41222=>"111111110",
  41223=>"111111100",
  41224=>"111110000",
  41225=>"000000111",
  41226=>"101100111",
  41227=>"000000110",
  41228=>"000000000",
  41229=>"000000100",
  41230=>"111111110",
  41231=>"000000000",
  41232=>"111000000",
  41233=>"101101001",
  41234=>"000000101",
  41235=>"001001111",
  41236=>"101001011",
  41237=>"111111000",
  41238=>"110000000",
  41239=>"000000000",
  41240=>"100111111",
  41241=>"101111111",
  41242=>"100000000",
  41243=>"000000000",
  41244=>"001000001",
  41245=>"111111111",
  41246=>"000000000",
  41247=>"101111000",
  41248=>"110100110",
  41249=>"000001111",
  41250=>"000000000",
  41251=>"111111111",
  41252=>"011111111",
  41253=>"111111111",
  41254=>"000000010",
  41255=>"000000101",
  41256=>"000111111",
  41257=>"000000111",
  41258=>"001111111",
  41259=>"111011000",
  41260=>"000000111",
  41261=>"111111111",
  41262=>"000111000",
  41263=>"111000000",
  41264=>"111111111",
  41265=>"001111111",
  41266=>"111111111",
  41267=>"100100111",
  41268=>"111010000",
  41269=>"010011000",
  41270=>"111011111",
  41271=>"111001000",
  41272=>"110000000",
  41273=>"111000000",
  41274=>"000000000",
  41275=>"000100111",
  41276=>"111111110",
  41277=>"111000110",
  41278=>"000000000",
  41279=>"111111000",
  41280=>"000000000",
  41281=>"100111110",
  41282=>"000000111",
  41283=>"111111111",
  41284=>"111111010",
  41285=>"100000111",
  41286=>"001111111",
  41287=>"000111010",
  41288=>"000000000",
  41289=>"111000000",
  41290=>"000100111",
  41291=>"110110110",
  41292=>"000100111",
  41293=>"111111111",
  41294=>"111100111",
  41295=>"000000110",
  41296=>"001001000",
  41297=>"100100000",
  41298=>"111111011",
  41299=>"000001000",
  41300=>"000111111",
  41301=>"001111111",
  41302=>"111111000",
  41303=>"111100000",
  41304=>"000000000",
  41305=>"000000000",
  41306=>"111010000",
  41307=>"001000011",
  41308=>"000000111",
  41309=>"000000000",
  41310=>"101101100",
  41311=>"001011111",
  41312=>"000000110",
  41313=>"000111111",
  41314=>"111110100",
  41315=>"001001000",
  41316=>"100100111",
  41317=>"000000101",
  41318=>"000000000",
  41319=>"011111111",
  41320=>"111111011",
  41321=>"111110000",
  41322=>"000011111",
  41323=>"110111011",
  41324=>"110111111",
  41325=>"011001111",
  41326=>"111001000",
  41327=>"011111010",
  41328=>"010000000",
  41329=>"111100110",
  41330=>"000100100",
  41331=>"111111111",
  41332=>"111111100",
  41333=>"000000001",
  41334=>"000000000",
  41335=>"010000000",
  41336=>"111111111",
  41337=>"001000000",
  41338=>"100111111",
  41339=>"000000000",
  41340=>"101000110",
  41341=>"001111110",
  41342=>"111111000",
  41343=>"111000000",
  41344=>"111001111",
  41345=>"100101111",
  41346=>"111100000",
  41347=>"000000000",
  41348=>"000000000",
  41349=>"111001111",
  41350=>"000000110",
  41351=>"000000111",
  41352=>"000000000",
  41353=>"000010111",
  41354=>"111100000",
  41355=>"111000000",
  41356=>"000011001",
  41357=>"000000100",
  41358=>"011111111",
  41359=>"010110111",
  41360=>"001000000",
  41361=>"000000001",
  41362=>"101000101",
  41363=>"111101111",
  41364=>"011000111",
  41365=>"000000000",
  41366=>"100101111",
  41367=>"100111111",
  41368=>"000000000",
  41369=>"001000110",
  41370=>"111111010",
  41371=>"110110110",
  41372=>"001001001",
  41373=>"000100111",
  41374=>"011000000",
  41375=>"111000000",
  41376=>"111111111",
  41377=>"000000110",
  41378=>"100111000",
  41379=>"111011001",
  41380=>"000000011",
  41381=>"000111100",
  41382=>"000000000",
  41383=>"000110111",
  41384=>"110000000",
  41385=>"000000000",
  41386=>"111111111",
  41387=>"100001000",
  41388=>"000000000",
  41389=>"000000000",
  41390=>"010000111",
  41391=>"111111100",
  41392=>"000000111",
  41393=>"000000000",
  41394=>"111111111",
  41395=>"111111101",
  41396=>"000000000",
  41397=>"000100111",
  41398=>"001000000",
  41399=>"000000111",
  41400=>"000000000",
  41401=>"000110111",
  41402=>"111101011",
  41403=>"000000110",
  41404=>"111011001",
  41405=>"111110111",
  41406=>"000000011",
  41407=>"010000000",
  41408=>"111111011",
  41409=>"000000010",
  41410=>"001000000",
  41411=>"000000000",
  41412=>"000001011",
  41413=>"100000000",
  41414=>"111001000",
  41415=>"011001111",
  41416=>"011000000",
  41417=>"010110000",
  41418=>"111101000",
  41419=>"100000111",
  41420=>"111001000",
  41421=>"101100011",
  41422=>"001011000",
  41423=>"000000010",
  41424=>"011011001",
  41425=>"110110111",
  41426=>"111111111",
  41427=>"000010100",
  41428=>"111111000",
  41429=>"111111111",
  41430=>"110111000",
  41431=>"000011110",
  41432=>"110000000",
  41433=>"001000000",
  41434=>"011011000",
  41435=>"001101101",
  41436=>"000000000",
  41437=>"100101111",
  41438=>"111111101",
  41439=>"001011000",
  41440=>"111011111",
  41441=>"111111000",
  41442=>"110100000",
  41443=>"000000010",
  41444=>"111001011",
  41445=>"100000111",
  41446=>"111000000",
  41447=>"111101101",
  41448=>"000110111",
  41449=>"000100111",
  41450=>"000000000",
  41451=>"000000000",
  41452=>"000000000",
  41453=>"001111111",
  41454=>"111011111",
  41455=>"111000111",
  41456=>"001000000",
  41457=>"101000110",
  41458=>"111011110",
  41459=>"000000000",
  41460=>"101000000",
  41461=>"101111111",
  41462=>"000000001",
  41463=>"100000000",
  41464=>"001111111",
  41465=>"100000000",
  41466=>"001001000",
  41467=>"111001001",
  41468=>"001100101",
  41469=>"111111011",
  41470=>"111000000",
  41471=>"100000110",
  41472=>"110111001",
  41473=>"110110110",
  41474=>"111100000",
  41475=>"000000000",
  41476=>"000000000",
  41477=>"100000000",
  41478=>"000000000",
  41479=>"111111111",
  41480=>"000010111",
  41481=>"111001001",
  41482=>"001001111",
  41483=>"000000001",
  41484=>"111000000",
  41485=>"000000000",
  41486=>"111111111",
  41487=>"111111111",
  41488=>"000000000",
  41489=>"000000000",
  41490=>"011011011",
  41491=>"000000000",
  41492=>"111111111",
  41493=>"111111000",
  41494=>"111000110",
  41495=>"011011011",
  41496=>"111111111",
  41497=>"100010111",
  41498=>"000000000",
  41499=>"110110110",
  41500=>"111001111",
  41501=>"111111111",
  41502=>"011010000",
  41503=>"000010010",
  41504=>"010000000",
  41505=>"011000000",
  41506=>"011011000",
  41507=>"000000000",
  41508=>"000000011",
  41509=>"000001011",
  41510=>"010011111",
  41511=>"101111111",
  41512=>"110011011",
  41513=>"000000000",
  41514=>"000000110",
  41515=>"000000000",
  41516=>"101111111",
  41517=>"000000000",
  41518=>"100111111",
  41519=>"111111111",
  41520=>"111110000",
  41521=>"000100111",
  41522=>"100100100",
  41523=>"000000000",
  41524=>"000111111",
  41525=>"111011011",
  41526=>"000000000",
  41527=>"000000100",
  41528=>"001000000",
  41529=>"000000000",
  41530=>"000000110",
  41531=>"111110101",
  41532=>"111111111",
  41533=>"111011011",
  41534=>"000000000",
  41535=>"111111111",
  41536=>"111000000",
  41537=>"111111111",
  41538=>"000000111",
  41539=>"100110000",
  41540=>"111111011",
  41541=>"000000000",
  41542=>"011001001",
  41543=>"000000000",
  41544=>"000000110",
  41545=>"111111111",
  41546=>"000000000",
  41547=>"000000000",
  41548=>"111111111",
  41549=>"111010010",
  41550=>"000000000",
  41551=>"000000000",
  41552=>"100000000",
  41553=>"110110000",
  41554=>"111101111",
  41555=>"111111011",
  41556=>"000000001",
  41557=>"100110110",
  41558=>"000000000",
  41559=>"000000000",
  41560=>"111111111",
  41561=>"000000101",
  41562=>"111111111",
  41563=>"011000011",
  41564=>"111011001",
  41565=>"111011000",
  41566=>"000101001",
  41567=>"000001011",
  41568=>"000000111",
  41569=>"111110111",
  41570=>"000000000",
  41571=>"000000000",
  41572=>"111111100",
  41573=>"111111111",
  41574=>"111111111",
  41575=>"111111111",
  41576=>"111111111",
  41577=>"111111111",
  41578=>"000000100",
  41579=>"111110000",
  41580=>"000000000",
  41581=>"111111000",
  41582=>"000000000",
  41583=>"111111010",
  41584=>"111111111",
  41585=>"111111111",
  41586=>"100100100",
  41587=>"111110000",
  41588=>"000000000",
  41589=>"000111100",
  41590=>"111111000",
  41591=>"001111111",
  41592=>"101111001",
  41593=>"110100000",
  41594=>"000000000",
  41595=>"000000000",
  41596=>"110110110",
  41597=>"011111111",
  41598=>"000000001",
  41599=>"000100110",
  41600=>"111111111",
  41601=>"111111111",
  41602=>"000000000",
  41603=>"001001000",
  41604=>"000000000",
  41605=>"111100111",
  41606=>"000000000",
  41607=>"000000000",
  41608=>"110000111",
  41609=>"111111111",
  41610=>"111111111",
  41611=>"111111111",
  41612=>"111111010",
  41613=>"111111100",
  41614=>"000000011",
  41615=>"000000000",
  41616=>"000010111",
  41617=>"010000000",
  41618=>"101000100",
  41619=>"100011011",
  41620=>"000000000",
  41621=>"000000000",
  41622=>"000000000",
  41623=>"000000000",
  41624=>"111000000",
  41625=>"000000000",
  41626=>"111011011",
  41627=>"111111111",
  41628=>"010000110",
  41629=>"111101101",
  41630=>"100110110",
  41631=>"101101111",
  41632=>"111111010",
  41633=>"111111111",
  41634=>"111000000",
  41635=>"111111010",
  41636=>"011011011",
  41637=>"111100000",
  41638=>"000000000",
  41639=>"011111111",
  41640=>"000010111",
  41641=>"010000010",
  41642=>"000000000",
  41643=>"101111111",
  41644=>"001000100",
  41645=>"001000111",
  41646=>"111111100",
  41647=>"000000000",
  41648=>"010110000",
  41649=>"100101111",
  41650=>"001111111",
  41651=>"110110000",
  41652=>"100101111",
  41653=>"000000001",
  41654=>"001011001",
  41655=>"101111110",
  41656=>"111111001",
  41657=>"000000001",
  41658=>"001000001",
  41659=>"010000000",
  41660=>"111110111",
  41661=>"110100111",
  41662=>"010111111",
  41663=>"001001111",
  41664=>"111110111",
  41665=>"001111111",
  41666=>"000000001",
  41667=>"000000000",
  41668=>"111110000",
  41669=>"000000000",
  41670=>"111111111",
  41671=>"000000111",
  41672=>"000000000",
  41673=>"000000000",
  41674=>"110010000",
  41675=>"111110010",
  41676=>"000100111",
  41677=>"010011000",
  41678=>"000000000",
  41679=>"000100111",
  41680=>"111111000",
  41681=>"011011011",
  41682=>"000000001",
  41683=>"111101111",
  41684=>"111111001",
  41685=>"111111111",
  41686=>"111011010",
  41687=>"000000000",
  41688=>"111111111",
  41689=>"001000000",
  41690=>"110000000",
  41691=>"000000000",
  41692=>"000111101",
  41693=>"100110111",
  41694=>"111010000",
  41695=>"000000000",
  41696=>"111111111",
  41697=>"110111111",
  41698=>"110010000",
  41699=>"111111000",
  41700=>"110000000",
  41701=>"111111111",
  41702=>"010111111",
  41703=>"111111111",
  41704=>"110111110",
  41705=>"111111111",
  41706=>"000000000",
  41707=>"111011010",
  41708=>"111111111",
  41709=>"111111111",
  41710=>"000000111",
  41711=>"111001000",
  41712=>"000100000",
  41713=>"111001000",
  41714=>"000000000",
  41715=>"011011011",
  41716=>"000000000",
  41717=>"111101000",
  41718=>"000000000",
  41719=>"000010000",
  41720=>"000100110",
  41721=>"000000010",
  41722=>"111111111",
  41723=>"011000000",
  41724=>"100100000",
  41725=>"000000000",
  41726=>"111111110",
  41727=>"111111111",
  41728=>"001001011",
  41729=>"011011001",
  41730=>"111111111",
  41731=>"101101111",
  41732=>"111111111",
  41733=>"000000000",
  41734=>"000000000",
  41735=>"000001111",
  41736=>"000000000",
  41737=>"111111111",
  41738=>"111110000",
  41739=>"010000000",
  41740=>"001000000",
  41741=>"111111111",
  41742=>"011000000",
  41743=>"000000000",
  41744=>"000000000",
  41745=>"001001000",
  41746=>"111101111",
  41747=>"111111111",
  41748=>"111111000",
  41749=>"111111111",
  41750=>"110100100",
  41751=>"000000000",
  41752=>"100000001",
  41753=>"111100000",
  41754=>"111111111",
  41755=>"010000000",
  41756=>"011011011",
  41757=>"010000000",
  41758=>"000000000",
  41759=>"111000000",
  41760=>"011000000",
  41761=>"000000000",
  41762=>"000000000",
  41763=>"111111000",
  41764=>"111111001",
  41765=>"000000011",
  41766=>"000000000",
  41767=>"000000000",
  41768=>"000000110",
  41769=>"000000000",
  41770=>"111111100",
  41771=>"111111111",
  41772=>"000010010",
  41773=>"000000000",
  41774=>"111111111",
  41775=>"000001111",
  41776=>"000000000",
  41777=>"111111111",
  41778=>"111000000",
  41779=>"111111110",
  41780=>"011111011",
  41781=>"000000000",
  41782=>"000000110",
  41783=>"111111111",
  41784=>"000000000",
  41785=>"010000001",
  41786=>"110110111",
  41787=>"110000110",
  41788=>"110000100",
  41789=>"100001111",
  41790=>"110110000",
  41791=>"111110100",
  41792=>"000100000",
  41793=>"111111111",
  41794=>"011001001",
  41795=>"111111111",
  41796=>"111111111",
  41797=>"000000000",
  41798=>"000000011",
  41799=>"011001001",
  41800=>"111011000",
  41801=>"000000000",
  41802=>"111101101",
  41803=>"011011010",
  41804=>"111111011",
  41805=>"111111111",
  41806=>"100000000",
  41807=>"000110110",
  41808=>"010010000",
  41809=>"000000000",
  41810=>"111000000",
  41811=>"000000000",
  41812=>"000000111",
  41813=>"011111111",
  41814=>"111000000",
  41815=>"111011111",
  41816=>"100111111",
  41817=>"111111111",
  41818=>"000110111",
  41819=>"111111111",
  41820=>"111111011",
  41821=>"000000000",
  41822=>"010011111",
  41823=>"111111111",
  41824=>"000000100",
  41825=>"000000000",
  41826=>"111111011",
  41827=>"000000000",
  41828=>"000000000",
  41829=>"000000000",
  41830=>"000000000",
  41831=>"011001000",
  41832=>"001001000",
  41833=>"000000000",
  41834=>"110111101",
  41835=>"100000000",
  41836=>"100000000",
  41837=>"000001111",
  41838=>"101001111",
  41839=>"000000000",
  41840=>"111111111",
  41841=>"111111111",
  41842=>"000110111",
  41843=>"111111111",
  41844=>"111111000",
  41845=>"011001001",
  41846=>"111100100",
  41847=>"110110100",
  41848=>"000000111",
  41849=>"000000000",
  41850=>"111111001",
  41851=>"011000010",
  41852=>"000001000",
  41853=>"111111111",
  41854=>"000000000",
  41855=>"000000000",
  41856=>"110100110",
  41857=>"000110111",
  41858=>"000000000",
  41859=>"110000000",
  41860=>"110111111",
  41861=>"000111110",
  41862=>"111111111",
  41863=>"010000001",
  41864=>"111111111",
  41865=>"111111111",
  41866=>"000000111",
  41867=>"111111111",
  41868=>"100100111",
  41869=>"111001111",
  41870=>"000000000",
  41871=>"111111111",
  41872=>"000100111",
  41873=>"000000000",
  41874=>"110000000",
  41875=>"111111111",
  41876=>"111111011",
  41877=>"000000000",
  41878=>"010110110",
  41879=>"101001000",
  41880=>"000000000",
  41881=>"111000000",
  41882=>"000000000",
  41883=>"111101100",
  41884=>"000000110",
  41885=>"000000000",
  41886=>"000000110",
  41887=>"010000000",
  41888=>"010000000",
  41889=>"011000000",
  41890=>"111111111",
  41891=>"111111111",
  41892=>"000100111",
  41893=>"011000000",
  41894=>"111111000",
  41895=>"100000000",
  41896=>"110000000",
  41897=>"011000100",
  41898=>"001000000",
  41899=>"001111111",
  41900=>"111000000",
  41901=>"110000010",
  41902=>"111101100",
  41903=>"111111111",
  41904=>"101100100",
  41905=>"111111111",
  41906=>"100110111",
  41907=>"110111001",
  41908=>"000001101",
  41909=>"000000000",
  41910=>"111111111",
  41911=>"111111101",
  41912=>"000111111",
  41913=>"000000000",
  41914=>"000000000",
  41915=>"111111111",
  41916=>"111111111",
  41917=>"001011111",
  41918=>"000000000",
  41919=>"011001011",
  41920=>"000100100",
  41921=>"111101111",
  41922=>"011011000",
  41923=>"011011111",
  41924=>"111111111",
  41925=>"001001011",
  41926=>"000011000",
  41927=>"010111011",
  41928=>"011001000",
  41929=>"000100111",
  41930=>"001001111",
  41931=>"000000000",
  41932=>"101001000",
  41933=>"000000000",
  41934=>"111010000",
  41935=>"000110110",
  41936=>"000000001",
  41937=>"111110100",
  41938=>"000000000",
  41939=>"011000000",
  41940=>"000000000",
  41941=>"011011000",
  41942=>"000000000",
  41943=>"100000010",
  41944=>"111111111",
  41945=>"001000000",
  41946=>"000111110",
  41947=>"000000000",
  41948=>"001110110",
  41949=>"111111111",
  41950=>"011110100",
  41951=>"001001011",
  41952=>"111111000",
  41953=>"000001111",
  41954=>"111111111",
  41955=>"111111111",
  41956=>"111110011",
  41957=>"100000000",
  41958=>"110100100",
  41959=>"000000000",
  41960=>"100000101",
  41961=>"110110111",
  41962=>"000000000",
  41963=>"000100100",
  41964=>"111111111",
  41965=>"000000000",
  41966=>"110100111",
  41967=>"000000000",
  41968=>"110111111",
  41969=>"111110111",
  41970=>"111111111",
  41971=>"111111111",
  41972=>"011111111",
  41973=>"000110010",
  41974=>"111111111",
  41975=>"101111111",
  41976=>"000010110",
  41977=>"000100111",
  41978=>"100100011",
  41979=>"010000000",
  41980=>"011100110",
  41981=>"111111111",
  41982=>"001001111",
  41983=>"000111111",
  41984=>"000111100",
  41985=>"111110110",
  41986=>"000000111",
  41987=>"001001001",
  41988=>"111111111",
  41989=>"001001000",
  41990=>"000001111",
  41991=>"000000000",
  41992=>"001100000",
  41993=>"000000000",
  41994=>"001111111",
  41995=>"000110111",
  41996=>"000000000",
  41997=>"111111111",
  41998=>"000000001",
  41999=>"111000011",
  42000=>"011000000",
  42001=>"101001000",
  42002=>"111111111",
  42003=>"001111111",
  42004=>"111111111",
  42005=>"110000111",
  42006=>"110000001",
  42007=>"110110110",
  42008=>"001111111",
  42009=>"001001100",
  42010=>"000111010",
  42011=>"000001000",
  42012=>"111011111",
  42013=>"111111111",
  42014=>"000100000",
  42015=>"111111111",
  42016=>"110110110",
  42017=>"001001011",
  42018=>"111111111",
  42019=>"000000000",
  42020=>"000000000",
  42021=>"101000111",
  42022=>"101000000",
  42023=>"010000000",
  42024=>"011011111",
  42025=>"010111011",
  42026=>"000100100",
  42027=>"111111111",
  42028=>"110111111",
  42029=>"011110010",
  42030=>"000000110",
  42031=>"000000000",
  42032=>"100110111",
  42033=>"111111111",
  42034=>"000011111",
  42035=>"111111111",
  42036=>"000010111",
  42037=>"010011111",
  42038=>"111111111",
  42039=>"110000000",
  42040=>"111100111",
  42041=>"100110111",
  42042=>"111100110",
  42043=>"111111111",
  42044=>"100000000",
  42045=>"111111111",
  42046=>"000000000",
  42047=>"100000000",
  42048=>"111111111",
  42049=>"000010000",
  42050=>"000100001",
  42051=>"000000000",
  42052=>"111111111",
  42053=>"101100100",
  42054=>"100000000",
  42055=>"111111111",
  42056=>"000000000",
  42057=>"111111000",
  42058=>"111111111",
  42059=>"111110111",
  42060=>"110011111",
  42061=>"111000001",
  42062=>"000000000",
  42063=>"000000000",
  42064=>"111101111",
  42065=>"111011000",
  42066=>"111111111",
  42067=>"010111110",
  42068=>"101000100",
  42069=>"011100111",
  42070=>"000110000",
  42071=>"100100100",
  42072=>"000000000",
  42073=>"000000000",
  42074=>"101111010",
  42075=>"100100110",
  42076=>"000000000",
  42077=>"110110111",
  42078=>"000000010",
  42079=>"000100101",
  42080=>"001111111",
  42081=>"000001000",
  42082=>"000000000",
  42083=>"000000000",
  42084=>"111000100",
  42085=>"100000100",
  42086=>"000000000",
  42087=>"110111000",
  42088=>"000000010",
  42089=>"111111101",
  42090=>"010111111",
  42091=>"000000111",
  42092=>"000000000",
  42093=>"011111111",
  42094=>"110000111",
  42095=>"111111111",
  42096=>"000111111",
  42097=>"000001111",
  42098=>"000000000",
  42099=>"000000100",
  42100=>"010010100",
  42101=>"010000101",
  42102=>"100110110",
  42103=>"001000000",
  42104=>"111111111",
  42105=>"000100100",
  42106=>"000000001",
  42107=>"111111111",
  42108=>"111111111",
  42109=>"100000001",
  42110=>"000111111",
  42111=>"000000000",
  42112=>"111111110",
  42113=>"110000000",
  42114=>"000000000",
  42115=>"111111111",
  42116=>"011111111",
  42117=>"111000000",
  42118=>"001100100",
  42119=>"111111111",
  42120=>"000000101",
  42121=>"111111111",
  42122=>"000000000",
  42123=>"111101000",
  42124=>"000000000",
  42125=>"000000000",
  42126=>"000000000",
  42127=>"100110110",
  42128=>"111111011",
  42129=>"111111011",
  42130=>"001000100",
  42131=>"000000110",
  42132=>"111111111",
  42133=>"100000000",
  42134=>"010000100",
  42135=>"100000110",
  42136=>"000111111",
  42137=>"000000000",
  42138=>"100100111",
  42139=>"011111111",
  42140=>"100110111",
  42141=>"111111100",
  42142=>"000100100",
  42143=>"000110111",
  42144=>"110000110",
  42145=>"111111000",
  42146=>"000010001",
  42147=>"000000000",
  42148=>"000000001",
  42149=>"110110110",
  42150=>"111101111",
  42151=>"100110100",
  42152=>"000010000",
  42153=>"111111101",
  42154=>"000000000",
  42155=>"000101001",
  42156=>"000100110",
  42157=>"000000111",
  42158=>"111111111",
  42159=>"110000110",
  42160=>"000011000",
  42161=>"000100001",
  42162=>"110010010",
  42163=>"000000000",
  42164=>"001000000",
  42165=>"001001111",
  42166=>"110000000",
  42167=>"110101100",
  42168=>"111110111",
  42169=>"100000000",
  42170=>"111000011",
  42171=>"000000000",
  42172=>"111111111",
  42173=>"000000111",
  42174=>"111111111",
  42175=>"111110111",
  42176=>"110100111",
  42177=>"010110111",
  42178=>"110110100",
  42179=>"000000000",
  42180=>"000011000",
  42181=>"000000000",
  42182=>"110111110",
  42183=>"111111111",
  42184=>"111011110",
  42185=>"111110111",
  42186=>"000000000",
  42187=>"111011111",
  42188=>"001011100",
  42189=>"100100111",
  42190=>"110110111",
  42191=>"001000000",
  42192=>"101001001",
  42193=>"000000000",
  42194=>"111111111",
  42195=>"000000000",
  42196=>"111001001",
  42197=>"111111111",
  42198=>"000000111",
  42199=>"000000000",
  42200=>"111011000",
  42201=>"100100001",
  42202=>"111000011",
  42203=>"001000011",
  42204=>"000000000",
  42205=>"111111111",
  42206=>"100100111",
  42207=>"111111110",
  42208=>"011011011",
  42209=>"011111000",
  42210=>"000000100",
  42211=>"111111111",
  42212=>"111000000",
  42213=>"000111111",
  42214=>"000000000",
  42215=>"000000001",
  42216=>"000000000",
  42217=>"011011111",
  42218=>"000100111",
  42219=>"000110111",
  42220=>"010000001",
  42221=>"110000000",
  42222=>"000111111",
  42223=>"111001011",
  42224=>"111111111",
  42225=>"111111111",
  42226=>"000000000",
  42227=>"000000000",
  42228=>"000000000",
  42229=>"100000110",
  42230=>"111111101",
  42231=>"000000000",
  42232=>"000000000",
  42233=>"111111111",
  42234=>"110001001",
  42235=>"111111111",
  42236=>"111111001",
  42237=>"011011001",
  42238=>"000000111",
  42239=>"000000111",
  42240=>"000000000",
  42241=>"111011011",
  42242=>"000001101",
  42243=>"101101000",
  42244=>"000000000",
  42245=>"000000000",
  42246=>"000000111",
  42247=>"000001001",
  42248=>"000111110",
  42249=>"000000101",
  42250=>"001001111",
  42251=>"111111111",
  42252=>"110000000",
  42253=>"111111011",
  42254=>"111111111",
  42255=>"111111011",
  42256=>"111111111",
  42257=>"111101101",
  42258=>"011111111",
  42259=>"011111110",
  42260=>"101100000",
  42261=>"000001011",
  42262=>"100100100",
  42263=>"000000000",
  42264=>"110011011",
  42265=>"111111111",
  42266=>"110111111",
  42267=>"111000000",
  42268=>"111111111",
  42269=>"000000000",
  42270=>"101111111",
  42271=>"100101001",
  42272=>"110110111",
  42273=>"111111111",
  42274=>"000000000",
  42275=>"101100100",
  42276=>"000000000",
  42277=>"100110000",
  42278=>"000000000",
  42279=>"010000111",
  42280=>"000000111",
  42281=>"000000000",
  42282=>"111010100",
  42283=>"001111111",
  42284=>"101000100",
  42285=>"111111001",
  42286=>"111111000",
  42287=>"000000110",
  42288=>"011001001",
  42289=>"000000001",
  42290=>"111111100",
  42291=>"000001111",
  42292=>"000000000",
  42293=>"001001101",
  42294=>"000000000",
  42295=>"111001001",
  42296=>"110010000",
  42297=>"000100111",
  42298=>"111100111",
  42299=>"111111111",
  42300=>"000000111",
  42301=>"000110110",
  42302=>"000000000",
  42303=>"111000011",
  42304=>"000111111",
  42305=>"110000000",
  42306=>"000000000",
  42307=>"000000000",
  42308=>"111101000",
  42309=>"110000000",
  42310=>"110111111",
  42311=>"000000000",
  42312=>"000000000",
  42313=>"110000000",
  42314=>"001001000",
  42315=>"000000000",
  42316=>"001000100",
  42317=>"111111000",
  42318=>"111000000",
  42319=>"111111000",
  42320=>"001111111",
  42321=>"000000000",
  42322=>"000110000",
  42323=>"110110110",
  42324=>"000011000",
  42325=>"011011001",
  42326=>"010000110",
  42327=>"000000000",
  42328=>"000000000",
  42329=>"000001111",
  42330=>"111111111",
  42331=>"110111111",
  42332=>"010110111",
  42333=>"101001000",
  42334=>"110111111",
  42335=>"000000100",
  42336=>"000011000",
  42337=>"111111111",
  42338=>"000110000",
  42339=>"111111111",
  42340=>"111011111",
  42341=>"000100111",
  42342=>"111111111",
  42343=>"100100100",
  42344=>"100000000",
  42345=>"000111111",
  42346=>"111111111",
  42347=>"000110110",
  42348=>"110110111",
  42349=>"000000000",
  42350=>"000101000",
  42351=>"000001001",
  42352=>"000000011",
  42353=>"001001111",
  42354=>"000000011",
  42355=>"111100111",
  42356=>"000000011",
  42357=>"000000111",
  42358=>"001111010",
  42359=>"000110000",
  42360=>"000000111",
  42361=>"000000000",
  42362=>"111000000",
  42363=>"111110100",
  42364=>"010000111",
  42365=>"000000000",
  42366=>"111111111",
  42367=>"111111000",
  42368=>"100110111",
  42369=>"111111110",
  42370=>"110100011",
  42371=>"000000000",
  42372=>"000100111",
  42373=>"110110000",
  42374=>"000000000",
  42375=>"001111010",
  42376=>"110111111",
  42377=>"000101111",
  42378=>"000100110",
  42379=>"000100111",
  42380=>"000000000",
  42381=>"000101110",
  42382=>"111001111",
  42383=>"000000001",
  42384=>"111111111",
  42385=>"111111110",
  42386=>"111111111",
  42387=>"110110000",
  42388=>"001111111",
  42389=>"111100111",
  42390=>"000010000",
  42391=>"000001001",
  42392=>"000000000",
  42393=>"001010111",
  42394=>"111111111",
  42395=>"111111111",
  42396=>"110111111",
  42397=>"000000101",
  42398=>"000001011",
  42399=>"111100000",
  42400=>"011100111",
  42401=>"000000001",
  42402=>"010000000",
  42403=>"000011000",
  42404=>"000010000",
  42405=>"000000000",
  42406=>"111101000",
  42407=>"000000000",
  42408=>"010010000",
  42409=>"110110000",
  42410=>"110111000",
  42411=>"111111111",
  42412=>"100111000",
  42413=>"000010110",
  42414=>"111111000",
  42415=>"111001001",
  42416=>"100110011",
  42417=>"111001000",
  42418=>"011111111",
  42419=>"000100000",
  42420=>"000000000",
  42421=>"100111111",
  42422=>"110110100",
  42423=>"000000000",
  42424=>"000000010",
  42425=>"000000000",
  42426=>"110001001",
  42427=>"111111111",
  42428=>"110111111",
  42429=>"000000000",
  42430=>"000000000",
  42431=>"000000011",
  42432=>"100100111",
  42433=>"000000111",
  42434=>"000000011",
  42435=>"100000000",
  42436=>"000000100",
  42437=>"100110110",
  42438=>"000011111",
  42439=>"000011000",
  42440=>"000100000",
  42441=>"111100100",
  42442=>"000000110",
  42443=>"111111111",
  42444=>"000010111",
  42445=>"000000000",
  42446=>"111110000",
  42447=>"000000000",
  42448=>"000000000",
  42449=>"111111111",
  42450=>"100000000",
  42451=>"111111111",
  42452=>"111111101",
  42453=>"111111111",
  42454=>"000000111",
  42455=>"000000000",
  42456=>"001111000",
  42457=>"010000000",
  42458=>"111111111",
  42459=>"110111000",
  42460=>"110100110",
  42461=>"000011000",
  42462=>"110000011",
  42463=>"111000001",
  42464=>"000000011",
  42465=>"001001111",
  42466=>"111111100",
  42467=>"101111111",
  42468=>"111111111",
  42469=>"001000011",
  42470=>"000100111",
  42471=>"111100000",
  42472=>"011101100",
  42473=>"000000000",
  42474=>"111111111",
  42475=>"111111111",
  42476=>"111111111",
  42477=>"000000100",
  42478=>"111111111",
  42479=>"100000000",
  42480=>"100000111",
  42481=>"100100111",
  42482=>"000000000",
  42483=>"111111111",
  42484=>"011011111",
  42485=>"111101100",
  42486=>"000000000",
  42487=>"001000011",
  42488=>"110110111",
  42489=>"000011011",
  42490=>"111101111",
  42491=>"000000110",
  42492=>"110100100",
  42493=>"010111000",
  42494=>"101101111",
  42495=>"111001001",
  42496=>"000011001",
  42497=>"001111011",
  42498=>"111111111",
  42499=>"100100100",
  42500=>"111111000",
  42501=>"100111111",
  42502=>"000000000",
  42503=>"111111111",
  42504=>"000100100",
  42505=>"000000000",
  42506=>"111111111",
  42507=>"000000000",
  42508=>"000000110",
  42509=>"000000000",
  42510=>"111111111",
  42511=>"111111111",
  42512=>"101001001",
  42513=>"000000000",
  42514=>"000000000",
  42515=>"110110000",
  42516=>"111111111",
  42517=>"000000000",
  42518=>"111111111",
  42519=>"100000000",
  42520=>"001001101",
  42521=>"000101101",
  42522=>"000000100",
  42523=>"100100111",
  42524=>"111111101",
  42525=>"000000000",
  42526=>"000000000",
  42527=>"000000000",
  42528=>"111000000",
  42529=>"111111111",
  42530=>"100000000",
  42531=>"100001111",
  42532=>"111111111",
  42533=>"111111111",
  42534=>"111101111",
  42535=>"111111001",
  42536=>"111111000",
  42537=>"000000101",
  42538=>"111111001",
  42539=>"011001011",
  42540=>"111101111",
  42541=>"100111111",
  42542=>"111111111",
  42543=>"111000010",
  42544=>"111111111",
  42545=>"000000000",
  42546=>"000100100",
  42547=>"111111110",
  42548=>"000000000",
  42549=>"000100100",
  42550=>"101111111",
  42551=>"111111000",
  42552=>"000000000",
  42553=>"111111001",
  42554=>"111111000",
  42555=>"000000000",
  42556=>"111111111",
  42557=>"110110100",
  42558=>"000110110",
  42559=>"111101101",
  42560=>"100111111",
  42561=>"010110110",
  42562=>"111111101",
  42563=>"111111111",
  42564=>"000000001",
  42565=>"111111111",
  42566=>"011001000",
  42567=>"111011011",
  42568=>"001011111",
  42569=>"101101111",
  42570=>"000000000",
  42571=>"011011000",
  42572=>"001111111",
  42573=>"111011111",
  42574=>"111111100",
  42575=>"000000110",
  42576=>"001001000",
  42577=>"111110110",
  42578=>"111111011",
  42579=>"100100000",
  42580=>"000000010",
  42581=>"110111001",
  42582=>"011000000",
  42583=>"111111111",
  42584=>"111111111",
  42585=>"111001101",
  42586=>"111111111",
  42587=>"000000000",
  42588=>"111111111",
  42589=>"111111111",
  42590=>"111000000",
  42591=>"000000000",
  42592=>"110000000",
  42593=>"111110110",
  42594=>"000000100",
  42595=>"111111111",
  42596=>"111111101",
  42597=>"000000000",
  42598=>"111111111",
  42599=>"111011111",
  42600=>"100110111",
  42601=>"111111111",
  42602=>"111111000",
  42603=>"000000000",
  42604=>"001000011",
  42605=>"101100000",
  42606=>"101000111",
  42607=>"111000000",
  42608=>"000000000",
  42609=>"000000000",
  42610=>"111111111",
  42611=>"111111111",
  42612=>"111111001",
  42613=>"000000000",
  42614=>"000001111",
  42615=>"001000000",
  42616=>"111111111",
  42617=>"000000000",
  42618=>"111110000",
  42619=>"101101100",
  42620=>"110110110",
  42621=>"111111111",
  42622=>"100000000",
  42623=>"111111111",
  42624=>"111111111",
  42625=>"000000000",
  42626=>"101101100",
  42627=>"011011000",
  42628=>"100000110",
  42629=>"000000000",
  42630=>"111111111",
  42631=>"110000000",
  42632=>"000000000",
  42633=>"111110111",
  42634=>"111111011",
  42635=>"110110000",
  42636=>"111111111",
  42637=>"000000111",
  42638=>"000000010",
  42639=>"110110000",
  42640=>"011111111",
  42641=>"000000010",
  42642=>"000010101",
  42643=>"111001001",
  42644=>"001000000",
  42645=>"011011111",
  42646=>"011111111",
  42647=>"000000000",
  42648=>"111111111",
  42649=>"111111111",
  42650=>"111111100",
  42651=>"111111111",
  42652=>"111111001",
  42653=>"101001001",
  42654=>"010000110",
  42655=>"000100100",
  42656=>"111111100",
  42657=>"000011111",
  42658=>"001000000",
  42659=>"111001000",
  42660=>"000101001",
  42661=>"000000000",
  42662=>"010110110",
  42663=>"000000000",
  42664=>"111111111",
  42665=>"111111111",
  42666=>"111001111",
  42667=>"111111111",
  42668=>"111111111",
  42669=>"001011110",
  42670=>"000100100",
  42671=>"100000000",
  42672=>"111111111",
  42673=>"100010000",
  42674=>"000000000",
  42675=>"000010000",
  42676=>"000000000",
  42677=>"111100000",
  42678=>"001000000",
  42679=>"000010000",
  42680=>"111111100",
  42681=>"000000110",
  42682=>"011111111",
  42683=>"000000100",
  42684=>"111111000",
  42685=>"001001000",
  42686=>"100000000",
  42687=>"111111111",
  42688=>"110100110",
  42689=>"000000000",
  42690=>"111111111",
  42691=>"001101111",
  42692=>"111000000",
  42693=>"111111111",
  42694=>"100100100",
  42695=>"001101101",
  42696=>"000010000",
  42697=>"111111111",
  42698=>"111111001",
  42699=>"000001001",
  42700=>"100000000",
  42701=>"000000000",
  42702=>"011010000",
  42703=>"010000000",
  42704=>"111010000",
  42705=>"100100100",
  42706=>"000000010",
  42707=>"000000000",
  42708=>"000000111",
  42709=>"101001001",
  42710=>"111111111",
  42711=>"001000000",
  42712=>"111111111",
  42713=>"111111011",
  42714=>"000000000",
  42715=>"000000000",
  42716=>"001101001",
  42717=>"000000000",
  42718=>"001011000",
  42719=>"100000000",
  42720=>"001000000",
  42721=>"000000000",
  42722=>"000000000",
  42723=>"100000100",
  42724=>"000000000",
  42725=>"001000000",
  42726=>"010111010",
  42727=>"000000000",
  42728=>"111110000",
  42729=>"001000000",
  42730=>"001001001",
  42731=>"000100111",
  42732=>"111111000",
  42733=>"111111111",
  42734=>"011011111",
  42735=>"111100100",
  42736=>"111100000",
  42737=>"111111100",
  42738=>"000000000",
  42739=>"010000000",
  42740=>"000000000",
  42741=>"000000000",
  42742=>"101111111",
  42743=>"111111111",
  42744=>"000000000",
  42745=>"111111111",
  42746=>"111111111",
  42747=>"011000000",
  42748=>"000000001",
  42749=>"000100000",
  42750=>"000000000",
  42751=>"110000000",
  42752=>"111111111",
  42753=>"000000001",
  42754=>"111111111",
  42755=>"000000010",
  42756=>"111110000",
  42757=>"001000000",
  42758=>"100000000",
  42759=>"111110110",
  42760=>"000000100",
  42761=>"000011000",
  42762=>"111111111",
  42763=>"000000000",
  42764=>"100110100",
  42765=>"110111111",
  42766=>"111111101",
  42767=>"100110000",
  42768=>"000000000",
  42769=>"111111111",
  42770=>"001000000",
  42771=>"111111111",
  42772=>"000000000",
  42773=>"000000001",
  42774=>"000000111",
  42775=>"111111111",
  42776=>"000000000",
  42777=>"001111111",
  42778=>"111111111",
  42779=>"000000100",
  42780=>"001101011",
  42781=>"000000000",
  42782=>"111111111",
  42783=>"000000000",
  42784=>"101110000",
  42785=>"111111011",
  42786=>"111110111",
  42787=>"000100111",
  42788=>"011011111",
  42789=>"001110111",
  42790=>"000010011",
  42791=>"110000000",
  42792=>"001001111",
  42793=>"000000000",
  42794=>"110110110",
  42795=>"000000000",
  42796=>"000000000",
  42797=>"100100000",
  42798=>"110000111",
  42799=>"001000101",
  42800=>"011001011",
  42801=>"111111111",
  42802=>"110110111",
  42803=>"111111111",
  42804=>"111111111",
  42805=>"000000000",
  42806=>"101111111",
  42807=>"001111111",
  42808=>"000111111",
  42809=>"111111111",
  42810=>"000000000",
  42811=>"110110110",
  42812=>"111111111",
  42813=>"000000000",
  42814=>"111111111",
  42815=>"111111111",
  42816=>"001000000",
  42817=>"111011111",
  42818=>"111111111",
  42819=>"111101111",
  42820=>"111111111",
  42821=>"111111111",
  42822=>"000000000",
  42823=>"000000000",
  42824=>"111101101",
  42825=>"111111111",
  42826=>"111011000",
  42827=>"100100100",
  42828=>"001000000",
  42829=>"111111110",
  42830=>"000000000",
  42831=>"111111110",
  42832=>"000000000",
  42833=>"000100100",
  42834=>"111101111",
  42835=>"000001111",
  42836=>"111101111",
  42837=>"001001011",
  42838=>"000000000",
  42839=>"000000000",
  42840=>"111111111",
  42841=>"111111111",
  42842=>"111111111",
  42843=>"000000000",
  42844=>"111111111",
  42845=>"111111001",
  42846=>"000000000",
  42847=>"001001001",
  42848=>"111111111",
  42849=>"011111000",
  42850=>"000000100",
  42851=>"001000001",
  42852=>"000000000",
  42853=>"111111011",
  42854=>"000111111",
  42855=>"001001111",
  42856=>"111111111",
  42857=>"000000110",
  42858=>"111111111",
  42859=>"101000000",
  42860=>"000001001",
  42861=>"001111000",
  42862=>"000000000",
  42863=>"111111111",
  42864=>"111101111",
  42865=>"010000000",
  42866=>"111111111",
  42867=>"000000000",
  42868=>"111100000",
  42869=>"111111110",
  42870=>"111111111",
  42871=>"110110000",
  42872=>"111100111",
  42873=>"000000000",
  42874=>"100000000",
  42875=>"000000000",
  42876=>"000000000",
  42877=>"111111111",
  42878=>"111111111",
  42879=>"111111111",
  42880=>"000001000",
  42881=>"100101101",
  42882=>"111111111",
  42883=>"111111111",
  42884=>"111111001",
  42885=>"111111110",
  42886=>"000000000",
  42887=>"111111111",
  42888=>"100000001",
  42889=>"111111111",
  42890=>"101111111",
  42891=>"111111000",
  42892=>"111111111",
  42893=>"000000110",
  42894=>"011111110",
  42895=>"000000000",
  42896=>"000000001",
  42897=>"000000001",
  42898=>"011111110",
  42899=>"111111111",
  42900=>"111111000",
  42901=>"000000010",
  42902=>"111111111",
  42903=>"000000000",
  42904=>"111101000",
  42905=>"000000000",
  42906=>"111111111",
  42907=>"111111111",
  42908=>"000000000",
  42909=>"000000000",
  42910=>"000000000",
  42911=>"000000111",
  42912=>"111111111",
  42913=>"110010110",
  42914=>"000000110",
  42915=>"111111111",
  42916=>"100100100",
  42917=>"111111001",
  42918=>"111011011",
  42919=>"000000100",
  42920=>"000000000",
  42921=>"000000101",
  42922=>"000000000",
  42923=>"000110110",
  42924=>"111101101",
  42925=>"000000000",
  42926=>"111101111",
  42927=>"111111001",
  42928=>"001111001",
  42929=>"111111110",
  42930=>"010000000",
  42931=>"111111000",
  42932=>"000001000",
  42933=>"000000000",
  42934=>"110111111",
  42935=>"111111111",
  42936=>"111111111",
  42937=>"111111111",
  42938=>"000000000",
  42939=>"111001000",
  42940=>"110011000",
  42941=>"111111111",
  42942=>"110111100",
  42943=>"100000000",
  42944=>"011000001",
  42945=>"100100111",
  42946=>"000000000",
  42947=>"111101100",
  42948=>"110111000",
  42949=>"011110111",
  42950=>"000011000",
  42951=>"000000000",
  42952=>"111111111",
  42953=>"000000000",
  42954=>"001011111",
  42955=>"000000111",
  42956=>"000111000",
  42957=>"111111111",
  42958=>"111111111",
  42959=>"010110010",
  42960=>"001000000",
  42961=>"111111000",
  42962=>"111111111",
  42963=>"111111111",
  42964=>"110110110",
  42965=>"001000000",
  42966=>"000100100",
  42967=>"000111111",
  42968=>"000000001",
  42969=>"110011111",
  42970=>"011000000",
  42971=>"111010000",
  42972=>"000100000",
  42973=>"111111111",
  42974=>"111111111",
  42975=>"000000001",
  42976=>"000000000",
  42977=>"000000100",
  42978=>"000110000",
  42979=>"000010100",
  42980=>"001000110",
  42981=>"001000111",
  42982=>"111100000",
  42983=>"111111111",
  42984=>"000000000",
  42985=>"111111111",
  42986=>"000000111",
  42987=>"111011000",
  42988=>"110110110",
  42989=>"000000100",
  42990=>"111000000",
  42991=>"110111111",
  42992=>"000000000",
  42993=>"000000111",
  42994=>"000000000",
  42995=>"111111111",
  42996=>"000000000",
  42997=>"111111111",
  42998=>"111001000",
  42999=>"111011001",
  43000=>"111111111",
  43001=>"011001111",
  43002=>"111111110",
  43003=>"111111110",
  43004=>"110110100",
  43005=>"000001100",
  43006=>"000000000",
  43007=>"111111011",
  43008=>"000100110",
  43009=>"000000100",
  43010=>"111111111",
  43011=>"111010011",
  43012=>"100011111",
  43013=>"110100111",
  43014=>"000000000",
  43015=>"111011001",
  43016=>"111000111",
  43017=>"000000000",
  43018=>"111111111",
  43019=>"111111111",
  43020=>"110111111",
  43021=>"111111111",
  43022=>"111101111",
  43023=>"111111111",
  43024=>"111011001",
  43025=>"011111111",
  43026=>"100000000",
  43027=>"111111111",
  43028=>"001011111",
  43029=>"000000111",
  43030=>"000000000",
  43031=>"011011011",
  43032=>"110101111",
  43033=>"111111111",
  43034=>"011000000",
  43035=>"000000001",
  43036=>"000000000",
  43037=>"000000000",
  43038=>"110110000",
  43039=>"100000100",
  43040=>"000000000",
  43041=>"110111111",
  43042=>"000001000",
  43043=>"111111111",
  43044=>"111111001",
  43045=>"111111111",
  43046=>"111111111",
  43047=>"010110111",
  43048=>"000001010",
  43049=>"000111111",
  43050=>"001101100",
  43051=>"000101101",
  43052=>"001111111",
  43053=>"000000000",
  43054=>"111111111",
  43055=>"000000101",
  43056=>"001001000",
  43057=>"001001111",
  43058=>"111111011",
  43059=>"000110111",
  43060=>"000010011",
  43061=>"000000000",
  43062=>"000000001",
  43063=>"000001011",
  43064=>"011111100",
  43065=>"111100000",
  43066=>"000111110",
  43067=>"000000000",
  43068=>"111101111",
  43069=>"111010000",
  43070=>"111111111",
  43071=>"101000101",
  43072=>"111111111",
  43073=>"101101101",
  43074=>"000001000",
  43075=>"000000000",
  43076=>"000000000",
  43077=>"000000100",
  43078=>"111111010",
  43079=>"000000000",
  43080=>"111011101",
  43081=>"001000011",
  43082=>"010111111",
  43083=>"110110111",
  43084=>"000000101",
  43085=>"111111000",
  43086=>"000000000",
  43087=>"111111111",
  43088=>"100000000",
  43089=>"011011000",
  43090=>"011000000",
  43091=>"110111000",
  43092=>"000000000",
  43093=>"000000101",
  43094=>"111111111",
  43095=>"000000000",
  43096=>"111111111",
  43097=>"111100111",
  43098=>"111111111",
  43099=>"111101100",
  43100=>"000001000",
  43101=>"011011000",
  43102=>"111111111",
  43103=>"110110010",
  43104=>"111111111",
  43105=>"111110001",
  43106=>"111000000",
  43107=>"111111111",
  43108=>"111000111",
  43109=>"000000011",
  43110=>"000000000",
  43111=>"111111111",
  43112=>"111111111",
  43113=>"000000000",
  43114=>"000010111",
  43115=>"000000011",
  43116=>"011111011",
  43117=>"100000000",
  43118=>"111110110",
  43119=>"111111111",
  43120=>"000000100",
  43121=>"111011010",
  43122=>"100110100",
  43123=>"000000000",
  43124=>"000000000",
  43125=>"110111010",
  43126=>"111111111",
  43127=>"011111111",
  43128=>"111111101",
  43129=>"101001000",
  43130=>"111111100",
  43131=>"011011000",
  43132=>"111111111",
  43133=>"111111111",
  43134=>"111001111",
  43135=>"000100111",
  43136=>"100001111",
  43137=>"111111111",
  43138=>"101001111",
  43139=>"011101000",
  43140=>"001111111",
  43141=>"001000000",
  43142=>"111111111",
  43143=>"000000001",
  43144=>"000000100",
  43145=>"000110111",
  43146=>"111101101",
  43147=>"000000000",
  43148=>"111111111",
  43149=>"111111111",
  43150=>"001000111",
  43151=>"100000000",
  43152=>"000000000",
  43153=>"000000100",
  43154=>"111111111",
  43155=>"001001000",
  43156=>"001101001",
  43157=>"010011001",
  43158=>"000100100",
  43159=>"111111001",
  43160=>"001001111",
  43161=>"111000000",
  43162=>"111001110",
  43163=>"000000000",
  43164=>"011111111",
  43165=>"101100100",
  43166=>"000000000",
  43167=>"000011111",
  43168=>"111111111",
  43169=>"001001000",
  43170=>"110011001",
  43171=>"000000110",
  43172=>"111111111",
  43173=>"000000101",
  43174=>"111111000",
  43175=>"000000000",
  43176=>"111111111",
  43177=>"111001111",
  43178=>"110111001",
  43179=>"000000000",
  43180=>"111111111",
  43181=>"000011111",
  43182=>"000001111",
  43183=>"111111111",
  43184=>"110111111",
  43185=>"110110101",
  43186=>"011011000",
  43187=>"000000000",
  43188=>"101000100",
  43189=>"000001000",
  43190=>"111100000",
  43191=>"100111110",
  43192=>"000000000",
  43193=>"000000000",
  43194=>"111001111",
  43195=>"000000000",
  43196=>"000000111",
  43197=>"000001111",
  43198=>"100100100",
  43199=>"111111111",
  43200=>"111100110",
  43201=>"000000000",
  43202=>"100111011",
  43203=>"000000000",
  43204=>"000000000",
  43205=>"110101101",
  43206=>"111111111",
  43207=>"001111011",
  43208=>"111111111",
  43209=>"111111010",
  43210=>"111111011",
  43211=>"111011001",
  43212=>"001011011",
  43213=>"000011011",
  43214=>"000000100",
  43215=>"111100000",
  43216=>"110110111",
  43217=>"111101100",
  43218=>"111111111",
  43219=>"000100110",
  43220=>"010001001",
  43221=>"000000010",
  43222=>"000000000",
  43223=>"110111111",
  43224=>"000000110",
  43225=>"011011111",
  43226=>"110000000",
  43227=>"111111101",
  43228=>"111000100",
  43229=>"010000000",
  43230=>"000000000",
  43231=>"010110111",
  43232=>"111111111",
  43233=>"111101111",
  43234=>"111111100",
  43235=>"000001000",
  43236=>"100000000",
  43237=>"110011000",
  43238=>"101111001",
  43239=>"110000111",
  43240=>"111111111",
  43241=>"000000100",
  43242=>"001001000",
  43243=>"001001111",
  43244=>"000000000",
  43245=>"110111111",
  43246=>"111111111",
  43247=>"111010000",
  43248=>"111111111",
  43249=>"000000011",
  43250=>"000000000",
  43251=>"000011011",
  43252=>"000000000",
  43253=>"000011011",
  43254=>"011111111",
  43255=>"111001000",
  43256=>"001011000",
  43257=>"000110000",
  43258=>"000001111",
  43259=>"111011011",
  43260=>"100000000",
  43261=>"100110111",
  43262=>"100110000",
  43263=>"111110000",
  43264=>"001000100",
  43265=>"011000000",
  43266=>"111111111",
  43267=>"000000000",
  43268=>"011110111",
  43269=>"001000000",
  43270=>"101000000",
  43271=>"111101001",
  43272=>"001011100",
  43273=>"111000101",
  43274=>"001111111",
  43275=>"000011000",
  43276=>"111000010",
  43277=>"111111111",
  43278=>"011011111",
  43279=>"011111011",
  43280=>"000000111",
  43281=>"000000000",
  43282=>"111011111",
  43283=>"000000101",
  43284=>"111111001",
  43285=>"000111111",
  43286=>"000000000",
  43287=>"000111111",
  43288=>"100100000",
  43289=>"110000000",
  43290=>"100001001",
  43291=>"111100000",
  43292=>"111001101",
  43293=>"000000000",
  43294=>"100111111",
  43295=>"110010000",
  43296=>"111111111",
  43297=>"111111101",
  43298=>"000000000",
  43299=>"011011000",
  43300=>"100100000",
  43301=>"111111001",
  43302=>"111111011",
  43303=>"000100100",
  43304=>"100000000",
  43305=>"111011000",
  43306=>"110111111",
  43307=>"000110000",
  43308=>"000000000",
  43309=>"000100100",
  43310=>"000000111",
  43311=>"100001001",
  43312=>"110111000",
  43313=>"101000000",
  43314=>"110000000",
  43315=>"111000100",
  43316=>"111111111",
  43317=>"011000110",
  43318=>"111111011",
  43319=>"111101001",
  43320=>"111111000",
  43321=>"111000000",
  43322=>"100000000",
  43323=>"111111111",
  43324=>"000000000",
  43325=>"000000010",
  43326=>"101001101",
  43327=>"000000000",
  43328=>"011001000",
  43329=>"000000000",
  43330=>"111111111",
  43331=>"000000110",
  43332=>"000001111",
  43333=>"111111000",
  43334=>"000000000",
  43335=>"000000000",
  43336=>"011000000",
  43337=>"000000111",
  43338=>"100111111",
  43339=>"000100000",
  43340=>"000001001",
  43341=>"011001101",
  43342=>"000000000",
  43343=>"010111011",
  43344=>"110010000",
  43345=>"000000000",
  43346=>"100101000",
  43347=>"101111111",
  43348=>"000001000",
  43349=>"111111111",
  43350=>"100000000",
  43351=>"011000000",
  43352=>"111111101",
  43353=>"111011000",
  43354=>"111111111",
  43355=>"011101110",
  43356=>"111001000",
  43357=>"101111111",
  43358=>"000001100",
  43359=>"000001011",
  43360=>"000100111",
  43361=>"000000000",
  43362=>"001001001",
  43363=>"001111111",
  43364=>"100010000",
  43365=>"000000000",
  43366=>"011011111",
  43367=>"000111111",
  43368=>"011111010",
  43369=>"110111111",
  43370=>"000100000",
  43371=>"111111111",
  43372=>"110110000",
  43373=>"000000000",
  43374=>"000111111",
  43375=>"110111001",
  43376=>"111111111",
  43377=>"111111111",
  43378=>"000000111",
  43379=>"111111111",
  43380=>"111111111",
  43381=>"000000000",
  43382=>"000000000",
  43383=>"111111111",
  43384=>"000000000",
  43385=>"111111100",
  43386=>"111111111",
  43387=>"100110111",
  43388=>"000000000",
  43389=>"001001001",
  43390=>"111110000",
  43391=>"111111111",
  43392=>"000000011",
  43393=>"111111111",
  43394=>"000000001",
  43395=>"000000000",
  43396=>"100000000",
  43397=>"000000010",
  43398=>"110100000",
  43399=>"111101111",
  43400=>"100100111",
  43401=>"111110000",
  43402=>"000000011",
  43403=>"111111000",
  43404=>"101001111",
  43405=>"000001110",
  43406=>"111111111",
  43407=>"100000000",
  43408=>"011001001",
  43409=>"100111111",
  43410=>"111101100",
  43411=>"000000000",
  43412=>"000010000",
  43413=>"000001011",
  43414=>"100000000",
  43415=>"000100100",
  43416=>"000000000",
  43417=>"111111100",
  43418=>"110000101",
  43419=>"000000000",
  43420=>"000000111",
  43421=>"111010011",
  43422=>"101110111",
  43423=>"100111111",
  43424=>"000000000",
  43425=>"010110110",
  43426=>"000011111",
  43427=>"111111000",
  43428=>"000000000",
  43429=>"110111111",
  43430=>"111111111",
  43431=>"000000000",
  43432=>"011011111",
  43433=>"110111111",
  43434=>"000000011",
  43435=>"111111000",
  43436=>"000011011",
  43437=>"111011011",
  43438=>"000100000",
  43439=>"111001111",
  43440=>"101000111",
  43441=>"100111111",
  43442=>"110111111",
  43443=>"011111010",
  43444=>"000000001",
  43445=>"111000000",
  43446=>"110000001",
  43447=>"111100000",
  43448=>"110111100",
  43449=>"111111111",
  43450=>"000111101",
  43451=>"000011111",
  43452=>"001000000",
  43453=>"001001001",
  43454=>"111111111",
  43455=>"011011011",
  43456=>"111000110",
  43457=>"111000000",
  43458=>"000000000",
  43459=>"011111111",
  43460=>"111011111",
  43461=>"011001001",
  43462=>"000000100",
  43463=>"111111110",
  43464=>"111111111",
  43465=>"001111111",
  43466=>"000000001",
  43467=>"111111110",
  43468=>"111111111",
  43469=>"000001011",
  43470=>"110101101",
  43471=>"011000000",
  43472=>"000000100",
  43473=>"111111001",
  43474=>"000011111",
  43475=>"000001001",
  43476=>"001000000",
  43477=>"100000000",
  43478=>"111011001",
  43479=>"011001001",
  43480=>"000000000",
  43481=>"011000000",
  43482=>"010001011",
  43483=>"111011110",
  43484=>"101000010",
  43485=>"111111011",
  43486=>"101101111",
  43487=>"000010000",
  43488=>"011011000",
  43489=>"000000000",
  43490=>"000001000",
  43491=>"000000001",
  43492=>"101101111",
  43493=>"101111111",
  43494=>"100000000",
  43495=>"000000000",
  43496=>"111111111",
  43497=>"000000000",
  43498=>"010111111",
  43499=>"111111111",
  43500=>"001110110",
  43501=>"000010010",
  43502=>"000000001",
  43503=>"111000001",
  43504=>"111111111",
  43505=>"111111111",
  43506=>"000001111",
  43507=>"110110100",
  43508=>"111111111",
  43509=>"000000001",
  43510=>"100000000",
  43511=>"000010111",
  43512=>"000000000",
  43513=>"001001011",
  43514=>"110000000",
  43515=>"111111000",
  43516=>"000000000",
  43517=>"111111111",
  43518=>"000000000",
  43519=>"111111011",
  43520=>"011000000",
  43521=>"101000000",
  43522=>"000000000",
  43523=>"000000000",
  43524=>"101000010",
  43525=>"100000000",
  43526=>"000000111",
  43527=>"000000000",
  43528=>"000000101",
  43529=>"001001111",
  43530=>"111110000",
  43531=>"000000000",
  43532=>"110110010",
  43533=>"111001001",
  43534=>"111000001",
  43535=>"000000011",
  43536=>"000001111",
  43537=>"010111001",
  43538=>"000000101",
  43539=>"000001111",
  43540=>"111111111",
  43541=>"100000110",
  43542=>"111100100",
  43543=>"011011111",
  43544=>"100000000",
  43545=>"000010011",
  43546=>"000000011",
  43547=>"000000000",
  43548=>"001000000",
  43549=>"000000100",
  43550=>"110111110",
  43551=>"011011001",
  43552=>"000000000",
  43553=>"111111111",
  43554=>"011001001",
  43555=>"111111000",
  43556=>"000100111",
  43557=>"111111010",
  43558=>"111000000",
  43559=>"111111111",
  43560=>"111111111",
  43561=>"001000111",
  43562=>"111111111",
  43563=>"111000000",
  43564=>"000100111",
  43565=>"101111111",
  43566=>"000000110",
  43567=>"110110000",
  43568=>"000000111",
  43569=>"110111111",
  43570=>"011111000",
  43571=>"000000000",
  43572=>"111111100",
  43573=>"100010000",
  43574=>"111111111",
  43575=>"111110110",
  43576=>"000001011",
  43577=>"110000100",
  43578=>"100111111",
  43579=>"110110000",
  43580=>"000000000",
  43581=>"111000000",
  43582=>"000000000",
  43583=>"000000111",
  43584=>"000000000",
  43585=>"000000010",
  43586=>"000011111",
  43587=>"111111000",
  43588=>"000001001",
  43589=>"000111111",
  43590=>"000000101",
  43591=>"100000000",
  43592=>"111111111",
  43593=>"000000000",
  43594=>"111110000",
  43595=>"011100111",
  43596=>"000000001",
  43597=>"100000000",
  43598=>"101000000",
  43599=>"111000000",
  43600=>"111110111",
  43601=>"111100110",
  43602=>"010000010",
  43603=>"000000000",
  43604=>"000000000",
  43605=>"111111110",
  43606=>"111000110",
  43607=>"010010000",
  43608=>"000000000",
  43609=>"111100111",
  43610=>"111111111",
  43611=>"011011110",
  43612=>"011111111",
  43613=>"001000101",
  43614=>"000011111",
  43615=>"101111000",
  43616=>"000000000",
  43617=>"111111111",
  43618=>"111000000",
  43619=>"111111000",
  43620=>"001001111",
  43621=>"000000000",
  43622=>"110110110",
  43623=>"111001000",
  43624=>"000000000",
  43625=>"111101111",
  43626=>"110110111",
  43627=>"000111100",
  43628=>"001000110",
  43629=>"111111011",
  43630=>"011000000",
  43631=>"000001001",
  43632=>"111110111",
  43633=>"100011011",
  43634=>"001001111",
  43635=>"000001000",
  43636=>"000000000",
  43637=>"000000000",
  43638=>"001101000",
  43639=>"100111111",
  43640=>"001000000",
  43641=>"000110111",
  43642=>"000000000",
  43643=>"111001101",
  43644=>"110110100",
  43645=>"000110111",
  43646=>"100100000",
  43647=>"000000011",
  43648=>"111000001",
  43649=>"100100111",
  43650=>"110110111",
  43651=>"111111011",
  43652=>"001011001",
  43653=>"000100000",
  43654=>"101111010",
  43655=>"111000000",
  43656=>"111001001",
  43657=>"111111111",
  43658=>"111011000",
  43659=>"000100101",
  43660=>"000101101",
  43661=>"001000110",
  43662=>"111111111",
  43663=>"000000111",
  43664=>"000110111",
  43665=>"000111011",
  43666=>"111100101",
  43667=>"000110110",
  43668=>"000000001",
  43669=>"000001000",
  43670=>"101000100",
  43671=>"000000101",
  43672=>"000000111",
  43673=>"100100000",
  43674=>"000000000",
  43675=>"111001000",
  43676=>"001111100",
  43677=>"000000000",
  43678=>"111010111",
  43679=>"000000010",
  43680=>"100000000",
  43681=>"001001000",
  43682=>"111000000",
  43683=>"001001011",
  43684=>"101000100",
  43685=>"000000011",
  43686=>"000000000",
  43687=>"111111111",
  43688=>"100000000",
  43689=>"111000000",
  43690=>"110111111",
  43691=>"100001111",
  43692=>"010011011",
  43693=>"000001000",
  43694=>"000100111",
  43695=>"000000000",
  43696=>"111000111",
  43697=>"011111111",
  43698=>"110011111",
  43699=>"000000000",
  43700=>"000010000",
  43701=>"111100100",
  43702=>"111111111",
  43703=>"000000111",
  43704=>"111111101",
  43705=>"000110110",
  43706=>"000000000",
  43707=>"110100111",
  43708=>"000000000",
  43709=>"111111111",
  43710=>"011000100",
  43711=>"000000000",
  43712=>"011111111",
  43713=>"110000010",
  43714=>"111111111",
  43715=>"111111110",
  43716=>"111111111",
  43717=>"111111111",
  43718=>"000111111",
  43719=>"000000001",
  43720=>"001000011",
  43721=>"000000111",
  43722=>"000000100",
  43723=>"100101101",
  43724=>"000000000",
  43725=>"011110100",
  43726=>"110111111",
  43727=>"010110100",
  43728=>"100000000",
  43729=>"000000000",
  43730=>"000000000",
  43731=>"000110111",
  43732=>"000000000",
  43733=>"110000101",
  43734=>"111111111",
  43735=>"101101000",
  43736=>"001000000",
  43737=>"000000100",
  43738=>"111111110",
  43739=>"001000110",
  43740=>"101001001",
  43741=>"111001000",
  43742=>"111111111",
  43743=>"011000110",
  43744=>"111011000",
  43745=>"000111000",
  43746=>"011000000",
  43747=>"000111111",
  43748=>"000111111",
  43749=>"110110111",
  43750=>"000000100",
  43751=>"000100110",
  43752=>"111100100",
  43753=>"100000000",
  43754=>"000000001",
  43755=>"111000000",
  43756=>"111111000",
  43757=>"000110111",
  43758=>"011111111",
  43759=>"000000000",
  43760=>"100110110",
  43761=>"111111111",
  43762=>"000111001",
  43763=>"111001000",
  43764=>"010111111",
  43765=>"011011000",
  43766=>"000011000",
  43767=>"000000100",
  43768=>"000000000",
  43769=>"111111001",
  43770=>"111000000",
  43771=>"111101001",
  43772=>"100110111",
  43773=>"110011011",
  43774=>"111000101",
  43775=>"000000000",
  43776=>"110000111",
  43777=>"011011000",
  43778=>"000010000",
  43779=>"000000001",
  43780=>"100110001",
  43781=>"111000010",
  43782=>"111111100",
  43783=>"111000101",
  43784=>"000000000",
  43785=>"000000000",
  43786=>"000000000",
  43787=>"000000101",
  43788=>"111010000",
  43789=>"001000000",
  43790=>"000000001",
  43791=>"001000000",
  43792=>"111000000",
  43793=>"111111111",
  43794=>"000000111",
  43795=>"000000100",
  43796=>"000011111",
  43797=>"001000000",
  43798=>"000011001",
  43799=>"101000000",
  43800=>"011111111",
  43801=>"000000000",
  43802=>"110001111",
  43803=>"010010111",
  43804=>"111111111",
  43805=>"111111000",
  43806=>"000000100",
  43807=>"111011001",
  43808=>"111000101",
  43809=>"111111111",
  43810=>"111100111",
  43811=>"111111001",
  43812=>"111001111",
  43813=>"110000111",
  43814=>"000000111",
  43815=>"001000000",
  43816=>"000000001",
  43817=>"000000011",
  43818=>"111111111",
  43819=>"100000000",
  43820=>"111111111",
  43821=>"011011111",
  43822=>"000011000",
  43823=>"110111110",
  43824=>"111111111",
  43825=>"111011111",
  43826=>"000000000",
  43827=>"000110111",
  43828=>"100000000",
  43829=>"110111000",
  43830=>"000000001",
  43831=>"000000000",
  43832=>"110000000",
  43833=>"000000100",
  43834=>"110100100",
  43835=>"111111011",
  43836=>"011000110",
  43837=>"000000000",
  43838=>"000000000",
  43839=>"000000010",
  43840=>"111000000",
  43841=>"111111001",
  43842=>"110110110",
  43843=>"000000000",
  43844=>"000001111",
  43845=>"111111000",
  43846=>"000000110",
  43847=>"111111110",
  43848=>"111011000",
  43849=>"010000000",
  43850=>"111101001",
  43851=>"011111011",
  43852=>"000000100",
  43853=>"000010000",
  43854=>"000000111",
  43855=>"000000011",
  43856=>"100100100",
  43857=>"001000100",
  43858=>"111011001",
  43859=>"111100100",
  43860=>"000110000",
  43861=>"001001001",
  43862=>"111111111",
  43863=>"111111111",
  43864=>"111111010",
  43865=>"000000010",
  43866=>"111110110",
  43867=>"111111111",
  43868=>"100000111",
  43869=>"000000111",
  43870=>"000000000",
  43871=>"011011011",
  43872=>"000000000",
  43873=>"001101111",
  43874=>"101111011",
  43875=>"111111011",
  43876=>"100000000",
  43877=>"000000111",
  43878=>"101101100",
  43879=>"000100100",
  43880=>"110110110",
  43881=>"111110000",
  43882=>"000000000",
  43883=>"110111000",
  43884=>"000110111",
  43885=>"111111111",
  43886=>"000111010",
  43887=>"111011000",
  43888=>"111111000",
  43889=>"110111111",
  43890=>"000010010",
  43891=>"111111011",
  43892=>"010110111",
  43893=>"100110110",
  43894=>"001001001",
  43895=>"111010000",
  43896=>"111111111",
  43897=>"101001000",
  43898=>"110110111",
  43899=>"111000000",
  43900=>"000000001",
  43901=>"000000000",
  43902=>"111000000",
  43903=>"010000000",
  43904=>"110000000",
  43905=>"000001111",
  43906=>"000111111",
  43907=>"101000000",
  43908=>"000000000",
  43909=>"000001000",
  43910=>"000111111",
  43911=>"001001100",
  43912=>"110111111",
  43913=>"111111011",
  43914=>"111111000",
  43915=>"101000100",
  43916=>"001001001",
  43917=>"001000110",
  43918=>"000110111",
  43919=>"010011000",
  43920=>"000000010",
  43921=>"101001000",
  43922=>"111111111",
  43923=>"000001001",
  43924=>"111101101",
  43925=>"000111111",
  43926=>"110111000",
  43927=>"000000000",
  43928=>"101001001",
  43929=>"110110010",
  43930=>"001101111",
  43931=>"111111110",
  43932=>"111101000",
  43933=>"000111110",
  43934=>"011110111",
  43935=>"000111111",
  43936=>"000000000",
  43937=>"010001111",
  43938=>"110000111",
  43939=>"111000100",
  43940=>"111001111",
  43941=>"111111111",
  43942=>"000101111",
  43943=>"111011111",
  43944=>"000000000",
  43945=>"001000001",
  43946=>"110011001",
  43947=>"111000000",
  43948=>"000000110",
  43949=>"111111111",
  43950=>"110000111",
  43951=>"011000111",
  43952=>"000000000",
  43953=>"000111011",
  43954=>"011001000",
  43955=>"100000000",
  43956=>"111100100",
  43957=>"111001001",
  43958=>"000110111",
  43959=>"110100011",
  43960=>"000000111",
  43961=>"100100101",
  43962=>"000000000",
  43963=>"000100111",
  43964=>"111111011",
  43965=>"111111110",
  43966=>"100000000",
  43967=>"111111011",
  43968=>"001001111",
  43969=>"111000000",
  43970=>"000000000",
  43971=>"000000100",
  43972=>"111001111",
  43973=>"110000000",
  43974=>"000000111",
  43975=>"111101000",
  43976=>"110000000",
  43977=>"011111011",
  43978=>"111110111",
  43979=>"111000000",
  43980=>"000000000",
  43981=>"000000000",
  43982=>"111000000",
  43983=>"010000000",
  43984=>"101111111",
  43985=>"111111011",
  43986=>"001000000",
  43987=>"000000000",
  43988=>"000001111",
  43989=>"100111111",
  43990=>"001000000",
  43991=>"111111001",
  43992=>"111000001",
  43993=>"101001000",
  43994=>"000000000",
  43995=>"011111111",
  43996=>"000011011",
  43997=>"000000000",
  43998=>"000000000",
  43999=>"000000111",
  44000=>"111111111",
  44001=>"111111001",
  44002=>"011000000",
  44003=>"000000100",
  44004=>"111000000",
  44005=>"000000000",
  44006=>"111101111",
  44007=>"111000000",
  44008=>"111001101",
  44009=>"000000000",
  44010=>"000010111",
  44011=>"000000000",
  44012=>"000001001",
  44013=>"000000001",
  44014=>"001001111",
  44015=>"111001111",
  44016=>"111111000",
  44017=>"111001111",
  44018=>"000000001",
  44019=>"111110110",
  44020=>"000000011",
  44021=>"111111111",
  44022=>"110111000",
  44023=>"000111111",
  44024=>"110111100",
  44025=>"011010110",
  44026=>"010011011",
  44027=>"000000011",
  44028=>"000001011",
  44029=>"111111111",
  44030=>"000000000",
  44031=>"000000110",
  44032=>"000000000",
  44033=>"101000010",
  44034=>"111000010",
  44035=>"111111110",
  44036=>"000000000",
  44037=>"111110110",
  44038=>"100111111",
  44039=>"111111111",
  44040=>"001000010",
  44041=>"111000000",
  44042=>"111111111",
  44043=>"110001001",
  44044=>"111111111",
  44045=>"111000011",
  44046=>"000000000",
  44047=>"000000000",
  44048=>"001001000",
  44049=>"111001001",
  44050=>"000001000",
  44051=>"111111111",
  44052=>"000000000",
  44053=>"110111100",
  44054=>"111111111",
  44055=>"111111111",
  44056=>"111001001",
  44057=>"100000000",
  44058=>"000000000",
  44059=>"111111111",
  44060=>"111111111",
  44061=>"111011111",
  44062=>"111101101",
  44063=>"001000000",
  44064=>"110111111",
  44065=>"110110000",
  44066=>"000000001",
  44067=>"111111110",
  44068=>"100100000",
  44069=>"000001111",
  44070=>"111111111",
  44071=>"000111111",
  44072=>"000000000",
  44073=>"110110000",
  44074=>"001101111",
  44075=>"000000000",
  44076=>"000000000",
  44077=>"100000000",
  44078=>"000001000",
  44079=>"000000000",
  44080=>"011010111",
  44081=>"010011111",
  44082=>"111111101",
  44083=>"000111111",
  44084=>"111111001",
  44085=>"011001001",
  44086=>"000100000",
  44087=>"111111100",
  44088=>"000001011",
  44089=>"111001000",
  44090=>"000001000",
  44091=>"001001011",
  44092=>"111111111",
  44093=>"000000000",
  44094=>"111000000",
  44095=>"000000000",
  44096=>"100000000",
  44097=>"111111111",
  44098=>"111111000",
  44099=>"111111111",
  44100=>"111111111",
  44101=>"110111111",
  44102=>"000000000",
  44103=>"111111111",
  44104=>"011011000",
  44105=>"000000000",
  44106=>"111111011",
  44107=>"111111111",
  44108=>"100110111",
  44109=>"000100000",
  44110=>"110000010",
  44111=>"111111111",
  44112=>"000000011",
  44113=>"110000000",
  44114=>"011000000",
  44115=>"111111111",
  44116=>"000100000",
  44117=>"010011011",
  44118=>"001001000",
  44119=>"111111111",
  44120=>"000000000",
  44121=>"111110111",
  44122=>"111111111",
  44123=>"011001001",
  44124=>"111111111",
  44125=>"000000001",
  44126=>"000000000",
  44127=>"111111110",
  44128=>"111111111",
  44129=>"111111110",
  44130=>"010000000",
  44131=>"111111111",
  44132=>"000000100",
  44133=>"011000000",
  44134=>"111000000",
  44135=>"001000000",
  44136=>"000000100",
  44137=>"100100111",
  44138=>"001111111",
  44139=>"001001000",
  44140=>"011111111",
  44141=>"111111000",
  44142=>"000001111",
  44143=>"111111000",
  44144=>"111111010",
  44145=>"001001001",
  44146=>"010111111",
  44147=>"100000000",
  44148=>"000000000",
  44149=>"111111111",
  44150=>"001001000",
  44151=>"111111111",
  44152=>"111100110",
  44153=>"110110111",
  44154=>"111111001",
  44155=>"111111111",
  44156=>"000000000",
  44157=>"111001000",
  44158=>"000000000",
  44159=>"100000000",
  44160=>"000111111",
  44161=>"011011001",
  44162=>"000000000",
  44163=>"001011100",
  44164=>"111111101",
  44165=>"111111000",
  44166=>"110111111",
  44167=>"111101000",
  44168=>"111011000",
  44169=>"010111111",
  44170=>"111111111",
  44171=>"000100110",
  44172=>"001011111",
  44173=>"000001111",
  44174=>"110111111",
  44175=>"000001000",
  44176=>"111111111",
  44177=>"000000100",
  44178=>"111101011",
  44179=>"010010110",
  44180=>"110110000",
  44181=>"110100100",
  44182=>"000000001",
  44183=>"000100110",
  44184=>"111000110",
  44185=>"000000000",
  44186=>"000000000",
  44187=>"111111111",
  44188=>"100000000",
  44189=>"111110111",
  44190=>"111111001",
  44191=>"100100000",
  44192=>"000000001",
  44193=>"111111111",
  44194=>"001111111",
  44195=>"111001001",
  44196=>"111111011",
  44197=>"111111111",
  44198=>"111111111",
  44199=>"001000101",
  44200=>"110111000",
  44201=>"000000000",
  44202=>"001001000",
  44203=>"111101001",
  44204=>"111011111",
  44205=>"001011111",
  44206=>"101001000",
  44207=>"000000000",
  44208=>"000000111",
  44209=>"000001111",
  44210=>"111110111",
  44211=>"111100100",
  44212=>"011000110",
  44213=>"001011011",
  44214=>"000000000",
  44215=>"000000000",
  44216=>"100100111",
  44217=>"000000101",
  44218=>"000110110",
  44219=>"000000110",
  44220=>"000010010",
  44221=>"111111111",
  44222=>"000000000",
  44223=>"111111001",
  44224=>"000000000",
  44225=>"000100000",
  44226=>"111011001",
  44227=>"000000000",
  44228=>"110000000",
  44229=>"111111000",
  44230=>"111110000",
  44231=>"000000000",
  44232=>"001000000",
  44233=>"001111011",
  44234=>"000000000",
  44235=>"000000000",
  44236=>"000000000",
  44237=>"111111111",
  44238=>"001011111",
  44239=>"111111111",
  44240=>"111110000",
  44241=>"101100100",
  44242=>"111000000",
  44243=>"010010000",
  44244=>"100100111",
  44245=>"111011111",
  44246=>"000000000",
  44247=>"111111000",
  44248=>"011011111",
  44249=>"000000000",
  44250=>"000000001",
  44251=>"000011111",
  44252=>"000111111",
  44253=>"100101111",
  44254=>"111111110",
  44255=>"110100110",
  44256=>"100000000",
  44257=>"010000011",
  44258=>"111111110",
  44259=>"000010001",
  44260=>"010010000",
  44261=>"100111111",
  44262=>"100111111",
  44263=>"111111001",
  44264=>"000011111",
  44265=>"111111111",
  44266=>"000010111",
  44267=>"000001111",
  44268=>"111100000",
  44269=>"011011111",
  44270=>"111111111",
  44271=>"111101100",
  44272=>"000000100",
  44273=>"111111111",
  44274=>"000000000",
  44275=>"000000111",
  44276=>"000111101",
  44277=>"011001011",
  44278=>"001001001",
  44279=>"100000100",
  44280=>"111111011",
  44281=>"000000000",
  44282=>"000000000",
  44283=>"001001100",
  44284=>"100110000",
  44285=>"001001100",
  44286=>"111111111",
  44287=>"000001000",
  44288=>"101111000",
  44289=>"111110100",
  44290=>"111110110",
  44291=>"011111110",
  44292=>"000000001",
  44293=>"100000000",
  44294=>"111111000",
  44295=>"000111111",
  44296=>"000000000",
  44297=>"111111111",
  44298=>"000001011",
  44299=>"111111110",
  44300=>"111111111",
  44301=>"000000000",
  44302=>"000000000",
  44303=>"000000000",
  44304=>"000000000",
  44305=>"000000000",
  44306=>"000000000",
  44307=>"011001001",
  44308=>"000000000",
  44309=>"111111111",
  44310=>"000001010",
  44311=>"111110110",
  44312=>"111001000",
  44313=>"111110110",
  44314=>"000000000",
  44315=>"110000000",
  44316=>"111111111",
  44317=>"111001100",
  44318=>"111111110",
  44319=>"110110000",
  44320=>"110111111",
  44321=>"000111011",
  44322=>"000000000",
  44323=>"000000000",
  44324=>"000000010",
  44325=>"111111111",
  44326=>"110110110",
  44327=>"000010000",
  44328=>"011000110",
  44329=>"000000000",
  44330=>"111111111",
  44331=>"111110000",
  44332=>"000110110",
  44333=>"100100110",
  44334=>"111001111",
  44335=>"101111001",
  44336=>"100000000",
  44337=>"111111011",
  44338=>"000010111",
  44339=>"011011010",
  44340=>"110111111",
  44341=>"000000000",
  44342=>"110000000",
  44343=>"000000000",
  44344=>"000000000",
  44345=>"000111111",
  44346=>"000000000",
  44347=>"001000000",
  44348=>"000111000",
  44349=>"000010111",
  44350=>"111000010",
  44351=>"111111111",
  44352=>"111111111",
  44353=>"111010010",
  44354=>"111111111",
  44355=>"101111111",
  44356=>"000000000",
  44357=>"111111111",
  44358=>"111111110",
  44359=>"111001111",
  44360=>"000000000",
  44361=>"000000001",
  44362=>"110111110",
  44363=>"111111111",
  44364=>"000000100",
  44365=>"000100000",
  44366=>"011111111",
  44367=>"000000000",
  44368=>"111111001",
  44369=>"000000000",
  44370=>"000000000",
  44371=>"000100100",
  44372=>"111111111",
  44373=>"000100000",
  44374=>"000000010",
  44375=>"000000000",
  44376=>"000000000",
  44377=>"000000111",
  44378=>"010010111",
  44379=>"001101000",
  44380=>"100000100",
  44381=>"000000111",
  44382=>"111110111",
  44383=>"111111011",
  44384=>"111101111",
  44385=>"000000000",
  44386=>"111111111",
  44387=>"000000100",
  44388=>"000000000",
  44389=>"111111000",
  44390=>"000001111",
  44391=>"001001111",
  44392=>"100110011",
  44393=>"000000000",
  44394=>"100101101",
  44395=>"000000000",
  44396=>"001000100",
  44397=>"000000000",
  44398=>"010000000",
  44399=>"000000010",
  44400=>"111011111",
  44401=>"111111111",
  44402=>"000000100",
  44403=>"100110111",
  44404=>"000000000",
  44405=>"100100100",
  44406=>"111111011",
  44407=>"001000111",
  44408=>"111110110",
  44409=>"100100000",
  44410=>"111110011",
  44411=>"111111111",
  44412=>"000100111",
  44413=>"001000001",
  44414=>"100110100",
  44415=>"000000000",
  44416=>"000000000",
  44417=>"111111011",
  44418=>"100110110",
  44419=>"000000000",
  44420=>"000001101",
  44421=>"000000000",
  44422=>"111111111",
  44423=>"110010110",
  44424=>"111111111",
  44425=>"100100100",
  44426=>"111111100",
  44427=>"111111101",
  44428=>"000000000",
  44429=>"100100111",
  44430=>"000000000",
  44431=>"111111111",
  44432=>"110111111",
  44433=>"000000000",
  44434=>"000000010",
  44435=>"111000000",
  44436=>"000000111",
  44437=>"000010000",
  44438=>"000000010",
  44439=>"001001001",
  44440=>"011011011",
  44441=>"111011101",
  44442=>"011001111",
  44443=>"001111111",
  44444=>"000000000",
  44445=>"111011111",
  44446=>"000000000",
  44447=>"000000111",
  44448=>"011011000",
  44449=>"011011011",
  44450=>"000001001",
  44451=>"000111111",
  44452=>"001011000",
  44453=>"110110111",
  44454=>"000000111",
  44455=>"000000001",
  44456=>"000000000",
  44457=>"000111011",
  44458=>"111011001",
  44459=>"000000000",
  44460=>"000000000",
  44461=>"000111111",
  44462=>"011010010",
  44463=>"111111111",
  44464=>"010111111",
  44465=>"001111000",
  44466=>"111000111",
  44467=>"000000000",
  44468=>"100100111",
  44469=>"000100101",
  44470=>"000000000",
  44471=>"000000000",
  44472=>"000000000",
  44473=>"111100111",
  44474=>"011000000",
  44475=>"000000000",
  44476=>"111101000",
  44477=>"111000000",
  44478=>"100000100",
  44479=>"111011011",
  44480=>"111111111",
  44481=>"000000111",
  44482=>"000000000",
  44483=>"111111100",
  44484=>"000001001",
  44485=>"111111111",
  44486=>"000100100",
  44487=>"000000000",
  44488=>"000001101",
  44489=>"000110110",
  44490=>"000000000",
  44491=>"000000111",
  44492=>"111110110",
  44493=>"000000111",
  44494=>"000000000",
  44495=>"100000111",
  44496=>"001001001",
  44497=>"111111111",
  44498=>"000000111",
  44499=>"000000000",
  44500=>"110110100",
  44501=>"011001000",
  44502=>"110110000",
  44503=>"110000000",
  44504=>"001111100",
  44505=>"100100000",
  44506=>"000000000",
  44507=>"000111111",
  44508=>"110000000",
  44509=>"000000000",
  44510=>"111001111",
  44511=>"111111111",
  44512=>"111111111",
  44513=>"000000000",
  44514=>"111101111",
  44515=>"000000000",
  44516=>"000000000",
  44517=>"111111100",
  44518=>"111011000",
  44519=>"000010111",
  44520=>"000000000",
  44521=>"111111011",
  44522=>"111111000",
  44523=>"000000000",
  44524=>"000000000",
  44525=>"000000000",
  44526=>"101101111",
  44527=>"111110000",
  44528=>"000000100",
  44529=>"000000001",
  44530=>"100100000",
  44531=>"001001001",
  44532=>"000000000",
  44533=>"000000000",
  44534=>"110110110",
  44535=>"111111111",
  44536=>"111000000",
  44537=>"110100000",
  44538=>"111111111",
  44539=>"000111111",
  44540=>"000000000",
  44541=>"010011000",
  44542=>"000000000",
  44543=>"011011011",
  44544=>"100110000",
  44545=>"000000000",
  44546=>"001000000",
  44547=>"111000000",
  44548=>"001010011",
  44549=>"000001000",
  44550=>"000000001",
  44551=>"111111000",
  44552=>"000000000",
  44553=>"110111100",
  44554=>"011111011",
  44555=>"111111101",
  44556=>"000000000",
  44557=>"001111111",
  44558=>"010000000",
  44559=>"111111111",
  44560=>"011000000",
  44561=>"111110011",
  44562=>"001001111",
  44563=>"000100000",
  44564=>"101111101",
  44565=>"111111000",
  44566=>"011111111",
  44567=>"001000100",
  44568=>"111000000",
  44569=>"001001000",
  44570=>"000001111",
  44571=>"100101110",
  44572=>"000000011",
  44573=>"001001100",
  44574=>"000001011",
  44575=>"111000111",
  44576=>"001111111",
  44577=>"111010000",
  44578=>"100000001",
  44579=>"111111000",
  44580=>"111000000",
  44581=>"000000000",
  44582=>"111111111",
  44583=>"111000010",
  44584=>"010001001",
  44585=>"000100100",
  44586=>"011001001",
  44587=>"000110010",
  44588=>"000000000",
  44589=>"000000100",
  44590=>"000111000",
  44591=>"011001000",
  44592=>"000000111",
  44593=>"000000111",
  44594=>"110110000",
  44595=>"111101111",
  44596=>"010000111",
  44597=>"110000000",
  44598=>"001000000",
  44599=>"000111000",
  44600=>"001011111",
  44601=>"111111111",
  44602=>"000011011",
  44603=>"000000000",
  44604=>"000000111",
  44605=>"111011001",
  44606=>"011111111",
  44607=>"000110000",
  44608=>"111110110",
  44609=>"011000100",
  44610=>"110110000",
  44611=>"100110111",
  44612=>"000000000",
  44613=>"111100111",
  44614=>"111111010",
  44615=>"110110111",
  44616=>"111111011",
  44617=>"000111000",
  44618=>"111001001",
  44619=>"111000000",
  44620=>"000000000",
  44621=>"111101111",
  44622=>"010000000",
  44623=>"010011001",
  44624=>"101111011",
  44625=>"110111110",
  44626=>"111111111",
  44627=>"111111110",
  44628=>"111100101",
  44629=>"111110110",
  44630=>"000110110",
  44631=>"011010111",
  44632=>"111011001",
  44633=>"000000000",
  44634=>"000000001",
  44635=>"100000000",
  44636=>"111000000",
  44637=>"010111010",
  44638=>"001111000",
  44639=>"111000001",
  44640=>"000000000",
  44641=>"111111111",
  44642=>"000000000",
  44643=>"000000111",
  44644=>"100000100",
  44645=>"111111111",
  44646=>"000000000",
  44647=>"100100101",
  44648=>"001000001",
  44649=>"110111000",
  44650=>"000110000",
  44651=>"111110101",
  44652=>"100001000",
  44653=>"111111111",
  44654=>"000000000",
  44655=>"111111100",
  44656=>"000000000",
  44657=>"110000000",
  44658=>"010110010",
  44659=>"000000000",
  44660=>"001011011",
  44661=>"001001000",
  44662=>"010111010",
  44663=>"111111010",
  44664=>"000000100",
  44665=>"011011000",
  44666=>"111100110",
  44667=>"000000001",
  44668=>"000111111",
  44669=>"101000000",
  44670=>"111111111",
  44671=>"000000100",
  44672=>"111111111",
  44673=>"011110111",
  44674=>"000111111",
  44675=>"110110111",
  44676=>"000000000",
  44677=>"111111000",
  44678=>"110101111",
  44679=>"001001000",
  44680=>"000001011",
  44681=>"011011000",
  44682=>"011000000",
  44683=>"000010010",
  44684=>"000011001",
  44685=>"110111010",
  44686=>"000000010",
  44687=>"000000010",
  44688=>"110111000",
  44689=>"010110111",
  44690=>"011000000",
  44691=>"000011011",
  44692=>"110111101",
  44693=>"111111011",
  44694=>"001001001",
  44695=>"000001111",
  44696=>"000101100",
  44697=>"101111111",
  44698=>"101000111",
  44699=>"001000000",
  44700=>"111111111",
  44701=>"000000000",
  44702=>"100100000",
  44703=>"011011000",
  44704=>"100000111",
  44705=>"000010000",
  44706=>"000001111",
  44707=>"000000011",
  44708=>"001000000",
  44709=>"000000010",
  44710=>"000000000",
  44711=>"011011110",
  44712=>"000100001",
  44713=>"111111001",
  44714=>"000100000",
  44715=>"010000000",
  44716=>"111101000",
  44717=>"000000001",
  44718=>"110000000",
  44719=>"000000000",
  44720=>"000010000",
  44721=>"111111101",
  44722=>"111011011",
  44723=>"011000000",
  44724=>"010001100",
  44725=>"111111111",
  44726=>"111001111",
  44727=>"000000000",
  44728=>"111111111",
  44729=>"001000101",
  44730=>"011011001",
  44731=>"000000111",
  44732=>"111000111",
  44733=>"000000111",
  44734=>"111111111",
  44735=>"000000000",
  44736=>"000000100",
  44737=>"111111111",
  44738=>"000000011",
  44739=>"000000000",
  44740=>"110111000",
  44741=>"101000111",
  44742=>"111100101",
  44743=>"011111111",
  44744=>"000001001",
  44745=>"111110111",
  44746=>"110000001",
  44747=>"011001111",
  44748=>"110111000",
  44749=>"000000001",
  44750=>"000000111",
  44751=>"000000000",
  44752=>"011011011",
  44753=>"001110011",
  44754=>"011011001",
  44755=>"101000111",
  44756=>"000000000",
  44757=>"011011011",
  44758=>"011001111",
  44759=>"000101001",
  44760=>"000000000",
  44761=>"000110111",
  44762=>"110111111",
  44763=>"000000000",
  44764=>"000001010",
  44765=>"011011011",
  44766=>"001001111",
  44767=>"000000000",
  44768=>"010111010",
  44769=>"111111111",
  44770=>"111011111",
  44771=>"000000000",
  44772=>"000000000",
  44773=>"000000001",
  44774=>"000000001",
  44775=>"101111001",
  44776=>"111000011",
  44777=>"111001101",
  44778=>"010100001",
  44779=>"100000100",
  44780=>"111111111",
  44781=>"111111111",
  44782=>"000000111",
  44783=>"111111011",
  44784=>"111111001",
  44785=>"000000000",
  44786=>"000000000",
  44787=>"110010110",
  44788=>"011000001",
  44789=>"111001110",
  44790=>"101101101",
  44791=>"100111111",
  44792=>"101000001",
  44793=>"000100000",
  44794=>"110111111",
  44795=>"000000001",
  44796=>"110101111",
  44797=>"100100110",
  44798=>"111000000",
  44799=>"000110110",
  44800=>"000000010",
  44801=>"111011111",
  44802=>"000000111",
  44803=>"011111111",
  44804=>"000111000",
  44805=>"000001001",
  44806=>"110111011",
  44807=>"111111000",
  44808=>"100111111",
  44809=>"111111100",
  44810=>"111001111",
  44811=>"111111111",
  44812=>"111111111",
  44813=>"111111110",
  44814=>"111111111",
  44815=>"000000111",
  44816=>"100000001",
  44817=>"011000000",
  44818=>"000000000",
  44819=>"000000001",
  44820=>"111001000",
  44821=>"000111111",
  44822=>"000011011",
  44823=>"000000000",
  44824=>"111110001",
  44825=>"111000111",
  44826=>"000000000",
  44827=>"000010000",
  44828=>"101111111",
  44829=>"111001000",
  44830=>"000010000",
  44831=>"000011011",
  44832=>"011001000",
  44833=>"000001000",
  44834=>"011000000",
  44835=>"111111111",
  44836=>"000000110",
  44837=>"110000110",
  44838=>"000111111",
  44839=>"110001001",
  44840=>"000000000",
  44841=>"000000000",
  44842=>"011011101",
  44843=>"000000000",
  44844=>"111100111",
  44845=>"011001000",
  44846=>"111000000",
  44847=>"001000000",
  44848=>"101100100",
  44849=>"101000000",
  44850=>"100011111",
  44851=>"000111000",
  44852=>"000000111",
  44853=>"000000000",
  44854=>"111111111",
  44855=>"011000000",
  44856=>"000000000",
  44857=>"111101000",
  44858=>"011010000",
  44859=>"111111011",
  44860=>"011000011",
  44861=>"001011001",
  44862=>"011111011",
  44863=>"111111110",
  44864=>"000001111",
  44865=>"111110000",
  44866=>"001011111",
  44867=>"110110110",
  44868=>"000110111",
  44869=>"100000100",
  44870=>"111100111",
  44871=>"001011000",
  44872=>"111000011",
  44873=>"111000000",
  44874=>"000000000",
  44875=>"100100101",
  44876=>"111111000",
  44877=>"111101000",
  44878=>"000110111",
  44879=>"001111001",
  44880=>"101001001",
  44881=>"110111000",
  44882=>"110100111",
  44883=>"000000111",
  44884=>"111110111",
  44885=>"111111111",
  44886=>"111011011",
  44887=>"000000000",
  44888=>"000000000",
  44889=>"000000000",
  44890=>"100000000",
  44891=>"110110000",
  44892=>"000000000",
  44893=>"000001000",
  44894=>"000000000",
  44895=>"001100000",
  44896=>"011010000",
  44897=>"111000000",
  44898=>"110110110",
  44899=>"101000101",
  44900=>"000000111",
  44901=>"000000000",
  44902=>"000000000",
  44903=>"000111011",
  44904=>"011001001",
  44905=>"111100101",
  44906=>"111111000",
  44907=>"001100100",
  44908=>"111111111",
  44909=>"011011011",
  44910=>"001000111",
  44911=>"000001000",
  44912=>"100110111",
  44913=>"000000000",
  44914=>"111111111",
  44915=>"111001001",
  44916=>"000000000",
  44917=>"000010000",
  44918=>"001000001",
  44919=>"111100110",
  44920=>"111000000",
  44921=>"111111111",
  44922=>"111000111",
  44923=>"110111111",
  44924=>"111111110",
  44925=>"000000000",
  44926=>"100000000",
  44927=>"001000001",
  44928=>"111111111",
  44929=>"100100111",
  44930=>"000111111",
  44931=>"000000000",
  44932=>"000000111",
  44933=>"000000000",
  44934=>"111100000",
  44935=>"000001001",
  44936=>"110000000",
  44937=>"011111111",
  44938=>"010111111",
  44939=>"000000000",
  44940=>"001001111",
  44941=>"010011111",
  44942=>"000000010",
  44943=>"100000000",
  44944=>"100000100",
  44945=>"010111000",
  44946=>"010111001",
  44947=>"001000001",
  44948=>"111111010",
  44949=>"000000110",
  44950=>"001101000",
  44951=>"100000011",
  44952=>"111111010",
  44953=>"000111001",
  44954=>"111000000",
  44955=>"111111111",
  44956=>"000100000",
  44957=>"010011001",
  44958=>"000100111",
  44959=>"111111111",
  44960=>"100100100",
  44961=>"010011000",
  44962=>"111110101",
  44963=>"000100001",
  44964=>"100110100",
  44965=>"110111010",
  44966=>"110111010",
  44967=>"000111111",
  44968=>"000000000",
  44969=>"000100110",
  44970=>"111001111",
  44971=>"000000000",
  44972=>"100100111",
  44973=>"000100000",
  44974=>"101111111",
  44975=>"000000000",
  44976=>"111111011",
  44977=>"000000000",
  44978=>"111011000",
  44979=>"001001001",
  44980=>"000011001",
  44981=>"011000000",
  44982=>"111111111",
  44983=>"111111110",
  44984=>"001001001",
  44985=>"001111111",
  44986=>"001111111",
  44987=>"111111011",
  44988=>"111111111",
  44989=>"111001000",
  44990=>"111001001",
  44991=>"010011011",
  44992=>"000000100",
  44993=>"000000011",
  44994=>"011011000",
  44995=>"111111000",
  44996=>"111111000",
  44997=>"101101001",
  44998=>"000000000",
  44999=>"111111111",
  45000=>"000000000",
  45001=>"111010011",
  45002=>"010111000",
  45003=>"110110100",
  45004=>"001100000",
  45005=>"001001000",
  45006=>"011111011",
  45007=>"111111000",
  45008=>"011111011",
  45009=>"111111111",
  45010=>"111111001",
  45011=>"000001111",
  45012=>"110110111",
  45013=>"011010000",
  45014=>"111111111",
  45015=>"011000010",
  45016=>"000000000",
  45017=>"100010110",
  45018=>"111111011",
  45019=>"001111000",
  45020=>"001000000",
  45021=>"001111011",
  45022=>"111110000",
  45023=>"001001011",
  45024=>"000000110",
  45025=>"000000000",
  45026=>"001000000",
  45027=>"000000000",
  45028=>"011111111",
  45029=>"011001011",
  45030=>"001000000",
  45031=>"000000111",
  45032=>"101101111",
  45033=>"001111111",
  45034=>"100100111",
  45035=>"001000000",
  45036=>"111111111",
  45037=>"001011111",
  45038=>"110110110",
  45039=>"000000000",
  45040=>"000000000",
  45041=>"111111001",
  45042=>"111011111",
  45043=>"000000001",
  45044=>"111001111",
  45045=>"001111000",
  45046=>"111111111",
  45047=>"011000001",
  45048=>"000000000",
  45049=>"001001001",
  45050=>"111011011",
  45051=>"000000000",
  45052=>"010011000",
  45053=>"000000101",
  45054=>"000000000",
  45055=>"000000111",
  45056=>"110111110",
  45057=>"010010010",
  45058=>"111000000",
  45059=>"111111111",
  45060=>"001011111",
  45061=>"111111000",
  45062=>"000000000",
  45063=>"000001101",
  45064=>"011011001",
  45065=>"100000000",
  45066=>"000001001",
  45067=>"111001000",
  45068=>"001101001",
  45069=>"101001001",
  45070=>"101100001",
  45071=>"100000000",
  45072=>"111101111",
  45073=>"000010111",
  45074=>"000011110",
  45075=>"111000100",
  45076=>"000000000",
  45077=>"111111111",
  45078=>"000000000",
  45079=>"011111111",
  45080=>"000001001",
  45081=>"101100000",
  45082=>"001010111",
  45083=>"000111000",
  45084=>"000001111",
  45085=>"000000000",
  45086=>"100110110",
  45087=>"000000000",
  45088=>"010010000",
  45089=>"111100000",
  45090=>"111110010",
  45091=>"110011001",
  45092=>"110000000",
  45093=>"000100111",
  45094=>"111111111",
  45095=>"001101111",
  45096=>"000000000",
  45097=>"010010010",
  45098=>"001000000",
  45099=>"000000000",
  45100=>"100100100",
  45101=>"011001001",
  45102=>"001000000",
  45103=>"111111111",
  45104=>"111111111",
  45105=>"001001101",
  45106=>"011001001",
  45107=>"000010000",
  45108=>"001001101",
  45109=>"000000000",
  45110=>"001010000",
  45111=>"000010110",
  45112=>"000110111",
  45113=>"111111101",
  45114=>"111001000",
  45115=>"001000111",
  45116=>"101101101",
  45117=>"101101111",
  45118=>"111111111",
  45119=>"001001111",
  45120=>"011011000",
  45121=>"110010000",
  45122=>"101001000",
  45123=>"111111111",
  45124=>"000100100",
  45125=>"010000100",
  45126=>"010000000",
  45127=>"111111111",
  45128=>"000000000",
  45129=>"111111111",
  45130=>"111111110",
  45131=>"001000000",
  45132=>"110110000",
  45133=>"111111111",
  45134=>"000100100",
  45135=>"101000101",
  45136=>"000000000",
  45137=>"101111111",
  45138=>"000000000",
  45139=>"000100100",
  45140=>"001000101",
  45141=>"000000010",
  45142=>"000111111",
  45143=>"101101111",
  45144=>"000110100",
  45145=>"000000000",
  45146=>"010111010",
  45147=>"111110100",
  45148=>"010011010",
  45149=>"111111111",
  45150=>"000001111",
  45151=>"111100000",
  45152=>"010110010",
  45153=>"000000000",
  45154=>"000000111",
  45155=>"001101000",
  45156=>"010000000",
  45157=>"111000101",
  45158=>"111111111",
  45159=>"000111111",
  45160=>"101111111",
  45161=>"011001100",
  45162=>"010010010",
  45163=>"100000100",
  45164=>"010110110",
  45165=>"100001111",
  45166=>"110111111",
  45167=>"110110110",
  45168=>"111011010",
  45169=>"000010111",
  45170=>"100100101",
  45171=>"100100101",
  45172=>"111000000",
  45173=>"000000000",
  45174=>"000000000",
  45175=>"101101101",
  45176=>"111000000",
  45177=>"101101111",
  45178=>"000000000",
  45179=>"000000000",
  45180=>"100110110",
  45181=>"111110010",
  45182=>"001001001",
  45183=>"000000000",
  45184=>"101001000",
  45185=>"001000111",
  45186=>"111000011",
  45187=>"000000010",
  45188=>"101101001",
  45189=>"111100101",
  45190=>"110110110",
  45191=>"000100100",
  45192=>"001001001",
  45193=>"000000000",
  45194=>"001001000",
  45195=>"010010110",
  45196=>"001001101",
  45197=>"111110011",
  45198=>"010000101",
  45199=>"011001111",
  45200=>"000000000",
  45201=>"000100111",
  45202=>"000000000",
  45203=>"111111111",
  45204=>"110110010",
  45205=>"111111001",
  45206=>"111011111",
  45207=>"101000000",
  45208=>"001001111",
  45209=>"000000100",
  45210=>"001001111",
  45211=>"000000000",
  45212=>"111111010",
  45213=>"000000110",
  45214=>"101101111",
  45215=>"110100000",
  45216=>"010010010",
  45217=>"001111111",
  45218=>"000010110",
  45219=>"111111111",
  45220=>"001001001",
  45221=>"111000000",
  45222=>"110111111",
  45223=>"000111111",
  45224=>"111101111",
  45225=>"000000101",
  45226=>"000010000",
  45227=>"000000110",
  45228=>"000000001",
  45229=>"110110110",
  45230=>"110111110",
  45231=>"011010011",
  45232=>"000010000",
  45233=>"000100000",
  45234=>"111111111",
  45235=>"000000101",
  45236=>"111111000",
  45237=>"000000001",
  45238=>"100101111",
  45239=>"010011010",
  45240=>"001101100",
  45241=>"001001001",
  45242=>"001100001",
  45243=>"110110111",
  45244=>"111101111",
  45245=>"000000000",
  45246=>"000000000",
  45247=>"111010011",
  45248=>"011011010",
  45249=>"000010010",
  45250=>"011001000",
  45251=>"010010000",
  45252=>"000000111",
  45253=>"111111111",
  45254=>"110000000",
  45255=>"110111010",
  45256=>"010010010",
  45257=>"000000000",
  45258=>"000000100",
  45259=>"000000011",
  45260=>"111111000",
  45261=>"110111111",
  45262=>"101000110",
  45263=>"101100111",
  45264=>"101100100",
  45265=>"110110110",
  45266=>"000010110",
  45267=>"000000001",
  45268=>"000000000",
  45269=>"000000000",
  45270=>"001001111",
  45271=>"000000001",
  45272=>"111111000",
  45273=>"001101111",
  45274=>"000000000",
  45275=>"010010010",
  45276=>"111111111",
  45277=>"011001111",
  45278=>"111111111",
  45279=>"000001001",
  45280=>"001001001",
  45281=>"000101000",
  45282=>"110000000",
  45283=>"010000000",
  45284=>"000000000",
  45285=>"111111111",
  45286=>"110111111",
  45287=>"000000111",
  45288=>"111011010",
  45289=>"001000000",
  45290=>"000000000",
  45291=>"101101111",
  45292=>"000000001",
  45293=>"000000110",
  45294=>"110111111",
  45295=>"000000000",
  45296=>"000010000",
  45297=>"111111111",
  45298=>"111111111",
  45299=>"001001001",
  45300=>"000000000",
  45301=>"111111010",
  45302=>"011011011",
  45303=>"101101111",
  45304=>"111000000",
  45305=>"010110111",
  45306=>"111000000",
  45307=>"000110000",
  45308=>"000101001",
  45309=>"011001011",
  45310=>"010010010",
  45311=>"001001101",
  45312=>"111111100",
  45313=>"001001000",
  45314=>"001000100",
  45315=>"000000000",
  45316=>"001000000",
  45317=>"000001000",
  45318=>"101101101",
  45319=>"000111110",
  45320=>"001101101",
  45321=>"101001101",
  45322=>"101000001",
  45323=>"101101111",
  45324=>"000010000",
  45325=>"101111111",
  45326=>"000001111",
  45327=>"101111111",
  45328=>"000000000",
  45329=>"000000000",
  45330=>"101001101",
  45331=>"110010000",
  45332=>"110000000",
  45333=>"100000000",
  45334=>"001100000",
  45335=>"000000000",
  45336=>"000001000",
  45337=>"001001000",
  45338=>"100111111",
  45339=>"010010011",
  45340=>"000011111",
  45341=>"000000100",
  45342=>"111110000",
  45343=>"001000011",
  45344=>"001011011",
  45345=>"000000011",
  45346=>"000110011",
  45347=>"011011111",
  45348=>"000010010",
  45349=>"111111111",
  45350=>"111111101",
  45351=>"001000100",
  45352=>"101000000",
  45353=>"000000000",
  45354=>"111110111",
  45355=>"101101101",
  45356=>"011000101",
  45357=>"110010111",
  45358=>"010000111",
  45359=>"101000100",
  45360=>"110110110",
  45361=>"011001111",
  45362=>"111011000",
  45363=>"000110111",
  45364=>"010010000",
  45365=>"010010010",
  45366=>"011001011",
  45367=>"101111111",
  45368=>"011111111",
  45369=>"111001000",
  45370=>"000000101",
  45371=>"111111000",
  45372=>"111111111",
  45373=>"111100000",
  45374=>"000000100",
  45375=>"111110010",
  45376=>"000000000",
  45377=>"111111111",
  45378=>"011011001",
  45379=>"001000001",
  45380=>"101001001",
  45381=>"100001001",
  45382=>"000000000",
  45383=>"111000000",
  45384=>"100101111",
  45385=>"000010110",
  45386=>"000100000",
  45387=>"011011011",
  45388=>"000000000",
  45389=>"010000000",
  45390=>"000000000",
  45391=>"000001001",
  45392=>"011011011",
  45393=>"110000000",
  45394=>"111111111",
  45395=>"110110010",
  45396=>"000000000",
  45397=>"001011001",
  45398=>"000001101",
  45399=>"100110100",
  45400=>"101101111",
  45401=>"111111111",
  45402=>"110000000",
  45403=>"000000101",
  45404=>"001001011",
  45405=>"000000000",
  45406=>"000000000",
  45407=>"000000110",
  45408=>"001001000",
  45409=>"000000000",
  45410=>"011011011",
  45411=>"101001001",
  45412=>"000010000",
  45413=>"000000000",
  45414=>"111111110",
  45415=>"100010111",
  45416=>"000110110",
  45417=>"000000000",
  45418=>"111111110",
  45419=>"111011001",
  45420=>"110110000",
  45421=>"000000001",
  45422=>"000000000",
  45423=>"000000000",
  45424=>"000000000",
  45425=>"000000000",
  45426=>"010110110",
  45427=>"111101000",
  45428=>"111111111",
  45429=>"101001001",
  45430=>"011011111",
  45431=>"110100101",
  45432=>"111101101",
  45433=>"110111011",
  45434=>"110100000",
  45435=>"010110110",
  45436=>"111101101",
  45437=>"110110011",
  45438=>"111110010",
  45439=>"110000000",
  45440=>"110110000",
  45441=>"110110010",
  45442=>"011111011",
  45443=>"000000101",
  45444=>"111111111",
  45445=>"000000000",
  45446=>"100100000",
  45447=>"000000000",
  45448=>"001001001",
  45449=>"000000000",
  45450=>"100100111",
  45451=>"000110100",
  45452=>"000000111",
  45453=>"000110110",
  45454=>"000000100",
  45455=>"101101101",
  45456=>"010010000",
  45457=>"100100000",
  45458=>"000000110",
  45459=>"111111110",
  45460=>"010010111",
  45461=>"000010010",
  45462=>"000000001",
  45463=>"011000000",
  45464=>"000011011",
  45465=>"100110110",
  45466=>"101000000",
  45467=>"011011111",
  45468=>"111111111",
  45469=>"011010110",
  45470=>"001000000",
  45471=>"000000100",
  45472=>"000110111",
  45473=>"001001000",
  45474=>"011001000",
  45475=>"010000000",
  45476=>"111110100",
  45477=>"010111011",
  45478=>"000000000",
  45479=>"111111111",
  45480=>"000000000",
  45481=>"110000000",
  45482=>"010010011",
  45483=>"000000000",
  45484=>"111111101",
  45485=>"110111111",
  45486=>"110110111",
  45487=>"110111011",
  45488=>"011001101",
  45489=>"001000000",
  45490=>"000011011",
  45491=>"000000000",
  45492=>"111111011",
  45493=>"000000000",
  45494=>"111111111",
  45495=>"011101101",
  45496=>"000000111",
  45497=>"010010000",
  45498=>"001000110",
  45499=>"001001000",
  45500=>"001111111",
  45501=>"110100000",
  45502=>"000001000",
  45503=>"000000011",
  45504=>"000000000",
  45505=>"111000001",
  45506=>"001001001",
  45507=>"000000000",
  45508=>"000000000",
  45509=>"100100101",
  45510=>"010010010",
  45511=>"100101101",
  45512=>"000001000",
  45513=>"011010000",
  45514=>"101001101",
  45515=>"000000110",
  45516=>"000000000",
  45517=>"111110110",
  45518=>"110110110",
  45519=>"110000100",
  45520=>"111010010",
  45521=>"000000001",
  45522=>"110110010",
  45523=>"011011000",
  45524=>"011011011",
  45525=>"001011011",
  45526=>"000000101",
  45527=>"100100111",
  45528=>"111011111",
  45529=>"000000001",
  45530=>"000000010",
  45531=>"010110110",
  45532=>"000001011",
  45533=>"011111011",
  45534=>"111111111",
  45535=>"110110010",
  45536=>"000000000",
  45537=>"111000000",
  45538=>"000000000",
  45539=>"011011000",
  45540=>"000010010",
  45541=>"000000000",
  45542=>"111001011",
  45543=>"000000000",
  45544=>"110110110",
  45545=>"111011000",
  45546=>"000011011",
  45547=>"001001000",
  45548=>"011010011",
  45549=>"111011000",
  45550=>"111010000",
  45551=>"101001111",
  45552=>"000000101",
  45553=>"111110111",
  45554=>"111111100",
  45555=>"111111111",
  45556=>"111010000",
  45557=>"000010010",
  45558=>"000000000",
  45559=>"110100000",
  45560=>"111111111",
  45561=>"000000000",
  45562=>"011011111",
  45563=>"101000000",
  45564=>"001111111",
  45565=>"111111111",
  45566=>"010010010",
  45567=>"111111111",
  45568=>"000000000",
  45569=>"100000000",
  45570=>"101100101",
  45571=>"110111110",
  45572=>"000000000",
  45573=>"111000101",
  45574=>"011011000",
  45575=>"111111111",
  45576=>"000000011",
  45577=>"000110111",
  45578=>"111001000",
  45579=>"111100000",
  45580=>"101101001",
  45581=>"111111111",
  45582=>"011011001",
  45583=>"000000001",
  45584=>"111001001",
  45585=>"111111111",
  45586=>"000000000",
  45587=>"111111111",
  45588=>"000000000",
  45589=>"111111111",
  45590=>"000000101",
  45591=>"111111110",
  45592=>"000000111",
  45593=>"100100101",
  45594=>"000100111",
  45595=>"100100110",
  45596=>"000001011",
  45597=>"111111111",
  45598=>"011111011",
  45599=>"011111011",
  45600=>"010000000",
  45601=>"000111111",
  45602=>"001001001",
  45603=>"111001001",
  45604=>"000000111",
  45605=>"110111000",
  45606=>"111111111",
  45607=>"000110110",
  45608=>"000000000",
  45609=>"111111111",
  45610=>"000000101",
  45611=>"111111111",
  45612=>"111111101",
  45613=>"100000000",
  45614=>"000000111",
  45615=>"111111111",
  45616=>"000000100",
  45617=>"000000001",
  45618=>"011000000",
  45619=>"000000000",
  45620=>"000000001",
  45621=>"100100111",
  45622=>"111111100",
  45623=>"111111110",
  45624=>"011000000",
  45625=>"010111111",
  45626=>"000110111",
  45627=>"001011011",
  45628=>"101001111",
  45629=>"000000001",
  45630=>"011111100",
  45631=>"100000100",
  45632=>"111111111",
  45633=>"011011010",
  45634=>"111111111",
  45635=>"000000000",
  45636=>"111011001",
  45637=>"000100100",
  45638=>"100111011",
  45639=>"111111111",
  45640=>"000000000",
  45641=>"111100111",
  45642=>"111111111",
  45643=>"000000011",
  45644=>"000000101",
  45645=>"110110111",
  45646=>"000000110",
  45647=>"110111010",
  45648=>"110110111",
  45649=>"111001000",
  45650=>"111111111",
  45651=>"000000001",
  45652=>"000000000",
  45653=>"111111111",
  45654=>"100000000",
  45655=>"111111111",
  45656=>"100100100",
  45657=>"000000000",
  45658=>"000000000",
  45659=>"000100010",
  45660=>"000001001",
  45661=>"000000000",
  45662=>"000000000",
  45663=>"000000000",
  45664=>"000000111",
  45665=>"111111000",
  45666=>"111111001",
  45667=>"000000000",
  45668=>"000001111",
  45669=>"000000111",
  45670=>"000111000",
  45671=>"111010000",
  45672=>"000000000",
  45673=>"111001001",
  45674=>"111011011",
  45675=>"111001000",
  45676=>"000100100",
  45677=>"111111111",
  45678=>"000000010",
  45679=>"110111111",
  45680=>"000110110",
  45681=>"000000000",
  45682=>"010011000",
  45683=>"111110110",
  45684=>"000110000",
  45685=>"000000000",
  45686=>"011000010",
  45687=>"111001111",
  45688=>"000000000",
  45689=>"001000000",
  45690=>"001111111",
  45691=>"100000111",
  45692=>"110110110",
  45693=>"110100110",
  45694=>"111111000",
  45695=>"100111111",
  45696=>"101111111",
  45697=>"111111000",
  45698=>"111110010",
  45699=>"000000100",
  45700=>"010000111",
  45701=>"011000000",
  45702=>"110110000",
  45703=>"000010000",
  45704=>"110111110",
  45705=>"111111011",
  45706=>"010111111",
  45707=>"111111110",
  45708=>"000000000",
  45709=>"000000000",
  45710=>"111111111",
  45711=>"001001000",
  45712=>"000110010",
  45713=>"000000000",
  45714=>"011000000",
  45715=>"000000000",
  45716=>"011000000",
  45717=>"100000100",
  45718=>"100111111",
  45719=>"111001000",
  45720=>"011000100",
  45721=>"111111111",
  45722=>"101110111",
  45723=>"101111111",
  45724=>"110110111",
  45725=>"000000111",
  45726=>"011001001",
  45727=>"011001000",
  45728=>"001000000",
  45729=>"110110000",
  45730=>"000111110",
  45731=>"011000101",
  45732=>"111111000",
  45733=>"110110100",
  45734=>"001111000",
  45735=>"000001011",
  45736=>"000000000",
  45737=>"111001011",
  45738=>"001000000",
  45739=>"010000000",
  45740=>"011011000",
  45741=>"100100000",
  45742=>"000000000",
  45743=>"011000111",
  45744=>"111111111",
  45745=>"000001011",
  45746=>"110111010",
  45747=>"011000000",
  45748=>"000000001",
  45749=>"111111111",
  45750=>"000110110",
  45751=>"000011001",
  45752=>"100101100",
  45753=>"001001001",
  45754=>"000000001",
  45755=>"110000000",
  45756=>"101000000",
  45757=>"000000001",
  45758=>"001111000",
  45759=>"111111111",
  45760=>"110100100",
  45761=>"001110110",
  45762=>"111101101",
  45763=>"111000000",
  45764=>"000000111",
  45765=>"000111111",
  45766=>"000111111",
  45767=>"000100111",
  45768=>"110000111",
  45769=>"111111010",
  45770=>"001000001",
  45771=>"000111111",
  45772=>"111111001",
  45773=>"000000011",
  45774=>"000000011",
  45775=>"000000000",
  45776=>"111111111",
  45777=>"111110000",
  45778=>"010000000",
  45779=>"010111111",
  45780=>"110111111",
  45781=>"100001001",
  45782=>"000000001",
  45783=>"111111101",
  45784=>"010000100",
  45785=>"110000000",
  45786=>"111111111",
  45787=>"000001111",
  45788=>"110111110",
  45789=>"110110000",
  45790=>"111111111",
  45791=>"111111101",
  45792=>"001000000",
  45793=>"000000000",
  45794=>"111111111",
  45795=>"000000111",
  45796=>"111101001",
  45797=>"100110110",
  45798=>"110110011",
  45799=>"000001011",
  45800=>"000000001",
  45801=>"111101101",
  45802=>"000000000",
  45803=>"011000000",
  45804=>"000000000",
  45805=>"111110000",
  45806=>"111111111",
  45807=>"111010000",
  45808=>"111111011",
  45809=>"000000000",
  45810=>"000010000",
  45811=>"110110000",
  45812=>"000000000",
  45813=>"110100000",
  45814=>"011111111",
  45815=>"100111000",
  45816=>"111110000",
  45817=>"000000000",
  45818=>"000001001",
  45819=>"111111111",
  45820=>"111111111",
  45821=>"111111000",
  45822=>"000000001",
  45823=>"010011011",
  45824=>"000000001",
  45825=>"100000000",
  45826=>"111111111",
  45827=>"110100111",
  45828=>"000110000",
  45829=>"000101111",
  45830=>"000000000",
  45831=>"001001001",
  45832=>"111111111",
  45833=>"111011011",
  45834=>"111111001",
  45835=>"000010010",
  45836=>"010000110",
  45837=>"000000000",
  45838=>"000110000",
  45839=>"000001000",
  45840=>"000001001",
  45841=>"110111110",
  45842=>"111100111",
  45843=>"001001001",
  45844=>"111111110",
  45845=>"100100000",
  45846=>"000000000",
  45847=>"001110110",
  45848=>"100101101",
  45849=>"001001000",
  45850=>"000000001",
  45851=>"110000111",
  45852=>"000001000",
  45853=>"000001000",
  45854=>"000000000",
  45855=>"000000110",
  45856=>"110100111",
  45857=>"111111000",
  45858=>"111111111",
  45859=>"110101111",
  45860=>"110000000",
  45861=>"111110110",
  45862=>"111111000",
  45863=>"000000001",
  45864=>"000000000",
  45865=>"111111010",
  45866=>"111111110",
  45867=>"001000000",
  45868=>"111101111",
  45869=>"001101111",
  45870=>"111111011",
  45871=>"010000000",
  45872=>"111111011",
  45873=>"111111110",
  45874=>"111011001",
  45875=>"111111000",
  45876=>"001000000",
  45877=>"110111110",
  45878=>"110100000",
  45879=>"011010000",
  45880=>"000000000",
  45881=>"111111111",
  45882=>"000100001",
  45883=>"010111111",
  45884=>"001001001",
  45885=>"111111000",
  45886=>"001001000",
  45887=>"000000000",
  45888=>"000000111",
  45889=>"000001111",
  45890=>"000000011",
  45891=>"111111111",
  45892=>"111111001",
  45893=>"111001000",
  45894=>"110111111",
  45895=>"110110000",
  45896=>"111111111",
  45897=>"100000000",
  45898=>"011000000",
  45899=>"000000000",
  45900=>"110000000",
  45901=>"111111111",
  45902=>"011111111",
  45903=>"000000000",
  45904=>"000000000",
  45905=>"001001001",
  45906=>"101110000",
  45907=>"000000111",
  45908=>"111010000",
  45909=>"011011011",
  45910=>"000000111",
  45911=>"110111000",
  45912=>"110111010",
  45913=>"111111000",
  45914=>"001001111",
  45915=>"111111100",
  45916=>"001001001",
  45917=>"000100000",
  45918=>"110111000",
  45919=>"000000101",
  45920=>"000000001",
  45921=>"001000001",
  45922=>"111111100",
  45923=>"000000101",
  45924=>"000001001",
  45925=>"000000000",
  45926=>"100100111",
  45927=>"111111000",
  45928=>"000000011",
  45929=>"000111111",
  45930=>"000001001",
  45931=>"111111111",
  45932=>"110111111",
  45933=>"000000011",
  45934=>"111011111",
  45935=>"000000000",
  45936=>"001111001",
  45937=>"000000001",
  45938=>"000110110",
  45939=>"100110100",
  45940=>"000111111",
  45941=>"000000001",
  45942=>"010000011",
  45943=>"000101011",
  45944=>"000000000",
  45945=>"111111000",
  45946=>"111111110",
  45947=>"000000000",
  45948=>"111111111",
  45949=>"001000000",
  45950=>"111000000",
  45951=>"111111101",
  45952=>"100111001",
  45953=>"000000000",
  45954=>"001011111",
  45955=>"101101101",
  45956=>"000000111",
  45957=>"010110000",
  45958=>"111111111",
  45959=>"110111111",
  45960=>"001000000",
  45961=>"010010111",
  45962=>"000111111",
  45963=>"100111111",
  45964=>"101100100",
  45965=>"000111111",
  45966=>"000110000",
  45967=>"000000101",
  45968=>"000000100",
  45969=>"111111110",
  45970=>"000101111",
  45971=>"000000000",
  45972=>"000000000",
  45973=>"000010010",
  45974=>"101000000",
  45975=>"111110000",
  45976=>"111111111",
  45977=>"111000001",
  45978=>"111001111",
  45979=>"111111111",
  45980=>"111111110",
  45981=>"100000000",
  45982=>"110100101",
  45983=>"111000000",
  45984=>"000000000",
  45985=>"000000111",
  45986=>"111111010",
  45987=>"111011000",
  45988=>"111001000",
  45989=>"000010011",
  45990=>"111111111",
  45991=>"000000000",
  45992=>"111011111",
  45993=>"111011001",
  45994=>"000001011",
  45995=>"110110111",
  45996=>"101100100",
  45997=>"110100111",
  45998=>"000000000",
  45999=>"000000100",
  46000=>"001000000",
  46001=>"111111000",
  46002=>"111001000",
  46003=>"000000000",
  46004=>"111000000",
  46005=>"000000000",
  46006=>"111001001",
  46007=>"000000001",
  46008=>"000000011",
  46009=>"111111111",
  46010=>"101100000",
  46011=>"110000000",
  46012=>"111000000",
  46013=>"110111111",
  46014=>"001011000",
  46015=>"100001001",
  46016=>"000000000",
  46017=>"000000000",
  46018=>"000000000",
  46019=>"110111000",
  46020=>"101101111",
  46021=>"011001000",
  46022=>"001001000",
  46023=>"000000101",
  46024=>"011000000",
  46025=>"010010000",
  46026=>"000100000",
  46027=>"101000000",
  46028=>"111011000",
  46029=>"111111000",
  46030=>"011111100",
  46031=>"011011000",
  46032=>"000000000",
  46033=>"111111111",
  46034=>"111111000",
  46035=>"000000111",
  46036=>"111111011",
  46037=>"000000111",
  46038=>"110000111",
  46039=>"001001000",
  46040=>"000101111",
  46041=>"000010110",
  46042=>"000000111",
  46043=>"111111001",
  46044=>"101111111",
  46045=>"000000001",
  46046=>"000000100",
  46047=>"000000000",
  46048=>"111111011",
  46049=>"011011011",
  46050=>"000000111",
  46051=>"000000111",
  46052=>"111101001",
  46053=>"000000001",
  46054=>"000000010",
  46055=>"100100101",
  46056=>"111100100",
  46057=>"000000000",
  46058=>"000000000",
  46059=>"000001001",
  46060=>"111111110",
  46061=>"100110000",
  46062=>"000000111",
  46063=>"111000000",
  46064=>"011011000",
  46065=>"000111111",
  46066=>"011111011",
  46067=>"001111001",
  46068=>"000000000",
  46069=>"000000000",
  46070=>"111111011",
  46071=>"000001001",
  46072=>"000011010",
  46073=>"000000000",
  46074=>"101000000",
  46075=>"111111111",
  46076=>"100100110",
  46077=>"001101001",
  46078=>"010011111",
  46079=>"000000001",
  46080=>"000110110",
  46081=>"111111111",
  46082=>"101000000",
  46083=>"001101101",
  46084=>"110100000",
  46085=>"001111000",
  46086=>"000000000",
  46087=>"111101110",
  46088=>"110111000",
  46089=>"000100110",
  46090=>"000010000",
  46091=>"100010000",
  46092=>"100101001",
  46093=>"000000111",
  46094=>"000100110",
  46095=>"111111111",
  46096=>"000000100",
  46097=>"000000000",
  46098=>"110111011",
  46099=>"011000000",
  46100=>"100110110",
  46101=>"000000011",
  46102=>"001000000",
  46103=>"000010000",
  46104=>"110010000",
  46105=>"001011110",
  46106=>"000111100",
  46107=>"000010110",
  46108=>"111111100",
  46109=>"111111000",
  46110=>"111111001",
  46111=>"000000001",
  46112=>"111111011",
  46113=>"011000000",
  46114=>"110111111",
  46115=>"000000000",
  46116=>"111111101",
  46117=>"010110111",
  46118=>"001000101",
  46119=>"010011000",
  46120=>"000000111",
  46121=>"000000000",
  46122=>"111111111",
  46123=>"000000000",
  46124=>"000000111",
  46125=>"000100111",
  46126=>"000000000",
  46127=>"001011111",
  46128=>"101111111",
  46129=>"000000011",
  46130=>"000000000",
  46131=>"111111111",
  46132=>"111111101",
  46133=>"110110110",
  46134=>"111111111",
  46135=>"000000000",
  46136=>"011000111",
  46137=>"001111111",
  46138=>"000000000",
  46139=>"000100111",
  46140=>"000000100",
  46141=>"111111111",
  46142=>"000000000",
  46143=>"111111111",
  46144=>"011010000",
  46145=>"101001001",
  46146=>"100000001",
  46147=>"011111111",
  46148=>"000000000",
  46149=>"000110110",
  46150=>"000000100",
  46151=>"111111111",
  46152=>"011011011",
  46153=>"111111111",
  46154=>"011000000",
  46155=>"111110101",
  46156=>"001000000",
  46157=>"000000001",
  46158=>"000000000",
  46159=>"111111111",
  46160=>"111001000",
  46161=>"000000100",
  46162=>"000000000",
  46163=>"111111101",
  46164=>"001011111",
  46165=>"100110111",
  46166=>"110110100",
  46167=>"111111111",
  46168=>"000000100",
  46169=>"101100101",
  46170=>"000000010",
  46171=>"000000010",
  46172=>"000110111",
  46173=>"000001101",
  46174=>"011011111",
  46175=>"111011000",
  46176=>"001101110",
  46177=>"000111000",
  46178=>"000000110",
  46179=>"000000000",
  46180=>"111111100",
  46181=>"111111011",
  46182=>"001001000",
  46183=>"010110110",
  46184=>"111111000",
  46185=>"111111111",
  46186=>"000000111",
  46187=>"001000111",
  46188=>"100111001",
  46189=>"000000000",
  46190=>"111111111",
  46191=>"111111111",
  46192=>"000000000",
  46193=>"011001111",
  46194=>"000001011",
  46195=>"111111111",
  46196=>"010111111",
  46197=>"000010111",
  46198=>"001111111",
  46199=>"010010000",
  46200=>"011001001",
  46201=>"000000000",
  46202=>"000000000",
  46203=>"000000000",
  46204=>"111000000",
  46205=>"000010000",
  46206=>"010000111",
  46207=>"000001000",
  46208=>"000000000",
  46209=>"111110111",
  46210=>"000111100",
  46211=>"111111110",
  46212=>"001111111",
  46213=>"110000000",
  46214=>"011000110",
  46215=>"001000101",
  46216=>"100100110",
  46217=>"000000000",
  46218=>"110100000",
  46219=>"000000000",
  46220=>"110110110",
  46221=>"100111110",
  46222=>"000000000",
  46223=>"000000000",
  46224=>"111101111",
  46225=>"111111001",
  46226=>"000000111",
  46227=>"100000000",
  46228=>"000000001",
  46229=>"000010000",
  46230=>"000011111",
  46231=>"100000100",
  46232=>"000000000",
  46233=>"001001111",
  46234=>"111110100",
  46235=>"000000000",
  46236=>"111111111",
  46237=>"111011000",
  46238=>"011001000",
  46239=>"000000010",
  46240=>"000000000",
  46241=>"111111111",
  46242=>"111111111",
  46243=>"000000000",
  46244=>"011000000",
  46245=>"111011111",
  46246=>"111000000",
  46247=>"001000000",
  46248=>"000010000",
  46249=>"111011111",
  46250=>"000001111",
  46251=>"001001101",
  46252=>"000000010",
  46253=>"000111111",
  46254=>"111111111",
  46255=>"100111101",
  46256=>"000000111",
  46257=>"110110111",
  46258=>"111111111",
  46259=>"101000000",
  46260=>"111111000",
  46261=>"111110011",
  46262=>"111001011",
  46263=>"111111111",
  46264=>"000000000",
  46265=>"111111111",
  46266=>"110100000",
  46267=>"011010111",
  46268=>"000000000",
  46269=>"000110110",
  46270=>"000111111",
  46271=>"111111111",
  46272=>"111111111",
  46273=>"000000001",
  46274=>"111110000",
  46275=>"001000000",
  46276=>"000010110",
  46277=>"000000000",
  46278=>"000011101",
  46279=>"011011001",
  46280=>"001001111",
  46281=>"000000000",
  46282=>"011011000",
  46283=>"111111111",
  46284=>"000000000",
  46285=>"000110110",
  46286=>"111111010",
  46287=>"000111001",
  46288=>"000000000",
  46289=>"000100000",
  46290=>"000000000",
  46291=>"000000000",
  46292=>"111111111",
  46293=>"010011111",
  46294=>"000000000",
  46295=>"011100100",
  46296=>"111110110",
  46297=>"111111100",
  46298=>"000011111",
  46299=>"111111111",
  46300=>"000000000",
  46301=>"000000000",
  46302=>"111111111",
  46303=>"111111111",
  46304=>"111000100",
  46305=>"001001001",
  46306=>"111111111",
  46307=>"001000000",
  46308=>"111111111",
  46309=>"000000000",
  46310=>"000010011",
  46311=>"000000110",
  46312=>"000000000",
  46313=>"100110100",
  46314=>"111111111",
  46315=>"000111111",
  46316=>"000111111",
  46317=>"101000111",
  46318=>"111000101",
  46319=>"000000000",
  46320=>"000010010",
  46321=>"111111111",
  46322=>"110111111",
  46323=>"111010001",
  46324=>"111111111",
  46325=>"000000000",
  46326=>"100110110",
  46327=>"111000000",
  46328=>"000000000",
  46329=>"000000000",
  46330=>"111111011",
  46331=>"111111111",
  46332=>"111111111",
  46333=>"011011100",
  46334=>"000000000",
  46335=>"000000000",
  46336=>"010110000",
  46337=>"001000000",
  46338=>"111011000",
  46339=>"011000000",
  46340=>"000010010",
  46341=>"111111111",
  46342=>"000000000",
  46343=>"000000100",
  46344=>"111111001",
  46345=>"111111111",
  46346=>"000000000",
  46347=>"111111110",
  46348=>"100000001",
  46349=>"000000011",
  46350=>"011111100",
  46351=>"110111111",
  46352=>"000001011",
  46353=>"111111111",
  46354=>"000001001",
  46355=>"110010111",
  46356=>"000000000",
  46357=>"000000000",
  46358=>"100000100",
  46359=>"010010000",
  46360=>"111111100",
  46361=>"110111111",
  46362=>"000010000",
  46363=>"000000000",
  46364=>"110110110",
  46365=>"000111110",
  46366=>"000000000",
  46367=>"111111111",
  46368=>"011011001",
  46369=>"111111011",
  46370=>"000100110",
  46371=>"001000000",
  46372=>"000001101",
  46373=>"100000111",
  46374=>"001001011",
  46375=>"111101111",
  46376=>"111011111",
  46377=>"011011001",
  46378=>"100110111",
  46379=>"100000000",
  46380=>"000000001",
  46381=>"010000100",
  46382=>"000000000",
  46383=>"000000000",
  46384=>"111111111",
  46385=>"111111111",
  46386=>"000000001",
  46387=>"111110110",
  46388=>"000110111",
  46389=>"011001011",
  46390=>"101111001",
  46391=>"000010000",
  46392=>"001000000",
  46393=>"111000011",
  46394=>"011011011",
  46395=>"110111001",
  46396=>"010010000",
  46397=>"000000100",
  46398=>"000000000",
  46399=>"010010010",
  46400=>"111110111",
  46401=>"011011111",
  46402=>"000101111",
  46403=>"000010010",
  46404=>"110111111",
  46405=>"111111111",
  46406=>"000000000",
  46407=>"111111111",
  46408=>"001001001",
  46409=>"000000000",
  46410=>"111111111",
  46411=>"110111011",
  46412=>"000000000",
  46413=>"000101111",
  46414=>"000000000",
  46415=>"111111111",
  46416=>"000000000",
  46417=>"011001001",
  46418=>"111111111",
  46419=>"000111111",
  46420=>"110100000",
  46421=>"011011011",
  46422=>"111111111",
  46423=>"111100100",
  46424=>"101100110",
  46425=>"111000000",
  46426=>"000000000",
  46427=>"100000000",
  46428=>"000000000",
  46429=>"000000000",
  46430=>"101000010",
  46431=>"000011101",
  46432=>"000000000",
  46433=>"001001101",
  46434=>"111110110",
  46435=>"000000001",
  46436=>"000000111",
  46437=>"000000011",
  46438=>"111111111",
  46439=>"000000000",
  46440=>"001100100",
  46441=>"111111111",
  46442=>"000001000",
  46443=>"000000001",
  46444=>"111001001",
  46445=>"111000110",
  46446=>"000000000",
  46447=>"111011011",
  46448=>"000000000",
  46449=>"000000000",
  46450=>"111000000",
  46451=>"111111001",
  46452=>"000000000",
  46453=>"111111111",
  46454=>"000000000",
  46455=>"001001000",
  46456=>"000000000",
  46457=>"000000000",
  46458=>"000000111",
  46459=>"010010011",
  46460=>"000000100",
  46461=>"111111111",
  46462=>"000000000",
  46463=>"111111111",
  46464=>"011010010",
  46465=>"010110111",
  46466=>"000011011",
  46467=>"000110110",
  46468=>"000100100",
  46469=>"000000000",
  46470=>"000001111",
  46471=>"000000000",
  46472=>"000000000",
  46473=>"011011011",
  46474=>"000000000",
  46475=>"111111100",
  46476=>"101000000",
  46477=>"010010110",
  46478=>"111111111",
  46479=>"111111111",
  46480=>"000000000",
  46481=>"000111111",
  46482=>"000111100",
  46483=>"000000000",
  46484=>"000110010",
  46485=>"000000010",
  46486=>"010000000",
  46487=>"010001001",
  46488=>"000000000",
  46489=>"010010000",
  46490=>"111010000",
  46491=>"111011111",
  46492=>"110000000",
  46493=>"000000000",
  46494=>"000111111",
  46495=>"111111100",
  46496=>"000000000",
  46497=>"111111101",
  46498=>"000000000",
  46499=>"111011111",
  46500=>"010111000",
  46501=>"001000001",
  46502=>"000000000",
  46503=>"000010000",
  46504=>"000000000",
  46505=>"000000000",
  46506=>"010000000",
  46507=>"111000001",
  46508=>"111111111",
  46509=>"100100000",
  46510=>"010110000",
  46511=>"111001001",
  46512=>"000111111",
  46513=>"000011011",
  46514=>"100000111",
  46515=>"000000001",
  46516=>"001000000",
  46517=>"000001001",
  46518=>"000110111",
  46519=>"111111100",
  46520=>"011111110",
  46521=>"110111111",
  46522=>"111100110",
  46523=>"000010011",
  46524=>"001111111",
  46525=>"110111100",
  46526=>"101111101",
  46527=>"000000010",
  46528=>"111001101",
  46529=>"000000000",
  46530=>"111011001",
  46531=>"000100110",
  46532=>"001111111",
  46533=>"011011101",
  46534=>"000001001",
  46535=>"001001101",
  46536=>"000100110",
  46537=>"011110111",
  46538=>"111001000",
  46539=>"000111111",
  46540=>"111101100",
  46541=>"000000000",
  46542=>"000100100",
  46543=>"100111111",
  46544=>"100111100",
  46545=>"011110111",
  46546=>"000000000",
  46547=>"000100111",
  46548=>"000100100",
  46549=>"000100111",
  46550=>"000000000",
  46551=>"111111111",
  46552=>"111111111",
  46553=>"000000001",
  46554=>"000000011",
  46555=>"111110000",
  46556=>"001001011",
  46557=>"111101011",
  46558=>"111111010",
  46559=>"011111011",
  46560=>"000000000",
  46561=>"111111111",
  46562=>"100110010",
  46563=>"110001000",
  46564=>"111111001",
  46565=>"111111110",
  46566=>"000000100",
  46567=>"000000011",
  46568=>"000000110",
  46569=>"111000000",
  46570=>"000000000",
  46571=>"111111111",
  46572=>"111111111",
  46573=>"011001001",
  46574=>"100100111",
  46575=>"010000110",
  46576=>"000000000",
  46577=>"000000111",
  46578=>"000000000",
  46579=>"101111101",
  46580=>"000011111",
  46581=>"001000100",
  46582=>"000000000",
  46583=>"010011111",
  46584=>"001000000",
  46585=>"000000001",
  46586=>"100000000",
  46587=>"000000000",
  46588=>"011011000",
  46589=>"000000101",
  46590=>"010110000",
  46591=>"100000000",
  46592=>"000000000",
  46593=>"101110110",
  46594=>"111110101",
  46595=>"000000000",
  46596=>"011111111",
  46597=>"000000000",
  46598=>"010000000",
  46599=>"100100110",
  46600=>"111111111",
  46601=>"110111111",
  46602=>"000000000",
  46603=>"001000000",
  46604=>"100110001",
  46605=>"111001111",
  46606=>"000111110",
  46607=>"001001111",
  46608=>"010111000",
  46609=>"000000011",
  46610=>"011011000",
  46611=>"000000000",
  46612=>"000001011",
  46613=>"001001111",
  46614=>"110110111",
  46615=>"111011001",
  46616=>"111110100",
  46617=>"000000000",
  46618=>"111111111",
  46619=>"111111111",
  46620=>"000111010",
  46621=>"000010010",
  46622=>"111011011",
  46623=>"010111111",
  46624=>"001000000",
  46625=>"111111111",
  46626=>"101101111",
  46627=>"000000001",
  46628=>"111110000",
  46629=>"111111011",
  46630=>"111111111",
  46631=>"000101111",
  46632=>"110000111",
  46633=>"001001111",
  46634=>"110111111",
  46635=>"000000000",
  46636=>"001111111",
  46637=>"000000000",
  46638=>"111111110",
  46639=>"001111111",
  46640=>"001101101",
  46641=>"000000000",
  46642=>"001011111",
  46643=>"100100100",
  46644=>"000000000",
  46645=>"000010011",
  46646=>"000110111",
  46647=>"000000010",
  46648=>"001001101",
  46649=>"001001101",
  46650=>"111111110",
  46651=>"000000000",
  46652=>"111000000",
  46653=>"010011111",
  46654=>"111101001",
  46655=>"010011010",
  46656=>"111111111",
  46657=>"111000000",
  46658=>"010111110",
  46659=>"000000000",
  46660=>"011001011",
  46661=>"000000000",
  46662=>"111000000",
  46663=>"100111111",
  46664=>"011111011",
  46665=>"111000000",
  46666=>"000000011",
  46667=>"001111111",
  46668=>"111111100",
  46669=>"110010000",
  46670=>"111100100",
  46671=>"111111111",
  46672=>"111111111",
  46673=>"010000100",
  46674=>"111111000",
  46675=>"011010111",
  46676=>"000000000",
  46677=>"000111110",
  46678=>"111101000",
  46679=>"111000000",
  46680=>"111111111",
  46681=>"000000000",
  46682=>"010000000",
  46683=>"100110100",
  46684=>"001000001",
  46685=>"001001111",
  46686=>"110111011",
  46687=>"001011011",
  46688=>"011000000",
  46689=>"111111111",
  46690=>"101101111",
  46691=>"101000111",
  46692=>"101100000",
  46693=>"001000110",
  46694=>"011111111",
  46695=>"010000000",
  46696=>"111100111",
  46697=>"000000101",
  46698=>"000000110",
  46699=>"000010110",
  46700=>"011011001",
  46701=>"111000000",
  46702=>"111111000",
  46703=>"000111111",
  46704=>"000111111",
  46705=>"000011111",
  46706=>"100111111",
  46707=>"000111111",
  46708=>"000000000",
  46709=>"000011011",
  46710=>"000111000",
  46711=>"000000000",
  46712=>"101101111",
  46713=>"101001101",
  46714=>"111111111",
  46715=>"111111111",
  46716=>"111110111",
  46717=>"110110111",
  46718=>"111111111",
  46719=>"011111001",
  46720=>"100100000",
  46721=>"000111111",
  46722=>"100100000",
  46723=>"111100100",
  46724=>"111111110",
  46725=>"000000100",
  46726=>"010110110",
  46727=>"000000000",
  46728=>"100000000",
  46729=>"011111111",
  46730=>"011001111",
  46731=>"111101100",
  46732=>"001101111",
  46733=>"101000000",
  46734=>"110011111",
  46735=>"001001100",
  46736=>"000100111",
  46737=>"111111101",
  46738=>"001000000",
  46739=>"001000000",
  46740=>"001111111",
  46741=>"111100111",
  46742=>"000100100",
  46743=>"000100111",
  46744=>"111111111",
  46745=>"011000000",
  46746=>"000010111",
  46747=>"101111111",
  46748=>"000000000",
  46749=>"111110110",
  46750=>"000000000",
  46751=>"111001000",
  46752=>"000000000",
  46753=>"111101000",
  46754=>"000001101",
  46755=>"001000110",
  46756=>"111111011",
  46757=>"110101111",
  46758=>"101001101",
  46759=>"011000111",
  46760=>"001001111",
  46761=>"001001111",
  46762=>"000000000",
  46763=>"111111010",
  46764=>"000000110",
  46765=>"110100100",
  46766=>"111111111",
  46767=>"001010111",
  46768=>"001001101",
  46769=>"011111011",
  46770=>"111111011",
  46771=>"111111111",
  46772=>"000000001",
  46773=>"011111000",
  46774=>"000111111",
  46775=>"111111001",
  46776=>"111111111",
  46777=>"111111111",
  46778=>"100111000",
  46779=>"101001001",
  46780=>"000000011",
  46781=>"111001000",
  46782=>"000000110",
  46783=>"001000100",
  46784=>"101000000",
  46785=>"100000100",
  46786=>"000000000",
  46787=>"000000000",
  46788=>"000000000",
  46789=>"000000000",
  46790=>"010110110",
  46791=>"000000100",
  46792=>"001000111",
  46793=>"111111000",
  46794=>"001000001",
  46795=>"000000111",
  46796=>"110110110",
  46797=>"111111100",
  46798=>"001000001",
  46799=>"111000000",
  46800=>"111111111",
  46801=>"111000010",
  46802=>"100000000",
  46803=>"000000000",
  46804=>"001000001",
  46805=>"111111111",
  46806=>"000000001",
  46807=>"000000000",
  46808=>"000001101",
  46809=>"111111101",
  46810=>"111100000",
  46811=>"000000000",
  46812=>"000000000",
  46813=>"111111010",
  46814=>"000000000",
  46815=>"000111111",
  46816=>"111111111",
  46817=>"000000000",
  46818=>"000000000",
  46819=>"011111000",
  46820=>"001001001",
  46821=>"111111111",
  46822=>"000111111",
  46823=>"111111001",
  46824=>"000000000",
  46825=>"001001101",
  46826=>"111111110",
  46827=>"011101101",
  46828=>"000010011",
  46829=>"011111111",
  46830=>"111111001",
  46831=>"111111000",
  46832=>"110110000",
  46833=>"000000000",
  46834=>"111110111",
  46835=>"101111011",
  46836=>"000000110",
  46837=>"110100110",
  46838=>"111111010",
  46839=>"000000000",
  46840=>"111000000",
  46841=>"001001001",
  46842=>"111111111",
  46843=>"111111111",
  46844=>"110110110",
  46845=>"100110111",
  46846=>"111111111",
  46847=>"110111111",
  46848=>"000001001",
  46849=>"100100110",
  46850=>"000000000",
  46851=>"111111111",
  46852=>"111111000",
  46853=>"111111000",
  46854=>"111111111",
  46855=>"100111111",
  46856=>"001111111",
  46857=>"101001001",
  46858=>"110111100",
  46859=>"111110100",
  46860=>"000000110",
  46861=>"000100000",
  46862=>"111111111",
  46863=>"111000000",
  46864=>"111101001",
  46865=>"000001101",
  46866=>"110110010",
  46867=>"000000000",
  46868=>"110000000",
  46869=>"000011111",
  46870=>"001001001",
  46871=>"000110110",
  46872=>"111100110",
  46873=>"111111001",
  46874=>"000000111",
  46875=>"001000000",
  46876=>"111111101",
  46877=>"000000000",
  46878=>"011111000",
  46879=>"111100000",
  46880=>"111111111",
  46881=>"111111100",
  46882=>"001100100",
  46883=>"001110110",
  46884=>"111111111",
  46885=>"000010011",
  46886=>"111001100",
  46887=>"000000000",
  46888=>"001000000",
  46889=>"000001111",
  46890=>"111000000",
  46891=>"100100110",
  46892=>"111111111",
  46893=>"101011111",
  46894=>"100100111",
  46895=>"111111111",
  46896=>"001001001",
  46897=>"111000000",
  46898=>"000101001",
  46899=>"011111100",
  46900=>"111101111",
  46901=>"000001001",
  46902=>"001000000",
  46903=>"000001111",
  46904=>"000000000",
  46905=>"000000000",
  46906=>"111011000",
  46907=>"000000000",
  46908=>"001001111",
  46909=>"110111010",
  46910=>"000000000",
  46911=>"001101101",
  46912=>"000101111",
  46913=>"100000011",
  46914=>"001111111",
  46915=>"111000000",
  46916=>"101111111",
  46917=>"001001101",
  46918=>"000000001",
  46919=>"110110111",
  46920=>"111101101",
  46921=>"111101000",
  46922=>"001001001",
  46923=>"101000100",
  46924=>"011011001",
  46925=>"000100111",
  46926=>"110110110",
  46927=>"011011111",
  46928=>"000010110",
  46929=>"100000000",
  46930=>"001001011",
  46931=>"000000111",
  46932=>"000000001",
  46933=>"011001011",
  46934=>"111111111",
  46935=>"111111111",
  46936=>"111111000",
  46937=>"111111111",
  46938=>"000000111",
  46939=>"010110111",
  46940=>"111001000",
  46941=>"000001111",
  46942=>"111111111",
  46943=>"000000001",
  46944=>"000000111",
  46945=>"000100111",
  46946=>"110110100",
  46947=>"000000000",
  46948=>"000000100",
  46949=>"000000000",
  46950=>"110100000",
  46951=>"110110110",
  46952=>"110000001",
  46953=>"000000111",
  46954=>"000000000",
  46955=>"110110110",
  46956=>"000010000",
  46957=>"111111110",
  46958=>"111111011",
  46959=>"111001000",
  46960=>"101111111",
  46961=>"101001001",
  46962=>"000000010",
  46963=>"000110111",
  46964=>"101111111",
  46965=>"000011111",
  46966=>"001000101",
  46967=>"001001111",
  46968=>"000000101",
  46969=>"011011111",
  46970=>"000000101",
  46971=>"010110010",
  46972=>"000001111",
  46973=>"111111000",
  46974=>"000000111",
  46975=>"000000000",
  46976=>"110000110",
  46977=>"001100100",
  46978=>"000000011",
  46979=>"000000000",
  46980=>"111111100",
  46981=>"111111111",
  46982=>"111111111",
  46983=>"111111001",
  46984=>"111101001",
  46985=>"100111111",
  46986=>"000010110",
  46987=>"000101111",
  46988=>"101000111",
  46989=>"111111111",
  46990=>"010000001",
  46991=>"000000000",
  46992=>"000000000",
  46993=>"000000001",
  46994=>"001001001",
  46995=>"000000001",
  46996=>"111110110",
  46997=>"111111111",
  46998=>"110001001",
  46999=>"011011011",
  47000=>"000000111",
  47001=>"011000000",
  47002=>"100111111",
  47003=>"001111111",
  47004=>"000000111",
  47005=>"111010000",
  47006=>"101111000",
  47007=>"000001001",
  47008=>"111111001",
  47009=>"110110111",
  47010=>"000111111",
  47011=>"000000000",
  47012=>"010011000",
  47013=>"100000001",
  47014=>"101101111",
  47015=>"000000000",
  47016=>"101000010",
  47017=>"111111001",
  47018=>"001001100",
  47019=>"000000000",
  47020=>"000000000",
  47021=>"000010111",
  47022=>"000001111",
  47023=>"001001111",
  47024=>"011000000",
  47025=>"000111111",
  47026=>"111111111",
  47027=>"000000000",
  47028=>"111000000",
  47029=>"000000000",
  47030=>"111111111",
  47031=>"010001111",
  47032=>"001000000",
  47033=>"001111111",
  47034=>"000000110",
  47035=>"111100000",
  47036=>"110110000",
  47037=>"100000101",
  47038=>"000000000",
  47039=>"011011011",
  47040=>"001000000",
  47041=>"111111110",
  47042=>"000111111",
  47043=>"111111110",
  47044=>"111111110",
  47045=>"001001011",
  47046=>"000001111",
  47047=>"000000000",
  47048=>"110110101",
  47049=>"000111111",
  47050=>"111111111",
  47051=>"010111111",
  47052=>"111000001",
  47053=>"110111111",
  47054=>"111110111",
  47055=>"000001111",
  47056=>"111111001",
  47057=>"000110010",
  47058=>"111000100",
  47059=>"001000111",
  47060=>"000100000",
  47061=>"111011010",
  47062=>"111111111",
  47063=>"111010111",
  47064=>"101111101",
  47065=>"000000001",
  47066=>"111111111",
  47067=>"111100000",
  47068=>"000010011",
  47069=>"000001111",
  47070=>"100100110",
  47071=>"000000110",
  47072=>"111111111",
  47073=>"101100101",
  47074=>"000111111",
  47075=>"000000011",
  47076=>"011111111",
  47077=>"000000000",
  47078=>"000011111",
  47079=>"000000000",
  47080=>"111100111",
  47081=>"000000010",
  47082=>"111001000",
  47083=>"111000000",
  47084=>"000000111",
  47085=>"101100100",
  47086=>"111101111",
  47087=>"111111111",
  47088=>"111111010",
  47089=>"001001000",
  47090=>"111011011",
  47091=>"101111111",
  47092=>"010110110",
  47093=>"011001001",
  47094=>"111111111",
  47095=>"111001101",
  47096=>"110000100",
  47097=>"000110100",
  47098=>"000000000",
  47099=>"000001001",
  47100=>"111111000",
  47101=>"001001000",
  47102=>"000010000",
  47103=>"000000001",
  47104=>"001111111",
  47105=>"001001111",
  47106=>"011111111",
  47107=>"100100101",
  47108=>"111100000",
  47109=>"000001001",
  47110=>"011110000",
  47111=>"111111111",
  47112=>"000000111",
  47113=>"111111111",
  47114=>"101111111",
  47115=>"000101111",
  47116=>"101111111",
  47117=>"111111000",
  47118=>"000000000",
  47119=>"111000000",
  47120=>"011011000",
  47121=>"111111111",
  47122=>"111111000",
  47123=>"111000000",
  47124=>"110111111",
  47125=>"000000110",
  47126=>"000000000",
  47127=>"001101111",
  47128=>"001000000",
  47129=>"101101000",
  47130=>"011001111",
  47131=>"000011001",
  47132=>"010111000",
  47133=>"000000000",
  47134=>"100100100",
  47135=>"110011011",
  47136=>"000100111",
  47137=>"110000000",
  47138=>"000000000",
  47139=>"111111111",
  47140=>"000000000",
  47141=>"100111111",
  47142=>"000000000",
  47143=>"000100110",
  47144=>"111101111",
  47145=>"000000000",
  47146=>"000000111",
  47147=>"000111111",
  47148=>"111111110",
  47149=>"111111110",
  47150=>"111111111",
  47151=>"100000001",
  47152=>"111101001",
  47153=>"111111000",
  47154=>"011100101",
  47155=>"111111111",
  47156=>"000111000",
  47157=>"101000000",
  47158=>"000000000",
  47159=>"000000100",
  47160=>"111111111",
  47161=>"101101111",
  47162=>"100001000",
  47163=>"000000111",
  47164=>"000100111",
  47165=>"111110111",
  47166=>"111111110",
  47167=>"000000000",
  47168=>"111111100",
  47169=>"000000000",
  47170=>"111111111",
  47171=>"000111100",
  47172=>"111111001",
  47173=>"001111111",
  47174=>"000001111",
  47175=>"111111000",
  47176=>"000000000",
  47177=>"000000111",
  47178=>"000111111",
  47179=>"111111111",
  47180=>"111100000",
  47181=>"000000000",
  47182=>"111001111",
  47183=>"100110110",
  47184=>"100111101",
  47185=>"111111111",
  47186=>"000000001",
  47187=>"001001111",
  47188=>"000110010",
  47189=>"100110111",
  47190=>"111101000",
  47191=>"000100000",
  47192=>"111111111",
  47193=>"011101111",
  47194=>"000001001",
  47195=>"110110110",
  47196=>"111111000",
  47197=>"001000000",
  47198=>"111111011",
  47199=>"011111111",
  47200=>"111000000",
  47201=>"111111100",
  47202=>"111111001",
  47203=>"111111000",
  47204=>"101001011",
  47205=>"111111011",
  47206=>"111000000",
  47207=>"111011000",
  47208=>"000111000",
  47209=>"000111111",
  47210=>"000000001",
  47211=>"111111111",
  47212=>"000001011",
  47213=>"000000011",
  47214=>"000000111",
  47215=>"111010000",
  47216=>"000010011",
  47217=>"000001111",
  47218=>"101100100",
  47219=>"111001111",
  47220=>"001011011",
  47221=>"101000000",
  47222=>"000011111",
  47223=>"000000000",
  47224=>"111101001",
  47225=>"000000000",
  47226=>"111000001",
  47227=>"000011111",
  47228=>"000001001",
  47229=>"101001001",
  47230=>"111111000",
  47231=>"011000000",
  47232=>"001000001",
  47233=>"111111111",
  47234=>"011000000",
  47235=>"110101001",
  47236=>"101000000",
  47237=>"000000000",
  47238=>"111111010",
  47239=>"001111110",
  47240=>"111110110",
  47241=>"001001001",
  47242=>"111111000",
  47243=>"011111111",
  47244=>"111100101",
  47245=>"000111111",
  47246=>"011011011",
  47247=>"111111000",
  47248=>"001101100",
  47249=>"000111111",
  47250=>"000000000",
  47251=>"100000000",
  47252=>"000011111",
  47253=>"111111111",
  47254=>"000000000",
  47255=>"001001101",
  47256=>"111111011",
  47257=>"000000110",
  47258=>"111111100",
  47259=>"001111111",
  47260=>"111100111",
  47261=>"011011000",
  47262=>"000000001",
  47263=>"000111000",
  47264=>"000011011",
  47265=>"011111111",
  47266=>"000000100",
  47267=>"000000100",
  47268=>"111111111",
  47269=>"111111000",
  47270=>"111100000",
  47271=>"111110000",
  47272=>"111111001",
  47273=>"101001111",
  47274=>"000000001",
  47275=>"101100000",
  47276=>"100111111",
  47277=>"001000000",
  47278=>"110000000",
  47279=>"000111000",
  47280=>"000111000",
  47281=>"111011000",
  47282=>"100100000",
  47283=>"111111000",
  47284=>"111011000",
  47285=>"100100000",
  47286=>"111111000",
  47287=>"111111111",
  47288=>"111101001",
  47289=>"111010111",
  47290=>"100100100",
  47291=>"110100101",
  47292=>"000111111",
  47293=>"100110111",
  47294=>"000011111",
  47295=>"000000000",
  47296=>"000100101",
  47297=>"000000000",
  47298=>"000000000",
  47299=>"000000000",
  47300=>"000000000",
  47301=>"000000000",
  47302=>"001000000",
  47303=>"100100111",
  47304=>"000000001",
  47305=>"101001111",
  47306=>"111111100",
  47307=>"100000100",
  47308=>"100100011",
  47309=>"000000000",
  47310=>"111101000",
  47311=>"000000000",
  47312=>"011001000",
  47313=>"010001111",
  47314=>"111111111",
  47315=>"000000111",
  47316=>"101101000",
  47317=>"100111111",
  47318=>"001111000",
  47319=>"100000011",
  47320=>"000011111",
  47321=>"111111011",
  47322=>"011111001",
  47323=>"000000000",
  47324=>"111111111",
  47325=>"000100111",
  47326=>"000000001",
  47327=>"001001000",
  47328=>"101111111",
  47329=>"000000000",
  47330=>"111111000",
  47331=>"111100001",
  47332=>"000000000",
  47333=>"111011000",
  47334=>"000111111",
  47335=>"111111100",
  47336=>"000100111",
  47337=>"111111110",
  47338=>"110110000",
  47339=>"001011111",
  47340=>"111111100",
  47341=>"000000011",
  47342=>"111000011",
  47343=>"001101111",
  47344=>"111011111",
  47345=>"111110111",
  47346=>"100111110",
  47347=>"100111110",
  47348=>"001111001",
  47349=>"110110100",
  47350=>"001001001",
  47351=>"110010111",
  47352=>"011111111",
  47353=>"000000000",
  47354=>"111111001",
  47355=>"011011000",
  47356=>"111111100",
  47357=>"000000000",
  47358=>"001000000",
  47359=>"000000000",
  47360=>"000000111",
  47361=>"101111111",
  47362=>"000111111",
  47363=>"001111111",
  47364=>"000000001",
  47365=>"000000001",
  47366=>"001000000",
  47367=>"001101000",
  47368=>"110110111",
  47369=>"111110100",
  47370=>"000111110",
  47371=>"111111111",
  47372=>"110100000",
  47373=>"001000011",
  47374=>"100100000",
  47375=>"011111111",
  47376=>"000010111",
  47377=>"000100101",
  47378=>"001111000",
  47379=>"000000001",
  47380=>"000110111",
  47381=>"111111111",
  47382=>"001011111",
  47383=>"000110111",
  47384=>"111100000",
  47385=>"000101001",
  47386=>"000000000",
  47387=>"011000100",
  47388=>"101000000",
  47389=>"111111111",
  47390=>"000101111",
  47391=>"111111101",
  47392=>"000001001",
  47393=>"000000000",
  47394=>"000000000",
  47395=>"000001001",
  47396=>"110000111",
  47397=>"000100001",
  47398=>"110100100",
  47399=>"000000000",
  47400=>"111111111",
  47401=>"100101000",
  47402=>"000001111",
  47403=>"000000000",
  47404=>"000000110",
  47405=>"110110100",
  47406=>"111110111",
  47407=>"000011111",
  47408=>"100111110",
  47409=>"000000000",
  47410=>"000001101",
  47411=>"000000001",
  47412=>"000000010",
  47413=>"111101111",
  47414=>"111111111",
  47415=>"101101111",
  47416=>"011111000",
  47417=>"000000000",
  47418=>"001111111",
  47419=>"000010000",
  47420=>"100100111",
  47421=>"000101000",
  47422=>"101101101",
  47423=>"110000111",
  47424=>"100000101",
  47425=>"110100000",
  47426=>"000001001",
  47427=>"000000111",
  47428=>"111111001",
  47429=>"100001001",
  47430=>"000000000",
  47431=>"001001000",
  47432=>"111100000",
  47433=>"011001011",
  47434=>"111001111",
  47435=>"001111011",
  47436=>"001001101",
  47437=>"111001000",
  47438=>"111111111",
  47439=>"011001000",
  47440=>"111110100",
  47441=>"011111001",
  47442=>"111000000",
  47443=>"011111111",
  47444=>"100100111",
  47445=>"011001001",
  47446=>"111100001",
  47447=>"111111000",
  47448=>"000110111",
  47449=>"111111111",
  47450=>"111111111",
  47451=>"000010011",
  47452=>"000000011",
  47453=>"111101000",
  47454=>"000011111",
  47455=>"111100000",
  47456=>"000000000",
  47457=>"000110100",
  47458=>"000000000",
  47459=>"001101111",
  47460=>"111101000",
  47461=>"110111111",
  47462=>"100110100",
  47463=>"001110111",
  47464=>"111111110",
  47465=>"000011011",
  47466=>"111000000",
  47467=>"000001001",
  47468=>"111110110",
  47469=>"000000000",
  47470=>"000010110",
  47471=>"100101111",
  47472=>"111000000",
  47473=>"111111111",
  47474=>"000000001",
  47475=>"110100000",
  47476=>"111010111",
  47477=>"000100000",
  47478=>"001000100",
  47479=>"111110010",
  47480=>"111111111",
  47481=>"000000111",
  47482=>"111011000",
  47483=>"000100100",
  47484=>"000000111",
  47485=>"000000000",
  47486=>"111111111",
  47487=>"111111111",
  47488=>"001001101",
  47489=>"111111111",
  47490=>"110010011",
  47491=>"000011111",
  47492=>"001011011",
  47493=>"010010010",
  47494=>"010000000",
  47495=>"000000111",
  47496=>"111111111",
  47497=>"001111111",
  47498=>"000011111",
  47499=>"000011011",
  47500=>"111111111",
  47501=>"100111110",
  47502=>"000111000",
  47503=>"111100000",
  47504=>"000011111",
  47505=>"000010001",
  47506=>"001011011",
  47507=>"000010111",
  47508=>"111111111",
  47509=>"001010000",
  47510=>"101101100",
  47511=>"001001000",
  47512=>"000000001",
  47513=>"111001001",
  47514=>"110111000",
  47515=>"001001111",
  47516=>"101101111",
  47517=>"000000100",
  47518=>"100000000",
  47519=>"011000000",
  47520=>"011000000",
  47521=>"111100100",
  47522=>"000111110",
  47523=>"000000000",
  47524=>"000000001",
  47525=>"000000000",
  47526=>"111111111",
  47527=>"111001011",
  47528=>"011011111",
  47529=>"000011011",
  47530=>"100101111",
  47531=>"001000000",
  47532=>"000000001",
  47533=>"001001000",
  47534=>"111111111",
  47535=>"111111000",
  47536=>"111100000",
  47537=>"000100010",
  47538=>"111011001",
  47539=>"001000000",
  47540=>"000000000",
  47541=>"000000101",
  47542=>"001000100",
  47543=>"001101001",
  47544=>"111111111",
  47545=>"100110111",
  47546=>"101111111",
  47547=>"010000110",
  47548=>"001011000",
  47549=>"000000000",
  47550=>"101111111",
  47551=>"100110101",
  47552=>"100000000",
  47553=>"001001111",
  47554=>"000000010",
  47555=>"011111111",
  47556=>"101101010",
  47557=>"111111001",
  47558=>"111111111",
  47559=>"000000001",
  47560=>"111111111",
  47561=>"111010011",
  47562=>"000000001",
  47563=>"111001001",
  47564=>"000011011",
  47565=>"000000000",
  47566=>"000000000",
  47567=>"000000000",
  47568=>"111110110",
  47569=>"100111111",
  47570=>"111111110",
  47571=>"000001111",
  47572=>"101110000",
  47573=>"111001001",
  47574=>"111011001",
  47575=>"010111011",
  47576=>"101001000",
  47577=>"001000011",
  47578=>"000101111",
  47579=>"111000000",
  47580=>"000000110",
  47581=>"000100100",
  47582=>"111101001",
  47583=>"110110010",
  47584=>"000000110",
  47585=>"010011001",
  47586=>"000100111",
  47587=>"111100100",
  47588=>"000100000",
  47589=>"111111111",
  47590=>"111011000",
  47591=>"000111111",
  47592=>"000000110",
  47593=>"111111111",
  47594=>"001111111",
  47595=>"100100000",
  47596=>"001000111",
  47597=>"111111110",
  47598=>"000000000",
  47599=>"111110110",
  47600=>"000000100",
  47601=>"001001111",
  47602=>"111111000",
  47603=>"000111111",
  47604=>"111100000",
  47605=>"000000111",
  47606=>"000111111",
  47607=>"111111111",
  47608=>"011011111",
  47609=>"000110010",
  47610=>"111001001",
  47611=>"010111111",
  47612=>"000000000",
  47613=>"111111101",
  47614=>"000000000",
  47615=>"111111111",
  47616=>"011001000",
  47617=>"001001000",
  47618=>"001000000",
  47619=>"000000000",
  47620=>"111001000",
  47621=>"111111001",
  47622=>"000000000",
  47623=>"111111111",
  47624=>"000000000",
  47625=>"001001000",
  47626=>"111111111",
  47627=>"110101001",
  47628=>"110010011",
  47629=>"111111111",
  47630=>"000011111",
  47631=>"010010000",
  47632=>"110000111",
  47633=>"110000000",
  47634=>"110111111",
  47635=>"011011111",
  47636=>"000000111",
  47637=>"000011111",
  47638=>"110100100",
  47639=>"100100111",
  47640=>"000100000",
  47641=>"000000110",
  47642=>"000000000",
  47643=>"011001000",
  47644=>"000000000",
  47645=>"111001111",
  47646=>"000011011",
  47647=>"111111000",
  47648=>"011011000",
  47649=>"111111111",
  47650=>"000001111",
  47651=>"111111100",
  47652=>"000000101",
  47653=>"000001000",
  47654=>"111111110",
  47655=>"001111010",
  47656=>"011011000",
  47657=>"000101001",
  47658=>"001001001",
  47659=>"100011001",
  47660=>"000000001",
  47661=>"111111111",
  47662=>"000000100",
  47663=>"000111111",
  47664=>"000000110",
  47665=>"110111111",
  47666=>"100111101",
  47667=>"000000000",
  47668=>"011010110",
  47669=>"111001001",
  47670=>"110101101",
  47671=>"101101011",
  47672=>"000000000",
  47673=>"000000001",
  47674=>"111001100",
  47675=>"000110110",
  47676=>"000000101",
  47677=>"000000000",
  47678=>"000000000",
  47679=>"111111111",
  47680=>"111000000",
  47681=>"001011000",
  47682=>"111111001",
  47683=>"000011111",
  47684=>"111101100",
  47685=>"000000100",
  47686=>"000000000",
  47687=>"111111111",
  47688=>"011000000",
  47689=>"000001001",
  47690=>"111111110",
  47691=>"000000000",
  47692=>"010010000",
  47693=>"110011000",
  47694=>"111100110",
  47695=>"000001001",
  47696=>"000000001",
  47697=>"011111111",
  47698=>"000000000",
  47699=>"011011111",
  47700=>"111000110",
  47701=>"110110110",
  47702=>"011000000",
  47703=>"111101000",
  47704=>"111110111",
  47705=>"000000000",
  47706=>"111000000",
  47707=>"011111011",
  47708=>"000000000",
  47709=>"001001000",
  47710=>"000001000",
  47711=>"111111111",
  47712=>"011001000",
  47713=>"001111111",
  47714=>"000110110",
  47715=>"111111001",
  47716=>"111111110",
  47717=>"000011111",
  47718=>"111101111",
  47719=>"101001001",
  47720=>"000000111",
  47721=>"010000000",
  47722=>"111111111",
  47723=>"111111111",
  47724=>"000001000",
  47725=>"000110111",
  47726=>"001011000",
  47727=>"001001011",
  47728=>"110110000",
  47729=>"001101111",
  47730=>"001001001",
  47731=>"001101111",
  47732=>"101110111",
  47733=>"000000000",
  47734=>"000000001",
  47735=>"000001111",
  47736=>"000000100",
  47737=>"010111111",
  47738=>"100000011",
  47739=>"000100111",
  47740=>"001011011",
  47741=>"110011111",
  47742=>"000000000",
  47743=>"111111000",
  47744=>"001001101",
  47745=>"111000110",
  47746=>"010010000",
  47747=>"111101111",
  47748=>"000100101",
  47749=>"000000000",
  47750=>"011111000",
  47751=>"111111111",
  47752=>"111111100",
  47753=>"000111111",
  47754=>"011011111",
  47755=>"111111000",
  47756=>"000110111",
  47757=>"111111111",
  47758=>"100100011",
  47759=>"110000100",
  47760=>"111100110",
  47761=>"111000000",
  47762=>"001001001",
  47763=>"000000110",
  47764=>"111110100",
  47765=>"110111111",
  47766=>"000001111",
  47767=>"000000000",
  47768=>"000000001",
  47769=>"111111111",
  47770=>"000000000",
  47771=>"000000000",
  47772=>"000010000",
  47773=>"001101101",
  47774=>"111111111",
  47775=>"000110010",
  47776=>"110100110",
  47777=>"011000000",
  47778=>"000000000",
  47779=>"000000000",
  47780=>"101001000",
  47781=>"000000000",
  47782=>"010000000",
  47783=>"111110111",
  47784=>"000000000",
  47785=>"111100100",
  47786=>"111111111",
  47787=>"111010010",
  47788=>"100100100",
  47789=>"110111111",
  47790=>"111000101",
  47791=>"000000111",
  47792=>"000100111",
  47793=>"000000111",
  47794=>"110110110",
  47795=>"000000111",
  47796=>"011011110",
  47797=>"000000111",
  47798=>"000000000",
  47799=>"111111110",
  47800=>"111101000",
  47801=>"111111111",
  47802=>"110000000",
  47803=>"110011001",
  47804=>"000111011",
  47805=>"100100100",
  47806=>"000000000",
  47807=>"000001101",
  47808=>"111111111",
  47809=>"110110000",
  47810=>"111111111",
  47811=>"000000000",
  47812=>"111001001",
  47813=>"000000000",
  47814=>"101011111",
  47815=>"000001000",
  47816=>"000000010",
  47817=>"111001000",
  47818=>"011111001",
  47819=>"010000000",
  47820=>"000000000",
  47821=>"000000000",
  47822=>"000000111",
  47823=>"110000111",
  47824=>"000100000",
  47825=>"001011111",
  47826=>"111111111",
  47827=>"000000000",
  47828=>"111111111",
  47829=>"011001000",
  47830=>"111111111",
  47831=>"000000000",
  47832=>"000000000",
  47833=>"110111111",
  47834=>"011111111",
  47835=>"000000000",
  47836=>"001000100",
  47837=>"001001000",
  47838=>"011000010",
  47839=>"000001000",
  47840=>"011011001",
  47841=>"001000000",
  47842=>"111001111",
  47843=>"110000000",
  47844=>"000000100",
  47845=>"111111010",
  47846=>"110010010",
  47847=>"111111100",
  47848=>"111111111",
  47849=>"000000101",
  47850=>"000000001",
  47851=>"111111111",
  47852=>"111001011",
  47853=>"001001111",
  47854=>"000111111",
  47855=>"111100000",
  47856=>"000000110",
  47857=>"000000000",
  47858=>"111111111",
  47859=>"111001111",
  47860=>"111111110",
  47861=>"111111111",
  47862=>"011011010",
  47863=>"111011111",
  47864=>"111101111",
  47865=>"111111111",
  47866=>"111111011",
  47867=>"000000000",
  47868=>"100111101",
  47869=>"000001000",
  47870=>"110111111",
  47871=>"000000000",
  47872=>"111111111",
  47873=>"001111011",
  47874=>"110110110",
  47875=>"001011000",
  47876=>"001111111",
  47877=>"111000000",
  47878=>"111111111",
  47879=>"000000000",
  47880=>"000101111",
  47881=>"110110111",
  47882=>"010111010",
  47883=>"001111110",
  47884=>"110110100",
  47885=>"111111001",
  47886=>"111111111",
  47887=>"000000000",
  47888=>"000110111",
  47889=>"111000100",
  47890=>"000000000",
  47891=>"011111100",
  47892=>"000100100",
  47893=>"000000000",
  47894=>"110100100",
  47895=>"000001111",
  47896=>"100100110",
  47897=>"000000111",
  47898=>"100000000",
  47899=>"000111010",
  47900=>"100100100",
  47901=>"111010000",
  47902=>"111111111",
  47903=>"111101000",
  47904=>"100000101",
  47905=>"000000000",
  47906=>"111111111",
  47907=>"001000000",
  47908=>"000001011",
  47909=>"100001011",
  47910=>"011111111",
  47911=>"000000000",
  47912=>"111001000",
  47913=>"111110110",
  47914=>"011101100",
  47915=>"111111111",
  47916=>"111111111",
  47917=>"111111101",
  47918=>"111111010",
  47919=>"100100110",
  47920=>"111111111",
  47921=>"100000011",
  47922=>"000101101",
  47923=>"111111111",
  47924=>"010000011",
  47925=>"111101000",
  47926=>"000000001",
  47927=>"000001000",
  47928=>"001000011",
  47929=>"001111111",
  47930=>"000000000",
  47931=>"111100001",
  47932=>"000000000",
  47933=>"100100110",
  47934=>"001101111",
  47935=>"100111110",
  47936=>"000111111",
  47937=>"111111111",
  47938=>"000000100",
  47939=>"000000000",
  47940=>"000100000",
  47941=>"000111111",
  47942=>"110111111",
  47943=>"111111111",
  47944=>"011111111",
  47945=>"000000000",
  47946=>"000001101",
  47947=>"010100110",
  47948=>"111111111",
  47949=>"001011010",
  47950=>"000001011",
  47951=>"110100100",
  47952=>"111111110",
  47953=>"001001100",
  47954=>"111110000",
  47955=>"111111110",
  47956=>"111111001",
  47957=>"000001001",
  47958=>"111110110",
  47959=>"011001111",
  47960=>"111111001",
  47961=>"110111000",
  47962=>"111111111",
  47963=>"001000001",
  47964=>"000100000",
  47965=>"111111111",
  47966=>"011000000",
  47967=>"001001000",
  47968=>"100000000",
  47969=>"111111101",
  47970=>"100000000",
  47971=>"000000000",
  47972=>"110001111",
  47973=>"111111111",
  47974=>"001000000",
  47975=>"000001001",
  47976=>"101001000",
  47977=>"011001000",
  47978=>"000000000",
  47979=>"000000000",
  47980=>"110111111",
  47981=>"111001101",
  47982=>"000000001",
  47983=>"000000111",
  47984=>"001011001",
  47985=>"000000000",
  47986=>"111111111",
  47987=>"000110111",
  47988=>"110110110",
  47989=>"100100100",
  47990=>"110111011",
  47991=>"001011011",
  47992=>"000000000",
  47993=>"000000000",
  47994=>"000000000",
  47995=>"000000000",
  47996=>"100111111",
  47997=>"000011111",
  47998=>"000000000",
  47999=>"000000000",
  48000=>"110111000",
  48001=>"000110000",
  48002=>"100110111",
  48003=>"000010000",
  48004=>"111111010",
  48005=>"111111000",
  48006=>"100110111",
  48007=>"000001111",
  48008=>"111111000",
  48009=>"000000000",
  48010=>"011111011",
  48011=>"000000011",
  48012=>"101101111",
  48013=>"111101100",
  48014=>"011100100",
  48015=>"111111111",
  48016=>"110110110",
  48017=>"111101000",
  48018=>"000101111",
  48019=>"000000101",
  48020=>"000000000",
  48021=>"111010010",
  48022=>"111101101",
  48023=>"101101111",
  48024=>"000000011",
  48025=>"000000000",
  48026=>"000000000",
  48027=>"101111111",
  48028=>"110110010",
  48029=>"110111011",
  48030=>"111110110",
  48031=>"110000011",
  48032=>"000000100",
  48033=>"001111011",
  48034=>"111100100",
  48035=>"100000100",
  48036=>"000100111",
  48037=>"011111011",
  48038=>"111111000",
  48039=>"001111111",
  48040=>"111111001",
  48041=>"000001001",
  48042=>"000000100",
  48043=>"111111111",
  48044=>"000000000",
  48045=>"011111111",
  48046=>"000001111",
  48047=>"011111110",
  48048=>"000000001",
  48049=>"000000000",
  48050=>"111111111",
  48051=>"000001001",
  48052=>"110000000",
  48053=>"000001111",
  48054=>"111111111",
  48055=>"110110000",
  48056=>"000000000",
  48057=>"000000000",
  48058=>"011111111",
  48059=>"110111111",
  48060=>"000000111",
  48061=>"100111111",
  48062=>"110100111",
  48063=>"111001001",
  48064=>"001101111",
  48065=>"111111110",
  48066=>"111111111",
  48067=>"000000000",
  48068=>"111111101",
  48069=>"111110110",
  48070=>"000001100",
  48071=>"111111111",
  48072=>"010000001",
  48073=>"011011001",
  48074=>"001000000",
  48075=>"000000000",
  48076=>"000111111",
  48077=>"000000000",
  48078=>"110110000",
  48079=>"100000011",
  48080=>"001000111",
  48081=>"000001111",
  48082=>"111111111",
  48083=>"000000111",
  48084=>"100111001",
  48085=>"110111111",
  48086=>"001011001",
  48087=>"011000111",
  48088=>"100111111",
  48089=>"010000001",
  48090=>"000100100",
  48091=>"111111111",
  48092=>"000000110",
  48093=>"000100110",
  48094=>"001000000",
  48095=>"111111001",
  48096=>"001000101",
  48097=>"000000000",
  48098=>"000000000",
  48099=>"111111111",
  48100=>"100000100",
  48101=>"000010111",
  48102=>"000000100",
  48103=>"000000111",
  48104=>"100100000",
  48105=>"000000000",
  48106=>"010111111",
  48107=>"111111111",
  48108=>"001001101",
  48109=>"011000111",
  48110=>"011010000",
  48111=>"110000001",
  48112=>"110000110",
  48113=>"111111001",
  48114=>"111101101",
  48115=>"000000000",
  48116=>"101000011",
  48117=>"111011011",
  48118=>"111111111",
  48119=>"110111111",
  48120=>"010000000",
  48121=>"110000100",
  48122=>"100101111",
  48123=>"000000000",
  48124=>"000111000",
  48125=>"000000000",
  48126=>"010000000",
  48127=>"000011111",
  48128=>"000000000",
  48129=>"000000111",
  48130=>"101101000",
  48131=>"111111111",
  48132=>"000000100",
  48133=>"000000000",
  48134=>"100101111",
  48135=>"111001100",
  48136=>"111111001",
  48137=>"111100000",
  48138=>"000011110",
  48139=>"100111111",
  48140=>"000000000",
  48141=>"110111111",
  48142=>"111111000",
  48143=>"000000000",
  48144=>"111111111",
  48145=>"111111110",
  48146=>"111111111",
  48147=>"111001011",
  48148=>"111011111",
  48149=>"111001001",
  48150=>"000000000",
  48151=>"111111110",
  48152=>"111111110",
  48153=>"000110111",
  48154=>"111101000",
  48155=>"010111111",
  48156=>"000100111",
  48157=>"000000111",
  48158=>"011111111",
  48159=>"000000000",
  48160=>"111111011",
  48161=>"111110111",
  48162=>"110110100",
  48163=>"110111000",
  48164=>"000000000",
  48165=>"011111111",
  48166=>"111110000",
  48167=>"111111000",
  48168=>"000000011",
  48169=>"111111000",
  48170=>"001111111",
  48171=>"001010110",
  48172=>"100000000",
  48173=>"110111111",
  48174=>"001111111",
  48175=>"110111110",
  48176=>"000000000",
  48177=>"000000000",
  48178=>"000000010",
  48179=>"111011000",
  48180=>"000111010",
  48181=>"000000100",
  48182=>"001000110",
  48183=>"001110000",
  48184=>"111111000",
  48185=>"000110011",
  48186=>"111111000",
  48187=>"111101000",
  48188=>"111101000",
  48189=>"000000100",
  48190=>"000000000",
  48191=>"001001111",
  48192=>"000010110",
  48193=>"111101000",
  48194=>"101101111",
  48195=>"111110010",
  48196=>"110110111",
  48197=>"000111110",
  48198=>"111011011",
  48199=>"000101100",
  48200=>"000111101",
  48201=>"111000011",
  48202=>"000000000",
  48203=>"101000000",
  48204=>"111010010",
  48205=>"000000001",
  48206=>"000001111",
  48207=>"000010110",
  48208=>"000000011",
  48209=>"000000000",
  48210=>"000000000",
  48211=>"111111000",
  48212=>"000011110",
  48213=>"000000011",
  48214=>"110000000",
  48215=>"000000000",
  48216=>"111111000",
  48217=>"111000000",
  48218=>"000100000",
  48219=>"001011011",
  48220=>"000000111",
  48221=>"111111011",
  48222=>"111010000",
  48223=>"000010010",
  48224=>"010000000",
  48225=>"111111010",
  48226=>"100000000",
  48227=>"000000000",
  48228=>"111111111",
  48229=>"111111000",
  48230=>"000000111",
  48231=>"000000111",
  48232=>"111100111",
  48233=>"111000000",
  48234=>"111000111",
  48235=>"000000000",
  48236=>"000110000",
  48237=>"111111010",
  48238=>"111000001",
  48239=>"000000000",
  48240=>"110111011",
  48241=>"000001101",
  48242=>"111111000",
  48243=>"000000101",
  48244=>"000010110",
  48245=>"111001001",
  48246=>"000000000",
  48247=>"000000000",
  48248=>"100010000",
  48249=>"111111111",
  48250=>"000000000",
  48251=>"000000000",
  48252=>"110111111",
  48253=>"010111111",
  48254=>"111000000",
  48255=>"111111000",
  48256=>"111011000",
  48257=>"101000000",
  48258=>"111111111",
  48259=>"111100001",
  48260=>"100111010",
  48261=>"111101111",
  48262=>"011001111",
  48263=>"000010111",
  48264=>"111111111",
  48265=>"001110110",
  48266=>"111010000",
  48267=>"000000000",
  48268=>"111111000",
  48269=>"111010011",
  48270=>"111111000",
  48271=>"111111110",
  48272=>"000111111",
  48273=>"000111111",
  48274=>"000000000",
  48275=>"010000110",
  48276=>"110110000",
  48277=>"000000111",
  48278=>"111000000",
  48279=>"000000000",
  48280=>"111101000",
  48281=>"000000000",
  48282=>"000000100",
  48283=>"101000001",
  48284=>"000110010",
  48285=>"000000111",
  48286=>"111111111",
  48287=>"000000000",
  48288=>"000000000",
  48289=>"011011111",
  48290=>"000000010",
  48291=>"000111111",
  48292=>"100111100",
  48293=>"111111000",
  48294=>"111111000",
  48295=>"010111111",
  48296=>"011010110",
  48297=>"110010000",
  48298=>"101101000",
  48299=>"000011111",
  48300=>"000110111",
  48301=>"000000100",
  48302=>"000000110",
  48303=>"000000000",
  48304=>"111111111",
  48305=>"110111010",
  48306=>"110111111",
  48307=>"100100000",
  48308=>"000111101",
  48309=>"000000100",
  48310=>"000110000",
  48311=>"011111110",
  48312=>"000000100",
  48313=>"100111111",
  48314=>"000000111",
  48315=>"000010010",
  48316=>"001000000",
  48317=>"111110111",
  48318=>"111000111",
  48319=>"111111100",
  48320=>"000000010",
  48321=>"001000000",
  48322=>"001111111",
  48323=>"100101001",
  48324=>"111001000",
  48325=>"101111011",
  48326=>"001000111",
  48327=>"000000000",
  48328=>"111111000",
  48329=>"000000110",
  48330=>"001111110",
  48331=>"000000111",
  48332=>"111111010",
  48333=>"110110010",
  48334=>"100110111",
  48335=>"000011111",
  48336=>"111100110",
  48337=>"000100000",
  48338=>"001000111",
  48339=>"000000100",
  48340=>"000010000",
  48341=>"110111111",
  48342=>"101101001",
  48343=>"011011111",
  48344=>"000110110",
  48345=>"111111111",
  48346=>"111111111",
  48347=>"111101000",
  48348=>"000000010",
  48349=>"111111001",
  48350=>"100110000",
  48351=>"000110000",
  48352=>"001001011",
  48353=>"001001000",
  48354=>"000000011",
  48355=>"000000000",
  48356=>"111000111",
  48357=>"000000110",
  48358=>"111111111",
  48359=>"000000111",
  48360=>"111011111",
  48361=>"111111111",
  48362=>"111011000",
  48363=>"111000000",
  48364=>"000101111",
  48365=>"000111101",
  48366=>"101111111",
  48367=>"001000000",
  48368=>"100110000",
  48369=>"011011010",
  48370=>"111000111",
  48371=>"010111001",
  48372=>"000000011",
  48373=>"001001001",
  48374=>"000000000",
  48375=>"000000011",
  48376=>"001111110",
  48377=>"000010111",
  48378=>"001111011",
  48379=>"110111111",
  48380=>"001011000",
  48381=>"011011011",
  48382=>"000000110",
  48383=>"000000000",
  48384=>"000000000",
  48385=>"001001001",
  48386=>"111111100",
  48387=>"110110000",
  48388=>"000000001",
  48389=>"001001111",
  48390=>"000000000",
  48391=>"000110111",
  48392=>"110110010",
  48393=>"000000000",
  48394=>"000000010",
  48395=>"111111000",
  48396=>"111111111",
  48397=>"000011001",
  48398=>"111110000",
  48399=>"000000001",
  48400=>"000001101",
  48401=>"001010111",
  48402=>"000001000",
  48403=>"000000000",
  48404=>"011111111",
  48405=>"101100000",
  48406=>"000000111",
  48407=>"000110111",
  48408=>"011011010",
  48409=>"111111011",
  48410=>"101111100",
  48411=>"011011001",
  48412=>"011011100",
  48413=>"100010000",
  48414=>"111111111",
  48415=>"111011111",
  48416=>"101101000",
  48417=>"001001110",
  48418=>"111011001",
  48419=>"000001001",
  48420=>"111111000",
  48421=>"110110000",
  48422=>"000000011",
  48423=>"001001100",
  48424=>"000000000",
  48425=>"010110010",
  48426=>"010011100",
  48427=>"000101000",
  48428=>"001111111",
  48429=>"010010110",
  48430=>"111111000",
  48431=>"000000000",
  48432=>"111111111",
  48433=>"110100010",
  48434=>"111111110",
  48435=>"111111000",
  48436=>"011001000",
  48437=>"000111111",
  48438=>"000010000",
  48439=>"001000000",
  48440=>"000000000",
  48441=>"101000111",
  48442=>"011111100",
  48443=>"101000001",
  48444=>"000100110",
  48445=>"110111111",
  48446=>"000110110",
  48447=>"000000000",
  48448=>"111111000",
  48449=>"111111000",
  48450=>"000010000",
  48451=>"001000001",
  48452=>"111111111",
  48453=>"111011011",
  48454=>"000000111",
  48455=>"100100111",
  48456=>"000111111",
  48457=>"000000010",
  48458=>"111111100",
  48459=>"110110010",
  48460=>"000100100",
  48461=>"111000000",
  48462=>"100110100",
  48463=>"011011011",
  48464=>"000100110",
  48465=>"000000000",
  48466=>"000010110",
  48467=>"001000001",
  48468=>"100101111",
  48469=>"011011011",
  48470=>"000010111",
  48471=>"111111111",
  48472=>"000001000",
  48473=>"111101000",
  48474=>"111111111",
  48475=>"111111001",
  48476=>"111000000",
  48477=>"011011111",
  48478=>"000001011",
  48479=>"011000000",
  48480=>"000001000",
  48481=>"000000000",
  48482=>"010011011",
  48483=>"101000000",
  48484=>"000000101",
  48485=>"000000000",
  48486=>"100100111",
  48487=>"000100100",
  48488=>"000111110",
  48489=>"110111111",
  48490=>"001111111",
  48491=>"101001001",
  48492=>"000000100",
  48493=>"000000000",
  48494=>"000000000",
  48495=>"000000000",
  48496=>"000110010",
  48497=>"111111000",
  48498=>"100111111",
  48499=>"000111111",
  48500=>"101111001",
  48501=>"000000000",
  48502=>"100111000",
  48503=>"100000000",
  48504=>"111111111",
  48505=>"111111111",
  48506=>"000000110",
  48507=>"000110010",
  48508=>"111111000",
  48509=>"111110100",
  48510=>"101101000",
  48511=>"000000000",
  48512=>"111101000",
  48513=>"111111000",
  48514=>"000111111",
  48515=>"111000001",
  48516=>"000000000",
  48517=>"111111001",
  48518=>"111111111",
  48519=>"100000111",
  48520=>"111111000",
  48521=>"000100100",
  48522=>"110000000",
  48523=>"001001111",
  48524=>"000111111",
  48525=>"000110110",
  48526=>"111111001",
  48527=>"000000000",
  48528=>"000000000",
  48529=>"110110110",
  48530=>"111111001",
  48531=>"000001001",
  48532=>"000101111",
  48533=>"000111000",
  48534=>"000110000",
  48535=>"000111000",
  48536=>"110000000",
  48537=>"000100110",
  48538=>"111111111",
  48539=>"111111001",
  48540=>"100000000",
  48541=>"000011111",
  48542=>"000110111",
  48543=>"010000000",
  48544=>"000000000",
  48545=>"111100100",
  48546=>"111111111",
  48547=>"010110101",
  48548=>"111111111",
  48549=>"000111000",
  48550=>"011000000",
  48551=>"000000111",
  48552=>"000000000",
  48553=>"000000000",
  48554=>"000000000",
  48555=>"000010110",
  48556=>"000000000",
  48557=>"000000001",
  48558=>"000000001",
  48559=>"000000110",
  48560=>"000000000",
  48561=>"001101111",
  48562=>"000000111",
  48563=>"000000110",
  48564=>"111110111",
  48565=>"111111000",
  48566=>"111111110",
  48567=>"000100111",
  48568=>"111000000",
  48569=>"100000000",
  48570=>"000111111",
  48571=>"010111111",
  48572=>"001000111",
  48573=>"111011000",
  48574=>"111001000",
  48575=>"000110110",
  48576=>"000000110",
  48577=>"111101111",
  48578=>"111101111",
  48579=>"001001000",
  48580=>"000000001",
  48581=>"000000000",
  48582=>"110110000",
  48583=>"110100100",
  48584=>"000110100",
  48585=>"000010000",
  48586=>"000000000",
  48587=>"000000000",
  48588=>"111000011",
  48589=>"000000100",
  48590=>"111111110",
  48591=>"000000001",
  48592=>"000101111",
  48593=>"110110011",
  48594=>"000000001",
  48595=>"111000000",
  48596=>"000100110",
  48597=>"000000101",
  48598=>"100110000",
  48599=>"000001011",
  48600=>"001111111",
  48601=>"000000000",
  48602=>"111111000",
  48603=>"111010010",
  48604=>"000110111",
  48605=>"111111000",
  48606=>"111111110",
  48607=>"000111011",
  48608=>"100100101",
  48609=>"000000000",
  48610=>"111111000",
  48611=>"000000100",
  48612=>"110111111",
  48613=>"001001000",
  48614=>"111111111",
  48615=>"101111111",
  48616=>"001000000",
  48617=>"000000000",
  48618=>"000111111",
  48619=>"111111010",
  48620=>"111111111",
  48621=>"000010000",
  48622=>"111101000",
  48623=>"100110010",
  48624=>"000110110",
  48625=>"000000010",
  48626=>"000100111",
  48627=>"000001001",
  48628=>"000000100",
  48629=>"011011001",
  48630=>"100110110",
  48631=>"111111001",
  48632=>"111111110",
  48633=>"100000000",
  48634=>"111001001",
  48635=>"110111000",
  48636=>"001111111",
  48637=>"101000000",
  48638=>"000000111",
  48639=>"000000111",
  48640=>"000111000",
  48641=>"111111000",
  48642=>"001000111",
  48643=>"000100100",
  48644=>"110111111",
  48645=>"111111011",
  48646=>"110111000",
  48647=>"111000000",
  48648=>"000000100",
  48649=>"100111110",
  48650=>"011001001",
  48651=>"110111111",
  48652=>"011111110",
  48653=>"101001011",
  48654=>"001010000",
  48655=>"110110010",
  48656=>"000000001",
  48657=>"000011111",
  48658=>"000000000",
  48659=>"000000000",
  48660=>"111111111",
  48661=>"111111111",
  48662=>"000000000",
  48663=>"110110111",
  48664=>"000001011",
  48665=>"000101001",
  48666=>"111111111",
  48667=>"011100001",
  48668=>"000000001",
  48669=>"000110010",
  48670=>"111011111",
  48671=>"111111000",
  48672=>"001001000",
  48673=>"000111010",
  48674=>"000000111",
  48675=>"111111110",
  48676=>"000000100",
  48677=>"011111101",
  48678=>"000000001",
  48679=>"000110000",
  48680=>"000000001",
  48681=>"001000000",
  48682=>"111111111",
  48683=>"101000000",
  48684=>"101101111",
  48685=>"110011111",
  48686=>"111111111",
  48687=>"001000100",
  48688=>"111111110",
  48689=>"001001100",
  48690=>"000000100",
  48691=>"001010000",
  48692=>"100001000",
  48693=>"100110000",
  48694=>"000000000",
  48695=>"110110111",
  48696=>"111110111",
  48697=>"000000110",
  48698=>"111101111",
  48699=>"000000011",
  48700=>"001000000",
  48701=>"000000111",
  48702=>"111111011",
  48703=>"111011000",
  48704=>"000000000",
  48705=>"011110110",
  48706=>"000000111",
  48707=>"110111000",
  48708=>"001000000",
  48709=>"111001001",
  48710=>"100101111",
  48711=>"111111111",
  48712=>"000000000",
  48713=>"001100110",
  48714=>"111111111",
  48715=>"000000111",
  48716=>"011011111",
  48717=>"111100100",
  48718=>"111111011",
  48719=>"000000000",
  48720=>"111011011",
  48721=>"000000000",
  48722=>"111011001",
  48723=>"000000000",
  48724=>"000110000",
  48725=>"101000000",
  48726=>"001001101",
  48727=>"000000111",
  48728=>"001111111",
  48729=>"010100100",
  48730=>"001001000",
  48731=>"111111101",
  48732=>"000000000",
  48733=>"110110110",
  48734=>"111111111",
  48735=>"111111101",
  48736=>"010010000",
  48737=>"111011111",
  48738=>"000000100",
  48739=>"001001001",
  48740=>"000000000",
  48741=>"111101111",
  48742=>"100100101",
  48743=>"100110110",
  48744=>"000010000",
  48745=>"000000111",
  48746=>"101000000",
  48747=>"000001100",
  48748=>"110110100",
  48749=>"111111111",
  48750=>"001101001",
  48751=>"000000000",
  48752=>"001001110",
  48753=>"000000100",
  48754=>"000000000",
  48755=>"111001001",
  48756=>"111011000",
  48757=>"110110000",
  48758=>"000000111",
  48759=>"000000000",
  48760=>"110110110",
  48761=>"001001101",
  48762=>"010000000",
  48763=>"100001001",
  48764=>"100110111",
  48765=>"101111001",
  48766=>"110010000",
  48767=>"000000000",
  48768=>"001000111",
  48769=>"111101111",
  48770=>"100000100",
  48771=>"011001001",
  48772=>"000000111",
  48773=>"101000000",
  48774=>"000000000",
  48775=>"000111111",
  48776=>"000000111",
  48777=>"000000000",
  48778=>"010001111",
  48779=>"110101000",
  48780=>"011010110",
  48781=>"110111010",
  48782=>"110110010",
  48783=>"001011000",
  48784=>"111101111",
  48785=>"011011011",
  48786=>"000000000",
  48787=>"011011011",
  48788=>"001000000",
  48789=>"110110000",
  48790=>"111101111",
  48791=>"001101000",
  48792=>"000000000",
  48793=>"111111110",
  48794=>"001101111",
  48795=>"111111111",
  48796=>"100000011",
  48797=>"000111111",
  48798=>"111001001",
  48799=>"111111111",
  48800=>"101000001",
  48801=>"110000000",
  48802=>"111111111",
  48803=>"111111001",
  48804=>"000000000",
  48805=>"110000000",
  48806=>"001000101",
  48807=>"010001000",
  48808=>"111111111",
  48809=>"010111110",
  48810=>"111100000",
  48811=>"110010100",
  48812=>"111000000",
  48813=>"110111000",
  48814=>"111011000",
  48815=>"000000011",
  48816=>"110010000",
  48817=>"000000000",
  48818=>"110110111",
  48819=>"000000001",
  48820=>"001011000",
  48821=>"111101111",
  48822=>"110111010",
  48823=>"011111001",
  48824=>"111100110",
  48825=>"001000000",
  48826=>"000001001",
  48827=>"110110000",
  48828=>"001000111",
  48829=>"001001001",
  48830=>"001000100",
  48831=>"001110111",
  48832=>"000000000",
  48833=>"111001111",
  48834=>"000011111",
  48835=>"000000001",
  48836=>"001001111",
  48837=>"110111111",
  48838=>"101000000",
  48839=>"000000001",
  48840=>"110110000",
  48841=>"000010111",
  48842=>"111111111",
  48843=>"000000000",
  48844=>"111001000",
  48845=>"110111000",
  48846=>"101110110",
  48847=>"010111111",
  48848=>"000000000",
  48849=>"111011110",
  48850=>"010000000",
  48851=>"111111111",
  48852=>"111011111",
  48853=>"111111111",
  48854=>"000000000",
  48855=>"001000101",
  48856=>"111111001",
  48857=>"000111001",
  48858=>"111110111",
  48859=>"000000000",
  48860=>"001001000",
  48861=>"111111111",
  48862=>"111111110",
  48863=>"000000011",
  48864=>"000000000",
  48865=>"000000001",
  48866=>"000100000",
  48867=>"001000011",
  48868=>"010110011",
  48869=>"100001001",
  48870=>"000110110",
  48871=>"010111011",
  48872=>"110110110",
  48873=>"000000000",
  48874=>"100110111",
  48875=>"000000101",
  48876=>"000000000",
  48877=>"000000110",
  48878=>"000110111",
  48879=>"000111111",
  48880=>"110110111",
  48881=>"111111111",
  48882=>"111111111",
  48883=>"000000110",
  48884=>"110110000",
  48885=>"100110000",
  48886=>"000011111",
  48887=>"111111000",
  48888=>"000000111",
  48889=>"110111000",
  48890=>"000000000",
  48891=>"111110110",
  48892=>"011001001",
  48893=>"010001001",
  48894=>"010000000",
  48895=>"110110000",
  48896=>"001000110",
  48897=>"110110110",
  48898=>"001000000",
  48899=>"000000111",
  48900=>"001111111",
  48901=>"000010011",
  48902=>"111110100",
  48903=>"110110110",
  48904=>"011000110",
  48905=>"011011011",
  48906=>"000000100",
  48907=>"000100111",
  48908=>"111111111",
  48909=>"000000000",
  48910=>"111111000",
  48911=>"000010000",
  48912=>"110110111",
  48913=>"110110111",
  48914=>"101001111",
  48915=>"000000000",
  48916=>"000000000",
  48917=>"000000011",
  48918=>"011110001",
  48919=>"110000000",
  48920=>"110111000",
  48921=>"111111000",
  48922=>"110100111",
  48923=>"000000001",
  48924=>"100110110",
  48925=>"111111111",
  48926=>"111111111",
  48927=>"110111011",
  48928=>"000000110",
  48929=>"000001111",
  48930=>"111111111",
  48931=>"111111111",
  48932=>"001000101",
  48933=>"111111111",
  48934=>"001111111",
  48935=>"111010111",
  48936=>"001101110",
  48937=>"000000000",
  48938=>"000110111",
  48939=>"011001101",
  48940=>"111110000",
  48941=>"000000000",
  48942=>"000000011",
  48943=>"000110010",
  48944=>"111111011",
  48945=>"110111111",
  48946=>"000000000",
  48947=>"000000000",
  48948=>"000101111",
  48949=>"011111011",
  48950=>"111111100",
  48951=>"000000011",
  48952=>"000000111",
  48953=>"111111111",
  48954=>"000110111",
  48955=>"111101111",
  48956=>"001001011",
  48957=>"111110000",
  48958=>"000110111",
  48959=>"010110000",
  48960=>"000001001",
  48961=>"000011001",
  48962=>"000000101",
  48963=>"001000110",
  48964=>"110000010",
  48965=>"001000000",
  48966=>"111111000",
  48967=>"111000000",
  48968=>"110100000",
  48969=>"000010111",
  48970=>"001011001",
  48971=>"000000000",
  48972=>"110000000",
  48973=>"001001001",
  48974=>"101001011",
  48975=>"001001010",
  48976=>"110111010",
  48977=>"011000100",
  48978=>"110011111",
  48979=>"000000100",
  48980=>"000100000",
  48981=>"011011011",
  48982=>"000000001",
  48983=>"001000000",
  48984=>"110110000",
  48985=>"111100000",
  48986=>"111011110",
  48987=>"011111100",
  48988=>"101111111",
  48989=>"111000001",
  48990=>"000110111",
  48991=>"111011011",
  48992=>"000001001",
  48993=>"111111110",
  48994=>"111111011",
  48995=>"000000000",
  48996=>"000000100",
  48997=>"000001001",
  48998=>"100110111",
  48999=>"000000000",
  49000=>"000000000",
  49001=>"000000110",
  49002=>"000000000",
  49003=>"000011011",
  49004=>"000000000",
  49005=>"000000000",
  49006=>"110111110",
  49007=>"000000000",
  49008=>"001001111",
  49009=>"000000000",
  49010=>"000001000",
  49011=>"011111011",
  49012=>"111111001",
  49013=>"111110100",
  49014=>"000000000",
  49015=>"000000111",
  49016=>"000000111",
  49017=>"111111010",
  49018=>"000000000",
  49019=>"110110000",
  49020=>"111010000",
  49021=>"000000000",
  49022=>"110111111",
  49023=>"010000100",
  49024=>"000000000",
  49025=>"110000000",
  49026=>"111111100",
  49027=>"001000111",
  49028=>"101111111",
  49029=>"100111111",
  49030=>"000100000",
  49031=>"111011000",
  49032=>"001000111",
  49033=>"101100000",
  49034=>"001000000",
  49035=>"111111111",
  49036=>"111000101",
  49037=>"001001001",
  49038=>"000000001",
  49039=>"001001111",
  49040=>"000000000",
  49041=>"110110110",
  49042=>"011010010",
  49043=>"110110100",
  49044=>"000100000",
  49045=>"000000000",
  49046=>"011011001",
  49047=>"011001000",
  49048=>"000001111",
  49049=>"100010010",
  49050=>"111111111",
  49051=>"001001000",
  49052=>"111100111",
  49053=>"110110000",
  49054=>"000000000",
  49055=>"000000111",
  49056=>"000000000",
  49057=>"001011000",
  49058=>"110011111",
  49059=>"100110110",
  49060=>"000000111",
  49061=>"000010010",
  49062=>"010000000",
  49063=>"100110100",
  49064=>"011011010",
  49065=>"110110101",
  49066=>"000010111",
  49067=>"000000001",
  49068=>"000000000",
  49069=>"000000000",
  49070=>"100110000",
  49071=>"100000100",
  49072=>"111111111",
  49073=>"111000000",
  49074=>"110111111",
  49075=>"001111111",
  49076=>"000000111",
  49077=>"111101110",
  49078=>"001110100",
  49079=>"111111111",
  49080=>"001000100",
  49081=>"000000010",
  49082=>"100000001",
  49083=>"100000000",
  49084=>"110010000",
  49085=>"110110111",
  49086=>"000000111",
  49087=>"000000000",
  49088=>"010110111",
  49089=>"001000101",
  49090=>"010011011",
  49091=>"110110110",
  49092=>"000011111",
  49093=>"000000011",
  49094=>"000000001",
  49095=>"001011000",
  49096=>"010000000",
  49097=>"000000000",
  49098=>"001001000",
  49099=>"111011010",
  49100=>"111010000",
  49101=>"110110000",
  49102=>"000000000",
  49103=>"100101000",
  49104=>"000000000",
  49105=>"111010011",
  49106=>"000111001",
  49107=>"111101111",
  49108=>"110110111",
  49109=>"111111000",
  49110=>"111111010",
  49111=>"001000001",
  49112=>"001000000",
  49113=>"111111011",
  49114=>"000000111",
  49115=>"111111111",
  49116=>"000011000",
  49117=>"000000000",
  49118=>"110110111",
  49119=>"000000000",
  49120=>"001011011",
  49121=>"100111111",
  49122=>"000111111",
  49123=>"000001000",
  49124=>"100111111",
  49125=>"111000000",
  49126=>"100000000",
  49127=>"111101111",
  49128=>"110111011",
  49129=>"000010000",
  49130=>"010101110",
  49131=>"000000011",
  49132=>"001001001",
  49133=>"000000000",
  49134=>"000000000",
  49135=>"110111111",
  49136=>"000000000",
  49137=>"110111011",
  49138=>"000011110",
  49139=>"110000110",
  49140=>"011110000",
  49141=>"110111000",
  49142=>"011001001",
  49143=>"100000000",
  49144=>"000110100",
  49145=>"000000000",
  49146=>"111111111",
  49147=>"111111111",
  49148=>"111000000",
  49149=>"001000000",
  49150=>"111011000",
  49151=>"000000010",
  49152=>"010010100",
  49153=>"100100100",
  49154=>"000000111",
  49155=>"110111111",
  49156=>"000000000",
  49157=>"111111111",
  49158=>"101101001",
  49159=>"000000000",
  49160=>"110000000",
  49161=>"111110110",
  49162=>"111100000",
  49163=>"001000000",
  49164=>"001000000",
  49165=>"011000000",
  49166=>"110111011",
  49167=>"000000000",
  49168=>"000100100",
  49169=>"000000101",
  49170=>"111111111",
  49171=>"000000000",
  49172=>"111111111",
  49173=>"001001111",
  49174=>"111111111",
  49175=>"111111110",
  49176=>"111111111",
  49177=>"011011001",
  49178=>"111000000",
  49179=>"100101111",
  49180=>"000000000",
  49181=>"110110111",
  49182=>"111111111",
  49183=>"101101101",
  49184=>"000110110",
  49185=>"111111000",
  49186=>"111111001",
  49187=>"110111111",
  49188=>"000000100",
  49189=>"110000000",
  49190=>"001111111",
  49191=>"000000000",
  49192=>"000100111",
  49193=>"111100000",
  49194=>"111111111",
  49195=>"000000000",
  49196=>"110111111",
  49197=>"000000000",
  49198=>"111111111",
  49199=>"000000000",
  49200=>"000000001",
  49201=>"000000000",
  49202=>"100000100",
  49203=>"001000000",
  49204=>"010011011",
  49205=>"110110110",
  49206=>"000000000",
  49207=>"111111111",
  49208=>"000000000",
  49209=>"010010000",
  49210=>"000000000",
  49211=>"000000000",
  49212=>"000000110",
  49213=>"000010000",
  49214=>"000001001",
  49215=>"000000000",
  49216=>"111111111",
  49217=>"101101101",
  49218=>"111111111",
  49219=>"111111111",
  49220=>"111111111",
  49221=>"011000000",
  49222=>"111111011",
  49223=>"000000000",
  49224=>"001000000",
  49225=>"000000000",
  49226=>"100000110",
  49227=>"110110111",
  49228=>"100100111",
  49229=>"011000000",
  49230=>"110111111",
  49231=>"000110111",
  49232=>"000000001",
  49233=>"111111110",
  49234=>"111111111",
  49235=>"110110100",
  49236=>"011011111",
  49237=>"111011000",
  49238=>"001011000",
  49239=>"000000100",
  49240=>"100110100",
  49241=>"111111111",
  49242=>"111111111",
  49243=>"111111011",
  49244=>"100000001",
  49245=>"000000000",
  49246=>"010001011",
  49247=>"110100000",
  49248=>"111011111",
  49249=>"000000011",
  49250=>"101100111",
  49251=>"111111010",
  49252=>"000000000",
  49253=>"111111111",
  49254=>"000010001",
  49255=>"100111101",
  49256=>"000000000",
  49257=>"011111111",
  49258=>"000100000",
  49259=>"000000000",
  49260=>"111111011",
  49261=>"000000000",
  49262=>"000000110",
  49263=>"110111111",
  49264=>"011011001",
  49265=>"111101101",
  49266=>"000001111",
  49267=>"000000000",
  49268=>"000000000",
  49269=>"000000000",
  49270=>"111111111",
  49271=>"000010000",
  49272=>"000100111",
  49273=>"000000000",
  49274=>"111001000",
  49275=>"000000000",
  49276=>"110110100",
  49277=>"000000000",
  49278=>"101011001",
  49279=>"111111011",
  49280=>"000000110",
  49281=>"000000111",
  49282=>"000100110",
  49283=>"000011011",
  49284=>"001101000",
  49285=>"000000000",
  49286=>"111110000",
  49287=>"000111111",
  49288=>"111111100",
  49289=>"000010110",
  49290=>"000011000",
  49291=>"111000101",
  49292=>"001101100",
  49293=>"111111110",
  49294=>"101100100",
  49295=>"011011000",
  49296=>"000000000",
  49297=>"111111000",
  49298=>"000001001",
  49299=>"111111011",
  49300=>"000111001",
  49301=>"111111000",
  49302=>"100000000",
  49303=>"100110100",
  49304=>"001001001",
  49305=>"111111111",
  49306=>"111101000",
  49307=>"100001001",
  49308=>"000000000",
  49309=>"001000001",
  49310=>"001010111",
  49311=>"111111111",
  49312=>"111111011",
  49313=>"111111111",
  49314=>"000000000",
  49315=>"000000000",
  49316=>"011010110",
  49317=>"000000110",
  49318=>"000000101",
  49319=>"001001001",
  49320=>"010010000",
  49321=>"111111111",
  49322=>"100110110",
  49323=>"111011011",
  49324=>"001000000",
  49325=>"110000001",
  49326=>"110111100",
  49327=>"001111111",
  49328=>"000000000",
  49329=>"000000010",
  49330=>"111111111",
  49331=>"000000000",
  49332=>"111001000",
  49333=>"111000100",
  49334=>"001000111",
  49335=>"111111111",
  49336=>"111011011",
  49337=>"100000000",
  49338=>"001000000",
  49339=>"111111000",
  49340=>"000000110",
  49341=>"000000101",
  49342=>"000000000",
  49343=>"000000000",
  49344=>"001001110",
  49345=>"000000000",
  49346=>"111111110",
  49347=>"111100111",
  49348=>"000001011",
  49349=>"111111001",
  49350=>"100000001",
  49351=>"000000000",
  49352=>"000000000",
  49353=>"111110111",
  49354=>"000000001",
  49355=>"000111110",
  49356=>"011011011",
  49357=>"001011111",
  49358=>"000011011",
  49359=>"011111011",
  49360=>"111010010",
  49361=>"000101000",
  49362=>"000010011",
  49363=>"111101111",
  49364=>"000000000",
  49365=>"000001001",
  49366=>"111100000",
  49367=>"100111111",
  49368=>"000000000",
  49369=>"000000000",
  49370=>"000000000",
  49371=>"001000000",
  49372=>"000000000",
  49373=>"001000000",
  49374=>"000000000",
  49375=>"111100001",
  49376=>"000000100",
  49377=>"111111111",
  49378=>"111100000",
  49379=>"000000000",
  49380=>"000000000",
  49381=>"110110000",
  49382=>"000000001",
  49383=>"000000111",
  49384=>"111111111",
  49385=>"111111111",
  49386=>"111110000",
  49387=>"111111101",
  49388=>"000000000",
  49389=>"000000000",
  49390=>"111111111",
  49391=>"111111111",
  49392=>"000010000",
  49393=>"000000000",
  49394=>"111000000",
  49395=>"000000100",
  49396=>"111100000",
  49397=>"111011010",
  49398=>"000011011",
  49399=>"111111110",
  49400=>"111111000",
  49401=>"000000000",
  49402=>"111111000",
  49403=>"000000000",
  49404=>"101111111",
  49405=>"000000001",
  49406=>"011111111",
  49407=>"100100111",
  49408=>"000001001",
  49409=>"111111111",
  49410=>"010111111",
  49411=>"011111000",
  49412=>"001101110",
  49413=>"100100110",
  49414=>"101110111",
  49415=>"111111111",
  49416=>"111111011",
  49417=>"000000000",
  49418=>"000011111",
  49419=>"000000000",
  49420=>"011111011",
  49421=>"111111100",
  49422=>"101001110",
  49423=>"000100000",
  49424=>"000000001",
  49425=>"001001000",
  49426=>"111000000",
  49427=>"000110111",
  49428=>"000000000",
  49429=>"000000000",
  49430=>"000000000",
  49431=>"000000000",
  49432=>"010111011",
  49433=>"110111111",
  49434=>"011011011",
  49435=>"001111111",
  49436=>"000010100",
  49437=>"111111000",
  49438=>"111111111",
  49439=>"111100010",
  49440=>"010011000",
  49441=>"000101111",
  49442=>"011000000",
  49443=>"111111111",
  49444=>"110010000",
  49445=>"001111111",
  49446=>"011000000",
  49447=>"000011011",
  49448=>"111111111",
  49449=>"111111010",
  49450=>"001000111",
  49451=>"111111111",
  49452=>"100110111",
  49453=>"110110111",
  49454=>"000001000",
  49455=>"000000000",
  49456=>"110110101",
  49457=>"000000000",
  49458=>"000000000",
  49459=>"000000000",
  49460=>"000000000",
  49461=>"001001001",
  49462=>"111110111",
  49463=>"001111111",
  49464=>"000000000",
  49465=>"000000000",
  49466=>"001000000",
  49467=>"100000100",
  49468=>"110111111",
  49469=>"101000000",
  49470=>"000000000",
  49471=>"000100000",
  49472=>"101101101",
  49473=>"011000000",
  49474=>"111111000",
  49475=>"110111111",
  49476=>"111110001",
  49477=>"000000000",
  49478=>"000000000",
  49479=>"101000000",
  49480=>"000000000",
  49481=>"000000000",
  49482=>"001100110",
  49483=>"110110100",
  49484=>"000011011",
  49485=>"100000000",
  49486=>"011000000",
  49487=>"111011001",
  49488=>"111100000",
  49489=>"000000100",
  49490=>"100100000",
  49491=>"011000000",
  49492=>"111111111",
  49493=>"011000001",
  49494=>"000000101",
  49495=>"001000000",
  49496=>"100100000",
  49497=>"111111111",
  49498=>"000011010",
  49499=>"110000001",
  49500=>"000000111",
  49501=>"000000000",
  49502=>"111110110",
  49503=>"111111111",
  49504=>"000110100",
  49505=>"111111111",
  49506=>"011001001",
  49507=>"111111111",
  49508=>"111111111",
  49509=>"011011011",
  49510=>"000000000",
  49511=>"000000000",
  49512=>"011111111",
  49513=>"001101110",
  49514=>"111111010",
  49515=>"110110111",
  49516=>"111111111",
  49517=>"001000011",
  49518=>"101101000",
  49519=>"000000000",
  49520=>"000000000",
  49521=>"110111000",
  49522=>"001100000",
  49523=>"011111111",
  49524=>"111111111",
  49525=>"000100111",
  49526=>"111011101",
  49527=>"000000000",
  49528=>"000110111",
  49529=>"001000010",
  49530=>"110010000",
  49531=>"111111011",
  49532=>"000000000",
  49533=>"010000000",
  49534=>"000000111",
  49535=>"111111111",
  49536=>"000111111",
  49537=>"110110111",
  49538=>"111111100",
  49539=>"111111111",
  49540=>"111111001",
  49541=>"100100000",
  49542=>"100000001",
  49543=>"101100100",
  49544=>"111111010",
  49545=>"111111111",
  49546=>"111001001",
  49547=>"100100100",
  49548=>"000000000",
  49549=>"000011011",
  49550=>"111111111",
  49551=>"000000000",
  49552=>"000000000",
  49553=>"100110111",
  49554=>"000000001",
  49555=>"111111111",
  49556=>"000000000",
  49557=>"000000000",
  49558=>"000000000",
  49559=>"111110000",
  49560=>"000000000",
  49561=>"000000011",
  49562=>"001001111",
  49563=>"100110000",
  49564=>"111111001",
  49565=>"111111111",
  49566=>"000000011",
  49567=>"000000000",
  49568=>"000000001",
  49569=>"100000000",
  49570=>"011110100",
  49571=>"111111101",
  49572=>"000110100",
  49573=>"000001001",
  49574=>"111110000",
  49575=>"000000000",
  49576=>"111111111",
  49577=>"111100100",
  49578=>"100100000",
  49579=>"000000000",
  49580=>"111100000",
  49581=>"111111001",
  49582=>"100101011",
  49583=>"111010000",
  49584=>"111010001",
  49585=>"000001000",
  49586=>"100000000",
  49587=>"000000000",
  49588=>"000000000",
  49589=>"111000000",
  49590=>"111111111",
  49591=>"111111111",
  49592=>"011111011",
  49593=>"101110000",
  49594=>"000111011",
  49595=>"111000000",
  49596=>"000000000",
  49597=>"000000100",
  49598=>"000000001",
  49599=>"111111111",
  49600=>"111111111",
  49601=>"000000000",
  49602=>"000000000",
  49603=>"111111111",
  49604=>"000000000",
  49605=>"000010111",
  49606=>"111111001",
  49607=>"100000001",
  49608=>"001001000",
  49609=>"111111111",
  49610=>"111100101",
  49611=>"111111100",
  49612=>"001001011",
  49613=>"000000000",
  49614=>"111111111",
  49615=>"010110111",
  49616=>"100110100",
  49617=>"011111111",
  49618=>"111110100",
  49619=>"000000000",
  49620=>"100000000",
  49621=>"000000000",
  49622=>"000000000",
  49623=>"100000100",
  49624=>"111111111",
  49625=>"111111010",
  49626=>"111000000",
  49627=>"000000000",
  49628=>"111111101",
  49629=>"111110100",
  49630=>"111111100",
  49631=>"111001001",
  49632=>"111111111",
  49633=>"110000000",
  49634=>"111111111",
  49635=>"111111111",
  49636=>"110111111",
  49637=>"101111111",
  49638=>"011001000",
  49639=>"100000110",
  49640=>"000110111",
  49641=>"111111111",
  49642=>"011000000",
  49643=>"000000000",
  49644=>"000000000",
  49645=>"001100100",
  49646=>"111111101",
  49647=>"000001001",
  49648=>"000000011",
  49649=>"111111111",
  49650=>"111111111",
  49651=>"100111111",
  49652=>"000110111",
  49653=>"111111111",
  49654=>"011111011",
  49655=>"011011111",
  49656=>"111111111",
  49657=>"010011001",
  49658=>"000000100",
  49659=>"000000000",
  49660=>"001000110",
  49661=>"011000000",
  49662=>"111111111",
  49663=>"000000010",
  49664=>"011001000",
  49665=>"111111111",
  49666=>"000000000",
  49667=>"111111111",
  49668=>"111000001",
  49669=>"111000000",
  49670=>"011000011",
  49671=>"111111111",
  49672=>"001111111",
  49673=>"111000000",
  49674=>"111000000",
  49675=>"000000000",
  49676=>"111111101",
  49677=>"000000100",
  49678=>"000000001",
  49679=>"000000001",
  49680=>"111001000",
  49681=>"110101000",
  49682=>"100000000",
  49683=>"111111111",
  49684=>"000011000",
  49685=>"100110100",
  49686=>"111111111",
  49687=>"111111111",
  49688=>"001111111",
  49689=>"111111111",
  49690=>"111111111",
  49691=>"110100001",
  49692=>"011111111",
  49693=>"111101101",
  49694=>"000001011",
  49695=>"000000000",
  49696=>"110110000",
  49697=>"000100111",
  49698=>"111111111",
  49699=>"000000000",
  49700=>"010000100",
  49701=>"001111111",
  49702=>"100100000",
  49703=>"000000010",
  49704=>"111111000",
  49705=>"000000000",
  49706=>"000111111",
  49707=>"000000000",
  49708=>"000000000",
  49709=>"111111111",
  49710=>"001001111",
  49711=>"000011000",
  49712=>"000000000",
  49713=>"111111111",
  49714=>"001001111",
  49715=>"000000000",
  49716=>"100100100",
  49717=>"001001101",
  49718=>"010011111",
  49719=>"110100000",
  49720=>"000000000",
  49721=>"101000000",
  49722=>"000010000",
  49723=>"000000000",
  49724=>"100100111",
  49725=>"001001000",
  49726=>"101111111",
  49727=>"011111111",
  49728=>"111101111",
  49729=>"000000000",
  49730=>"000000001",
  49731=>"000010000",
  49732=>"001000000",
  49733=>"111111111",
  49734=>"000000100",
  49735=>"100000000",
  49736=>"111111111",
  49737=>"100000000",
  49738=>"000000000",
  49739=>"000000000",
  49740=>"111111111",
  49741=>"111111111",
  49742=>"000000100",
  49743=>"000000000",
  49744=>"100100111",
  49745=>"100100101",
  49746=>"000100000",
  49747=>"000000000",
  49748=>"111100101",
  49749=>"000011111",
  49750=>"000010010",
  49751=>"000000000",
  49752=>"110100000",
  49753=>"000000000",
  49754=>"111111111",
  49755=>"001001001",
  49756=>"111111111",
  49757=>"000000000",
  49758=>"111111111",
  49759=>"100100100",
  49760=>"001000100",
  49761=>"100110111",
  49762=>"111110100",
  49763=>"000000000",
  49764=>"000000111",
  49765=>"000001001",
  49766=>"100100000",
  49767=>"000000000",
  49768=>"111111111",
  49769=>"000000111",
  49770=>"000000111",
  49771=>"111111110",
  49772=>"111111111",
  49773=>"000110110",
  49774=>"000000000",
  49775=>"000100100",
  49776=>"000001001",
  49777=>"010000100",
  49778=>"100101111",
  49779=>"000111111",
  49780=>"111111100",
  49781=>"000001011",
  49782=>"001000000",
  49783=>"111111111",
  49784=>"111011111",
  49785=>"000101001",
  49786=>"000000000",
  49787=>"111111111",
  49788=>"001001011",
  49789=>"000010010",
  49790=>"010110110",
  49791=>"000111110",
  49792=>"000000000",
  49793=>"000000000",
  49794=>"001001000",
  49795=>"000001111",
  49796=>"000000000",
  49797=>"000000000",
  49798=>"100110111",
  49799=>"101100100",
  49800=>"000000000",
  49801=>"111111111",
  49802=>"000000101",
  49803=>"011011001",
  49804=>"111111111",
  49805=>"111111111",
  49806=>"101101101",
  49807=>"111111111",
  49808=>"011111111",
  49809=>"111101100",
  49810=>"111101000",
  49811=>"000010111",
  49812=>"000010010",
  49813=>"000000000",
  49814=>"111111111",
  49815=>"000001001",
  49816=>"111110000",
  49817=>"010000000",
  49818=>"111101000",
  49819=>"111101101",
  49820=>"100101100",
  49821=>"111111111",
  49822=>"010010000",
  49823=>"000000000",
  49824=>"000000000",
  49825=>"000000000",
  49826=>"111111111",
  49827=>"100100101",
  49828=>"011001111",
  49829=>"011011011",
  49830=>"101000111",
  49831=>"100100110",
  49832=>"111000000",
  49833=>"011011000",
  49834=>"000000000",
  49835=>"111101101",
  49836=>"001100000",
  49837=>"111111000",
  49838=>"111111111",
  49839=>"000011000",
  49840=>"000000000",
  49841=>"101111111",
  49842=>"111110111",
  49843=>"000000100",
  49844=>"010011011",
  49845=>"011011001",
  49846=>"111010000",
  49847=>"001001101",
  49848=>"001011111",
  49849=>"100000000",
  49850=>"111000111",
  49851=>"111110000",
  49852=>"000111111",
  49853=>"000010111",
  49854=>"000000000",
  49855=>"111011000",
  49856=>"000000110",
  49857=>"001010000",
  49858=>"111110000",
  49859=>"000000000",
  49860=>"111111111",
  49861=>"000000000",
  49862=>"111000000",
  49863=>"111011000",
  49864=>"111111110",
  49865=>"100111111",
  49866=>"010110000",
  49867=>"000001101",
  49868=>"001111100",
  49869=>"000000000",
  49870=>"000000000",
  49871=>"000001111",
  49872=>"111001000",
  49873=>"111111100",
  49874=>"111000000",
  49875=>"000110000",
  49876=>"111111111",
  49877=>"000000000",
  49878=>"110000000",
  49879=>"011111000",
  49880=>"111111100",
  49881=>"000000110",
  49882=>"000000100",
  49883=>"111111111",
  49884=>"100111000",
  49885=>"110111111",
  49886=>"000001111",
  49887=>"000000010",
  49888=>"111001001",
  49889=>"100000000",
  49890=>"000000000",
  49891=>"011000000",
  49892=>"111011011",
  49893=>"100110100",
  49894=>"000111111",
  49895=>"111111110",
  49896=>"111111100",
  49897=>"110010111",
  49898=>"011111101",
  49899=>"001011110",
  49900=>"111011000",
  49901=>"000000000",
  49902=>"111001000",
  49903=>"000000000",
  49904=>"011111111",
  49905=>"111101111",
  49906=>"111000000",
  49907=>"000000111",
  49908=>"011111111",
  49909=>"111000100",
  49910=>"111111001",
  49911=>"000000110",
  49912=>"000010000",
  49913=>"000000000",
  49914=>"000000000",
  49915=>"111111111",
  49916=>"001111111",
  49917=>"011000110",
  49918=>"111111111",
  49919=>"010110100",
  49920=>"000000011",
  49921=>"111011000",
  49922=>"111111111",
  49923=>"000000101",
  49924=>"000000111",
  49925=>"000011011",
  49926=>"000000000",
  49927=>"010010011",
  49928=>"100100000",
  49929=>"111111111",
  49930=>"111000000",
  49931=>"111001011",
  49932=>"111111101",
  49933=>"111111111",
  49934=>"000010011",
  49935=>"100001111",
  49936=>"000001001",
  49937=>"110000000",
  49938=>"111111111",
  49939=>"011001111",
  49940=>"011111111",
  49941=>"111111111",
  49942=>"111011110",
  49943=>"111110000",
  49944=>"001001111",
  49945=>"011000000",
  49946=>"000111111",
  49947=>"011110000",
  49948=>"101101111",
  49949=>"000000000",
  49950=>"010010010",
  49951=>"110000000",
  49952=>"001001001",
  49953=>"110110011",
  49954=>"011011111",
  49955=>"000010000",
  49956=>"011001001",
  49957=>"110110000",
  49958=>"111111011",
  49959=>"011000011",
  49960=>"111100100",
  49961=>"111111111",
  49962=>"111101000",
  49963=>"111111000",
  49964=>"000100111",
  49965=>"110110111",
  49966=>"000101111",
  49967=>"110110111",
  49968=>"111111101",
  49969=>"000011111",
  49970=>"000000000",
  49971=>"001000000",
  49972=>"111111111",
  49973=>"111111000",
  49974=>"111111000",
  49975=>"010011011",
  49976=>"100000111",
  49977=>"010111111",
  49978=>"110110000",
  49979=>"000001111",
  49980=>"000000000",
  49981=>"000000111",
  49982=>"011001111",
  49983=>"000011011",
  49984=>"000000111",
  49985=>"010011111",
  49986=>"111111111",
  49987=>"000100000",
  49988=>"110111000",
  49989=>"000000000",
  49990=>"000000000",
  49991=>"111111111",
  49992=>"000100110",
  49993=>"001000000",
  49994=>"001001010",
  49995=>"011110100",
  49996=>"000000000",
  49997=>"111111111",
  49998=>"000000000",
  49999=>"000001001",
  50000=>"011011011",
  50001=>"011010010",
  50002=>"000100000",
  50003=>"100100001",
  50004=>"000000100",
  50005=>"010011010",
  50006=>"111110000",
  50007=>"111111111",
  50008=>"111111111",
  50009=>"111000100",
  50010=>"101001111",
  50011=>"001101110",
  50012=>"000000000",
  50013=>"111111110",
  50014=>"000000000",
  50015=>"110100000",
  50016=>"100111111",
  50017=>"101101100",
  50018=>"100100100",
  50019=>"000000110",
  50020=>"000000100",
  50021=>"000000000",
  50022=>"100100000",
  50023=>"110000000",
  50024=>"110010001",
  50025=>"101111101",
  50026=>"101100111",
  50027=>"111111111",
  50028=>"111111111",
  50029=>"010000001",
  50030=>"000000000",
  50031=>"000000101",
  50032=>"111111111",
  50033=>"111001000",
  50034=>"000100100",
  50035=>"110100111",
  50036=>"000000000",
  50037=>"011010111",
  50038=>"111001001",
  50039=>"100110100",
  50040=>"111111111",
  50041=>"001110000",
  50042=>"100100111",
  50043=>"111001001",
  50044=>"000000000",
  50045=>"000001011",
  50046=>"000000000",
  50047=>"111110000",
  50048=>"100110110",
  50049=>"111111101",
  50050=>"111111111",
  50051=>"000000000",
  50052=>"000000000",
  50053=>"000000000",
  50054=>"111111111",
  50055=>"001001001",
  50056=>"111101111",
  50057=>"110110111",
  50058=>"101100100",
  50059=>"010010010",
  50060=>"111111111",
  50061=>"100110111",
  50062=>"010000000",
  50063=>"100111000",
  50064=>"001000000",
  50065=>"000000000",
  50066=>"000000000",
  50067=>"001000001",
  50068=>"111111111",
  50069=>"111001000",
  50070=>"010000010",
  50071=>"011001111",
  50072=>"111001000",
  50073=>"111111000",
  50074=>"000100000",
  50075=>"110110111",
  50076=>"000000111",
  50077=>"001000001",
  50078=>"000000111",
  50079=>"000000000",
  50080=>"000011001",
  50081=>"001001111",
  50082=>"001110110",
  50083=>"011011101",
  50084=>"000000010",
  50085=>"101000001",
  50086=>"111111111",
  50087=>"111110100",
  50088=>"111110100",
  50089=>"000000000",
  50090=>"111000000",
  50091=>"111111111",
  50092=>"000010000",
  50093=>"000000000",
  50094=>"000000000",
  50095=>"111011011",
  50096=>"111100111",
  50097=>"000000000",
  50098=>"001000110",
  50099=>"000110110",
  50100=>"111101100",
  50101=>"011011010",
  50102=>"110110010",
  50103=>"000000111",
  50104=>"000110111",
  50105=>"111111111",
  50106=>"101101101",
  50107=>"000000000",
  50108=>"011111110",
  50109=>"000110110",
  50110=>"111110110",
  50111=>"111011011",
  50112=>"000111110",
  50113=>"100111111",
  50114=>"000000000",
  50115=>"100000000",
  50116=>"000000110",
  50117=>"011001001",
  50118=>"001111111",
  50119=>"111111000",
  50120=>"111111111",
  50121=>"000000010",
  50122=>"000000000",
  50123=>"111110000",
  50124=>"000000111",
  50125=>"001111101",
  50126=>"001111101",
  50127=>"001000010",
  50128=>"001001111",
  50129=>"111110000",
  50130=>"000000000",
  50131=>"000000001",
  50132=>"001011001",
  50133=>"111111111",
  50134=>"111111110",
  50135=>"101001011",
  50136=>"001000111",
  50137=>"111001001",
  50138=>"111000000",
  50139=>"011011000",
  50140=>"111100101",
  50141=>"000010110",
  50142=>"000000100",
  50143=>"011011011",
  50144=>"111111111",
  50145=>"100100100",
  50146=>"011001111",
  50147=>"100110110",
  50148=>"000000000",
  50149=>"110111001",
  50150=>"000100100",
  50151=>"000000000",
  50152=>"000110010",
  50153=>"000000000",
  50154=>"001011000",
  50155=>"000000111",
  50156=>"011111111",
  50157=>"000000001",
  50158=>"101111111",
  50159=>"111111100",
  50160=>"111110111",
  50161=>"000000000",
  50162=>"111111111",
  50163=>"000001001",
  50164=>"000100100",
  50165=>"000000111",
  50166=>"000000000",
  50167=>"011001101",
  50168=>"110111111",
  50169=>"011111111",
  50170=>"000000000",
  50171=>"000000000",
  50172=>"001110110",
  50173=>"001001000",
  50174=>"001001100",
  50175=>"110111111",
  50176=>"001111000",
  50177=>"111111100",
  50178=>"000000101",
  50179=>"111111111",
  50180=>"111111111",
  50181=>"011011000",
  50182=>"000000000",
  50183=>"111111001",
  50184=>"111001001",
  50185=>"111111111",
  50186=>"000000000",
  50187=>"111110111",
  50188=>"010000000",
  50189=>"100000000",
  50190=>"000000000",
  50191=>"000000000",
  50192=>"000000100",
  50193=>"111111111",
  50194=>"111111111",
  50195=>"000000000",
  50196=>"000000000",
  50197=>"000000000",
  50198=>"000000000",
  50199=>"000001000",
  50200=>"011111101",
  50201=>"110101000",
  50202=>"111111011",
  50203=>"000111111",
  50204=>"101001001",
  50205=>"000000000",
  50206=>"001001001",
  50207=>"111111001",
  50208=>"111111110",
  50209=>"000000011",
  50210=>"111111111",
  50211=>"000000000",
  50212=>"011000110",
  50213=>"111111111",
  50214=>"000000000",
  50215=>"111000000",
  50216=>"111110000",
  50217=>"000000000",
  50218=>"110100000",
  50219=>"111110111",
  50220=>"000000000",
  50221=>"000000001",
  50222=>"000000000",
  50223=>"000000000",
  50224=>"001001100",
  50225=>"000000000",
  50226=>"011011000",
  50227=>"011000000",
  50228=>"100100000",
  50229=>"011111111",
  50230=>"100100000",
  50231=>"011111100",
  50232=>"011011000",
  50233=>"000111111",
  50234=>"111111111",
  50235=>"000000000",
  50236=>"000000000",
  50237=>"111111111",
  50238=>"100011111",
  50239=>"000111111",
  50240=>"111111111",
  50241=>"111010000",
  50242=>"111010010",
  50243=>"111011111",
  50244=>"000000111",
  50245=>"111110110",
  50246=>"000000000",
  50247=>"000000011",
  50248=>"011011000",
  50249=>"000001111",
  50250=>"111111010",
  50251=>"011000011",
  50252=>"000000000",
  50253=>"100111111",
  50254=>"001111111",
  50255=>"100111111",
  50256=>"111111110",
  50257=>"000000100",
  50258=>"100000000",
  50259=>"001001010",
  50260=>"111111111",
  50261=>"110111111",
  50262=>"111111100",
  50263=>"000000101",
  50264=>"100101101",
  50265=>"001000111",
  50266=>"011000000",
  50267=>"111011000",
  50268=>"010000000",
  50269=>"011011111",
  50270=>"000000000",
  50271=>"000000000",
  50272=>"000111111",
  50273=>"111111111",
  50274=>"100100000",
  50275=>"000000000",
  50276=>"111111000",
  50277=>"000010011",
  50278=>"111111000",
  50279=>"111111111",
  50280=>"000000111",
  50281=>"011111111",
  50282=>"011011010",
  50283=>"101111000",
  50284=>"000110110",
  50285=>"111110111",
  50286=>"111000000",
  50287=>"100100111",
  50288=>"111111000",
  50289=>"111111111",
  50290=>"001011000",
  50291=>"000000000",
  50292=>"101000111",
  50293=>"011111110",
  50294=>"011000000",
  50295=>"000000000",
  50296=>"000000000",
  50297=>"000000111",
  50298=>"111111111",
  50299=>"111111111",
  50300=>"000000000",
  50301=>"000000011",
  50302=>"100000000",
  50303=>"000000000",
  50304=>"000000000",
  50305=>"111111000",
  50306=>"000000000",
  50307=>"000110010",
  50308=>"100111111",
  50309=>"110111000",
  50310=>"001000000",
  50311=>"111001000",
  50312=>"111111111",
  50313=>"010000000",
  50314=>"000000111",
  50315=>"000010111",
  50316=>"111111111",
  50317=>"111111111",
  50318=>"000001101",
  50319=>"001000111",
  50320=>"111111000",
  50321=>"000000000",
  50322=>"100000000",
  50323=>"000000001",
  50324=>"111001000",
  50325=>"110111101",
  50326=>"111111111",
  50327=>"000000001",
  50328=>"010000000",
  50329=>"111111111",
  50330=>"001000000",
  50331=>"111111000",
  50332=>"001001100",
  50333=>"111101000",
  50334=>"001000100",
  50335=>"111111111",
  50336=>"000010111",
  50337=>"001111111",
  50338=>"111111111",
  50339=>"111000000",
  50340=>"101000100",
  50341=>"000000000",
  50342=>"111111111",
  50343=>"110100110",
  50344=>"111111111",
  50345=>"110111000",
  50346=>"111111111",
  50347=>"111111111",
  50348=>"111111000",
  50349=>"101001001",
  50350=>"000100011",
  50351=>"000000000",
  50352=>"011011000",
  50353=>"011110100",
  50354=>"110010010",
  50355=>"111111111",
  50356=>"000000000",
  50357=>"111111110",
  50358=>"111100110",
  50359=>"000000000",
  50360=>"011000000",
  50361=>"001000000",
  50362=>"110000000",
  50363=>"011001000",
  50364=>"000000010",
  50365=>"111011000",
  50366=>"111111111",
  50367=>"111111010",
  50368=>"111111010",
  50369=>"000000000",
  50370=>"010011011",
  50371=>"000111111",
  50372=>"101001001",
  50373=>"110000000",
  50374=>"111111000",
  50375=>"001001111",
  50376=>"111111111",
  50377=>"000000000",
  50378=>"000000000",
  50379=>"111000000",
  50380=>"000100111",
  50381=>"000000000",
  50382=>"110111011",
  50383=>"111111110",
  50384=>"111011000",
  50385=>"000000000",
  50386=>"111111111",
  50387=>"000000000",
  50388=>"111111000",
  50389=>"000000000",
  50390=>"000000000",
  50391=>"010111111",
  50392=>"111111110",
  50393=>"010010011",
  50394=>"000000011",
  50395=>"000000000",
  50396=>"000000111",
  50397=>"000000000",
  50398=>"000000000",
  50399=>"111100000",
  50400=>"111111111",
  50401=>"111111111",
  50402=>"111111000",
  50403=>"011111111",
  50404=>"000000000",
  50405=>"110100100",
  50406=>"000010010",
  50407=>"111111111",
  50408=>"000000011",
  50409=>"000000101",
  50410=>"110101101",
  50411=>"000100110",
  50412=>"000110100",
  50413=>"000000000",
  50414=>"000111111",
  50415=>"011011111",
  50416=>"000000000",
  50417=>"011010000",
  50418=>"111111111",
  50419=>"000000111",
  50420=>"011000000",
  50421=>"111111111",
  50422=>"111111111",
  50423=>"000000000",
  50424=>"001110000",
  50425=>"111111111",
  50426=>"000010011",
  50427=>"111111111",
  50428=>"000000000",
  50429=>"000000000",
  50430=>"011111001",
  50431=>"111111111",
  50432=>"000000000",
  50433=>"000000000",
  50434=>"000000000",
  50435=>"000000000",
  50436=>"000000000",
  50437=>"111001000",
  50438=>"000000000",
  50439=>"011000000",
  50440=>"111111111",
  50441=>"111111111",
  50442=>"110100000",
  50443=>"000011011",
  50444=>"101001001",
  50445=>"001010111",
  50446=>"111111001",
  50447=>"111111111",
  50448=>"000000000",
  50449=>"111111111",
  50450=>"000000000",
  50451=>"000000111",
  50452=>"000000000",
  50453=>"000000001",
  50454=>"000100110",
  50455=>"000000100",
  50456=>"000000111",
  50457=>"011010110",
  50458=>"011011111",
  50459=>"111111111",
  50460=>"110110111",
  50461=>"111000000",
  50462=>"111111111",
  50463=>"100000000",
  50464=>"000110000",
  50465=>"111111111",
  50466=>"111111010",
  50467=>"110111111",
  50468=>"000100100",
  50469=>"011000000",
  50470=>"111101111",
  50471=>"000000000",
  50472=>"000000000",
  50473=>"000000000",
  50474=>"011100111",
  50475=>"000110111",
  50476=>"000000111",
  50477=>"000110000",
  50478=>"111111000",
  50479=>"000000000",
  50480=>"000110100",
  50481=>"111111111",
  50482=>"000111110",
  50483=>"111111111",
  50484=>"000000000",
  50485=>"111111000",
  50486=>"111000011",
  50487=>"000000111",
  50488=>"000000111",
  50489=>"000000011",
  50490=>"111011011",
  50491=>"111010010",
  50492=>"110110110",
  50493=>"000000001",
  50494=>"111100001",
  50495=>"110110111",
  50496=>"000111101",
  50497=>"110110111",
  50498=>"011111111",
  50499=>"111000000",
  50500=>"001000010",
  50501=>"111111111",
  50502=>"000000000",
  50503=>"111111111",
  50504=>"111110111",
  50505=>"000111111",
  50506=>"111111011",
  50507=>"000001010",
  50508=>"000000010",
  50509=>"111100110",
  50510=>"110100101",
  50511=>"000000000",
  50512=>"111110110",
  50513=>"111100000",
  50514=>"010011010",
  50515=>"100111110",
  50516=>"000110111",
  50517=>"000000000",
  50518=>"001001000",
  50519=>"000000000",
  50520=>"111111111",
  50521=>"000000000",
  50522=>"001000000",
  50523=>"111111000",
  50524=>"111111111",
  50525=>"101000100",
  50526=>"111111111",
  50527=>"110111101",
  50528=>"000001000",
  50529=>"000000000",
  50530=>"010111100",
  50531=>"111111111",
  50532=>"000000000",
  50533=>"000010000",
  50534=>"000000011",
  50535=>"000111111",
  50536=>"101111101",
  50537=>"000110111",
  50538=>"100000000",
  50539=>"000000000",
  50540=>"011111111",
  50541=>"111111101",
  50542=>"000000000",
  50543=>"111000000",
  50544=>"000000000",
  50545=>"111111111",
  50546=>"000000100",
  50547=>"111111111",
  50548=>"001000000",
  50549=>"000000000",
  50550=>"111111111",
  50551=>"111111111",
  50552=>"011111111",
  50553=>"111000000",
  50554=>"000000000",
  50555=>"000000000",
  50556=>"111000000",
  50557=>"000100111",
  50558=>"111111111",
  50559=>"010010011",
  50560=>"100000000",
  50561=>"100100100",
  50562=>"000000000",
  50563=>"000000000",
  50564=>"000000000",
  50565=>"000000110",
  50566=>"011111111",
  50567=>"000000000",
  50568=>"000001000",
  50569=>"011010111",
  50570=>"111111001",
  50571=>"010011000",
  50572=>"001001001",
  50573=>"111111000",
  50574=>"111111001",
  50575=>"000000000",
  50576=>"111111111",
  50577=>"000000000",
  50578=>"110010000",
  50579=>"111111111",
  50580=>"000000000",
  50581=>"000000000",
  50582=>"001000001",
  50583=>"000000100",
  50584=>"000001111",
  50585=>"101000000",
  50586=>"000000000",
  50587=>"101111111",
  50588=>"111111111",
  50589=>"000100100",
  50590=>"000000000",
  50591=>"000100110",
  50592=>"111111100",
  50593=>"110100000",
  50594=>"000110110",
  50595=>"011011101",
  50596=>"010110000",
  50597=>"000000000",
  50598=>"111010000",
  50599=>"111111111",
  50600=>"010000000",
  50601=>"011111111",
  50602=>"001000000",
  50603=>"000100111",
  50604=>"000000000",
  50605=>"000000001",
  50606=>"111111100",
  50607=>"111111111",
  50608=>"000000000",
  50609=>"111111110",
  50610=>"111000000",
  50611=>"000010000",
  50612=>"011111011",
  50613=>"111011111",
  50614=>"001100111",
  50615=>"111000110",
  50616=>"010001111",
  50617=>"000011111",
  50618=>"000111111",
  50619=>"000000111",
  50620=>"000111111",
  50621=>"000000000",
  50622=>"100111111",
  50623=>"000000000",
  50624=>"000110110",
  50625=>"111011001",
  50626=>"111111111",
  50627=>"000000000",
  50628=>"111111111",
  50629=>"011011000",
  50630=>"011011111",
  50631=>"000000001",
  50632=>"111000000",
  50633=>"100100000",
  50634=>"111111111",
  50635=>"111111111",
  50636=>"001111111",
  50637=>"000000000",
  50638=>"000000000",
  50639=>"100100101",
  50640=>"000001001",
  50641=>"011011010",
  50642=>"110110000",
  50643=>"111111110",
  50644=>"110110110",
  50645=>"001111111",
  50646=>"000100110",
  50647=>"001001011",
  50648=>"000000000",
  50649=>"111111111",
  50650=>"000000000",
  50651=>"101111001",
  50652=>"011000000",
  50653=>"111111111",
  50654=>"000000000",
  50655=>"000011000",
  50656=>"011011111",
  50657=>"000000000",
  50658=>"110111110",
  50659=>"010000000",
  50660=>"001011010",
  50661=>"001000000",
  50662=>"000000000",
  50663=>"110111111",
  50664=>"111111111",
  50665=>"111111010",
  50666=>"000000000",
  50667=>"000100110",
  50668=>"000001000",
  50669=>"011000000",
  50670=>"000000000",
  50671=>"110111110",
  50672=>"111011011",
  50673=>"111001100",
  50674=>"000000110",
  50675=>"011011000",
  50676=>"010000001",
  50677=>"100100000",
  50678=>"111111111",
  50679=>"001111111",
  50680=>"000000000",
  50681=>"000100100",
  50682=>"110111111",
  50683=>"110110110",
  50684=>"111111000",
  50685=>"100000111",
  50686=>"000000110",
  50687=>"000000000",
  50688=>"110100100",
  50689=>"110111011",
  50690=>"111111111",
  50691=>"000000000",
  50692=>"110110111",
  50693=>"110000110",
  50694=>"000000000",
  50695=>"101111111",
  50696=>"101001001",
  50697=>"000000000",
  50698=>"110011000",
  50699=>"000011111",
  50700=>"000000000",
  50701=>"100100110",
  50702=>"000000000",
  50703=>"000000000",
  50704=>"100000001",
  50705=>"000001000",
  50706=>"111111111",
  50707=>"100111111",
  50708=>"111111111",
  50709=>"000000000",
  50710=>"000000100",
  50711=>"111111111",
  50712=>"000100100",
  50713=>"111111001",
  50714=>"000001001",
  50715=>"011111111",
  50716=>"111111111",
  50717=>"011111101",
  50718=>"111111111",
  50719=>"111111111",
  50720=>"100100111",
  50721=>"111111111",
  50722=>"110000111",
  50723=>"111111111",
  50724=>"000000000",
  50725=>"111111101",
  50726=>"010000000",
  50727=>"111111110",
  50728=>"001111111",
  50729=>"010000000",
  50730=>"011111001",
  50731=>"111111111",
  50732=>"111111111",
  50733=>"011000000",
  50734=>"111111111",
  50735=>"100000000",
  50736=>"011011000",
  50737=>"011000001",
  50738=>"001000000",
  50739=>"111100100",
  50740=>"001111111",
  50741=>"000000000",
  50742=>"110000000",
  50743=>"000111011",
  50744=>"000000000",
  50745=>"101110111",
  50746=>"000001001",
  50747=>"111111111",
  50748=>"111000000",
  50749=>"000000000",
  50750=>"000000100",
  50751=>"010010111",
  50752=>"000101111",
  50753=>"000000000",
  50754=>"111111111",
  50755=>"110111111",
  50756=>"000000000",
  50757=>"110010000",
  50758=>"000011111",
  50759=>"000000000",
  50760=>"011001000",
  50761=>"000000000",
  50762=>"100100000",
  50763=>"000000000",
  50764=>"111111000",
  50765=>"111111111",
  50766=>"001110111",
  50767=>"111111111",
  50768=>"000000000",
  50769=>"111000000",
  50770=>"111111111",
  50771=>"100010011",
  50772=>"000011011",
  50773=>"111111000",
  50774=>"001001001",
  50775=>"000100100",
  50776=>"000000001",
  50777=>"000000000",
  50778=>"111111111",
  50779=>"011001000",
  50780=>"111001001",
  50781=>"111111010",
  50782=>"000000000",
  50783=>"111111111",
  50784=>"111001000",
  50785=>"111111111",
  50786=>"000000000",
  50787=>"000000010",
  50788=>"100000000",
  50789=>"000000000",
  50790=>"110001011",
  50791=>"000101111",
  50792=>"011111000",
  50793=>"111111111",
  50794=>"111100000",
  50795=>"111111011",
  50796=>"001011111",
  50797=>"000000000",
  50798=>"100111110",
  50799=>"000000000",
  50800=>"000000000",
  50801=>"000000100",
  50802=>"100000000",
  50803=>"111101100",
  50804=>"000000001",
  50805=>"110110110",
  50806=>"000000000",
  50807=>"111111111",
  50808=>"100100000",
  50809=>"000000000",
  50810=>"111111111",
  50811=>"111111111",
  50812=>"000000000",
  50813=>"111111111",
  50814=>"111111111",
  50815=>"010010010",
  50816=>"001011000",
  50817=>"110111111",
  50818=>"110111111",
  50819=>"011000000",
  50820=>"000000001",
  50821=>"100000000",
  50822=>"000110000",
  50823=>"111111111",
  50824=>"000000100",
  50825=>"000000000",
  50826=>"111111101",
  50827=>"111111111",
  50828=>"000000000",
  50829=>"000000101",
  50830=>"111111100",
  50831=>"000000000",
  50832=>"111101111",
  50833=>"000010000",
  50834=>"000000000",
  50835=>"000111111",
  50836=>"111110100",
  50837=>"000001011",
  50838=>"011001111",
  50839=>"000000000",
  50840=>"010010111",
  50841=>"000001001",
  50842=>"000000011",
  50843=>"001011000",
  50844=>"000000001",
  50845=>"000000000",
  50846=>"111111111",
  50847=>"000000000",
  50848=>"111111111",
  50849=>"001000000",
  50850=>"000000000",
  50851=>"000000000",
  50852=>"111000000",
  50853=>"010100101",
  50854=>"111111111",
  50855=>"111111110",
  50856=>"000001111",
  50857=>"100000000",
  50858=>"110100100",
  50859=>"000000111",
  50860=>"011011111",
  50861=>"111111111",
  50862=>"101101000",
  50863=>"000011011",
  50864=>"000000000",
  50865=>"111111111",
  50866=>"111010010",
  50867=>"111111000",
  50868=>"000000000",
  50869=>"110111111",
  50870=>"110110010",
  50871=>"001100111",
  50872=>"100000001",
  50873=>"000000000",
  50874=>"111110111",
  50875=>"111011111",
  50876=>"101101111",
  50877=>"000000110",
  50878=>"111111111",
  50879=>"111000000",
  50880=>"111110010",
  50881=>"000000000",
  50882=>"100000000",
  50883=>"111111000",
  50884=>"111111000",
  50885=>"111100000",
  50886=>"011011000",
  50887=>"111111011",
  50888=>"100000000",
  50889=>"001000000",
  50890=>"001000000",
  50891=>"111000100",
  50892=>"000100111",
  50893=>"000000000",
  50894=>"000001111",
  50895=>"111111111",
  50896=>"111000000",
  50897=>"000010010",
  50898=>"111111111",
  50899=>"101000100",
  50900=>"011000000",
  50901=>"111111111",
  50902=>"100000000",
  50903=>"111111101",
  50904=>"000000001",
  50905=>"100111111",
  50906=>"011111111",
  50907=>"111111000",
  50908=>"000110110",
  50909=>"101000000",
  50910=>"000000010",
  50911=>"000000000",
  50912=>"111111111",
  50913=>"000011111",
  50914=>"111111111",
  50915=>"111111111",
  50916=>"100100100",
  50917=>"011000000",
  50918=>"010000000",
  50919=>"111111111",
  50920=>"111101111",
  50921=>"111111111",
  50922=>"110111111",
  50923=>"000000000",
  50924=>"111111111",
  50925=>"000000000",
  50926=>"111000000",
  50927=>"001111111",
  50928=>"111101001",
  50929=>"100000000",
  50930=>"011111001",
  50931=>"010000011",
  50932=>"111111111",
  50933=>"111111111",
  50934=>"001100110",
  50935=>"001000000",
  50936=>"000000111",
  50937=>"111111111",
  50938=>"111100111",
  50939=>"111111011",
  50940=>"111111000",
  50941=>"111100000",
  50942=>"111111111",
  50943=>"101000000",
  50944=>"110110111",
  50945=>"101000000",
  50946=>"111101111",
  50947=>"111111001",
  50948=>"011000000",
  50949=>"111111011",
  50950=>"001001111",
  50951=>"111111111",
  50952=>"111111111",
  50953=>"001001101",
  50954=>"000000000",
  50955=>"111101111",
  50956=>"111111110",
  50957=>"000100000",
  50958=>"000000010",
  50959=>"111000000",
  50960=>"000000111",
  50961=>"111111101",
  50962=>"011111111",
  50963=>"010010001",
  50964=>"001001111",
  50965=>"111111111",
  50966=>"111111111",
  50967=>"010110000",
  50968=>"111101101",
  50969=>"001111111",
  50970=>"110010000",
  50971=>"000000000",
  50972=>"111000000",
  50973=>"000010000",
  50974=>"111111111",
  50975=>"111111111",
  50976=>"101000000",
  50977=>"000111111",
  50978=>"000000000",
  50979=>"100000100",
  50980=>"000011111",
  50981=>"000100110",
  50982=>"000110110",
  50983=>"000001000",
  50984=>"111010000",
  50985=>"010111111",
  50986=>"010000000",
  50987=>"000000000",
  50988=>"111111111",
  50989=>"111111100",
  50990=>"111010000",
  50991=>"000000000",
  50992=>"111111111",
  50993=>"000000000",
  50994=>"111111111",
  50995=>"111111000",
  50996=>"111111111",
  50997=>"111111011",
  50998=>"011000000",
  50999=>"111111111",
  51000=>"111111001",
  51001=>"111111111",
  51002=>"000000000",
  51003=>"111000000",
  51004=>"111110111",
  51005=>"111001000",
  51006=>"000000111",
  51007=>"000000111",
  51008=>"111111001",
  51009=>"111111111",
  51010=>"001001000",
  51011=>"111111111",
  51012=>"000000001",
  51013=>"111111111",
  51014=>"010110110",
  51015=>"110110010",
  51016=>"111110110",
  51017=>"000111111",
  51018=>"110101111",
  51019=>"011111111",
  51020=>"111011000",
  51021=>"000000000",
  51022=>"000000000",
  51023=>"000000000",
  51024=>"111111111",
  51025=>"111111111",
  51026=>"100100000",
  51027=>"111000111",
  51028=>"000010111",
  51029=>"000000001",
  51030=>"111111100",
  51031=>"111111111",
  51032=>"001001101",
  51033=>"000000000",
  51034=>"110111111",
  51035=>"111111111",
  51036=>"111111000",
  51037=>"000000000",
  51038=>"111111111",
  51039=>"011011111",
  51040=>"000000001",
  51041=>"001000000",
  51042=>"100111111",
  51043=>"110111111",
  51044=>"001000000",
  51045=>"000000000",
  51046=>"000001011",
  51047=>"000000000",
  51048=>"110111111",
  51049=>"000000001",
  51050=>"000000111",
  51051=>"000000000",
  51052=>"000000000",
  51053=>"111010000",
  51054=>"111111001",
  51055=>"000000100",
  51056=>"111111001",
  51057=>"111111111",
  51058=>"000000000",
  51059=>"000100011",
  51060=>"001000001",
  51061=>"000000000",
  51062=>"001011011",
  51063=>"000100101",
  51064=>"000100110",
  51065=>"000000011",
  51066=>"111111111",
  51067=>"010110111",
  51068=>"000011111",
  51069=>"111111111",
  51070=>"001000011",
  51071=>"111111100",
  51072=>"000000100",
  51073=>"000001001",
  51074=>"011001000",
  51075=>"000000111",
  51076=>"000100000",
  51077=>"110111111",
  51078=>"001001000",
  51079=>"001001011",
  51080=>"111111111",
  51081=>"011001011",
  51082=>"111111000",
  51083=>"001101000",
  51084=>"111111111",
  51085=>"000000000",
  51086=>"111111111",
  51087=>"000000000",
  51088=>"111111110",
  51089=>"000001011",
  51090=>"111111111",
  51091=>"111000100",
  51092=>"111111100",
  51093=>"000000000",
  51094=>"000000001",
  51095=>"000000011",
  51096=>"100101111",
  51097=>"111111000",
  51098=>"000000000",
  51099=>"110001001",
  51100=>"000110111",
  51101=>"010010111",
  51102=>"000000000",
  51103=>"000000000",
  51104=>"011111000",
  51105=>"100000000",
  51106=>"110110111",
  51107=>"000000111",
  51108=>"100111111",
  51109=>"000000000",
  51110=>"000010010",
  51111=>"111111111",
  51112=>"110010000",
  51113=>"000000100",
  51114=>"000001111",
  51115=>"000000000",
  51116=>"111111000",
  51117=>"111111111",
  51118=>"000000000",
  51119=>"000000000",
  51120=>"001100101",
  51121=>"000000000",
  51122=>"010010011",
  51123=>"000000000",
  51124=>"100000000",
  51125=>"111111111",
  51126=>"111111111",
  51127=>"111000000",
  51128=>"000000111",
  51129=>"100110111",
  51130=>"000011011",
  51131=>"000000011",
  51132=>"111111111",
  51133=>"111111111",
  51134=>"010000001",
  51135=>"100100111",
  51136=>"000101111",
  51137=>"011011000",
  51138=>"111000000",
  51139=>"001011000",
  51140=>"111100001",
  51141=>"111111001",
  51142=>"000100111",
  51143=>"110000000",
  51144=>"111111111",
  51145=>"101111011",
  51146=>"111111111",
  51147=>"000000000",
  51148=>"111111110",
  51149=>"000000000",
  51150=>"111111000",
  51151=>"011111111",
  51152=>"101000000",
  51153=>"111001000",
  51154=>"111110110",
  51155=>"111111111",
  51156=>"000000000",
  51157=>"110110000",
  51158=>"000100000",
  51159=>"000000011",
  51160=>"111110111",
  51161=>"100100100",
  51162=>"100000001",
  51163=>"000000100",
  51164=>"001001000",
  51165=>"110100100",
  51166=>"000000000",
  51167=>"001000000",
  51168=>"001000000",
  51169=>"111111111",
  51170=>"111111111",
  51171=>"100100000",
  51172=>"111000000",
  51173=>"000000000",
  51174=>"000000101",
  51175=>"000000000",
  51176=>"000000001",
  51177=>"111011111",
  51178=>"111111110",
  51179=>"110100000",
  51180=>"110110000",
  51181=>"010111110",
  51182=>"111000000",
  51183=>"011110001",
  51184=>"111110110",
  51185=>"000110111",
  51186=>"101000000",
  51187=>"111111111",
  51188=>"000000001",
  51189=>"111111000",
  51190=>"000111111",
  51191=>"110111111",
  51192=>"110110111",
  51193=>"111100111",
  51194=>"111111111",
  51195=>"000010000",
  51196=>"011111000",
  51197=>"010111111",
  51198=>"111111100",
  51199=>"100111111",
  51200=>"111110000",
  51201=>"000010010",
  51202=>"000000000",
  51203=>"111111101",
  51204=>"000000100",
  51205=>"000001000",
  51206=>"000000000",
  51207=>"000000000",
  51208=>"000000000",
  51209=>"000001001",
  51210=>"000011111",
  51211=>"001111110",
  51212=>"000010010",
  51213=>"111110000",
  51214=>"011011001",
  51215=>"000000000",
  51216=>"111111111",
  51217=>"000010111",
  51218=>"111111111",
  51219=>"111111111",
  51220=>"000010000",
  51221=>"000000000",
  51222=>"001000000",
  51223=>"001001000",
  51224=>"011111111",
  51225=>"111111001",
  51226=>"001100000",
  51227=>"011001001",
  51228=>"111111111",
  51229=>"011111011",
  51230=>"011001101",
  51231=>"111111111",
  51232=>"000000000",
  51233=>"111110000",
  51234=>"001001000",
  51235=>"000001001",
  51236=>"111111000",
  51237=>"111111111",
  51238=>"000000000",
  51239=>"000100001",
  51240=>"000000000",
  51241=>"000000000",
  51242=>"011111111",
  51243=>"000000000",
  51244=>"111111111",
  51245=>"111111111",
  51246=>"000000101",
  51247=>"100000000",
  51248=>"000111111",
  51249=>"001111111",
  51250=>"000000000",
  51251=>"011011011",
  51252=>"111011000",
  51253=>"100111000",
  51254=>"000000001",
  51255=>"000000110",
  51256=>"111111000",
  51257=>"110111111",
  51258=>"001111001",
  51259=>"001001000",
  51260=>"111110110",
  51261=>"111111110",
  51262=>"000011011",
  51263=>"000000000",
  51264=>"010010000",
  51265=>"011001000",
  51266=>"000000000",
  51267=>"000111111",
  51268=>"000000000",
  51269=>"110111111",
  51270=>"111111111",
  51271=>"000110111",
  51272=>"000001001",
  51273=>"001001001",
  51274=>"000100111",
  51275=>"000000111",
  51276=>"000000101",
  51277=>"000010111",
  51278=>"111111111",
  51279=>"000111111",
  51280=>"000000000",
  51281=>"000000000",
  51282=>"100000000",
  51283=>"110000000",
  51284=>"011011011",
  51285=>"011000000",
  51286=>"111111111",
  51287=>"111111111",
  51288=>"000000000",
  51289=>"111111000",
  51290=>"100101111",
  51291=>"111011001",
  51292=>"010000000",
  51293=>"000010111",
  51294=>"000000001",
  51295=>"111111111",
  51296=>"111100100",
  51297=>"011010010",
  51298=>"000000000",
  51299=>"000000000",
  51300=>"101101001",
  51301=>"000000110",
  51302=>"000001000",
  51303=>"111111111",
  51304=>"000110111",
  51305=>"111111101",
  51306=>"010011001",
  51307=>"000111111",
  51308=>"111111111",
  51309=>"111111111",
  51310=>"001000011",
  51311=>"111111111",
  51312=>"110110110",
  51313=>"000100111",
  51314=>"001101111",
  51315=>"000011001",
  51316=>"000000000",
  51317=>"001001000",
  51318=>"001000000",
  51319=>"000000011",
  51320=>"010111111",
  51321=>"101101101",
  51322=>"000001011",
  51323=>"111111000",
  51324=>"011000010",
  51325=>"111111111",
  51326=>"000000000",
  51327=>"000000000",
  51328=>"101111000",
  51329=>"000000001",
  51330=>"111111111",
  51331=>"111111111",
  51332=>"111111111",
  51333=>"000111101",
  51334=>"000100100",
  51335=>"100010000",
  51336=>"100000100",
  51337=>"000100100",
  51338=>"001001001",
  51339=>"111111100",
  51340=>"000000000",
  51341=>"000000000",
  51342=>"000100000",
  51343=>"111111111",
  51344=>"110000100",
  51345=>"011111111",
  51346=>"111111111",
  51347=>"000000000",
  51348=>"100111011",
  51349=>"000000000",
  51350=>"111000000",
  51351=>"000000000",
  51352=>"000011001",
  51353=>"111111110",
  51354=>"001001001",
  51355=>"111010000",
  51356=>"000000000",
  51357=>"110110000",
  51358=>"111111001",
  51359=>"111000111",
  51360=>"111111111",
  51361=>"011000000",
  51362=>"000011000",
  51363=>"110100111",
  51364=>"101111111",
  51365=>"000000000",
  51366=>"111111110",
  51367=>"011111111",
  51368=>"001010000",
  51369=>"111111111",
  51370=>"000000000",
  51371=>"111011111",
  51372=>"110000001",
  51373=>"111111011",
  51374=>"000001111",
  51375=>"000100101",
  51376=>"111000011",
  51377=>"101111001",
  51378=>"010110110",
  51379=>"010010110",
  51380=>"000000011",
  51381=>"111111111",
  51382=>"111111111",
  51383=>"110111100",
  51384=>"111001000",
  51385=>"111111111",
  51386=>"111111111",
  51387=>"110000000",
  51388=>"000000000",
  51389=>"110101001",
  51390=>"111111111",
  51391=>"000000000",
  51392=>"010011011",
  51393=>"001000001",
  51394=>"000000000",
  51395=>"101011011",
  51396=>"000110000",
  51397=>"010010000",
  51398=>"100000000",
  51399=>"111111101",
  51400=>"110110100",
  51401=>"000000000",
  51402=>"100000100",
  51403=>"111111111",
  51404=>"001001011",
  51405=>"000000001",
  51406=>"000000000",
  51407=>"000000000",
  51408=>"001000000",
  51409=>"000010111",
  51410=>"010011110",
  51411=>"111111111",
  51412=>"101101111",
  51413=>"000001001",
  51414=>"000000000",
  51415=>"111111111",
  51416=>"111111101",
  51417=>"001001100",
  51418=>"000000010",
  51419=>"011100000",
  51420=>"000011010",
  51421=>"111111111",
  51422=>"000000000",
  51423=>"110100000",
  51424=>"111111111",
  51425=>"000000011",
  51426=>"000000000",
  51427=>"111000000",
  51428=>"010100100",
  51429=>"111111110",
  51430=>"000000000",
  51431=>"101101111",
  51432=>"000000100",
  51433=>"110110000",
  51434=>"001000000",
  51435=>"111111111",
  51436=>"111111011",
  51437=>"000000000",
  51438=>"111111111",
  51439=>"110101111",
  51440=>"111111011",
  51441=>"110110100",
  51442=>"011100000",
  51443=>"111101000",
  51444=>"111111111",
  51445=>"001111111",
  51446=>"000100000",
  51447=>"000111111",
  51448=>"000110111",
  51449=>"111111111",
  51450=>"000000000",
  51451=>"001001111",
  51452=>"110110110",
  51453=>"100111111",
  51454=>"111010000",
  51455=>"000000000",
  51456=>"001001000",
  51457=>"000000000",
  51458=>"100011101",
  51459=>"000001001",
  51460=>"111111111",
  51461=>"000000000",
  51462=>"000000000",
  51463=>"111011111",
  51464=>"000000000",
  51465=>"000000000",
  51466=>"011011110",
  51467=>"001001000",
  51468=>"111011000",
  51469=>"001101111",
  51470=>"111111111",
  51471=>"111111001",
  51472=>"000001000",
  51473=>"000100000",
  51474=>"000000001",
  51475=>"111111011",
  51476=>"111111100",
  51477=>"111111011",
  51478=>"011111111",
  51479=>"111111111",
  51480=>"010000000",
  51481=>"111111001",
  51482=>"111011000",
  51483=>"111101111",
  51484=>"000100100",
  51485=>"000000000",
  51486=>"011011001",
  51487=>"011011011",
  51488=>"100111111",
  51489=>"001000000",
  51490=>"110110111",
  51491=>"000000000",
  51492=>"111000011",
  51493=>"111111101",
  51494=>"000001000",
  51495=>"000000011",
  51496=>"111111111",
  51497=>"000000000",
  51498=>"111011100",
  51499=>"111111111",
  51500=>"000000000",
  51501=>"010011100",
  51502=>"010011111",
  51503=>"111000001",
  51504=>"111111111",
  51505=>"000000011",
  51506=>"000000000",
  51507=>"000000000",
  51508=>"000000000",
  51509=>"001011011",
  51510=>"111111111",
  51511=>"110110100",
  51512=>"000000000",
  51513=>"111111111",
  51514=>"111101111",
  51515=>"000000000",
  51516=>"110110111",
  51517=>"000000111",
  51518=>"100000001",
  51519=>"000100110",
  51520=>"000000000",
  51521=>"000000000",
  51522=>"111111111",
  51523=>"001000000",
  51524=>"000101000",
  51525=>"101001001",
  51526=>"010000000",
  51527=>"111111011",
  51528=>"111111010",
  51529=>"000000110",
  51530=>"000000100",
  51531=>"000010000",
  51532=>"110111111",
  51533=>"110110010",
  51534=>"010000000",
  51535=>"111110110",
  51536=>"110110110",
  51537=>"101111111",
  51538=>"110110111",
  51539=>"111111000",
  51540=>"000000000",
  51541=>"011001001",
  51542=>"111111111",
  51543=>"111111111",
  51544=>"110110000",
  51545=>"111111111",
  51546=>"000100110",
  51547=>"111111111",
  51548=>"111111111",
  51549=>"000000000",
  51550=>"000000110",
  51551=>"000000110",
  51552=>"000000000",
  51553=>"010110000",
  51554=>"110100000",
  51555=>"111111111",
  51556=>"110010000",
  51557=>"000000000",
  51558=>"000000000",
  51559=>"111001000",
  51560=>"110110100",
  51561=>"100100000",
  51562=>"000000101",
  51563=>"000000110",
  51564=>"111111111",
  51565=>"000000000",
  51566=>"000111111",
  51567=>"111101111",
  51568=>"111111111",
  51569=>"111011001",
  51570=>"111111111",
  51571=>"000110111",
  51572=>"000000000",
  51573=>"100101001",
  51574=>"000000111",
  51575=>"100000001",
  51576=>"111111111",
  51577=>"111111111",
  51578=>"000000000",
  51579=>"111111111",
  51580=>"000000001",
  51581=>"111101100",
  51582=>"000000000",
  51583=>"111111111",
  51584=>"110110000",
  51585=>"111111111",
  51586=>"111111111",
  51587=>"000000000",
  51588=>"111111100",
  51589=>"001000000",
  51590=>"000000111",
  51591=>"100110111",
  51592=>"000000000",
  51593=>"110110111",
  51594=>"111111100",
  51595=>"001111111",
  51596=>"111111111",
  51597=>"111010110",
  51598=>"111111111",
  51599=>"000000000",
  51600=>"010010000",
  51601=>"101111111",
  51602=>"000011000",
  51603=>"111111111",
  51604=>"001001000",
  51605=>"000000000",
  51606=>"110000100",
  51607=>"100000000",
  51608=>"000000000",
  51609=>"000010100",
  51610=>"000000101",
  51611=>"111111111",
  51612=>"000000000",
  51613=>"000000000",
  51614=>"010000000",
  51615=>"111111111",
  51616=>"111101111",
  51617=>"111101111",
  51618=>"001111100",
  51619=>"111111111",
  51620=>"111111101",
  51621=>"000111001",
  51622=>"000000000",
  51623=>"011111111",
  51624=>"000000000",
  51625=>"111111111",
  51626=>"001001001",
  51627=>"001000000",
  51628=>"000000000",
  51629=>"000000000",
  51630=>"100101111",
  51631=>"000000000",
  51632=>"000000000",
  51633=>"000000000",
  51634=>"000000000",
  51635=>"000000000",
  51636=>"010100100",
  51637=>"111111111",
  51638=>"111111111",
  51639=>"000100000",
  51640=>"000000000",
  51641=>"110110111",
  51642=>"111110011",
  51643=>"111011001",
  51644=>"111100111",
  51645=>"000000000",
  51646=>"000000000",
  51647=>"100100111",
  51648=>"111101000",
  51649=>"000000100",
  51650=>"111111111",
  51651=>"110111111",
  51652=>"111111111",
  51653=>"111000101",
  51654=>"111111111",
  51655=>"000000111",
  51656=>"111011011",
  51657=>"000000000",
  51658=>"111111001",
  51659=>"000000000",
  51660=>"111000000",
  51661=>"111111111",
  51662=>"111111111",
  51663=>"111111111",
  51664=>"111100110",
  51665=>"111111111",
  51666=>"110110110",
  51667=>"000000000",
  51668=>"111100000",
  51669=>"100100001",
  51670=>"111111001",
  51671=>"000001011",
  51672=>"100000101",
  51673=>"111111110",
  51674=>"000000000",
  51675=>"111111110",
  51676=>"111111111",
  51677=>"110110000",
  51678=>"111110111",
  51679=>"101000101",
  51680=>"000000010",
  51681=>"010010010",
  51682=>"111111111",
  51683=>"111011001",
  51684=>"010011111",
  51685=>"111111111",
  51686=>"111111111",
  51687=>"000000000",
  51688=>"111111111",
  51689=>"000000001",
  51690=>"000000000",
  51691=>"001101111",
  51692=>"100110100",
  51693=>"011111110",
  51694=>"010011011",
  51695=>"111111111",
  51696=>"111111100",
  51697=>"000000000",
  51698=>"111111111",
  51699=>"000111011",
  51700=>"001010000",
  51701=>"000000000",
  51702=>"000000000",
  51703=>"111111110",
  51704=>"100100110",
  51705=>"010000000",
  51706=>"000011111",
  51707=>"011000000",
  51708=>"100000000",
  51709=>"000000001",
  51710=>"001000000",
  51711=>"101001111",
  51712=>"001011111",
  51713=>"000000000",
  51714=>"000000111",
  51715=>"000000000",
  51716=>"000000100",
  51717=>"110001111",
  51718=>"001001000",
  51719=>"110111111",
  51720=>"000001011",
  51721=>"110111111",
  51722=>"110000111",
  51723=>"101111011",
  51724=>"100100111",
  51725=>"001010010",
  51726=>"001001001",
  51727=>"000111111",
  51728=>"111001010",
  51729=>"000110011",
  51730=>"011101101",
  51731=>"111111111",
  51732=>"000100111",
  51733=>"010111000",
  51734=>"000000100",
  51735=>"000111111",
  51736=>"000000000",
  51737=>"110100000",
  51738=>"010110000",
  51739=>"101000000",
  51740=>"000000000",
  51741=>"101111111",
  51742=>"011111000",
  51743=>"100000000",
  51744=>"111101101",
  51745=>"111110110",
  51746=>"111111111",
  51747=>"101110100",
  51748=>"000000000",
  51749=>"111111111",
  51750=>"111001101",
  51751=>"001001011",
  51752=>"001001100",
  51753=>"000000000",
  51754=>"000001111",
  51755=>"111111101",
  51756=>"100000000",
  51757=>"111111111",
  51758=>"110110110",
  51759=>"100100110",
  51760=>"001000000",
  51761=>"000000001",
  51762=>"010011011",
  51763=>"000000000",
  51764=>"110110000",
  51765=>"011011011",
  51766=>"010110011",
  51767=>"000001000",
  51768=>"000001001",
  51769=>"001000110",
  51770=>"000000000",
  51771=>"010000010",
  51772=>"000000000",
  51773=>"110100111",
  51774=>"011111111",
  51775=>"000000000",
  51776=>"110110110",
  51777=>"110010110",
  51778=>"000000000",
  51779=>"010100000",
  51780=>"011111111",
  51781=>"110110000",
  51782=>"100000000",
  51783=>"100100111",
  51784=>"111111011",
  51785=>"101101101",
  51786=>"011111111",
  51787=>"100101111",
  51788=>"100100000",
  51789=>"001110010",
  51790=>"000000101",
  51791=>"111000000",
  51792=>"111111111",
  51793=>"111111111",
  51794=>"001101000",
  51795=>"000000000",
  51796=>"011111011",
  51797=>"000001001",
  51798=>"001001111",
  51799=>"111000010",
  51800=>"000000000",
  51801=>"101000101",
  51802=>"010111111",
  51803=>"111111111",
  51804=>"101111111",
  51805=>"000000111",
  51806=>"111110000",
  51807=>"111111111",
  51808=>"110110111",
  51809=>"110101110",
  51810=>"101111111",
  51811=>"000000011",
  51812=>"100001001",
  51813=>"111111111",
  51814=>"000000000",
  51815=>"000110011",
  51816=>"111111111",
  51817=>"001000000",
  51818=>"001111110",
  51819=>"000000111",
  51820=>"101111111",
  51821=>"111111000",
  51822=>"101011101",
  51823=>"111001000",
  51824=>"000000000",
  51825=>"011011101",
  51826=>"111111011",
  51827=>"000100111",
  51828=>"100000000",
  51829=>"000000001",
  51830=>"000000000",
  51831=>"000000000",
  51832=>"101001001",
  51833=>"001000000",
  51834=>"101101101",
  51835=>"111110111",
  51836=>"111111011",
  51837=>"011000011",
  51838=>"101101101",
  51839=>"010000000",
  51840=>"101000111",
  51841=>"000000111",
  51842=>"111010000",
  51843=>"010000111",
  51844=>"010000000",
  51845=>"001000101",
  51846=>"000000100",
  51847=>"000111110",
  51848=>"111111110",
  51849=>"000100000",
  51850=>"000000001",
  51851=>"111111111",
  51852=>"111000000",
  51853=>"000000000",
  51854=>"110111111",
  51855=>"000001001",
  51856=>"000100111",
  51857=>"110110110",
  51858=>"110110000",
  51859=>"111000000",
  51860=>"101001111",
  51861=>"111111001",
  51862=>"000000000",
  51863=>"111111111",
  51864=>"001111010",
  51865=>"111111111",
  51866=>"000101111",
  51867=>"101111111",
  51868=>"001001111",
  51869=>"001001100",
  51870=>"110001001",
  51871=>"101111111",
  51872=>"111101001",
  51873=>"000000000",
  51874=>"000100100",
  51875=>"000010010",
  51876=>"000001001",
  51877=>"001110110",
  51878=>"000000111",
  51879=>"111111100",
  51880=>"100101101",
  51881=>"000000110",
  51882=>"111000000",
  51883=>"110110000",
  51884=>"000000010",
  51885=>"000000010",
  51886=>"100111111",
  51887=>"101111111",
  51888=>"001000000",
  51889=>"000011011",
  51890=>"111111110",
  51891=>"000000000",
  51892=>"111011110",
  51893=>"001000000",
  51894=>"000000100",
  51895=>"000000000",
  51896=>"111111111",
  51897=>"111111111",
  51898=>"001000000",
  51899=>"101101000",
  51900=>"010000111",
  51901=>"111111011",
  51902=>"111000000",
  51903=>"000000111",
  51904=>"000000000",
  51905=>"100101110",
  51906=>"111111001",
  51907=>"000000000",
  51908=>"000001111",
  51909=>"000111111",
  51910=>"101111010",
  51911=>"000001000",
  51912=>"111111111",
  51913=>"111111101",
  51914=>"110000001",
  51915=>"000000111",
  51916=>"110000100",
  51917=>"100111111",
  51918=>"001000000",
  51919=>"000001000",
  51920=>"111111111",
  51921=>"111000001",
  51922=>"000001001",
  51923=>"010000000",
  51924=>"000000001",
  51925=>"111111111",
  51926=>"110110001",
  51927=>"111110110",
  51928=>"100111111",
  51929=>"100000001",
  51930=>"000000000",
  51931=>"101001111",
  51932=>"000000000",
  51933=>"110000000",
  51934=>"001101111",
  51935=>"111111010",
  51936=>"010011000",
  51937=>"000000010",
  51938=>"101101101",
  51939=>"111111111",
  51940=>"001001001",
  51941=>"100100100",
  51942=>"111000000",
  51943=>"001001001",
  51944=>"100011111",
  51945=>"001000000",
  51946=>"010111111",
  51947=>"011000100",
  51948=>"011111111",
  51949=>"110000000",
  51950=>"111000000",
  51951=>"111111101",
  51952=>"000111111",
  51953=>"000011111",
  51954=>"000000000",
  51955=>"000000111",
  51956=>"111101001",
  51957=>"110100110",
  51958=>"111111011",
  51959=>"110110000",
  51960=>"110110000",
  51961=>"101101000",
  51962=>"010000000",
  51963=>"110111110",
  51964=>"111111111",
  51965=>"100000001",
  51966=>"001001111",
  51967=>"111110001",
  51968=>"000001001",
  51969=>"100101111",
  51970=>"000000000",
  51971=>"000000000",
  51972=>"111111100",
  51973=>"000000100",
  51974=>"111110110",
  51975=>"000000101",
  51976=>"111111001",
  51977=>"111111101",
  51978=>"000000011",
  51979=>"001001000",
  51980=>"100000111",
  51981=>"010100001",
  51982=>"101111011",
  51983=>"100000000",
  51984=>"111101001",
  51985=>"001001000",
  51986=>"111010000",
  51987=>"000111011",
  51988=>"110110001",
  51989=>"111111111",
  51990=>"011011000",
  51991=>"000000000",
  51992=>"000111111",
  51993=>"111111011",
  51994=>"011111011",
  51995=>"000000011",
  51996=>"111111111",
  51997=>"111111010",
  51998=>"000000000",
  51999=>"000001111",
  52000=>"000000000",
  52001=>"000101111",
  52002=>"000101111",
  52003=>"000000000",
  52004=>"111100111",
  52005=>"010000000",
  52006=>"000001000",
  52007=>"000000111",
  52008=>"011111000",
  52009=>"000000000",
  52010=>"000000000",
  52011=>"000000111",
  52012=>"001001001",
  52013=>"101011111",
  52014=>"000000111",
  52015=>"001000000",
  52016=>"101101111",
  52017=>"011000111",
  52018=>"111000111",
  52019=>"111111101",
  52020=>"000000001",
  52021=>"100000001",
  52022=>"010110000",
  52023=>"101101100",
  52024=>"010110000",
  52025=>"111111011",
  52026=>"111111111",
  52027=>"110000000",
  52028=>"111111111",
  52029=>"110111000",
  52030=>"111111011",
  52031=>"101101111",
  52032=>"000000010",
  52033=>"000100100",
  52034=>"110110010",
  52035=>"111100100",
  52036=>"100110111",
  52037=>"001000111",
  52038=>"111111111",
  52039=>"101111111",
  52040=>"111111111",
  52041=>"000000101",
  52042=>"000000000",
  52043=>"100100110",
  52044=>"011011011",
  52045=>"111110010",
  52046=>"101001100",
  52047=>"110000100",
  52048=>"100100100",
  52049=>"001111011",
  52050=>"111000000",
  52051=>"001111111",
  52052=>"100100100",
  52053=>"000001001",
  52054=>"000000100",
  52055=>"000000000",
  52056=>"101101000",
  52057=>"000000100",
  52058=>"011010111",
  52059=>"101111111",
  52060=>"000000111",
  52061=>"111111111",
  52062=>"101100101",
  52063=>"001100100",
  52064=>"101001111",
  52065=>"000000001",
  52066=>"110111111",
  52067=>"100000100",
  52068=>"000100110",
  52069=>"010000000",
  52070=>"001111001",
  52071=>"100000000",
  52072=>"111001000",
  52073=>"111111111",
  52074=>"111000000",
  52075=>"110110110",
  52076=>"100111011",
  52077=>"000100000",
  52078=>"000000000",
  52079=>"111111111",
  52080=>"000001111",
  52081=>"111111111",
  52082=>"100101110",
  52083=>"000100100",
  52084=>"001010000",
  52085=>"111111111",
  52086=>"000000000",
  52087=>"111111111",
  52088=>"000101000",
  52089=>"110000000",
  52090=>"111010000",
  52091=>"000000000",
  52092=>"011111111",
  52093=>"111110000",
  52094=>"111001111",
  52095=>"000000000",
  52096=>"101000110",
  52097=>"001000010",
  52098=>"011011011",
  52099=>"001000000",
  52100=>"101101111",
  52101=>"111111111",
  52102=>"100000000",
  52103=>"111001000",
  52104=>"111111111",
  52105=>"000111111",
  52106=>"100000100",
  52107=>"101001101",
  52108=>"111101111",
  52109=>"000000010",
  52110=>"000000000",
  52111=>"000000000",
  52112=>"010001000",
  52113=>"111011111",
  52114=>"100000011",
  52115=>"001001000",
  52116=>"110111000",
  52117=>"000000000",
  52118=>"000000001",
  52119=>"011011010",
  52120=>"011111111",
  52121=>"111110110",
  52122=>"111111111",
  52123=>"000000000",
  52124=>"101101110",
  52125=>"010111111",
  52126=>"000000110",
  52127=>"000000000",
  52128=>"111111011",
  52129=>"100110110",
  52130=>"000100010",
  52131=>"111111111",
  52132=>"000000100",
  52133=>"100000000",
  52134=>"001001111",
  52135=>"111011111",
  52136=>"010010010",
  52137=>"110000000",
  52138=>"001100100",
  52139=>"000001001",
  52140=>"001000010",
  52141=>"000000000",
  52142=>"111111000",
  52143=>"000000100",
  52144=>"000000100",
  52145=>"000000000",
  52146=>"111000000",
  52147=>"010000000",
  52148=>"000000000",
  52149=>"111111111",
  52150=>"111000001",
  52151=>"001001000",
  52152=>"001011000",
  52153=>"010011011",
  52154=>"111000000",
  52155=>"001110000",
  52156=>"111111000",
  52157=>"100101111",
  52158=>"010110000",
  52159=>"111111001",
  52160=>"001001000",
  52161=>"110111110",
  52162=>"111111111",
  52163=>"000000000",
  52164=>"100100100",
  52165=>"001001001",
  52166=>"100111111",
  52167=>"110111111",
  52168=>"000100111",
  52169=>"100111000",
  52170=>"001001110",
  52171=>"110110111",
  52172=>"110000100",
  52173=>"110111111",
  52174=>"000100100",
  52175=>"010000000",
  52176=>"000000000",
  52177=>"010011011",
  52178=>"111001001",
  52179=>"001000111",
  52180=>"000110111",
  52181=>"000000000",
  52182=>"110111011",
  52183=>"000000011",
  52184=>"111111100",
  52185=>"000000001",
  52186=>"000001001",
  52187=>"101000000",
  52188=>"111110111",
  52189=>"001011011",
  52190=>"000000100",
  52191=>"011000010",
  52192=>"110110110",
  52193=>"001000111",
  52194=>"000111111",
  52195=>"110110111",
  52196=>"111110111",
  52197=>"111110000",
  52198=>"111111000",
  52199=>"000000000",
  52200=>"111111001",
  52201=>"000010000",
  52202=>"000000000",
  52203=>"110110111",
  52204=>"010010000",
  52205=>"100100100",
  52206=>"110010110",
  52207=>"111111111",
  52208=>"011110000",
  52209=>"000000000",
  52210=>"000000000",
  52211=>"111110111",
  52212=>"000000000",
  52213=>"111011111",
  52214=>"111111111",
  52215=>"011001000",
  52216=>"000000000",
  52217=>"100100000",
  52218=>"100100001",
  52219=>"111111011",
  52220=>"110010000",
  52221=>"001001001",
  52222=>"111111000",
  52223=>"111011111",
  52224=>"100000000",
  52225=>"000000000",
  52226=>"111000000",
  52227=>"000000000",
  52228=>"111111111",
  52229=>"000000111",
  52230=>"000111000",
  52231=>"111110110",
  52232=>"000000000",
  52233=>"001111111",
  52234=>"000000000",
  52235=>"000000000",
  52236=>"100100110",
  52237=>"000001011",
  52238=>"000110111",
  52239=>"000000000",
  52240=>"011000000",
  52241=>"000100111",
  52242=>"011111111",
  52243=>"000000000",
  52244=>"111111111",
  52245=>"111111110",
  52246=>"111000000",
  52247=>"111111000",
  52248=>"110110110",
  52249=>"011110010",
  52250=>"100000111",
  52251=>"000001011",
  52252=>"101001111",
  52253=>"111111101",
  52254=>"001000101",
  52255=>"111110000",
  52256=>"110110100",
  52257=>"110111110",
  52258=>"001000001",
  52259=>"111111111",
  52260=>"000000000",
  52261=>"000001000",
  52262=>"000000011",
  52263=>"111111111",
  52264=>"001101111",
  52265=>"111111000",
  52266=>"010000000",
  52267=>"111111111",
  52268=>"000000000",
  52269=>"000000000",
  52270=>"111110000",
  52271=>"001001001",
  52272=>"000000000",
  52273=>"000000000",
  52274=>"000000000",
  52275=>"000000000",
  52276=>"101101101",
  52277=>"011001000",
  52278=>"000101101",
  52279=>"110111111",
  52280=>"000000110",
  52281=>"001011111",
  52282=>"000001011",
  52283=>"111111000",
  52284=>"001000101",
  52285=>"001000000",
  52286=>"000000000",
  52287=>"110111111",
  52288=>"000000000",
  52289=>"000000001",
  52290=>"001001011",
  52291=>"111111111",
  52292=>"001101110",
  52293=>"110111011",
  52294=>"000000111",
  52295=>"111111110",
  52296=>"011111111",
  52297=>"111111111",
  52298=>"000000011",
  52299=>"000000001",
  52300=>"111111111",
  52301=>"111100000",
  52302=>"101000000",
  52303=>"110111011",
  52304=>"001011111",
  52305=>"001001011",
  52306=>"010111111",
  52307=>"000001101",
  52308=>"101101001",
  52309=>"001101111",
  52310=>"001001001",
  52311=>"110110110",
  52312=>"100100111",
  52313=>"101000101",
  52314=>"000010000",
  52315=>"001110000",
  52316=>"000000000",
  52317=>"101000100",
  52318=>"000000010",
  52319=>"111110100",
  52320=>"000000111",
  52321=>"000001000",
  52322=>"001011111",
  52323=>"101101001",
  52324=>"111110000",
  52325=>"010000000",
  52326=>"111111111",
  52327=>"000001111",
  52328=>"110100000",
  52329=>"111111001",
  52330=>"111010000",
  52331=>"111111111",
  52332=>"011001001",
  52333=>"000000000",
  52334=>"111111111",
  52335=>"111110010",
  52336=>"000000000",
  52337=>"001111111",
  52338=>"110111111",
  52339=>"111111110",
  52340=>"000000000",
  52341=>"111101000",
  52342=>"100101111",
  52343=>"111110000",
  52344=>"000000000",
  52345=>"111111111",
  52346=>"111111111",
  52347=>"000000000",
  52348=>"100100100",
  52349=>"111111110",
  52350=>"010000000",
  52351=>"000000000",
  52352=>"110111111",
  52353=>"001000000",
  52354=>"111111111",
  52355=>"011111001",
  52356=>"001000111",
  52357=>"111111111",
  52358=>"011111111",
  52359=>"111101001",
  52360=>"000101100",
  52361=>"000111111",
  52362=>"100000110",
  52363=>"000000101",
  52364=>"000111111",
  52365=>"000000000",
  52366=>"000001111",
  52367=>"000011000",
  52368=>"100000000",
  52369=>"000000101",
  52370=>"111111111",
  52371=>"111111111",
  52372=>"111111001",
  52373=>"110111111",
  52374=>"000001000",
  52375=>"011111011",
  52376=>"000000001",
  52377=>"010110000",
  52378=>"000111111",
  52379=>"000000000",
  52380=>"110111111",
  52381=>"000000001",
  52382=>"000000000",
  52383=>"111111111",
  52384=>"111111111",
  52385=>"101111100",
  52386=>"000000000",
  52387=>"000111111",
  52388=>"111111001",
  52389=>"110111111",
  52390=>"110100111",
  52391=>"100000001",
  52392=>"111111110",
  52393=>"111111111",
  52394=>"000000000",
  52395=>"000000000",
  52396=>"111111111",
  52397=>"100110101",
  52398=>"111000000",
  52399=>"001001001",
  52400=>"111111000",
  52401=>"111111110",
  52402=>"111111111",
  52403=>"111111001",
  52404=>"011011111",
  52405=>"110000000",
  52406=>"000010000",
  52407=>"110111110",
  52408=>"001001111",
  52409=>"111001000",
  52410=>"111111111",
  52411=>"000000000",
  52412=>"011000111",
  52413=>"101100111",
  52414=>"100011111",
  52415=>"000100100",
  52416=>"101111111",
  52417=>"011001011",
  52418=>"110110000",
  52419=>"111000000",
  52420=>"111111000",
  52421=>"111001000",
  52422=>"111111100",
  52423=>"000000000",
  52424=>"011111010",
  52425=>"000000001",
  52426=>"101001101",
  52427=>"011000111",
  52428=>"111111111",
  52429=>"000001111",
  52430=>"000001001",
  52431=>"000101110",
  52432=>"111111100",
  52433=>"111111111",
  52434=>"000001001",
  52435=>"010010000",
  52436=>"101001000",
  52437=>"001000110",
  52438=>"000000111",
  52439=>"111111111",
  52440=>"000000000",
  52441=>"111000000",
  52442=>"111101000",
  52443=>"111111111",
  52444=>"000111111",
  52445=>"000101111",
  52446=>"101001001",
  52447=>"011000001",
  52448=>"000000101",
  52449=>"010010000",
  52450=>"111111000",
  52451=>"001000100",
  52452=>"000110010",
  52453=>"001000100",
  52454=>"111111111",
  52455=>"000000111",
  52456=>"111111110",
  52457=>"101111111",
  52458=>"001001111",
  52459=>"000111000",
  52460=>"000000001",
  52461=>"100110111",
  52462=>"000000111",
  52463=>"000000000",
  52464=>"110111000",
  52465=>"000000000",
  52466=>"111111111",
  52467=>"100000001",
  52468=>"010011111",
  52469=>"110110110",
  52470=>"000000000",
  52471=>"111000010",
  52472=>"000000100",
  52473=>"111111111",
  52474=>"000001111",
  52475=>"111100100",
  52476=>"110110011",
  52477=>"110111110",
  52478=>"001000000",
  52479=>"000000100",
  52480=>"000000000",
  52481=>"001000000",
  52482=>"000000000",
  52483=>"010110010",
  52484=>"111111110",
  52485=>"000000111",
  52486=>"000000000",
  52487=>"000010111",
  52488=>"010000000",
  52489=>"000000001",
  52490=>"001001111",
  52491=>"001111111",
  52492=>"110000000",
  52493=>"111111111",
  52494=>"000000101",
  52495=>"111111111",
  52496=>"000100111",
  52497=>"001011101",
  52498=>"000000000",
  52499=>"001001001",
  52500=>"000000100",
  52501=>"111011011",
  52502=>"100100100",
  52503=>"111111111",
  52504=>"101111110",
  52505=>"000000000",
  52506=>"000001000",
  52507=>"111011010",
  52508=>"110111101",
  52509=>"001000000",
  52510=>"001001111",
  52511=>"111001001",
  52512=>"000100100",
  52513=>"000000000",
  52514=>"011011001",
  52515=>"100101101",
  52516=>"000111110",
  52517=>"111111000",
  52518=>"000000111",
  52519=>"000000111",
  52520=>"010011000",
  52521=>"000000000",
  52522=>"001001011",
  52523=>"000000111",
  52524=>"000010010",
  52525=>"011111111",
  52526=>"000111001",
  52527=>"000000100",
  52528=>"011000000",
  52529=>"111111110",
  52530=>"001000000",
  52531=>"111111001",
  52532=>"111101111",
  52533=>"111111011",
  52534=>"000011000",
  52535=>"111111111",
  52536=>"111011000",
  52537=>"000000000",
  52538=>"011000000",
  52539=>"111110001",
  52540=>"000000000",
  52541=>"000001001",
  52542=>"000000000",
  52543=>"000000000",
  52544=>"000011000",
  52545=>"111111000",
  52546=>"100100110",
  52547=>"011000000",
  52548=>"101001000",
  52549=>"010111111",
  52550=>"000010011",
  52551=>"001001001",
  52552=>"000000111",
  52553=>"000011000",
  52554=>"000100111",
  52555=>"001000100",
  52556=>"111111111",
  52557=>"111011000",
  52558=>"000000111",
  52559=>"011011111",
  52560=>"011011001",
  52561=>"011000111",
  52562=>"000000000",
  52563=>"001000000",
  52564=>"111111111",
  52565=>"011011011",
  52566=>"010000000",
  52567=>"000000001",
  52568=>"100111111",
  52569=>"000000000",
  52570=>"000000000",
  52571=>"000100110",
  52572=>"000000000",
  52573=>"000000000",
  52574=>"100100101",
  52575=>"001001001",
  52576=>"000000111",
  52577=>"111111101",
  52578=>"000000000",
  52579=>"000100110",
  52580=>"101111111",
  52581=>"001001001",
  52582=>"111001000",
  52583=>"000000001",
  52584=>"111111111",
  52585=>"111111000",
  52586=>"001000111",
  52587=>"100000001",
  52588=>"000000000",
  52589=>"001111111",
  52590=>"011011011",
  52591=>"000010000",
  52592=>"001101101",
  52593=>"000000000",
  52594=>"111000000",
  52595=>"111111001",
  52596=>"110010000",
  52597=>"111111111",
  52598=>"111111100",
  52599=>"000000000",
  52600=>"000000000",
  52601=>"000000110",
  52602=>"111000000",
  52603=>"000000000",
  52604=>"000011111",
  52605=>"111000000",
  52606=>"000000000",
  52607=>"001001111",
  52608=>"101111101",
  52609=>"111111001",
  52610=>"111110100",
  52611=>"000000000",
  52612=>"000010111",
  52613=>"010111000",
  52614=>"100100100",
  52615=>"101000111",
  52616=>"101001101",
  52617=>"011011111",
  52618=>"111111111",
  52619=>"000011010",
  52620=>"111111111",
  52621=>"000110100",
  52622=>"111111001",
  52623=>"111111111",
  52624=>"000000000",
  52625=>"001100110",
  52626=>"001001001",
  52627=>"001100111",
  52628=>"001111111",
  52629=>"000010000",
  52630=>"011111111",
  52631=>"001001111",
  52632=>"000000000",
  52633=>"000111111",
  52634=>"111110110",
  52635=>"101000101",
  52636=>"000000111",
  52637=>"010000000",
  52638=>"001011001",
  52639=>"000000001",
  52640=>"111111111",
  52641=>"000000000",
  52642=>"001000000",
  52643=>"000010000",
  52644=>"000100100",
  52645=>"111111011",
  52646=>"001001001",
  52647=>"000000111",
  52648=>"001001001",
  52649=>"111110111",
  52650=>"011000001",
  52651=>"001000000",
  52652=>"000000000",
  52653=>"001001000",
  52654=>"000000110",
  52655=>"110111111",
  52656=>"000000100",
  52657=>"111111001",
  52658=>"001000100",
  52659=>"000110111",
  52660=>"000101101",
  52661=>"111111101",
  52662=>"011101100",
  52663=>"000010000",
  52664=>"111111000",
  52665=>"000101000",
  52666=>"111111000",
  52667=>"011010100",
  52668=>"001111111",
  52669=>"111111111",
  52670=>"100000001",
  52671=>"100101101",
  52672=>"000000000",
  52673=>"000000000",
  52674=>"011000000",
  52675=>"111101101",
  52676=>"101111111",
  52677=>"011111111",
  52678=>"000001001",
  52679=>"111101001",
  52680=>"100100100",
  52681=>"010000000",
  52682=>"000000000",
  52683=>"001101111",
  52684=>"000000101",
  52685=>"001111111",
  52686=>"101001001",
  52687=>"110111111",
  52688=>"111001000",
  52689=>"001000101",
  52690=>"001001111",
  52691=>"111111111",
  52692=>"000001111",
  52693=>"100000000",
  52694=>"011001111",
  52695=>"001000100",
  52696=>"000100000",
  52697=>"000000111",
  52698=>"000000000",
  52699=>"111101101",
  52700=>"000000000",
  52701=>"000000000",
  52702=>"011000000",
  52703=>"001011011",
  52704=>"000000000",
  52705=>"000000000",
  52706=>"011011111",
  52707=>"000110110",
  52708=>"011011000",
  52709=>"000000000",
  52710=>"100000010",
  52711=>"010111111",
  52712=>"000001111",
  52713=>"111111111",
  52714=>"111000000",
  52715=>"111111010",
  52716=>"111101100",
  52717=>"101111111",
  52718=>"111111111",
  52719=>"001111111",
  52720=>"100000111",
  52721=>"000010000",
  52722=>"111110100",
  52723=>"000000000",
  52724=>"011011111",
  52725=>"000000000",
  52726=>"001000001",
  52727=>"000000001",
  52728=>"000000000",
  52729=>"001001001",
  52730=>"000000000",
  52731=>"101001111",
  52732=>"111010101",
  52733=>"100100100",
  52734=>"100100000",
  52735=>"010110100",
  52736=>"111111111",
  52737=>"111111010",
  52738=>"111111100",
  52739=>"100100111",
  52740=>"011000000",
  52741=>"000000000",
  52742=>"111101101",
  52743=>"111111111",
  52744=>"000001111",
  52745=>"000000111",
  52746=>"001000001",
  52747=>"101000101",
  52748=>"111101001",
  52749=>"011000011",
  52750=>"111111000",
  52751=>"101001011",
  52752=>"101110111",
  52753=>"100000000",
  52754=>"110000110",
  52755=>"111000101",
  52756=>"111111110",
  52757=>"001001111",
  52758=>"010000000",
  52759=>"111111110",
  52760=>"100000000",
  52761=>"111111110",
  52762=>"111011000",
  52763=>"111111011",
  52764=>"000000111",
  52765=>"101111011",
  52766=>"100110000",
  52767=>"111100110",
  52768=>"010000000",
  52769=>"111111111",
  52770=>"111111111",
  52771=>"001001000",
  52772=>"111001000",
  52773=>"000010000",
  52774=>"111111110",
  52775=>"001111000",
  52776=>"111011000",
  52777=>"000010000",
  52778=>"111111010",
  52779=>"111010111",
  52780=>"111100100",
  52781=>"000000000",
  52782=>"100100000",
  52783=>"110100101",
  52784=>"101101101",
  52785=>"101001111",
  52786=>"001111000",
  52787=>"100110000",
  52788=>"111111011",
  52789=>"111000000",
  52790=>"101111111",
  52791=>"010110111",
  52792=>"000000111",
  52793=>"110110001",
  52794=>"101001101",
  52795=>"000000000",
  52796=>"001100100",
  52797=>"111100000",
  52798=>"111010000",
  52799=>"101101111",
  52800=>"011000000",
  52801=>"011111000",
  52802=>"111101101",
  52803=>"111111000",
  52804=>"111101111",
  52805=>"111111111",
  52806=>"111111000",
  52807=>"111111111",
  52808=>"001111100",
  52809=>"111101101",
  52810=>"111111010",
  52811=>"001000011",
  52812=>"000000000",
  52813=>"111111001",
  52814=>"000000000",
  52815=>"011001101",
  52816=>"100111111",
  52817=>"000110000",
  52818=>"101001101",
  52819=>"100110110",
  52820=>"000000111",
  52821=>"000111111",
  52822=>"001000001",
  52823=>"010010000",
  52824=>"111111111",
  52825=>"000000001",
  52826=>"000000000",
  52827=>"111111000",
  52828=>"000110110",
  52829=>"111111111",
  52830=>"111111011",
  52831=>"001001001",
  52832=>"010000000",
  52833=>"000000000",
  52834=>"101101001",
  52835=>"111111010",
  52836=>"011001011",
  52837=>"001000100",
  52838=>"001011001",
  52839=>"000000101",
  52840=>"111011111",
  52841=>"000000111",
  52842=>"111110110",
  52843=>"000000000",
  52844=>"100100000",
  52845=>"101100111",
  52846=>"011111111",
  52847=>"000111111",
  52848=>"100111111",
  52849=>"100010110",
  52850=>"000011011",
  52851=>"001000001",
  52852=>"101101111",
  52853=>"111011111",
  52854=>"000000011",
  52855=>"001000101",
  52856=>"110010000",
  52857=>"111111011",
  52858=>"101001101",
  52859=>"000000111",
  52860=>"110110010",
  52861=>"110110100",
  52862=>"100000101",
  52863=>"110000001",
  52864=>"011001011",
  52865=>"101111111",
  52866=>"000000110",
  52867=>"011011111",
  52868=>"111101000",
  52869=>"110000100",
  52870=>"000000000",
  52871=>"000000010",
  52872=>"000000000",
  52873=>"000011011",
  52874=>"000111111",
  52875=>"111110111",
  52876=>"111001001",
  52877=>"111101101",
  52878=>"111111111",
  52879=>"111101101",
  52880=>"000000000",
  52881=>"100110111",
  52882=>"000001001",
  52883=>"111001001",
  52884=>"110110111",
  52885=>"000000000",
  52886=>"000000010",
  52887=>"101111100",
  52888=>"001011111",
  52889=>"111111111",
  52890=>"111111111",
  52891=>"001001001",
  52892=>"011111110",
  52893=>"001000011",
  52894=>"000000100",
  52895=>"111111001",
  52896=>"110000010",
  52897=>"001010000",
  52898=>"101101111",
  52899=>"000100000",
  52900=>"101001111",
  52901=>"000000000",
  52902=>"110110110",
  52903=>"110011000",
  52904=>"111101000",
  52905=>"000000001",
  52906=>"000110100",
  52907=>"001001011",
  52908=>"010010011",
  52909=>"111111011",
  52910=>"000110111",
  52911=>"000000001",
  52912=>"111011011",
  52913=>"001001001",
  52914=>"111100000",
  52915=>"000000000",
  52916=>"101100100",
  52917=>"001111111",
  52918=>"001000101",
  52919=>"000000010",
  52920=>"000000000",
  52921=>"001000111",
  52922=>"100100011",
  52923=>"111111001",
  52924=>"111111000",
  52925=>"010110011",
  52926=>"010000111",
  52927=>"111111111",
  52928=>"000000000",
  52929=>"000001000",
  52930=>"000000000",
  52931=>"000000000",
  52932=>"110000000",
  52933=>"111111000",
  52934=>"111110100",
  52935=>"110110010",
  52936=>"010010010",
  52937=>"001001111",
  52938=>"101000000",
  52939=>"000000011",
  52940=>"110110111",
  52941=>"010110010",
  52942=>"000000110",
  52943=>"101101100",
  52944=>"000000000",
  52945=>"000000010",
  52946=>"111010000",
  52947=>"101101111",
  52948=>"111111011",
  52949=>"000000000",
  52950=>"000010110",
  52951=>"010000001",
  52952=>"110110000",
  52953=>"000001001",
  52954=>"000000001",
  52955=>"000111111",
  52956=>"001001001",
  52957=>"001001100",
  52958=>"111111111",
  52959=>"001000000",
  52960=>"111000000",
  52961=>"011110111",
  52962=>"111111111",
  52963=>"110111001",
  52964=>"111100000",
  52965=>"011001001",
  52966=>"010010000",
  52967=>"000000001",
  52968=>"011111100",
  52969=>"100001001",
  52970=>"000010001",
  52971=>"111111000",
  52972=>"111111111",
  52973=>"111111010",
  52974=>"000111011",
  52975=>"111000000",
  52976=>"000111111",
  52977=>"000001111",
  52978=>"101000100",
  52979=>"011011001",
  52980=>"111010111",
  52981=>"110110000",
  52982=>"011111000",
  52983=>"100000000",
  52984=>"001001111",
  52985=>"110110000",
  52986=>"000001001",
  52987=>"000000010",
  52988=>"000000000",
  52989=>"111001111",
  52990=>"000000000",
  52991=>"101000000",
  52992=>"111111111",
  52993=>"001001001",
  52994=>"111111111",
  52995=>"000001011",
  52996=>"101001011",
  52997=>"011011011",
  52998=>"001000100",
  52999=>"000111111",
  53000=>"000000101",
  53001=>"000000011",
  53002=>"000000111",
  53003=>"100111111",
  53004=>"110100000",
  53005=>"000111111",
  53006=>"000000000",
  53007=>"000000000",
  53008=>"000001101",
  53009=>"000011110",
  53010=>"000000000",
  53011=>"111111001",
  53012=>"000100000",
  53013=>"111111000",
  53014=>"111110000",
  53015=>"111111111",
  53016=>"000110111",
  53017=>"001000000",
  53018=>"000000111",
  53019=>"010010000",
  53020=>"100011001",
  53021=>"111011000",
  53022=>"000010000",
  53023=>"111011001",
  53024=>"000100110",
  53025=>"111111010",
  53026=>"000001111",
  53027=>"011000000",
  53028=>"111111111",
  53029=>"001001001",
  53030=>"100110111",
  53031=>"100111111",
  53032=>"000000111",
  53033=>"111111111",
  53034=>"000000111",
  53035=>"000101111",
  53036=>"011111100",
  53037=>"100001000",
  53038=>"000000000",
  53039=>"011000000",
  53040=>"011000000",
  53041=>"000100101",
  53042=>"000000000",
  53043=>"000111111",
  53044=>"010110000",
  53045=>"110110100",
  53046=>"001111111",
  53047=>"111000001",
  53048=>"011111001",
  53049=>"011000000",
  53050=>"110111111",
  53051=>"001001000",
  53052=>"110111000",
  53053=>"111001101",
  53054=>"000000111",
  53055=>"000010000",
  53056=>"001101111",
  53057=>"100000101",
  53058=>"000001111",
  53059=>"111111010",
  53060=>"111001001",
  53061=>"111111011",
  53062=>"100000111",
  53063=>"111001111",
  53064=>"000001110",
  53065=>"000010000",
  53066=>"111110000",
  53067=>"111110000",
  53068=>"000000001",
  53069=>"000000001",
  53070=>"001001111",
  53071=>"000001100",
  53072=>"001000001",
  53073=>"001000000",
  53074=>"111111111",
  53075=>"110110010",
  53076=>"000000110",
  53077=>"001000000",
  53078=>"000000000",
  53079=>"111111111",
  53080=>"111110110",
  53081=>"011111000",
  53082=>"111110001",
  53083=>"001001111",
  53084=>"000111111",
  53085=>"111101001",
  53086=>"000000000",
  53087=>"000010000",
  53088=>"011111000",
  53089=>"000000000",
  53090=>"011011011",
  53091=>"111001011",
  53092=>"001111111",
  53093=>"001111000",
  53094=>"111000000",
  53095=>"101111111",
  53096=>"111011000",
  53097=>"111111011",
  53098=>"110111011",
  53099=>"011000000",
  53100=>"000111101",
  53101=>"111000011",
  53102=>"000000001",
  53103=>"011001001",
  53104=>"000100100",
  53105=>"000000000",
  53106=>"110111111",
  53107=>"111101100",
  53108=>"111001001",
  53109=>"001001001",
  53110=>"111001001",
  53111=>"001011111",
  53112=>"001000001",
  53113=>"111111010",
  53114=>"111111111",
  53115=>"110110000",
  53116=>"011010111",
  53117=>"110110111",
  53118=>"000000000",
  53119=>"000000000",
  53120=>"111000000",
  53121=>"000000110",
  53122=>"000111111",
  53123=>"011001111",
  53124=>"111110000",
  53125=>"010000011",
  53126=>"000111111",
  53127=>"111111111",
  53128=>"000000001",
  53129=>"111111111",
  53130=>"111111111",
  53131=>"000000000",
  53132=>"101101111",
  53133=>"110111000",
  53134=>"000001100",
  53135=>"001111111",
  53136=>"010010000",
  53137=>"001001111",
  53138=>"000000000",
  53139=>"110110100",
  53140=>"000000000",
  53141=>"000000110",
  53142=>"100000101",
  53143=>"001101111",
  53144=>"100111111",
  53145=>"010111111",
  53146=>"101000001",
  53147=>"111011000",
  53148=>"110110100",
  53149=>"111011111",
  53150=>"000000110",
  53151=>"000000000",
  53152=>"110110000",
  53153=>"000001001",
  53154=>"000001001",
  53155=>"000000000",
  53156=>"011011101",
  53157=>"011111000",
  53158=>"111111011",
  53159=>"000111011",
  53160=>"000000011",
  53161=>"001000000",
  53162=>"100100000",
  53163=>"000000000",
  53164=>"011111000",
  53165=>"000111111",
  53166=>"111111111",
  53167=>"111000001",
  53168=>"011001101",
  53169=>"000000000",
  53170=>"111111111",
  53171=>"111101000",
  53172=>"111111011",
  53173=>"111000111",
  53174=>"101100000",
  53175=>"000101111",
  53176=>"000111111",
  53177=>"110111110",
  53178=>"111001001",
  53179=>"000000111",
  53180=>"010000000",
  53181=>"101000001",
  53182=>"000000111",
  53183=>"001011011",
  53184=>"000000111",
  53185=>"000001001",
  53186=>"000001000",
  53187=>"001001000",
  53188=>"001001111",
  53189=>"111110110",
  53190=>"110110111",
  53191=>"000001111",
  53192=>"000001000",
  53193=>"101000000",
  53194=>"000001001",
  53195=>"110000000",
  53196=>"111000001",
  53197=>"110110111",
  53198=>"000010000",
  53199=>"000000000",
  53200=>"010000000",
  53201=>"000111111",
  53202=>"110110010",
  53203=>"011111000",
  53204=>"001001011",
  53205=>"111000000",
  53206=>"110010001",
  53207=>"100100111",
  53208=>"001001001",
  53209=>"000110110",
  53210=>"001001111",
  53211=>"100111111",
  53212=>"110000001",
  53213=>"111111110",
  53214=>"110100011",
  53215=>"100100100",
  53216=>"111111111",
  53217=>"110111111",
  53218=>"000000101",
  53219=>"111110110",
  53220=>"000000000",
  53221=>"000000111",
  53222=>"001001001",
  53223=>"110111111",
  53224=>"111100100",
  53225=>"001001000",
  53226=>"001111110",
  53227=>"000000000",
  53228=>"111010000",
  53229=>"110110000",
  53230=>"000100011",
  53231=>"111000000",
  53232=>"001000000",
  53233=>"111111000",
  53234=>"000000000",
  53235=>"000010000",
  53236=>"111111111",
  53237=>"000111010",
  53238=>"011011001",
  53239=>"110111110",
  53240=>"000000111",
  53241=>"010110000",
  53242=>"000000000",
  53243=>"100000100",
  53244=>"001000000",
  53245=>"000110111",
  53246=>"000000000",
  53247=>"111111111",
  53248=>"001000111",
  53249=>"000000000",
  53250=>"000000101",
  53251=>"000100100",
  53252=>"001001001",
  53253=>"001101101",
  53254=>"111111110",
  53255=>"111111111",
  53256=>"000000000",
  53257=>"111011000",
  53258=>"111111111",
  53259=>"000111111",
  53260=>"111111111",
  53261=>"111101110",
  53262=>"000011011",
  53263=>"111001000",
  53264=>"001001000",
  53265=>"111111110",
  53266=>"100111100",
  53267=>"100111111",
  53268=>"111111110",
  53269=>"110000000",
  53270=>"111000111",
  53271=>"001101101",
  53272=>"100110110",
  53273=>"001011011",
  53274=>"000000000",
  53275=>"001011000",
  53276=>"110110100",
  53277=>"110111111",
  53278=>"000001000",
  53279=>"000111111",
  53280=>"111111111",
  53281=>"000000000",
  53282=>"000000000",
  53283=>"111111111",
  53284=>"011000011",
  53285=>"000000001",
  53286=>"000000111",
  53287=>"100000111",
  53288=>"001000000",
  53289=>"000000111",
  53290=>"111011011",
  53291=>"111111000",
  53292=>"111111110",
  53293=>"111111100",
  53294=>"001001000",
  53295=>"100000001",
  53296=>"000000000",
  53297=>"111111111",
  53298=>"000111000",
  53299=>"000000000",
  53300=>"100111110",
  53301=>"001000000",
  53302=>"001001001",
  53303=>"011011000",
  53304=>"111000000",
  53305=>"000000000",
  53306=>"111011000",
  53307=>"000000000",
  53308=>"001000111",
  53309=>"101000101",
  53310=>"111001100",
  53311=>"000000000",
  53312=>"000011000",
  53313=>"110110110",
  53314=>"011011010",
  53315=>"000000111",
  53316=>"100111000",
  53317=>"000000000",
  53318=>"000000000",
  53319=>"111111100",
  53320=>"011000000",
  53321=>"000000000",
  53322=>"110100000",
  53323=>"111111111",
  53324=>"000111111",
  53325=>"111111010",
  53326=>"110100100",
  53327=>"111000100",
  53328=>"001001010",
  53329=>"110111111",
  53330=>"001011011",
  53331=>"000101101",
  53332=>"111101100",
  53333=>"000000000",
  53334=>"001000110",
  53335=>"111001001",
  53336=>"000011000",
  53337=>"111100000",
  53338=>"110001000",
  53339=>"111111111",
  53340=>"111111011",
  53341=>"111111000",
  53342=>"000000110",
  53343=>"100100000",
  53344=>"110110000",
  53345=>"000010001",
  53346=>"000000110",
  53347=>"111111110",
  53348=>"000000111",
  53349=>"100111111",
  53350=>"111111111",
  53351=>"000000000",
  53352=>"111000111",
  53353=>"111111111",
  53354=>"011011111",
  53355=>"000000000",
  53356=>"001001011",
  53357=>"111111010",
  53358=>"000000111",
  53359=>"000000000",
  53360=>"000000000",
  53361=>"000000000",
  53362=>"010110110",
  53363=>"100000000",
  53364=>"111101000",
  53365=>"011111001",
  53366=>"000111111",
  53367=>"101111111",
  53368=>"100101111",
  53369=>"000000110",
  53370=>"001111011",
  53371=>"111111111",
  53372=>"000011111",
  53373=>"010010000",
  53374=>"001001001",
  53375=>"011000000",
  53376=>"101001111",
  53377=>"111101001",
  53378=>"110001111",
  53379=>"000000000",
  53380=>"001111111",
  53381=>"111011111",
  53382=>"000000000",
  53383=>"111111111",
  53384=>"000000000",
  53385=>"111111011",
  53386=>"111110010",
  53387=>"111000000",
  53388=>"000000000",
  53389=>"000000101",
  53390=>"100000000",
  53391=>"111111111",
  53392=>"000000100",
  53393=>"111111000",
  53394=>"000000000",
  53395=>"000000000",
  53396=>"111111111",
  53397=>"001010000",
  53398=>"011000000",
  53399=>"000000000",
  53400=>"000000000",
  53401=>"001011111",
  53402=>"111111011",
  53403=>"111111110",
  53404=>"001000100",
  53405=>"001111110",
  53406=>"111101001",
  53407=>"111111111",
  53408=>"000000001",
  53409=>"000110000",
  53410=>"111011000",
  53411=>"111100000",
  53412=>"001000110",
  53413=>"000000000",
  53414=>"111111101",
  53415=>"000100111",
  53416=>"111111000",
  53417=>"001000000",
  53418=>"000000100",
  53419=>"111011000",
  53420=>"000110110",
  53421=>"000100000",
  53422=>"111000000",
  53423=>"101100000",
  53424=>"111111111",
  53425=>"011111100",
  53426=>"111111110",
  53427=>"111000000",
  53428=>"111011000",
  53429=>"001111111",
  53430=>"111000000",
  53431=>"111110111",
  53432=>"111110100",
  53433=>"111111111",
  53434=>"111000111",
  53435=>"101000111",
  53436=>"000011111",
  53437=>"000000100",
  53438=>"111111111",
  53439=>"101001001",
  53440=>"011011001",
  53441=>"111111000",
  53442=>"000011111",
  53443=>"000001001",
  53444=>"111100110",
  53445=>"110110111",
  53446=>"001001100",
  53447=>"001101000",
  53448=>"111110110",
  53449=>"000000000",
  53450=>"010000000",
  53451=>"111100111",
  53452=>"101111111",
  53453=>"110011000",
  53454=>"111111111",
  53455=>"000100111",
  53456=>"010111000",
  53457=>"001110111",
  53458=>"111110110",
  53459=>"000000000",
  53460=>"110110111",
  53461=>"000000100",
  53462=>"000000000",
  53463=>"011111110",
  53464=>"000000000",
  53465=>"011111111",
  53466=>"111000000",
  53467=>"000010111",
  53468=>"000111111",
  53469=>"000000010",
  53470=>"111011000",
  53471=>"111111111",
  53472=>"110110000",
  53473=>"110111000",
  53474=>"100111111",
  53475=>"100110000",
  53476=>"011011001",
  53477=>"100111111",
  53478=>"000111111",
  53479=>"001111111",
  53480=>"110000000",
  53481=>"111111111",
  53482=>"111110111",
  53483=>"000111111",
  53484=>"111011000",
  53485=>"111000101",
  53486=>"100000111",
  53487=>"111111101",
  53488=>"111111111",
  53489=>"000000000",
  53490=>"000000110",
  53491=>"000011011",
  53492=>"001000100",
  53493=>"000001000",
  53494=>"000100110",
  53495=>"000111111",
  53496=>"000111111",
  53497=>"100111001",
  53498=>"111111111",
  53499=>"000000111",
  53500=>"000001110",
  53501=>"000000000",
  53502=>"001111111",
  53503=>"111111111",
  53504=>"000000000",
  53505=>"111010100",
  53506=>"010000000",
  53507=>"010110111",
  53508=>"000110110",
  53509=>"111000000",
  53510=>"000000000",
  53511=>"000000000",
  53512=>"000000000",
  53513=>"010010000",
  53514=>"111000000",
  53515=>"111111110",
  53516=>"000111111",
  53517=>"111111111",
  53518=>"011000000",
  53519=>"100111101",
  53520=>"001111001",
  53521=>"111110000",
  53522=>"011001000",
  53523=>"000001000",
  53524=>"000111111",
  53525=>"000000111",
  53526=>"111011000",
  53527=>"111111101",
  53528=>"111000000",
  53529=>"110111010",
  53530=>"000000111",
  53531=>"001001000",
  53532=>"000100000",
  53533=>"000000000",
  53534=>"011000000",
  53535=>"111110101",
  53536=>"001001011",
  53537=>"111111111",
  53538=>"011000000",
  53539=>"000100110",
  53540=>"110000000",
  53541=>"111111111",
  53542=>"100101101",
  53543=>"111111111",
  53544=>"111111000",
  53545=>"111110000",
  53546=>"011111111",
  53547=>"111111111",
  53548=>"000100111",
  53549=>"111111111",
  53550=>"000000000",
  53551=>"111111111",
  53552=>"000000001",
  53553=>"111111111",
  53554=>"000000001",
  53555=>"000000110",
  53556=>"000111111",
  53557=>"100110100",
  53558=>"000000000",
  53559=>"111000000",
  53560=>"111111111",
  53561=>"000111111",
  53562=>"000000001",
  53563=>"111111111",
  53564=>"111100110",
  53565=>"100111101",
  53566=>"001000000",
  53567=>"001101111",
  53568=>"000000011",
  53569=>"000000001",
  53570=>"111111111",
  53571=>"111011000",
  53572=>"011111000",
  53573=>"001011001",
  53574=>"001101111",
  53575=>"111000101",
  53576=>"000000111",
  53577=>"111111000",
  53578=>"000000000",
  53579=>"000000001",
  53580=>"111111011",
  53581=>"000000000",
  53582=>"000000011",
  53583=>"000100000",
  53584=>"001111111",
  53585=>"000000011",
  53586=>"000000011",
  53587=>"011111111",
  53588=>"100110100",
  53589=>"000010000",
  53590=>"000110111",
  53591=>"000000111",
  53592=>"101100000",
  53593=>"111111100",
  53594=>"000011111",
  53595=>"111111111",
  53596=>"000000000",
  53597=>"100000000",
  53598=>"001001111",
  53599=>"111111000",
  53600=>"000000001",
  53601=>"111111111",
  53602=>"000000000",
  53603=>"111100101",
  53604=>"000000000",
  53605=>"111000111",
  53606=>"100000111",
  53607=>"001000000",
  53608=>"100110010",
  53609=>"111111011",
  53610=>"000000000",
  53611=>"000010110",
  53612=>"001001011",
  53613=>"101111111",
  53614=>"000111011",
  53615=>"111111111",
  53616=>"000000000",
  53617=>"011011111",
  53618=>"100110111",
  53619=>"000000011",
  53620=>"011111111",
  53621=>"001100111",
  53622=>"111111010",
  53623=>"001111011",
  53624=>"000000111",
  53625=>"000000110",
  53626=>"000000000",
  53627=>"111100000",
  53628=>"001101000",
  53629=>"111101000",
  53630=>"011101111",
  53631=>"111110110",
  53632=>"010001001",
  53633=>"001111000",
  53634=>"001000001",
  53635=>"111111110",
  53636=>"000111011",
  53637=>"111111111",
  53638=>"000111111",
  53639=>"011111000",
  53640=>"111000000",
  53641=>"110100100",
  53642=>"001000000",
  53643=>"111001111",
  53644=>"000111111",
  53645=>"111001001",
  53646=>"111111000",
  53647=>"111111111",
  53648=>"000000000",
  53649=>"111101110",
  53650=>"000110110",
  53651=>"111111011",
  53652=>"000001111",
  53653=>"011111010",
  53654=>"000000000",
  53655=>"001001001",
  53656=>"001011010",
  53657=>"001100111",
  53658=>"001000000",
  53659=>"111100011",
  53660=>"100111000",
  53661=>"000000011",
  53662=>"101101101",
  53663=>"000111111",
  53664=>"000000111",
  53665=>"001001001",
  53666=>"000001011",
  53667=>"001101111",
  53668=>"011001000",
  53669=>"110110000",
  53670=>"000000110",
  53671=>"111110100",
  53672=>"000010111",
  53673=>"000011111",
  53674=>"111111111",
  53675=>"111000001",
  53676=>"000000000",
  53677=>"001111011",
  53678=>"000000000",
  53679=>"101000000",
  53680=>"000000000",
  53681=>"000000000",
  53682=>"100000001",
  53683=>"110000000",
  53684=>"101101000",
  53685=>"111111111",
  53686=>"000100000",
  53687=>"011011000",
  53688=>"111111111",
  53689=>"111001000",
  53690=>"111111000",
  53691=>"111111000",
  53692=>"000000000",
  53693=>"000000000",
  53694=>"010111111",
  53695=>"111111101",
  53696=>"000000010",
  53697=>"000000000",
  53698=>"000000000",
  53699=>"111111111",
  53700=>"000000010",
  53701=>"000000000",
  53702=>"000101111",
  53703=>"000010110",
  53704=>"101010011",
  53705=>"011111000",
  53706=>"000000000",
  53707=>"111111011",
  53708=>"110111111",
  53709=>"100110110",
  53710=>"000000000",
  53711=>"100000000",
  53712=>"000000000",
  53713=>"111000000",
  53714=>"001111011",
  53715=>"000001111",
  53716=>"000010000",
  53717=>"010111111",
  53718=>"111111111",
  53719=>"110110101",
  53720=>"111000000",
  53721=>"111001101",
  53722=>"111111001",
  53723=>"000000111",
  53724=>"000010000",
  53725=>"001011000",
  53726=>"111110111",
  53727=>"000001011",
  53728=>"000000000",
  53729=>"111111000",
  53730=>"011000000",
  53731=>"100111100",
  53732=>"100000000",
  53733=>"011111011",
  53734=>"110111100",
  53735=>"001000000",
  53736=>"111000000",
  53737=>"111111111",
  53738=>"000000000",
  53739=>"000011111",
  53740=>"111111111",
  53741=>"101100101",
  53742=>"111110110",
  53743=>"101101001",
  53744=>"101100101",
  53745=>"000000100",
  53746=>"000100000",
  53747=>"000000000",
  53748=>"111000100",
  53749=>"011111111",
  53750=>"111000100",
  53751=>"000000100",
  53752=>"110111110",
  53753=>"101111101",
  53754=>"111111111",
  53755=>"111111000",
  53756=>"000000000",
  53757=>"000000000",
  53758=>"001010111",
  53759=>"100100000",
  53760=>"111111011",
  53761=>"000000000",
  53762=>"101000000",
  53763=>"111000000",
  53764=>"011011011",
  53765=>"111111111",
  53766=>"111111110",
  53767=>"000001111",
  53768=>"000011000",
  53769=>"011010111",
  53770=>"110100101",
  53771=>"001000100",
  53772=>"011111000",
  53773=>"110110111",
  53774=>"000000000",
  53775=>"000100111",
  53776=>"111111111",
  53777=>"000000010",
  53778=>"111111110",
  53779=>"111101000",
  53780=>"001000001",
  53781=>"111110110",
  53782=>"110111111",
  53783=>"110110110",
  53784=>"101001111",
  53785=>"100111000",
  53786=>"100000000",
  53787=>"111111111",
  53788=>"011000011",
  53789=>"000000000",
  53790=>"000100111",
  53791=>"000000111",
  53792=>"000000000",
  53793=>"100000000",
  53794=>"110110000",
  53795=>"111011011",
  53796=>"011000000",
  53797=>"111010000",
  53798=>"111001111",
  53799=>"000110000",
  53800=>"111011011",
  53801=>"000000000",
  53802=>"000100100",
  53803=>"111111110",
  53804=>"000000011",
  53805=>"111111111",
  53806=>"010011010",
  53807=>"000000110",
  53808=>"000000110",
  53809=>"000101111",
  53810=>"111111000",
  53811=>"000000000",
  53812=>"010110000",
  53813=>"000000110",
  53814=>"000000000",
  53815=>"011101101",
  53816=>"000000000",
  53817=>"000110111",
  53818=>"100111111",
  53819=>"000111111",
  53820=>"000000110",
  53821=>"000000010",
  53822=>"110110111",
  53823=>"000000000",
  53824=>"111111010",
  53825=>"011011000",
  53826=>"000010110",
  53827=>"111000000",
  53828=>"001000000",
  53829=>"000000100",
  53830=>"111000000",
  53831=>"111000000",
  53832=>"001001111",
  53833=>"010000011",
  53834=>"111111000",
  53835=>"101000111",
  53836=>"000000000",
  53837=>"001001000",
  53838=>"001111111",
  53839=>"000000100",
  53840=>"111111010",
  53841=>"110110000",
  53842=>"100000000",
  53843=>"001001000",
  53844=>"000000010",
  53845=>"111000000",
  53846=>"111111001",
  53847=>"000000000",
  53848=>"110100000",
  53849=>"100100100",
  53850=>"111111111",
  53851=>"011111111",
  53852=>"000100100",
  53853=>"100000111",
  53854=>"000000111",
  53855=>"000000000",
  53856=>"010111100",
  53857=>"111111010",
  53858=>"000000001",
  53859=>"000000000",
  53860=>"111000000",
  53861=>"111111000",
  53862=>"001000000",
  53863=>"111111111",
  53864=>"000000000",
  53865=>"111111111",
  53866=>"000010110",
  53867=>"000000000",
  53868=>"111111111",
  53869=>"000000001",
  53870=>"000000000",
  53871=>"011101001",
  53872=>"100110110",
  53873=>"000000001",
  53874=>"000000011",
  53875=>"010110110",
  53876=>"111111000",
  53877=>"000000110",
  53878=>"000000111",
  53879=>"111111111",
  53880=>"111001001",
  53881=>"111111011",
  53882=>"100000000",
  53883=>"111111001",
  53884=>"101001000",
  53885=>"101000000",
  53886=>"111111111",
  53887=>"000111111",
  53888=>"000111111",
  53889=>"001111111",
  53890=>"000010111",
  53891=>"111111010",
  53892=>"100111011",
  53893=>"000000000",
  53894=>"000001111",
  53895=>"000000000",
  53896=>"000000000",
  53897=>"000000000",
  53898=>"111110100",
  53899=>"111111000",
  53900=>"000110111",
  53901=>"000000000",
  53902=>"110111111",
  53903=>"111111111",
  53904=>"111000111",
  53905=>"000000111",
  53906=>"000001111",
  53907=>"000000000",
  53908=>"110000000",
  53909=>"000001001",
  53910=>"011000000",
  53911=>"000000000",
  53912=>"000000100",
  53913=>"000000111",
  53914=>"100111111",
  53915=>"001001001",
  53916=>"100111100",
  53917=>"000000000",
  53918=>"111111011",
  53919=>"110100000",
  53920=>"111111111",
  53921=>"000111111",
  53922=>"110000100",
  53923=>"111111011",
  53924=>"101111000",
  53925=>"111100100",
  53926=>"001000100",
  53927=>"000010000",
  53928=>"001111101",
  53929=>"100101000",
  53930=>"000000111",
  53931=>"000100110",
  53932=>"101100100",
  53933=>"111100000",
  53934=>"111111000",
  53935=>"111111100",
  53936=>"110000111",
  53937=>"100000111",
  53938=>"110111010",
  53939=>"000000000",
  53940=>"011000010",
  53941=>"111111111",
  53942=>"000101000",
  53943=>"000110111",
  53944=>"010000111",
  53945=>"111111011",
  53946=>"100000000",
  53947=>"110111011",
  53948=>"111111001",
  53949=>"000100111",
  53950=>"111111111",
  53951=>"000000000",
  53952=>"100100111",
  53953=>"101000111",
  53954=>"000000111",
  53955=>"000000001",
  53956=>"111111111",
  53957=>"000001000",
  53958=>"011001000",
  53959=>"111111110",
  53960=>"110110110",
  53961=>"110110111",
  53962=>"001001111",
  53963=>"000000000",
  53964=>"111000000",
  53965=>"000000000",
  53966=>"000000001",
  53967=>"111110000",
  53968=>"100000110",
  53969=>"001110110",
  53970=>"000000111",
  53971=>"111100100",
  53972=>"000000000",
  53973=>"100111000",
  53974=>"111111101",
  53975=>"111111111",
  53976=>"111010100",
  53977=>"000000111",
  53978=>"111111111",
  53979=>"000110111",
  53980=>"000000001",
  53981=>"111001011",
  53982=>"001000100",
  53983=>"001100111",
  53984=>"111111111",
  53985=>"111111111",
  53986=>"110111111",
  53987=>"000000000",
  53988=>"001100111",
  53989=>"100100110",
  53990=>"000000000",
  53991=>"101111111",
  53992=>"111111001",
  53993=>"000111011",
  53994=>"111000101",
  53995=>"001011111",
  53996=>"110000000",
  53997=>"111011001",
  53998=>"000100100",
  53999=>"111010000",
  54000=>"111110110",
  54001=>"000101111",
  54002=>"111111111",
  54003=>"000000011",
  54004=>"111111111",
  54005=>"000000000",
  54006=>"100101111",
  54007=>"000000001",
  54008=>"111111110",
  54009=>"011000000",
  54010=>"000000001",
  54011=>"100100100",
  54012=>"111111111",
  54013=>"011111000",
  54014=>"111110111",
  54015=>"100000000",
  54016=>"000000001",
  54017=>"001001111",
  54018=>"110000000",
  54019=>"111111000",
  54020=>"000000000",
  54021=>"000000000",
  54022=>"111001001",
  54023=>"101001001",
  54024=>"000000000",
  54025=>"010000011",
  54026=>"111111111",
  54027=>"111111000",
  54028=>"110100100",
  54029=>"011000000",
  54030=>"000001111",
  54031=>"010111111",
  54032=>"111111000",
  54033=>"010111111",
  54034=>"111111000",
  54035=>"000000001",
  54036=>"001001111",
  54037=>"000011000",
  54038=>"000110000",
  54039=>"111010011",
  54040=>"101100101",
  54041=>"100111111",
  54042=>"101110110",
  54043=>"111000000",
  54044=>"100110100",
  54045=>"110101011",
  54046=>"000100000",
  54047=>"000010110",
  54048=>"100100111",
  54049=>"000000111",
  54050=>"100100100",
  54051=>"111111111",
  54052=>"000011111",
  54053=>"000111100",
  54054=>"000000010",
  54055=>"111001111",
  54056=>"111111111",
  54057=>"110111010",
  54058=>"011111110",
  54059=>"101001101",
  54060=>"000111001",
  54061=>"001011011",
  54062=>"100111111",
  54063=>"110110110",
  54064=>"111101101",
  54065=>"001000001",
  54066=>"000000010",
  54067=>"111111000",
  54068=>"000000000",
  54069=>"000000001",
  54070=>"001111111",
  54071=>"110100000",
  54072=>"111111010",
  54073=>"111000000",
  54074=>"000000000",
  54075=>"011000111",
  54076=>"100100100",
  54077=>"111000100",
  54078=>"000000000",
  54079=>"100100100",
  54080=>"000000000",
  54081=>"110000000",
  54082=>"001100111",
  54083=>"001111111",
  54084=>"111111110",
  54085=>"100000000",
  54086=>"111111110",
  54087=>"000011000",
  54088=>"010110111",
  54089=>"001001001",
  54090=>"000000100",
  54091=>"110110110",
  54092=>"000100111",
  54093=>"000000110",
  54094=>"000010111",
  54095=>"000000100",
  54096=>"101100110",
  54097=>"000111111",
  54098=>"110000010",
  54099=>"011011011",
  54100=>"111011001",
  54101=>"001001001",
  54102=>"011000111",
  54103=>"010010000",
  54104=>"111111111",
  54105=>"111000000",
  54106=>"111111000",
  54107=>"111111110",
  54108=>"110110110",
  54109=>"111100111",
  54110=>"101111110",
  54111=>"111111111",
  54112=>"101101101",
  54113=>"111100000",
  54114=>"000111111",
  54115=>"111111000",
  54116=>"110110000",
  54117=>"001000001",
  54118=>"011111001",
  54119=>"111111010",
  54120=>"111111110",
  54121=>"111111110",
  54122=>"001001011",
  54123=>"110111010",
  54124=>"001001100",
  54125=>"000000000",
  54126=>"010111111",
  54127=>"000000000",
  54128=>"111000000",
  54129=>"111000111",
  54130=>"000000000",
  54131=>"001111111",
  54132=>"000000000",
  54133=>"000000001",
  54134=>"000010000",
  54135=>"111111111",
  54136=>"111111111",
  54137=>"111111000",
  54138=>"001000001",
  54139=>"011110000",
  54140=>"100000000",
  54141=>"101000000",
  54142=>"000000000",
  54143=>"001111101",
  54144=>"110111111",
  54145=>"100100111",
  54146=>"000000000",
  54147=>"000000000",
  54148=>"111111001",
  54149=>"010110111",
  54150=>"111001001",
  54151=>"100000000",
  54152=>"011000000",
  54153=>"010010000",
  54154=>"111111010",
  54155=>"010011000",
  54156=>"111111111",
  54157=>"111111111",
  54158=>"110111000",
  54159=>"000000111",
  54160=>"111111111",
  54161=>"111100000",
  54162=>"000000111",
  54163=>"000001011",
  54164=>"010000000",
  54165=>"010110000",
  54166=>"001001101",
  54167=>"000000110",
  54168=>"001001111",
  54169=>"000100111",
  54170=>"111111111",
  54171=>"111111000",
  54172=>"111111111",
  54173=>"011011111",
  54174=>"111000100",
  54175=>"110110111",
  54176=>"111101111",
  54177=>"010000100",
  54178=>"110111011",
  54179=>"000000000",
  54180=>"111111111",
  54181=>"111111111",
  54182=>"000000100",
  54183=>"001000000",
  54184=>"010010000",
  54185=>"000001111",
  54186=>"111111000",
  54187=>"001011000",
  54188=>"001001001",
  54189=>"010000001",
  54190=>"000011110",
  54191=>"000000000",
  54192=>"000000000",
  54193=>"111111000",
  54194=>"000111100",
  54195=>"000000110",
  54196=>"111111001",
  54197=>"111111010",
  54198=>"110000000",
  54199=>"000000000",
  54200=>"101100000",
  54201=>"111101001",
  54202=>"000000000",
  54203=>"110110110",
  54204=>"000000000",
  54205=>"111111111",
  54206=>"111101100",
  54207=>"111111111",
  54208=>"110010000",
  54209=>"111111111",
  54210=>"111111111",
  54211=>"000000001",
  54212=>"111101110",
  54213=>"111000000",
  54214=>"000000111",
  54215=>"000000000",
  54216=>"000000000",
  54217=>"100100000",
  54218=>"000000000",
  54219=>"111111111",
  54220=>"000000010",
  54221=>"000000111",
  54222=>"000000100",
  54223=>"001001100",
  54224=>"011100110",
  54225=>"111110000",
  54226=>"110111011",
  54227=>"011000001",
  54228=>"111111101",
  54229=>"001111111",
  54230=>"010111000",
  54231=>"110111000",
  54232=>"000110110",
  54233=>"111111111",
  54234=>"011001001",
  54235=>"111110000",
  54236=>"100111100",
  54237=>"111111111",
  54238=>"011000000",
  54239=>"101111111",
  54240=>"000010110",
  54241=>"000110110",
  54242=>"110000000",
  54243=>"000000101",
  54244=>"110000000",
  54245=>"001001001",
  54246=>"000111111",
  54247=>"001000000",
  54248=>"101001101",
  54249=>"110110111",
  54250=>"111111011",
  54251=>"111110110",
  54252=>"000000111",
  54253=>"000000000",
  54254=>"111111111",
  54255=>"100111111",
  54256=>"111100100",
  54257=>"110110110",
  54258=>"111110000",
  54259=>"000110111",
  54260=>"111111000",
  54261=>"011111001",
  54262=>"111111111",
  54263=>"111111111",
  54264=>"111111010",
  54265=>"100100100",
  54266=>"000000011",
  54267=>"001000000",
  54268=>"010110010",
  54269=>"111111000",
  54270=>"000010111",
  54271=>"100111111",
  54272=>"001100000",
  54273=>"000000000",
  54274=>"000000000",
  54275=>"000110110",
  54276=>"000000100",
  54277=>"001001101",
  54278=>"000000110",
  54279=>"111001000",
  54280=>"111000000",
  54281=>"000000000",
  54282=>"111100100",
  54283=>"100101001",
  54284=>"110000000",
  54285=>"111111101",
  54286=>"111001011",
  54287=>"000000000",
  54288=>"001001111",
  54289=>"000000110",
  54290=>"111101000",
  54291=>"111011001",
  54292=>"000000000",
  54293=>"000001111",
  54294=>"100000000",
  54295=>"111111001",
  54296=>"111011010",
  54297=>"110010000",
  54298=>"111000000",
  54299=>"011001000",
  54300=>"000000000",
  54301=>"000000000",
  54302=>"010111000",
  54303=>"111111000",
  54304=>"111001000",
  54305=>"111111000",
  54306=>"001000000",
  54307=>"111111110",
  54308=>"111001000",
  54309=>"111111110",
  54310=>"000001010",
  54311=>"010000000",
  54312=>"000000000",
  54313=>"000000000",
  54314=>"111111000",
  54315=>"000000111",
  54316=>"111111001",
  54317=>"000000111",
  54318=>"000000100",
  54319=>"100111111",
  54320=>"111101111",
  54321=>"110000000",
  54322=>"100110000",
  54323=>"000000000",
  54324=>"111111000",
  54325=>"000000000",
  54326=>"000100111",
  54327=>"111110100",
  54328=>"000100101",
  54329=>"111111000",
  54330=>"001011011",
  54331=>"111111101",
  54332=>"101100111",
  54333=>"000000000",
  54334=>"000000011",
  54335=>"000000011",
  54336=>"000001001",
  54337=>"000000000",
  54338=>"001001001",
  54339=>"011011111",
  54340=>"000010110",
  54341=>"000000110",
  54342=>"000000110",
  54343=>"000000000",
  54344=>"111111011",
  54345=>"011011111",
  54346=>"000101000",
  54347=>"001001000",
  54348=>"111110010",
  54349=>"001000000",
  54350=>"000000001",
  54351=>"111111111",
  54352=>"000001000",
  54353=>"111111111",
  54354=>"000100000",
  54355=>"001001011",
  54356=>"000000000",
  54357=>"000000000",
  54358=>"111111111",
  54359=>"000100000",
  54360=>"000000000",
  54361=>"000000011",
  54362=>"000000000",
  54363=>"001001100",
  54364=>"000000000",
  54365=>"111111010",
  54366=>"111111010",
  54367=>"010010100",
  54368=>"000000000",
  54369=>"100000100",
  54370=>"111111111",
  54371=>"111101100",
  54372=>"111110000",
  54373=>"000000000",
  54374=>"111111111",
  54375=>"111111111",
  54376=>"000001111",
  54377=>"111101111",
  54378=>"011000000",
  54379=>"011001000",
  54380=>"010110110",
  54381=>"000000000",
  54382=>"000000010",
  54383=>"000000000",
  54384=>"101000000",
  54385=>"001001111",
  54386=>"100111111",
  54387=>"111101000",
  54388=>"111111110",
  54389=>"111010000",
  54390=>"111100111",
  54391=>"000000111",
  54392=>"101001001",
  54393=>"111111000",
  54394=>"111000000",
  54395=>"000000000",
  54396=>"110111110",
  54397=>"000010000",
  54398=>"000000000",
  54399=>"000000111",
  54400=>"000000000",
  54401=>"000001111",
  54402=>"111111000",
  54403=>"111111000",
  54404=>"001001000",
  54405=>"111000101",
  54406=>"111111111",
  54407=>"000100111",
  54408=>"101111111",
  54409=>"111111111",
  54410=>"000110110",
  54411=>"100100100",
  54412=>"101101111",
  54413=>"000000000",
  54414=>"000100111",
  54415=>"111111111",
  54416=>"111001000",
  54417=>"000000000",
  54418=>"001000000",
  54419=>"110111110",
  54420=>"100000011",
  54421=>"111111111",
  54422=>"110111111",
  54423=>"111111001",
  54424=>"000000111",
  54425=>"000000000",
  54426=>"000000000",
  54427=>"110000000",
  54428=>"000000110",
  54429=>"001001111",
  54430=>"000100100",
  54431=>"000000111",
  54432=>"100000000",
  54433=>"001011001",
  54434=>"000000111",
  54435=>"010111111",
  54436=>"000000000",
  54437=>"111100111",
  54438=>"111000001",
  54439=>"111111011",
  54440=>"111010000",
  54441=>"000000100",
  54442=>"111100100",
  54443=>"001000111",
  54444=>"111001000",
  54445=>"111100001",
  54446=>"001001111",
  54447=>"111111111",
  54448=>"111111000",
  54449=>"111011011",
  54450=>"111111111",
  54451=>"000000000",
  54452=>"111111010",
  54453=>"111111011",
  54454=>"000000111",
  54455=>"000000111",
  54456=>"111000111",
  54457=>"111000000",
  54458=>"000000000",
  54459=>"111111100",
  54460=>"010111010",
  54461=>"111100000",
  54462=>"100000000",
  54463=>"001000000",
  54464=>"001111011",
  54465=>"111111010",
  54466=>"111111111",
  54467=>"000000000",
  54468=>"111111111",
  54469=>"111111101",
  54470=>"111111000",
  54471=>"101111011",
  54472=>"000001011",
  54473=>"111111001",
  54474=>"111111100",
  54475=>"110111010",
  54476=>"101001001",
  54477=>"100101111",
  54478=>"110000000",
  54479=>"111111000",
  54480=>"111111100",
  54481=>"000011111",
  54482=>"000000000",
  54483=>"000100000",
  54484=>"000000000",
  54485=>"011000000",
  54486=>"000100000",
  54487=>"111111111",
  54488=>"000000000",
  54489=>"100000000",
  54490=>"111100110",
  54491=>"000001001",
  54492=>"111110000",
  54493=>"000011001",
  54494=>"111111011",
  54495=>"100111111",
  54496=>"000000000",
  54497=>"000000110",
  54498=>"111111011",
  54499=>"000000000",
  54500=>"000110100",
  54501=>"010000000",
  54502=>"111111010",
  54503=>"111111111",
  54504=>"000000110",
  54505=>"000001000",
  54506=>"000001011",
  54507=>"000111111",
  54508=>"111111000",
  54509=>"000000000",
  54510=>"111111111",
  54511=>"000000000",
  54512=>"000001000",
  54513=>"110110110",
  54514=>"111111111",
  54515=>"000000101",
  54516=>"000000100",
  54517=>"001111001",
  54518=>"110110011",
  54519=>"000001111",
  54520=>"111111111",
  54521=>"001001000",
  54522=>"000000000",
  54523=>"000000101",
  54524=>"111111111",
  54525=>"011011110",
  54526=>"100000000",
  54527=>"111111111",
  54528=>"000000111",
  54529=>"001101111",
  54530=>"110000111",
  54531=>"111110000",
  54532=>"100100110",
  54533=>"000010010",
  54534=>"000000001",
  54535=>"011111000",
  54536=>"000110111",
  54537=>"000000111",
  54538=>"000000001",
  54539=>"001000001",
  54540=>"111000000",
  54541=>"000000000",
  54542=>"001000011",
  54543=>"000001001",
  54544=>"000111111",
  54545=>"000111101",
  54546=>"101000000",
  54547=>"111111111",
  54548=>"000111111",
  54549=>"111111111",
  54550=>"111100100",
  54551=>"000100111",
  54552=>"111111000",
  54553=>"110000000",
  54554=>"111111000",
  54555=>"110110000",
  54556=>"010011111",
  54557=>"000000000",
  54558=>"000000000",
  54559=>"000010111",
  54560=>"111111111",
  54561=>"111111111",
  54562=>"111111000",
  54563=>"011111111",
  54564=>"001000000",
  54565=>"111111000",
  54566=>"000011011",
  54567=>"011001001",
  54568=>"111010110",
  54569=>"111111110",
  54570=>"001001100",
  54571=>"000000111",
  54572=>"110111000",
  54573=>"000000100",
  54574=>"111011010",
  54575=>"000000000",
  54576=>"011011011",
  54577=>"111011000",
  54578=>"000000000",
  54579=>"110111111",
  54580=>"000000000",
  54581=>"111001011",
  54582=>"000000001",
  54583=>"111111111",
  54584=>"101111101",
  54585=>"001000001",
  54586=>"110000000",
  54587=>"111111111",
  54588=>"000111010",
  54589=>"000100110",
  54590=>"000110110",
  54591=>"000000000",
  54592=>"100000000",
  54593=>"000000000",
  54594=>"111010010",
  54595=>"000000101",
  54596=>"000110111",
  54597=>"111110000",
  54598=>"000000000",
  54599=>"111000000",
  54600=>"111011000",
  54601=>"110111000",
  54602=>"001111011",
  54603=>"100100111",
  54604=>"100000000",
  54605=>"000000000",
  54606=>"001001001",
  54607=>"000111011",
  54608=>"110110110",
  54609=>"010110110",
  54610=>"100100110",
  54611=>"000000111",
  54612=>"000000100",
  54613=>"011011001",
  54614=>"100000000",
  54615=>"001000111",
  54616=>"111110111",
  54617=>"000100111",
  54618=>"111111001",
  54619=>"000000000",
  54620=>"111111111",
  54621=>"111000111",
  54622=>"000000000",
  54623=>"111111010",
  54624=>"000100110",
  54625=>"100000000",
  54626=>"111111100",
  54627=>"000000100",
  54628=>"000110110",
  54629=>"000000000",
  54630=>"000000011",
  54631=>"000000000",
  54632=>"001001011",
  54633=>"011010100",
  54634=>"000000100",
  54635=>"111011111",
  54636=>"000001000",
  54637=>"100111111",
  54638=>"000000000",
  54639=>"100100100",
  54640=>"110111000",
  54641=>"010110110",
  54642=>"000111000",
  54643=>"011111111",
  54644=>"000000010",
  54645=>"110000000",
  54646=>"111110000",
  54647=>"100111111",
  54648=>"000000000",
  54649=>"000000000",
  54650=>"111111000",
  54651=>"000001001",
  54652=>"110110010",
  54653=>"111011000",
  54654=>"111111011",
  54655=>"000000000",
  54656=>"111111000",
  54657=>"000110111",
  54658=>"100000111",
  54659=>"000110010",
  54660=>"000000111",
  54661=>"111110000",
  54662=>"000001001",
  54663=>"000000111",
  54664=>"000010111",
  54665=>"111000000",
  54666=>"101101000",
  54667=>"111111000",
  54668=>"111111111",
  54669=>"001111001",
  54670=>"111111000",
  54671=>"000000110",
  54672=>"000000000",
  54673=>"000000111",
  54674=>"000101111",
  54675=>"011010110",
  54676=>"001001111",
  54677=>"000000000",
  54678=>"111111111",
  54679=>"000000000",
  54680=>"000111111",
  54681=>"110000000",
  54682=>"000000001",
  54683=>"000000111",
  54684=>"100100111",
  54685=>"111111111",
  54686=>"100000100",
  54687=>"111000000",
  54688=>"100000000",
  54689=>"111111000",
  54690=>"001001100",
  54691=>"010000000",
  54692=>"000100000",
  54693=>"000000000",
  54694=>"001001011",
  54695=>"000001011",
  54696=>"000000101",
  54697=>"111111001",
  54698=>"111011111",
  54699=>"000000111",
  54700=>"000000000",
  54701=>"100100011",
  54702=>"000000000",
  54703=>"111010010",
  54704=>"101101000",
  54705=>"100000000",
  54706=>"111111111",
  54707=>"111100000",
  54708=>"111111111",
  54709=>"001100110",
  54710=>"000000100",
  54711=>"111111001",
  54712=>"000000000",
  54713=>"111111111",
  54714=>"000000000",
  54715=>"111111011",
  54716=>"101111111",
  54717=>"110111000",
  54718=>"000000101",
  54719=>"100100100",
  54720=>"111111000",
  54721=>"010000100",
  54722=>"111111111",
  54723=>"010000111",
  54724=>"000001111",
  54725=>"111111110",
  54726=>"100101001",
  54727=>"000101101",
  54728=>"111000000",
  54729=>"001101101",
  54730=>"000101111",
  54731=>"110000000",
  54732=>"000000111",
  54733=>"001001001",
  54734=>"101101101",
  54735=>"000000000",
  54736=>"100100110",
  54737=>"011111011",
  54738=>"011011011",
  54739=>"111000000",
  54740=>"111111111",
  54741=>"000000000",
  54742=>"000000101",
  54743=>"001111111",
  54744=>"000000000",
  54745=>"000000000",
  54746=>"001011111",
  54747=>"111000000",
  54748=>"000000000",
  54749=>"001011111",
  54750=>"000000000",
  54751=>"100100000",
  54752=>"000001111",
  54753=>"001001000",
  54754=>"111111000",
  54755=>"111011000",
  54756=>"100110100",
  54757=>"111001000",
  54758=>"111111011",
  54759=>"000000011",
  54760=>"001000000",
  54761=>"000000100",
  54762=>"000010110",
  54763=>"101111111",
  54764=>"111111011",
  54765=>"011001011",
  54766=>"001001001",
  54767=>"111111001",
  54768=>"100101111",
  54769=>"111111111",
  54770=>"000001111",
  54771=>"000000101",
  54772=>"111111111",
  54773=>"000110110",
  54774=>"001000111",
  54775=>"000011001",
  54776=>"111111111",
  54777=>"001000010",
  54778=>"111000001",
  54779=>"011010000",
  54780=>"111110111",
  54781=>"000000001",
  54782=>"000011111",
  54783=>"111111111",
  54784=>"000001001",
  54785=>"001101101",
  54786=>"111100000",
  54787=>"111111111",
  54788=>"001101011",
  54789=>"011001001",
  54790=>"000011011",
  54791=>"111111111",
  54792=>"000000000",
  54793=>"111111111",
  54794=>"111111111",
  54795=>"000000111",
  54796=>"000000110",
  54797=>"000000000",
  54798=>"000100100",
  54799=>"000111001",
  54800=>"000000000",
  54801=>"001111111",
  54802=>"000000000",
  54803=>"111111111",
  54804=>"000000011",
  54805=>"010001000",
  54806=>"010000000",
  54807=>"101100100",
  54808=>"101000001",
  54809=>"101001011",
  54810=>"011011111",
  54811=>"111111100",
  54812=>"110000000",
  54813=>"001001000",
  54814=>"000011111",
  54815=>"000000001",
  54816=>"010000000",
  54817=>"000000111",
  54818=>"000000000",
  54819=>"111111111",
  54820=>"000000000",
  54821=>"000110000",
  54822=>"000000111",
  54823=>"000000011",
  54824=>"000100111",
  54825=>"000000000",
  54826=>"000000000",
  54827=>"111000100",
  54828=>"111111111",
  54829=>"111111111",
  54830=>"111000110",
  54831=>"000000000",
  54832=>"111111111",
  54833=>"000000000",
  54834=>"100110111",
  54835=>"110100100",
  54836=>"111111111",
  54837=>"111100110",
  54838=>"001000000",
  54839=>"101101111",
  54840=>"001011011",
  54841=>"000111111",
  54842=>"000000000",
  54843=>"000000000",
  54844=>"111111011",
  54845=>"000000000",
  54846=>"111111111",
  54847=>"101000101",
  54848=>"111111111",
  54849=>"011111100",
  54850=>"111111111",
  54851=>"011111000",
  54852=>"011000000",
  54853=>"000000110",
  54854=>"111111111",
  54855=>"000000000",
  54856=>"011111011",
  54857=>"000000000",
  54858=>"000000010",
  54859=>"001000000",
  54860=>"001000001",
  54861=>"000000000",
  54862=>"111100100",
  54863=>"100000000",
  54864=>"000000000",
  54865=>"111110000",
  54866=>"000001111",
  54867=>"001001111",
  54868=>"111100100",
  54869=>"001000000",
  54870=>"100110100",
  54871=>"111111101",
  54872=>"000000000",
  54873=>"111111011",
  54874=>"111111111",
  54875=>"000001001",
  54876=>"000110110",
  54877=>"000000111",
  54878=>"110111111",
  54879=>"110111111",
  54880=>"100000000",
  54881=>"011011111",
  54882=>"000000000",
  54883=>"111111111",
  54884=>"001111111",
  54885=>"110100111",
  54886=>"001011010",
  54887=>"000000000",
  54888=>"000000000",
  54889=>"001001111",
  54890=>"111111111",
  54891=>"001101000",
  54892=>"011011011",
  54893=>"010111111",
  54894=>"000111110",
  54895=>"000000000",
  54896=>"000111111",
  54897=>"000000000",
  54898=>"101100110",
  54899=>"000111111",
  54900=>"111111110",
  54901=>"000000000",
  54902=>"111000010",
  54903=>"000000000",
  54904=>"111111000",
  54905=>"000000111",
  54906=>"000100111",
  54907=>"111100100",
  54908=>"011011000",
  54909=>"100000000",
  54910=>"000011001",
  54911=>"001111111",
  54912=>"000011000",
  54913=>"010010010",
  54914=>"000000111",
  54915=>"111111100",
  54916=>"111000000",
  54917=>"111111000",
  54918=>"001001000",
  54919=>"000100110",
  54920=>"101001001",
  54921=>"111111111",
  54922=>"111111000",
  54923=>"001000000",
  54924=>"110011111",
  54925=>"000000000",
  54926=>"111010000",
  54927=>"110111110",
  54928=>"111111111",
  54929=>"100100111",
  54930=>"111001000",
  54931=>"110110000",
  54932=>"000000000",
  54933=>"000001111",
  54934=>"000000001",
  54935=>"001000000",
  54936=>"111111101",
  54937=>"111011111",
  54938=>"000000001",
  54939=>"101000100",
  54940=>"000000000",
  54941=>"111100101",
  54942=>"001000111",
  54943=>"011111011",
  54944=>"000000000",
  54945=>"011011011",
  54946=>"111111111",
  54947=>"000001000",
  54948=>"000000000",
  54949=>"111111111",
  54950=>"001000111",
  54951=>"101100111",
  54952=>"111011000",
  54953=>"000000100",
  54954=>"111111111",
  54955=>"111111111",
  54956=>"111111111",
  54957=>"101001000",
  54958=>"110010010",
  54959=>"001001000",
  54960=>"000011000",
  54961=>"111111100",
  54962=>"111111111",
  54963=>"111111111",
  54964=>"000000101",
  54965=>"001000000",
  54966=>"000000101",
  54967=>"111111000",
  54968=>"111111111",
  54969=>"111111000",
  54970=>"110110110",
  54971=>"100100000",
  54972=>"111111000",
  54973=>"100111111",
  54974=>"111000000",
  54975=>"000000111",
  54976=>"100000000",
  54977=>"011001000",
  54978=>"111111111",
  54979=>"000010110",
  54980=>"000000000",
  54981=>"000000000",
  54982=>"000000000",
  54983=>"100001111",
  54984=>"111110111",
  54985=>"111111111",
  54986=>"111111111",
  54987=>"000000000",
  54988=>"111111111",
  54989=>"111111111",
  54990=>"110100111",
  54991=>"111110000",
  54992=>"110111111",
  54993=>"000000000",
  54994=>"101101111",
  54995=>"000000000",
  54996=>"101001000",
  54997=>"111001100",
  54998=>"000000000",
  54999=>"101111111",
  55000=>"000001001",
  55001=>"100110010",
  55002=>"111001000",
  55003=>"001000000",
  55004=>"000000111",
  55005=>"001001001",
  55006=>"111111111",
  55007=>"000000011",
  55008=>"011111111",
  55009=>"000000000",
  55010=>"111111111",
  55011=>"111011000",
  55012=>"001000000",
  55013=>"000000001",
  55014=>"010010000",
  55015=>"111111111",
  55016=>"111000000",
  55017=>"001100100",
  55018=>"111110000",
  55019=>"000010001",
  55020=>"111111111",
  55021=>"000100111",
  55022=>"000000011",
  55023=>"110000111",
  55024=>"111010000",
  55025=>"000100000",
  55026=>"111001001",
  55027=>"010000000",
  55028=>"000010000",
  55029=>"001001111",
  55030=>"000000110",
  55031=>"001000000",
  55032=>"000000000",
  55033=>"000000000",
  55034=>"111111000",
  55035=>"111111111",
  55036=>"000000111",
  55037=>"101000001",
  55038=>"110000001",
  55039=>"000111111",
  55040=>"000010000",
  55041=>"001011111",
  55042=>"000000100",
  55043=>"010111111",
  55044=>"010111111",
  55045=>"111111100",
  55046=>"010011111",
  55047=>"111111011",
  55048=>"000000000",
  55049=>"111011000",
  55050=>"110000101",
  55051=>"000000111",
  55052=>"110000110",
  55053=>"111111111",
  55054=>"111111111",
  55055=>"111000000",
  55056=>"001001110",
  55057=>"111111111",
  55058=>"101101111",
  55059=>"111000000",
  55060=>"000000000",
  55061=>"111111111",
  55062=>"100100110",
  55063=>"111111000",
  55064=>"111111111",
  55065=>"000000000",
  55066=>"101110111",
  55067=>"000000000",
  55068=>"000000000",
  55069=>"111111001",
  55070=>"011010000",
  55071=>"000111111",
  55072=>"100100111",
  55073=>"111111111",
  55074=>"001001001",
  55075=>"111111111",
  55076=>"111101110",
  55077=>"000000110",
  55078=>"000000010",
  55079=>"111111111",
  55080=>"011111111",
  55081=>"000000000",
  55082=>"110100000",
  55083=>"111010011",
  55084=>"000001001",
  55085=>"011001001",
  55086=>"000110111",
  55087=>"100111000",
  55088=>"011111111",
  55089=>"111000000",
  55090=>"111111010",
  55091=>"010000111",
  55092=>"111111111",
  55093=>"000001000",
  55094=>"000000000",
  55095=>"000000000",
  55096=>"111111100",
  55097=>"001011011",
  55098=>"010110111",
  55099=>"000111000",
  55100=>"111111111",
  55101=>"111000111",
  55102=>"100110000",
  55103=>"000001111",
  55104=>"000001111",
  55105=>"100111111",
  55106=>"000000000",
  55107=>"111000000",
  55108=>"001001111",
  55109=>"101111101",
  55110=>"000000101",
  55111=>"000100110",
  55112=>"000100000",
  55113=>"000000001",
  55114=>"111101111",
  55115=>"000000010",
  55116=>"000000111",
  55117=>"111110111",
  55118=>"011111111",
  55119=>"100000100",
  55120=>"000000000",
  55121=>"011000001",
  55122=>"000000000",
  55123=>"000000000",
  55124=>"000000000",
  55125=>"100110110",
  55126=>"000001000",
  55127=>"111100111",
  55128=>"111110000",
  55129=>"000000000",
  55130=>"101101101",
  55131=>"111000000",
  55132=>"000000001",
  55133=>"000000000",
  55134=>"001101101",
  55135=>"111111111",
  55136=>"111101111",
  55137=>"111111111",
  55138=>"100111111",
  55139=>"000000000",
  55140=>"111111111",
  55141=>"000000100",
  55142=>"001111110",
  55143=>"111111111",
  55144=>"000100111",
  55145=>"000000000",
  55146=>"111111111",
  55147=>"111111111",
  55148=>"001001001",
  55149=>"111101100",
  55150=>"010000000",
  55151=>"111111111",
  55152=>"000000100",
  55153=>"111111110",
  55154=>"111111000",
  55155=>"000001001",
  55156=>"100100111",
  55157=>"000110111",
  55158=>"000000000",
  55159=>"000000000",
  55160=>"000000000",
  55161=>"000011000",
  55162=>"000000100",
  55163=>"110000100",
  55164=>"100000111",
  55165=>"111111010",
  55166=>"111110100",
  55167=>"000000000",
  55168=>"000001001",
  55169=>"000001101",
  55170=>"000000000",
  55171=>"110010000",
  55172=>"000011011",
  55173=>"110110110",
  55174=>"111000000",
  55175=>"000000000",
  55176=>"000111111",
  55177=>"011011011",
  55178=>"001001101",
  55179=>"111111101",
  55180=>"000000011",
  55181=>"100101100",
  55182=>"000100100",
  55183=>"111111000",
  55184=>"000000000",
  55185=>"000000111",
  55186=>"111000000",
  55187=>"111101011",
  55188=>"011000000",
  55189=>"000011011",
  55190=>"111110000",
  55191=>"001001000",
  55192=>"000000000",
  55193=>"111000110",
  55194=>"111111011",
  55195=>"000000000",
  55196=>"000000000",
  55197=>"111111110",
  55198=>"101000000",
  55199=>"000000000",
  55200=>"000000100",
  55201=>"000000110",
  55202=>"011111010",
  55203=>"111111111",
  55204=>"000000010",
  55205=>"111111111",
  55206=>"111100100",
  55207=>"111111111",
  55208=>"011011001",
  55209=>"000000100",
  55210=>"111110110",
  55211=>"000000010",
  55212=>"000101111",
  55213=>"000000000",
  55214=>"111111111",
  55215=>"110111111",
  55216=>"111111000",
  55217=>"111111010",
  55218=>"000000000",
  55219=>"111100101",
  55220=>"000010011",
  55221=>"011011010",
  55222=>"000010010",
  55223=>"111111111",
  55224=>"111011011",
  55225=>"111111111",
  55226=>"111111111",
  55227=>"000000000",
  55228=>"111111111",
  55229=>"010110010",
  55230=>"100100111",
  55231=>"110110000",
  55232=>"000000000",
  55233=>"000111111",
  55234=>"111111111",
  55235=>"110111111",
  55236=>"011010111",
  55237=>"111010111",
  55238=>"000000000",
  55239=>"001110111",
  55240=>"000000000",
  55241=>"000000000",
  55242=>"000000000",
  55243=>"111111111",
  55244=>"000011010",
  55245=>"001011111",
  55246=>"100000011",
  55247=>"000000000",
  55248=>"000000000",
  55249=>"000111111",
  55250=>"111111111",
  55251=>"000000100",
  55252=>"100000000",
  55253=>"111111111",
  55254=>"001001000",
  55255=>"000010001",
  55256=>"000111110",
  55257=>"111001101",
  55258=>"000000010",
  55259=>"111001111",
  55260=>"000000000",
  55261=>"000001111",
  55262=>"100100110",
  55263=>"000001001",
  55264=>"111111111",
  55265=>"100110111",
  55266=>"110111101",
  55267=>"000111111",
  55268=>"111111111",
  55269=>"111111001",
  55270=>"110110111",
  55271=>"111001000",
  55272=>"100100000",
  55273=>"000110101",
  55274=>"110000000",
  55275=>"111111111",
  55276=>"110110111",
  55277=>"111001001",
  55278=>"000000111",
  55279=>"001000000",
  55280=>"100000000",
  55281=>"111000100",
  55282=>"111100110",
  55283=>"101001111",
  55284=>"000000000",
  55285=>"111111111",
  55286=>"111101111",
  55287=>"000000000",
  55288=>"111011000",
  55289=>"110100110",
  55290=>"111111100",
  55291=>"111111111",
  55292=>"000000000",
  55293=>"111110111",
  55294=>"110111000",
  55295=>"000000000",
  55296=>"001001110",
  55297=>"000000100",
  55298=>"011001001",
  55299=>"111111001",
  55300=>"001100111",
  55301=>"000000000",
  55302=>"100000000",
  55303=>"011111111",
  55304=>"000000000",
  55305=>"011001011",
  55306=>"000101110",
  55307=>"001000100",
  55308=>"100100000",
  55309=>"100000001",
  55310=>"111111110",
  55311=>"110000100",
  55312=>"111110110",
  55313=>"111111111",
  55314=>"001000000",
  55315=>"000011111",
  55316=>"111111000",
  55317=>"000000111",
  55318=>"111000110",
  55319=>"110110000",
  55320=>"110011011",
  55321=>"100000001",
  55322=>"111111110",
  55323=>"100010010",
  55324=>"111001001",
  55325=>"100000000",
  55326=>"111111000",
  55327=>"111111000",
  55328=>"011111101",
  55329=>"101101001",
  55330=>"110000000",
  55331=>"110110110",
  55332=>"111000000",
  55333=>"000000011",
  55334=>"000000110",
  55335=>"000000111",
  55336=>"111111000",
  55337=>"000110111",
  55338=>"101001000",
  55339=>"000000110",
  55340=>"000000110",
  55341=>"000000000",
  55342=>"111111101",
  55343=>"000110111",
  55344=>"111111110",
  55345=>"001000000",
  55346=>"000000000",
  55347=>"000000000",
  55348=>"000000001",
  55349=>"111111111",
  55350=>"000110000",
  55351=>"011001001",
  55352=>"000000000",
  55353=>"000001111",
  55354=>"000000000",
  55355=>"111110000",
  55356=>"001001111",
  55357=>"110010000",
  55358=>"000000111",
  55359=>"111101111",
  55360=>"111111001",
  55361=>"111111111",
  55362=>"000000000",
  55363=>"111111000",
  55364=>"110110100",
  55365=>"000111111",
  55366=>"111011010",
  55367=>"001111111",
  55368=>"111000100",
  55369=>"011000000",
  55370=>"000000000",
  55371=>"111111111",
  55372=>"100100000",
  55373=>"111111110",
  55374=>"111000000",
  55375=>"111111111",
  55376=>"000000000",
  55377=>"111110110",
  55378=>"111110110",
  55379=>"100100000",
  55380=>"100101001",
  55381=>"110011011",
  55382=>"000010000",
  55383=>"100100101",
  55384=>"000000000",
  55385=>"001000000",
  55386=>"111111000",
  55387=>"111111111",
  55388=>"000000000",
  55389=>"111100100",
  55390=>"000000011",
  55391=>"111111111",
  55392=>"011000000",
  55393=>"110110000",
  55394=>"011011001",
  55395=>"000000110",
  55396=>"000000000",
  55397=>"000000111",
  55398=>"001001111",
  55399=>"000111101",
  55400=>"001001001",
  55401=>"101000000",
  55402=>"000000000",
  55403=>"111000000",
  55404=>"100000000",
  55405=>"000000000",
  55406=>"111111111",
  55407=>"010111111",
  55408=>"010110111",
  55409=>"000011111",
  55410=>"100100111",
  55411=>"000000000",
  55412=>"000000111",
  55413=>"111111110",
  55414=>"111111110",
  55415=>"111000000",
  55416=>"110000101",
  55417=>"001111111",
  55418=>"111110110",
  55419=>"000000010",
  55420=>"010011110",
  55421=>"000000000",
  55422=>"111111111",
  55423=>"110111111",
  55424=>"000000000",
  55425=>"111011111",
  55426=>"110000000",
  55427=>"111111111",
  55428=>"100111111",
  55429=>"111000000",
  55430=>"111011010",
  55431=>"111111110",
  55432=>"111000000",
  55433=>"000111111",
  55434=>"100000000",
  55435=>"000000100",
  55436=>"001111111",
  55437=>"000100000",
  55438=>"011000111",
  55439=>"001111110",
  55440=>"000000001",
  55441=>"001000000",
  55442=>"000001111",
  55443=>"111111000",
  55444=>"111111011",
  55445=>"110100000",
  55446=>"000001001",
  55447=>"111000001",
  55448=>"111000110",
  55449=>"011011000",
  55450=>"110000000",
  55451=>"011001001",
  55452=>"001000000",
  55453=>"001110100",
  55454=>"000001000",
  55455=>"111111111",
  55456=>"111111110",
  55457=>"011011011",
  55458=>"000000000",
  55459=>"111010000",
  55460=>"001101100",
  55461=>"111000000",
  55462=>"100100000",
  55463=>"000000011",
  55464=>"000000000",
  55465=>"111000000",
  55466=>"000000000",
  55467=>"111001111",
  55468=>"111111101",
  55469=>"110100101",
  55470=>"111111000",
  55471=>"111110000",
  55472=>"111111000",
  55473=>"000000000",
  55474=>"111001000",
  55475=>"000000000",
  55476=>"000111111",
  55477=>"100000100",
  55478=>"100000100",
  55479=>"000000000",
  55480=>"000000100",
  55481=>"000000000",
  55482=>"001111110",
  55483=>"111111110",
  55484=>"111010111",
  55485=>"111001000",
  55486=>"111000010",
  55487=>"111101001",
  55488=>"110000000",
  55489=>"000000000",
  55490=>"111011011",
  55491=>"000000101",
  55492=>"000000111",
  55493=>"101000111",
  55494=>"001111000",
  55495=>"000011111",
  55496=>"001000000",
  55497=>"000010111",
  55498=>"001011000",
  55499=>"000000001",
  55500=>"111001000",
  55501=>"111111000",
  55502=>"000100100",
  55503=>"111000000",
  55504=>"111000000",
  55505=>"000000000",
  55506=>"001001000",
  55507=>"000000011",
  55508=>"001001011",
  55509=>"110111000",
  55510=>"000111111",
  55511=>"010001000",
  55512=>"000100001",
  55513=>"111000000",
  55514=>"110111010",
  55515=>"000010000",
  55516=>"000000000",
  55517=>"001000000",
  55518=>"000110111",
  55519=>"000000110",
  55520=>"111111110",
  55521=>"111111111",
  55522=>"000011111",
  55523=>"000000000",
  55524=>"111111110",
  55525=>"111111011",
  55526=>"111111111",
  55527=>"111101110",
  55528=>"000000000",
  55529=>"000000100",
  55530=>"111100000",
  55531=>"000000000",
  55532=>"000000000",
  55533=>"000000011",
  55534=>"000111110",
  55535=>"000000000",
  55536=>"110111011",
  55537=>"111111111",
  55538=>"111000101",
  55539=>"101111110",
  55540=>"000000000",
  55541=>"111111111",
  55542=>"111011000",
  55543=>"011001111",
  55544=>"101001000",
  55545=>"000000000",
  55546=>"111001111",
  55547=>"111111000",
  55548=>"000000000",
  55549=>"001011011",
  55550=>"000000000",
  55551=>"101011111",
  55552=>"111111000",
  55553=>"000000100",
  55554=>"111111111",
  55555=>"000000110",
  55556=>"110111111",
  55557=>"000110111",
  55558=>"000111111",
  55559=>"000000000",
  55560=>"100000000",
  55561=>"101000000",
  55562=>"111111010",
  55563=>"111111000",
  55564=>"111011111",
  55565=>"011100101",
  55566=>"100110100",
  55567=>"111111111",
  55568=>"111111111",
  55569=>"001001000",
  55570=>"000001000",
  55571=>"111111000",
  55572=>"000000011",
  55573=>"000000001",
  55574=>"111111100",
  55575=>"000000101",
  55576=>"111111111",
  55577=>"000000000",
  55578=>"000000111",
  55579=>"000000000",
  55580=>"000001001",
  55581=>"000000000",
  55582=>"000000000",
  55583=>"000000010",
  55584=>"100100111",
  55585=>"111000000",
  55586=>"001011111",
  55587=>"111011000",
  55588=>"011110111",
  55589=>"100110110",
  55590=>"111111111",
  55591=>"000000000",
  55592=>"000000000",
  55593=>"010000110",
  55594=>"000000111",
  55595=>"000000111",
  55596=>"110000000",
  55597=>"000001011",
  55598=>"000111000",
  55599=>"000000101",
  55600=>"000011111",
  55601=>"101001111",
  55602=>"000000000",
  55603=>"010110111",
  55604=>"011001001",
  55605=>"101000100",
  55606=>"111111111",
  55607=>"000100111",
  55608=>"010110000",
  55609=>"000000001",
  55610=>"000000110",
  55611=>"111000010",
  55612=>"111111111",
  55613=>"111111000",
  55614=>"000000000",
  55615=>"000000111",
  55616=>"000000000",
  55617=>"001111101",
  55618=>"000000000",
  55619=>"111000000",
  55620=>"000111111",
  55621=>"111110110",
  55622=>"011000000",
  55623=>"100000000",
  55624=>"110000000",
  55625=>"010000010",
  55626=>"111110111",
  55627=>"000000001",
  55628=>"000000000",
  55629=>"111000000",
  55630=>"000000000",
  55631=>"100100111",
  55632=>"110111110",
  55633=>"000110110",
  55634=>"010111111",
  55635=>"000000000",
  55636=>"000001000",
  55637=>"011000000",
  55638=>"001111011",
  55639=>"111000111",
  55640=>"001000000",
  55641=>"000100110",
  55642=>"001100110",
  55643=>"111111111",
  55644=>"111100000",
  55645=>"000001011",
  55646=>"001000000",
  55647=>"110110000",
  55648=>"100111111",
  55649=>"000000000",
  55650=>"111111111",
  55651=>"111111000",
  55652=>"111111111",
  55653=>"111111111",
  55654=>"111001001",
  55655=>"111110110",
  55656=>"011001101",
  55657=>"000010000",
  55658=>"111111111",
  55659=>"000000011",
  55660=>"000000000",
  55661=>"000111111",
  55662=>"000000000",
  55663=>"000000000",
  55664=>"010000000",
  55665=>"111001000",
  55666=>"101111111",
  55667=>"111011011",
  55668=>"111110001",
  55669=>"110111111",
  55670=>"111111110",
  55671=>"000011111",
  55672=>"111111000",
  55673=>"000000111",
  55674=>"111010010",
  55675=>"110111011",
  55676=>"111101001",
  55677=>"111111110",
  55678=>"000000111",
  55679=>"111111111",
  55680=>"111111110",
  55681=>"101111101",
  55682=>"000111111",
  55683=>"000000110",
  55684=>"000111100",
  55685=>"000000011",
  55686=>"000000000",
  55687=>"000110111",
  55688=>"111010000",
  55689=>"000100000",
  55690=>"111100110",
  55691=>"000000001",
  55692=>"111111111",
  55693=>"011011111",
  55694=>"111111111",
  55695=>"000000100",
  55696=>"010000100",
  55697=>"000000000",
  55698=>"011001001",
  55699=>"111111111",
  55700=>"111001011",
  55701=>"000000000",
  55702=>"001100110",
  55703=>"000000100",
  55704=>"111111000",
  55705=>"101111110",
  55706=>"000000000",
  55707=>"001001011",
  55708=>"111111010",
  55709=>"011000000",
  55710=>"000001001",
  55711=>"100000100",
  55712=>"000110111",
  55713=>"110110111",
  55714=>"000000100",
  55715=>"000011111",
  55716=>"111111110",
  55717=>"111111111",
  55718=>"001000111",
  55719=>"111111011",
  55720=>"111110000",
  55721=>"000110111",
  55722=>"110000000",
  55723=>"001111111",
  55724=>"010001001",
  55725=>"111011100",
  55726=>"000000000",
  55727=>"000000111",
  55728=>"001001000",
  55729=>"011000000",
  55730=>"000000000",
  55731=>"100110110",
  55732=>"111110011",
  55733=>"000000000",
  55734=>"000000000",
  55735=>"100000001",
  55736=>"111101111",
  55737=>"000000000",
  55738=>"000000000",
  55739=>"001011111",
  55740=>"111111111",
  55741=>"000000001",
  55742=>"111111101",
  55743=>"111111101",
  55744=>"000100100",
  55745=>"111001111",
  55746=>"000000000",
  55747=>"001001000",
  55748=>"000110111",
  55749=>"100100111",
  55750=>"000000000",
  55751=>"000000100",
  55752=>"110110000",
  55753=>"111111111",
  55754=>"111000101",
  55755=>"000011001",
  55756=>"111000000",
  55757=>"000000101",
  55758=>"000110111",
  55759=>"110111111",
  55760=>"110000000",
  55761=>"101111011",
  55762=>"000000000",
  55763=>"000111111",
  55764=>"011111111",
  55765=>"111010000",
  55766=>"000000000",
  55767=>"011011000",
  55768=>"111100110",
  55769=>"010010010",
  55770=>"000000011",
  55771=>"000010010",
  55772=>"000000000",
  55773=>"100000010",
  55774=>"111111111",
  55775=>"111000000",
  55776=>"100000000",
  55777=>"000000011",
  55778=>"000000001",
  55779=>"111111000",
  55780=>"000000011",
  55781=>"000001000",
  55782=>"111001101",
  55783=>"000000000",
  55784=>"011001111",
  55785=>"111111100",
  55786=>"000000000",
  55787=>"101111110",
  55788=>"011111111",
  55789=>"101111011",
  55790=>"100111111",
  55791=>"000000010",
  55792=>"111111111",
  55793=>"000000111",
  55794=>"100111000",
  55795=>"000000000",
  55796=>"111110000",
  55797=>"010000000",
  55798=>"111111000",
  55799=>"111111100",
  55800=>"000000000",
  55801=>"000000001",
  55802=>"000000000",
  55803=>"111111011",
  55804=>"110110110",
  55805=>"111111110",
  55806=>"101000111",
  55807=>"111111001",
  55808=>"111111111",
  55809=>"000000000",
  55810=>"000000111",
  55811=>"111111000",
  55812=>"001001001",
  55813=>"011001100",
  55814=>"111111111",
  55815=>"111111101",
  55816=>"010000000",
  55817=>"111001001",
  55818=>"111111111",
  55819=>"000111111",
  55820=>"011011001",
  55821=>"100101111",
  55822=>"100100100",
  55823=>"000101101",
  55824=>"000000111",
  55825=>"011010110",
  55826=>"001000111",
  55827=>"111111111",
  55828=>"000111111",
  55829=>"110000000",
  55830=>"000000000",
  55831=>"011111111",
  55832=>"001000000",
  55833=>"111111111",
  55834=>"111111111",
  55835=>"111111100",
  55836=>"111111111",
  55837=>"000000111",
  55838=>"101100000",
  55839=>"000011111",
  55840=>"000000000",
  55841=>"111111111",
  55842=>"111111100",
  55843=>"000000000",
  55844=>"111111111",
  55845=>"000000111",
  55846=>"111111111",
  55847=>"100000000",
  55848=>"111111111",
  55849=>"000000000",
  55850=>"000101001",
  55851=>"111000000",
  55852=>"000000110",
  55853=>"111100000",
  55854=>"000000000",
  55855=>"100000000",
  55856=>"001001000",
  55857=>"101001001",
  55858=>"101101111",
  55859=>"110001000",
  55860=>"101110000",
  55861=>"000110111",
  55862=>"000001001",
  55863=>"000010111",
  55864=>"111111111",
  55865=>"111000111",
  55866=>"000000000",
  55867=>"111111110",
  55868=>"111111110",
  55869=>"101001001",
  55870=>"001001100",
  55871=>"000001111",
  55872=>"100111100",
  55873=>"101001111",
  55874=>"011001001",
  55875=>"111111000",
  55876=>"110110110",
  55877=>"011011010",
  55878=>"001000000",
  55879=>"111111111",
  55880=>"101111110",
  55881=>"000000000",
  55882=>"000000010",
  55883=>"111111000",
  55884=>"110111011",
  55885=>"000111111",
  55886=>"100000011",
  55887=>"010010000",
  55888=>"000000000",
  55889=>"101011011",
  55890=>"000010001",
  55891=>"010000000",
  55892=>"101001111",
  55893=>"000001000",
  55894=>"111011111",
  55895=>"010110010",
  55896=>"001001111",
  55897=>"000000000",
  55898=>"110110111",
  55899=>"000101110",
  55900=>"000000001",
  55901=>"000000001",
  55902=>"111111101",
  55903=>"000011001",
  55904=>"111111111",
  55905=>"110110111",
  55906=>"111111010",
  55907=>"100110110",
  55908=>"111100110",
  55909=>"000101111",
  55910=>"111010000",
  55911=>"111000001",
  55912=>"111110000",
  55913=>"000001001",
  55914=>"110000000",
  55915=>"110111111",
  55916=>"000101000",
  55917=>"000000100",
  55918=>"100100000",
  55919=>"111111111",
  55920=>"000010000",
  55921=>"111111000",
  55922=>"111010000",
  55923=>"010110010",
  55924=>"111101101",
  55925=>"011101111",
  55926=>"111111111",
  55927=>"001001001",
  55928=>"000100000",
  55929=>"000110011",
  55930=>"111000001",
  55931=>"000000000",
  55932=>"100100100",
  55933=>"001001110",
  55934=>"000001001",
  55935=>"110110000",
  55936=>"000000000",
  55937=>"000011001",
  55938=>"000000111",
  55939=>"100110110",
  55940=>"111111111",
  55941=>"111000000",
  55942=>"000001111",
  55943=>"111000000",
  55944=>"110010000",
  55945=>"000100111",
  55946=>"001001001",
  55947=>"110010000",
  55948=>"000001111",
  55949=>"111111110",
  55950=>"111000000",
  55951=>"000000000",
  55952=>"010000000",
  55953=>"101101001",
  55954=>"010110100",
  55955=>"110011001",
  55956=>"111101001",
  55957=>"000000000",
  55958=>"000000000",
  55959=>"000000000",
  55960=>"101000000",
  55961=>"001111111",
  55962=>"000000000",
  55963=>"111111111",
  55964=>"000010110",
  55965=>"000000111",
  55966=>"111110111",
  55967=>"001101111",
  55968=>"111111111",
  55969=>"000000000",
  55970=>"000100111",
  55971=>"000110000",
  55972=>"001011011",
  55973=>"111110111",
  55974=>"111111111",
  55975=>"000010001",
  55976=>"011111000",
  55977=>"101001011",
  55978=>"000000000",
  55979=>"101000000",
  55980=>"000000111",
  55981=>"111111111",
  55982=>"000101010",
  55983=>"011011111",
  55984=>"110010000",
  55985=>"110110101",
  55986=>"111111111",
  55987=>"000001001",
  55988=>"111101000",
  55989=>"010000000",
  55990=>"000000000",
  55991=>"000000000",
  55992=>"001001001",
  55993=>"100000000",
  55994=>"101001001",
  55995=>"000000100",
  55996=>"000000111",
  55997=>"111000000",
  55998=>"000000111",
  55999=>"000000000",
  56000=>"000110111",
  56001=>"001011111",
  56002=>"111111000",
  56003=>"000001111",
  56004=>"000000000",
  56005=>"000000111",
  56006=>"000000000",
  56007=>"101001101",
  56008=>"000010000",
  56009=>"000000001",
  56010=>"000000000",
  56011=>"001011000",
  56012=>"011110110",
  56013=>"110000000",
  56014=>"000000011",
  56015=>"000000000",
  56016=>"000110110",
  56017=>"000000000",
  56018=>"000000110",
  56019=>"001000000",
  56020=>"000000101",
  56021=>"110110100",
  56022=>"111110010",
  56023=>"111100110",
  56024=>"001111111",
  56025=>"111011000",
  56026=>"111111111",
  56027=>"000000001",
  56028=>"010110010",
  56029=>"000101000",
  56030=>"001001111",
  56031=>"000110110",
  56032=>"000111111",
  56033=>"111001001",
  56034=>"001000000",
  56035=>"000010010",
  56036=>"001011000",
  56037=>"001111001",
  56038=>"111111111",
  56039=>"001001000",
  56040=>"111110100",
  56041=>"111111111",
  56042=>"111111111",
  56043=>"101000000",
  56044=>"111110000",
  56045=>"110111111",
  56046=>"111111000",
  56047=>"001111000",
  56048=>"100000100",
  56049=>"000000000",
  56050=>"111111011",
  56051=>"000001001",
  56052=>"111101000",
  56053=>"001001000",
  56054=>"000111110",
  56055=>"001000000",
  56056=>"000000000",
  56057=>"000000000",
  56058=>"001001001",
  56059=>"111111111",
  56060=>"110110100",
  56061=>"011011001",
  56062=>"010111000",
  56063=>"111111111",
  56064=>"111111111",
  56065=>"001001001",
  56066=>"000000000",
  56067=>"001001000",
  56068=>"110010000",
  56069=>"101001000",
  56070=>"111111110",
  56071=>"000000100",
  56072=>"000000000",
  56073=>"000101000",
  56074=>"000010000",
  56075=>"000000011",
  56076=>"000000100",
  56077=>"110110010",
  56078=>"000000000",
  56079=>"000000000",
  56080=>"110000000",
  56081=>"111111111",
  56082=>"110000000",
  56083=>"000000000",
  56084=>"110110010",
  56085=>"111111100",
  56086=>"001011011",
  56087=>"000000101",
  56088=>"001111011",
  56089=>"111001101",
  56090=>"000111111",
  56091=>"000010110",
  56092=>"111111100",
  56093=>"000000000",
  56094=>"100110110",
  56095=>"011111000",
  56096=>"111011001",
  56097=>"100000001",
  56098=>"010010000",
  56099=>"111101111",
  56100=>"111001001",
  56101=>"001001000",
  56102=>"110111111",
  56103=>"011011001",
  56104=>"111111100",
  56105=>"000000000",
  56106=>"111010110",
  56107=>"000000101",
  56108=>"000010000",
  56109=>"110110000",
  56110=>"000001001",
  56111=>"100101000",
  56112=>"000000000",
  56113=>"111111111",
  56114=>"000110100",
  56115=>"010111011",
  56116=>"100000101",
  56117=>"011111100",
  56118=>"111000000",
  56119=>"000110110",
  56120=>"000000010",
  56121=>"111001001",
  56122=>"000001001",
  56123=>"110110111",
  56124=>"110110100",
  56125=>"011001001",
  56126=>"000001101",
  56127=>"010010010",
  56128=>"001001000",
  56129=>"110111001",
  56130=>"001001011",
  56131=>"111000000",
  56132=>"011111100",
  56133=>"111111111",
  56134=>"000000000",
  56135=>"001000000",
  56136=>"000000111",
  56137=>"110010000",
  56138=>"100000000",
  56139=>"001101100",
  56140=>"000111111",
  56141=>"010111111",
  56142=>"000100100",
  56143=>"101001101",
  56144=>"000000001",
  56145=>"100000000",
  56146=>"000000001",
  56147=>"000001101",
  56148=>"000000000",
  56149=>"011001001",
  56150=>"000010010",
  56151=>"000000000",
  56152=>"100000100",
  56153=>"011011011",
  56154=>"111011011",
  56155=>"001000100",
  56156=>"000010001",
  56157=>"001001001",
  56158=>"100000000",
  56159=>"000101110",
  56160=>"110111111",
  56161=>"000001101",
  56162=>"011000000",
  56163=>"111111111",
  56164=>"100110100",
  56165=>"000010000",
  56166=>"111011111",
  56167=>"111111100",
  56168=>"110111001",
  56169=>"111111001",
  56170=>"000100000",
  56171=>"100011111",
  56172=>"011011001",
  56173=>"000001000",
  56174=>"000000000",
  56175=>"000001111",
  56176=>"000000000",
  56177=>"000111111",
  56178=>"100000000",
  56179=>"100100001",
  56180=>"000000000",
  56181=>"011000000",
  56182=>"001000111",
  56183=>"111111111",
  56184=>"000100100",
  56185=>"101100111",
  56186=>"111111001",
  56187=>"000110111",
  56188=>"000000000",
  56189=>"010110001",
  56190=>"110110000",
  56191=>"101111101",
  56192=>"000000000",
  56193=>"110110111",
  56194=>"110111111",
  56195=>"000000000",
  56196=>"011010111",
  56197=>"010110010",
  56198=>"001001001",
  56199=>"010110110",
  56200=>"000000000",
  56201=>"111111010",
  56202=>"001000000",
  56203=>"111001111",
  56204=>"111110100",
  56205=>"110110110",
  56206=>"110110000",
  56207=>"000000001",
  56208=>"000000001",
  56209=>"000000000",
  56210=>"000000000",
  56211=>"011001001",
  56212=>"010010010",
  56213=>"010010000",
  56214=>"000001011",
  56215=>"001001001",
  56216=>"100101000",
  56217=>"111110000",
  56218=>"000000000",
  56219=>"000111111",
  56220=>"000000000",
  56221=>"000100000",
  56222=>"000000000",
  56223=>"000110110",
  56224=>"111111111",
  56225=>"011011011",
  56226=>"000000000",
  56227=>"000000001",
  56228=>"101001000",
  56229=>"110111110",
  56230=>"001000000",
  56231=>"000110111",
  56232=>"000010000",
  56233=>"010110110",
  56234=>"000001111",
  56235=>"000000000",
  56236=>"000000100",
  56237=>"000001001",
  56238=>"111101001",
  56239=>"111011000",
  56240=>"111111110",
  56241=>"000000001",
  56242=>"001001000",
  56243=>"000000000",
  56244=>"111111010",
  56245=>"001001000",
  56246=>"101111111",
  56247=>"011010000",
  56248=>"101011111",
  56249=>"110110111",
  56250=>"011011111",
  56251=>"001000111",
  56252=>"100111111",
  56253=>"000001000",
  56254=>"101000101",
  56255=>"001011011",
  56256=>"000000000",
  56257=>"101000000",
  56258=>"001001111",
  56259=>"000110100",
  56260=>"011000110",
  56261=>"110111111",
  56262=>"100101101",
  56263=>"111101000",
  56264=>"001000000",
  56265=>"000011111",
  56266=>"000001000",
  56267=>"000000000",
  56268=>"111000000",
  56269=>"111111101",
  56270=>"000110110",
  56271=>"000000000",
  56272=>"100110111",
  56273=>"000000000",
  56274=>"000000000",
  56275=>"111101001",
  56276=>"001011011",
  56277=>"000000100",
  56278=>"111010000",
  56279=>"100000001",
  56280=>"111111011",
  56281=>"010010000",
  56282=>"001111010",
  56283=>"001000000",
  56284=>"110111111",
  56285=>"100111111",
  56286=>"111111111",
  56287=>"000000001",
  56288=>"101000111",
  56289=>"110100000",
  56290=>"010111010",
  56291=>"110111110",
  56292=>"010011110",
  56293=>"101000101",
  56294=>"001000000",
  56295=>"000000001",
  56296=>"100100000",
  56297=>"000000000",
  56298=>"111000000",
  56299=>"000000000",
  56300=>"001111111",
  56301=>"001101101",
  56302=>"111000000",
  56303=>"001101101",
  56304=>"001001101",
  56305=>"000110111",
  56306=>"000000000",
  56307=>"100100100",
  56308=>"100100000",
  56309=>"111001001",
  56310=>"110110110",
  56311=>"101100111",
  56312=>"001001000",
  56313=>"100110111",
  56314=>"011001000",
  56315=>"000011011",
  56316=>"111100111",
  56317=>"001001001",
  56318=>"000001010",
  56319=>"111001001",
  56320=>"001001010",
  56321=>"000000000",
  56322=>"000000000",
  56323=>"001001111",
  56324=>"001111111",
  56325=>"010111010",
  56326=>"010111111",
  56327=>"111111111",
  56328=>"000000011",
  56329=>"000000000",
  56330=>"000000000",
  56331=>"000000000",
  56332=>"000000110",
  56333=>"110000111",
  56334=>"000011111",
  56335=>"010011111",
  56336=>"001001000",
  56337=>"000000000",
  56338=>"101100000",
  56339=>"000000000",
  56340=>"111111101",
  56341=>"111111000",
  56342=>"111111111",
  56343=>"000101001",
  56344=>"111001001",
  56345=>"100100111",
  56346=>"010110111",
  56347=>"000000000",
  56348=>"010011000",
  56349=>"111111000",
  56350=>"110100000",
  56351=>"110011100",
  56352=>"110111111",
  56353=>"000100000",
  56354=>"000110110",
  56355=>"111111110",
  56356=>"000001011",
  56357=>"011111111",
  56358=>"000000000",
  56359=>"000000000",
  56360=>"111111111",
  56361=>"000000111",
  56362=>"011001001",
  56363=>"111111000",
  56364=>"100000111",
  56365=>"010000010",
  56366=>"011011001",
  56367=>"000111111",
  56368=>"000000100",
  56369=>"000111111",
  56370=>"111111010",
  56371=>"000000000",
  56372=>"110110010",
  56373=>"110101110",
  56374=>"011000000",
  56375=>"101111111",
  56376=>"000000111",
  56377=>"001000000",
  56378=>"001111111",
  56379=>"111111101",
  56380=>"111111111",
  56381=>"000000111",
  56382=>"011111111",
  56383=>"100000100",
  56384=>"111001111",
  56385=>"011011011",
  56386=>"000000000",
  56387=>"000000010",
  56388=>"111100111",
  56389=>"111000100",
  56390=>"101000000",
  56391=>"111111100",
  56392=>"111001000",
  56393=>"111000000",
  56394=>"111111110",
  56395=>"101000000",
  56396=>"000000000",
  56397=>"110100111",
  56398=>"000000000",
  56399=>"000000111",
  56400=>"110111111",
  56401=>"111001000",
  56402=>"000000000",
  56403=>"000100110",
  56404=>"100000000",
  56405=>"111000001",
  56406=>"000000111",
  56407=>"000000000",
  56408=>"110111111",
  56409=>"111101001",
  56410=>"111111111",
  56411=>"011110110",
  56412=>"000111011",
  56413=>"000000000",
  56414=>"001000000",
  56415=>"111111111",
  56416=>"111111000",
  56417=>"010000000",
  56418=>"000000000",
  56419=>"000000000",
  56420=>"111111000",
  56421=>"100100101",
  56422=>"000100101",
  56423=>"111111111",
  56424=>"111111011",
  56425=>"111010110",
  56426=>"111111111",
  56427=>"000000000",
  56428=>"000111111",
  56429=>"111111000",
  56430=>"001000000",
  56431=>"110100000",
  56432=>"011111111",
  56433=>"000000111",
  56434=>"111111011",
  56435=>"111110111",
  56436=>"000000000",
  56437=>"000000000",
  56438=>"000000000",
  56439=>"000100000",
  56440=>"111000001",
  56441=>"111111111",
  56442=>"001000000",
  56443=>"000111111",
  56444=>"000000000",
  56445=>"000000101",
  56446=>"111001001",
  56447=>"000000000",
  56448=>"000000000",
  56449=>"111111001",
  56450=>"101100100",
  56451=>"001011111",
  56452=>"000000000",
  56453=>"000000111",
  56454=>"111111100",
  56455=>"010000111",
  56456=>"110100000",
  56457=>"000000000",
  56458=>"000000111",
  56459=>"111111111",
  56460=>"000010110",
  56461=>"111111111",
  56462=>"111001000",
  56463=>"111111111",
  56464=>"111001101",
  56465=>"000000111",
  56466=>"111111111",
  56467=>"000000111",
  56468=>"000000000",
  56469=>"111100000",
  56470=>"100101000",
  56471=>"000000000",
  56472=>"000000000",
  56473=>"000000000",
  56474=>"010111111",
  56475=>"111001001",
  56476=>"100000000",
  56477=>"011000000",
  56478=>"110111011",
  56479=>"111110110",
  56480=>"000000111",
  56481=>"001000000",
  56482=>"101001000",
  56483=>"100000110",
  56484=>"110111111",
  56485=>"001000000",
  56486=>"000000000",
  56487=>"011011101",
  56488=>"111110111",
  56489=>"000000100",
  56490=>"000000000",
  56491=>"000000100",
  56492=>"100101111",
  56493=>"111110100",
  56494=>"110111111",
  56495=>"111111111",
  56496=>"111011011",
  56497=>"110100111",
  56498=>"111111111",
  56499=>"000000000",
  56500=>"100010001",
  56501=>"000000000",
  56502=>"111111111",
  56503=>"111111110",
  56504=>"111100000",
  56505=>"111111000",
  56506=>"001001000",
  56507=>"100001000",
  56508=>"001101111",
  56509=>"000000000",
  56510=>"111100110",
  56511=>"111011000",
  56512=>"111011010",
  56513=>"101001001",
  56514=>"000000000",
  56515=>"011000000",
  56516=>"001001111",
  56517=>"101001000",
  56518=>"111111111",
  56519=>"010110110",
  56520=>"111111111",
  56521=>"111001111",
  56522=>"000000111",
  56523=>"100001000",
  56524=>"000000001",
  56525=>"111111110",
  56526=>"000000000",
  56527=>"000000000",
  56528=>"111010000",
  56529=>"111001110",
  56530=>"000011111",
  56531=>"111000000",
  56532=>"001001000",
  56533=>"000110111",
  56534=>"000000000",
  56535=>"000001111",
  56536=>"011010000",
  56537=>"000000001",
  56538=>"111111111",
  56539=>"000000111",
  56540=>"100100110",
  56541=>"000000000",
  56542=>"011000110",
  56543=>"100100111",
  56544=>"000000000",
  56545=>"011110110",
  56546=>"100000101",
  56547=>"000100101",
  56548=>"111111010",
  56549=>"111001001",
  56550=>"000000011",
  56551=>"101110111",
  56552=>"101001000",
  56553=>"111010000",
  56554=>"101000111",
  56555=>"100111111",
  56556=>"011011101",
  56557=>"000100111",
  56558=>"000001000",
  56559=>"111111100",
  56560=>"000000000",
  56561=>"111101111",
  56562=>"110111111",
  56563=>"000010111",
  56564=>"010010010",
  56565=>"111111111",
  56566=>"111101100",
  56567=>"111011111",
  56568=>"111111111",
  56569=>"100000000",
  56570=>"001010011",
  56571=>"111111000",
  56572=>"111111110",
  56573=>"000000100",
  56574=>"110111111",
  56575=>"000000000",
  56576=>"100000000",
  56577=>"111111000",
  56578=>"000000010",
  56579=>"000000000",
  56580=>"000010110",
  56581=>"011000100",
  56582=>"111110110",
  56583=>"000000110",
  56584=>"000000000",
  56585=>"000000000",
  56586=>"001011111",
  56587=>"110111111",
  56588=>"111111100",
  56589=>"001000000",
  56590=>"111111111",
  56591=>"111000010",
  56592=>"011011011",
  56593=>"000010111",
  56594=>"010000000",
  56595=>"000000000",
  56596=>"111000111",
  56597=>"111111101",
  56598=>"100110111",
  56599=>"100000000",
  56600=>"111111110",
  56601=>"011011111",
  56602=>"111111000",
  56603=>"100000000",
  56604=>"111111111",
  56605=>"111111011",
  56606=>"000000000",
  56607=>"000111110",
  56608=>"110111001",
  56609=>"111111001",
  56610=>"111000100",
  56611=>"000000111",
  56612=>"010110110",
  56613=>"000000100",
  56614=>"000111111",
  56615=>"111111000",
  56616=>"111111111",
  56617=>"111111111",
  56618=>"001010010",
  56619=>"101111011",
  56620=>"001000000",
  56621=>"000100110",
  56622=>"000000111",
  56623=>"011111110",
  56624=>"000111011",
  56625=>"100000001",
  56626=>"111000000",
  56627=>"010010110",
  56628=>"000000100",
  56629=>"000000011",
  56630=>"000000000",
  56631=>"101100000",
  56632=>"000010000",
  56633=>"000000111",
  56634=>"000000000",
  56635=>"000000001",
  56636=>"111101100",
  56637=>"001001101",
  56638=>"001001101",
  56639=>"100111011",
  56640=>"001000000",
  56641=>"001000001",
  56642=>"111111111",
  56643=>"001011001",
  56644=>"110110110",
  56645=>"111111011",
  56646=>"111001001",
  56647=>"000000111",
  56648=>"000100000",
  56649=>"000000000",
  56650=>"001110111",
  56651=>"000111011",
  56652=>"000000000",
  56653=>"111000000",
  56654=>"001111111",
  56655=>"001001000",
  56656=>"110101111",
  56657=>"111111111",
  56658=>"111111111",
  56659=>"111110100",
  56660=>"000000110",
  56661=>"011001011",
  56662=>"000010110",
  56663=>"111011011",
  56664=>"001001001",
  56665=>"111000000",
  56666=>"111111100",
  56667=>"111111010",
  56668=>"000000000",
  56669=>"000110111",
  56670=>"110000010",
  56671=>"101101011",
  56672=>"111111000",
  56673=>"111111000",
  56674=>"011011100",
  56675=>"111111111",
  56676=>"111111111",
  56677=>"000000000",
  56678=>"111111111",
  56679=>"001001011",
  56680=>"000100100",
  56681=>"111111111",
  56682=>"000000000",
  56683=>"111111100",
  56684=>"000000100",
  56685=>"111101000",
  56686=>"111111010",
  56687=>"000000100",
  56688=>"000100100",
  56689=>"100000000",
  56690=>"111001111",
  56691=>"000000010",
  56692=>"111011011",
  56693=>"000000000",
  56694=>"000000000",
  56695=>"111001001",
  56696=>"111111111",
  56697=>"110111010",
  56698=>"000000100",
  56699=>"100100110",
  56700=>"111111000",
  56701=>"000000000",
  56702=>"110110110",
  56703=>"100100000",
  56704=>"000011011",
  56705=>"000000100",
  56706=>"000001001",
  56707=>"111011111",
  56708=>"111000000",
  56709=>"111001001",
  56710=>"000000000",
  56711=>"001111000",
  56712=>"111111111",
  56713=>"111111111",
  56714=>"001000000",
  56715=>"010000001",
  56716=>"111111111",
  56717=>"000101101",
  56718=>"010110100",
  56719=>"000000111",
  56720=>"000000000",
  56721=>"111001000",
  56722=>"000011000",
  56723=>"000000100",
  56724=>"111111000",
  56725=>"000010010",
  56726=>"111001000",
  56727=>"001001111",
  56728=>"111111110",
  56729=>"101111110",
  56730=>"100001000",
  56731=>"000000111",
  56732=>"100000101",
  56733=>"000000111",
  56734=>"100100101",
  56735=>"000110110",
  56736=>"000000000",
  56737=>"000000001",
  56738=>"010010111",
  56739=>"111111111",
  56740=>"000000000",
  56741=>"111111011",
  56742=>"000000000",
  56743=>"011111111",
  56744=>"000001111",
  56745=>"000001001",
  56746=>"110111111",
  56747=>"000000110",
  56748=>"001000000",
  56749=>"101101111",
  56750=>"000100111",
  56751=>"111111110",
  56752=>"001111111",
  56753=>"010010010",
  56754=>"000010111",
  56755=>"000000000",
  56756=>"011011000",
  56757=>"000000100",
  56758=>"000000000",
  56759=>"111000001",
  56760=>"111111001",
  56761=>"111111000",
  56762=>"000110000",
  56763=>"111111111",
  56764=>"000000100",
  56765=>"111111111",
  56766=>"111111000",
  56767=>"111101101",
  56768=>"111111111",
  56769=>"111111111",
  56770=>"111000000",
  56771=>"111111111",
  56772=>"000000111",
  56773=>"000000100",
  56774=>"111111011",
  56775=>"111111000",
  56776=>"000000000",
  56777=>"111111000",
  56778=>"001111111",
  56779=>"000101101",
  56780=>"111111000",
  56781=>"111011100",
  56782=>"111001110",
  56783=>"111111110",
  56784=>"010111111",
  56785=>"110110100",
  56786=>"011000011",
  56787=>"111000001",
  56788=>"001011111",
  56789=>"000000000",
  56790=>"000000111",
  56791=>"000000011",
  56792=>"000000001",
  56793=>"110111111",
  56794=>"000100111",
  56795=>"111111011",
  56796=>"000000000",
  56797=>"000000000",
  56798=>"000000100",
  56799=>"000100000",
  56800=>"000000110",
  56801=>"111111100",
  56802=>"011010000",
  56803=>"000000110",
  56804=>"111111111",
  56805=>"111111101",
  56806=>"111111111",
  56807=>"000000100",
  56808=>"110110111",
  56809=>"111011011",
  56810=>"111111110",
  56811=>"000000000",
  56812=>"001010111",
  56813=>"001011100",
  56814=>"000000000",
  56815=>"111111111",
  56816=>"000000000",
  56817=>"110000000",
  56818=>"001000000",
  56819=>"000011011",
  56820=>"111111111",
  56821=>"110111111",
  56822=>"000000100",
  56823=>"000000110",
  56824=>"011011000",
  56825=>"111111111",
  56826=>"000000111",
  56827=>"111000000",
  56828=>"000000100",
  56829=>"101110111",
  56830=>"000000000",
  56831=>"000000000",
  56832=>"000000000",
  56833=>"111001000",
  56834=>"000000000",
  56835=>"000000011",
  56836=>"111111111",
  56837=>"000000001",
  56838=>"000000000",
  56839=>"111000100",
  56840=>"011111111",
  56841=>"011001001",
  56842=>"000000001",
  56843=>"000010001",
  56844=>"001000000",
  56845=>"010110000",
  56846=>"000000010",
  56847=>"101001111",
  56848=>"000000000",
  56849=>"110011111",
  56850=>"001101111",
  56851=>"111101000",
  56852=>"111111111",
  56853=>"000000000",
  56854=>"111111111",
  56855=>"111111111",
  56856=>"110111110",
  56857=>"101111011",
  56858=>"111001001",
  56859=>"100001001",
  56860=>"100000000",
  56861=>"111111001",
  56862=>"000000101",
  56863=>"010010010",
  56864=>"101101100",
  56865=>"110111010",
  56866=>"000000110",
  56867=>"000100001",
  56868=>"111111111",
  56869=>"000000111",
  56870=>"111101011",
  56871=>"111111110",
  56872=>"000000000",
  56873=>"111011011",
  56874=>"011001000",
  56875=>"110111111",
  56876=>"001001111",
  56877=>"111010111",
  56878=>"110000011",
  56879=>"111011001",
  56880=>"110110000",
  56881=>"000000001",
  56882=>"000110000",
  56883=>"011111011",
  56884=>"000000100",
  56885=>"000000000",
  56886=>"000000000",
  56887=>"011001001",
  56888=>"011000110",
  56889=>"000000000",
  56890=>"110111110",
  56891=>"111010000",
  56892=>"110100100",
  56893=>"000000110",
  56894=>"000000011",
  56895=>"111000000",
  56896=>"000000000",
  56897=>"000000000",
  56898=>"101111111",
  56899=>"111111111",
  56900=>"110111110",
  56901=>"110110100",
  56902=>"111000000",
  56903=>"111100000",
  56904=>"111111100",
  56905=>"000000000",
  56906=>"111111111",
  56907=>"111111100",
  56908=>"000000000",
  56909=>"000000111",
  56910=>"000111111",
  56911=>"000000000",
  56912=>"000000111",
  56913=>"010110111",
  56914=>"000011010",
  56915=>"101101100",
  56916=>"000111100",
  56917=>"010110000",
  56918=>"001000000",
  56919=>"111111010",
  56920=>"111010000",
  56921=>"100000000",
  56922=>"011011001",
  56923=>"001001000",
  56924=>"000000000",
  56925=>"000000000",
  56926=>"011010110",
  56927=>"100111000",
  56928=>"100001100",
  56929=>"111110000",
  56930=>"111001000",
  56931=>"100000000",
  56932=>"100000000",
  56933=>"111000000",
  56934=>"111001011",
  56935=>"111011000",
  56936=>"000000111",
  56937=>"000000100",
  56938=>"001000000",
  56939=>"111111111",
  56940=>"000110110",
  56941=>"111111111",
  56942=>"001101111",
  56943=>"010010000",
  56944=>"110111010",
  56945=>"000000100",
  56946=>"110100110",
  56947=>"000000000",
  56948=>"000000101",
  56949=>"011001000",
  56950=>"111111111",
  56951=>"000000001",
  56952=>"000110100",
  56953=>"111100000",
  56954=>"111001000",
  56955=>"000000111",
  56956=>"100110110",
  56957=>"000000011",
  56958=>"111110100",
  56959=>"110110011",
  56960=>"101101001",
  56961=>"000000111",
  56962=>"111111001",
  56963=>"111111100",
  56964=>"111101011",
  56965=>"111000100",
  56966=>"000000001",
  56967=>"111101101",
  56968=>"010000000",
  56969=>"010000011",
  56970=>"100111010",
  56971=>"111111001",
  56972=>"000000000",
  56973=>"000000000",
  56974=>"100100101",
  56975=>"000000000",
  56976=>"111011010",
  56977=>"110110010",
  56978=>"000000001",
  56979=>"111111111",
  56980=>"000000000",
  56981=>"111001000",
  56982=>"111111111",
  56983=>"000000000",
  56984=>"000011001",
  56985=>"000000000",
  56986=>"000000000",
  56987=>"111000000",
  56988=>"011011010",
  56989=>"000001001",
  56990=>"110111111",
  56991=>"000001011",
  56992=>"000000000",
  56993=>"000110111",
  56994=>"000000000",
  56995=>"000000010",
  56996=>"001001001",
  56997=>"010110110",
  56998=>"101000000",
  56999=>"010011111",
  57000=>"001001001",
  57001=>"000000000",
  57002=>"001000001",
  57003=>"110100000",
  57004=>"111111111",
  57005=>"101111111",
  57006=>"000000000",
  57007=>"110001000",
  57008=>"111110010",
  57009=>"000000110",
  57010=>"111111110",
  57011=>"110000000",
  57012=>"001001001",
  57013=>"000111111",
  57014=>"110111110",
  57015=>"011111111",
  57016=>"000000000",
  57017=>"101111111",
  57018=>"111001111",
  57019=>"000010110",
  57020=>"001000001",
  57021=>"110100111",
  57022=>"110110000",
  57023=>"011011001",
  57024=>"000000000",
  57025=>"111111100",
  57026=>"001011011",
  57027=>"000111111",
  57028=>"111111111",
  57029=>"001000000",
  57030=>"011111111",
  57031=>"111111111",
  57032=>"001001000",
  57033=>"000000000",
  57034=>"000000000",
  57035=>"111111111",
  57036=>"000110111",
  57037=>"000000001",
  57038=>"010010111",
  57039=>"111001001",
  57040=>"111111000",
  57041=>"111111111",
  57042=>"111000000",
  57043=>"000000010",
  57044=>"100000100",
  57045=>"000000110",
  57046=>"000001011",
  57047=>"000001010",
  57048=>"010010110",
  57049=>"010000000",
  57050=>"000000001",
  57051=>"110110110",
  57052=>"000000000",
  57053=>"000001111",
  57054=>"000000000",
  57055=>"111111000",
  57056=>"000000111",
  57057=>"010110000",
  57058=>"011010000",
  57059=>"011011111",
  57060=>"000101100",
  57061=>"000000000",
  57062=>"000000001",
  57063=>"111111111",
  57064=>"111001000",
  57065=>"111011000",
  57066=>"100100100",
  57067=>"001000000",
  57068=>"000000000",
  57069=>"011000000",
  57070=>"001000011",
  57071=>"111111000",
  57072=>"111110101",
  57073=>"111111000",
  57074=>"110000000",
  57075=>"000000000",
  57076=>"011000001",
  57077=>"001001000",
  57078=>"000000011",
  57079=>"000111111",
  57080=>"111111111",
  57081=>"001001111",
  57082=>"000000000",
  57083=>"000000000",
  57084=>"000000110",
  57085=>"100111000",
  57086=>"001000000",
  57087=>"000000001",
  57088=>"000000100",
  57089=>"011011011",
  57090=>"111111111",
  57091=>"111111011",
  57092=>"000000000",
  57093=>"100111111",
  57094=>"000000100",
  57095=>"111111111",
  57096=>"101111111",
  57097=>"000000111",
  57098=>"000111011",
  57099=>"111111111",
  57100=>"000000100",
  57101=>"111111111",
  57102=>"110110110",
  57103=>"000000000",
  57104=>"000011110",
  57105=>"100110000",
  57106=>"011000000",
  57107=>"010111111",
  57108=>"100001111",
  57109=>"111010010",
  57110=>"011111111",
  57111=>"111110000",
  57112=>"110100000",
  57113=>"010000011",
  57114=>"000000001",
  57115=>"011001000",
  57116=>"100110100",
  57117=>"111111111",
  57118=>"000000110",
  57119=>"001000000",
  57120=>"111111000",
  57121=>"000011111",
  57122=>"110000000",
  57123=>"111111111",
  57124=>"101001001",
  57125=>"000000001",
  57126=>"110100000",
  57127=>"000001111",
  57128=>"111111111",
  57129=>"011001001",
  57130=>"100000000",
  57131=>"011110110",
  57132=>"101111000",
  57133=>"000000100",
  57134=>"111111111",
  57135=>"000000000",
  57136=>"000000101",
  57137=>"000001011",
  57138=>"001000000",
  57139=>"000001111",
  57140=>"111101000",
  57141=>"100000111",
  57142=>"000001000",
  57143=>"000000100",
  57144=>"111011001",
  57145=>"000000111",
  57146=>"011011010",
  57147=>"111011111",
  57148=>"000001011",
  57149=>"000000000",
  57150=>"000000000",
  57151=>"000111100",
  57152=>"000000000",
  57153=>"000000000",
  57154=>"000000000",
  57155=>"000000000",
  57156=>"111111000",
  57157=>"000000000",
  57158=>"111001000",
  57159=>"111111111",
  57160=>"000001011",
  57161=>"110000000",
  57162=>"101001001",
  57163=>"111000000",
  57164=>"011001111",
  57165=>"000000000",
  57166=>"011000000",
  57167=>"101101000",
  57168=>"000000101",
  57169=>"000100100",
  57170=>"111111000",
  57171=>"111011011",
  57172=>"001001000",
  57173=>"011011011",
  57174=>"111111111",
  57175=>"000000101",
  57176=>"000000111",
  57177=>"111101100",
  57178=>"101101000",
  57179=>"100000000",
  57180=>"000000000",
  57181=>"000000000",
  57182=>"000000110",
  57183=>"111111110",
  57184=>"110000000",
  57185=>"000000000",
  57186=>"111100000",
  57187=>"101000101",
  57188=>"111111111",
  57189=>"001000000",
  57190=>"111001000",
  57191=>"111110100",
  57192=>"001001001",
  57193=>"000000001",
  57194=>"000000000",
  57195=>"000110111",
  57196=>"110111110",
  57197=>"100111111",
  57198=>"000001111",
  57199=>"010111100",
  57200=>"001001001",
  57201=>"000011010",
  57202=>"111111111",
  57203=>"110000100",
  57204=>"011011011",
  57205=>"100000000",
  57206=>"000000100",
  57207=>"000000000",
  57208=>"111101111",
  57209=>"011110110",
  57210=>"001000111",
  57211=>"011011011",
  57212=>"111011000",
  57213=>"111111110",
  57214=>"001001000",
  57215=>"000000101",
  57216=>"100100000",
  57217=>"000010000",
  57218=>"011010000",
  57219=>"110111111",
  57220=>"011000000",
  57221=>"000110110",
  57222=>"000111111",
  57223=>"000000111",
  57224=>"000000111",
  57225=>"100000000",
  57226=>"000000111",
  57227=>"000000000",
  57228=>"111100111",
  57229=>"011111110",
  57230=>"010110110",
  57231=>"011000000",
  57232=>"000000000",
  57233=>"111111000",
  57234=>"111111110",
  57235=>"000010011",
  57236=>"111111111",
  57237=>"010010000",
  57238=>"000000000",
  57239=>"111111110",
  57240=>"111111110",
  57241=>"000001001",
  57242=>"000000101",
  57243=>"111111010",
  57244=>"001011001",
  57245=>"000000000",
  57246=>"111001111",
  57247=>"000000000",
  57248=>"001011011",
  57249=>"010010000",
  57250=>"100100111",
  57251=>"000111111",
  57252=>"110000000",
  57253=>"111011111",
  57254=>"111111110",
  57255=>"000000000",
  57256=>"000000000",
  57257=>"100000000",
  57258=>"000100000",
  57259=>"111000000",
  57260=>"111001001",
  57261=>"001000000",
  57262=>"011111110",
  57263=>"111011000",
  57264=>"000100110",
  57265=>"011111001",
  57266=>"000111111",
  57267=>"000000111",
  57268=>"101111111",
  57269=>"000001100",
  57270=>"101000100",
  57271=>"111000000",
  57272=>"111000000",
  57273=>"000011001",
  57274=>"101101001",
  57275=>"000000001",
  57276=>"010111111",
  57277=>"000111111",
  57278=>"111000100",
  57279=>"111111101",
  57280=>"000111111",
  57281=>"111000111",
  57282=>"000000000",
  57283=>"111111000",
  57284=>"000000000",
  57285=>"011000100",
  57286=>"111111100",
  57287=>"000000000",
  57288=>"000000000",
  57289=>"000000001",
  57290=>"000000000",
  57291=>"111111111",
  57292=>"110111110",
  57293=>"111000000",
  57294=>"110001011",
  57295=>"111111110",
  57296=>"000100110",
  57297=>"000000111",
  57298=>"000111000",
  57299=>"000000000",
  57300=>"111111001",
  57301=>"001000011",
  57302=>"000000011",
  57303=>"000000000",
  57304=>"000000101",
  57305=>"000111111",
  57306=>"001001000",
  57307=>"011011111",
  57308=>"000000000",
  57309=>"111111111",
  57310=>"111111000",
  57311=>"000000110",
  57312=>"000000000",
  57313=>"001111111",
  57314=>"101000000",
  57315=>"111111111",
  57316=>"111111111",
  57317=>"000000000",
  57318=>"111011000",
  57319=>"111111011",
  57320=>"110001000",
  57321=>"000000111",
  57322=>"111001000",
  57323=>"000000000",
  57324=>"111101110",
  57325=>"110100000",
  57326=>"101000100",
  57327=>"000001111",
  57328=>"001111111",
  57329=>"000000001",
  57330=>"010111111",
  57331=>"111000000",
  57332=>"000000000",
  57333=>"000111111",
  57334=>"110111111",
  57335=>"111101001",
  57336=>"010010010",
  57337=>"100101111",
  57338=>"000001001",
  57339=>"010011000",
  57340=>"111111100",
  57341=>"000000000",
  57342=>"011000101",
  57343=>"000110111",
  57344=>"000000000",
  57345=>"111000000",
  57346=>"000000001",
  57347=>"100110110",
  57348=>"100110110",
  57349=>"000000000",
  57350=>"000001011",
  57351=>"111111111",
  57352=>"101001111",
  57353=>"000101111",
  57354=>"111111000",
  57355=>"011110111",
  57356=>"111111111",
  57357=>"011000000",
  57358=>"001100000",
  57359=>"111101011",
  57360=>"000001000",
  57361=>"111111111",
  57362=>"000000000",
  57363=>"000000000",
  57364=>"000001000",
  57365=>"000000000",
  57366=>"111111111",
  57367=>"011000000",
  57368=>"010000000",
  57369=>"110000000",
  57370=>"111111111",
  57371=>"000000000",
  57372=>"110111111",
  57373=>"111001001",
  57374=>"011111110",
  57375=>"000111010",
  57376=>"100000000",
  57377=>"111111111",
  57378=>"110110110",
  57379=>"111111111",
  57380=>"111001001",
  57381=>"111101001",
  57382=>"010100000",
  57383=>"000000100",
  57384=>"111111111",
  57385=>"111111000",
  57386=>"000000000",
  57387=>"000000000",
  57388=>"000000000",
  57389=>"000000000",
  57390=>"001111111",
  57391=>"000000000",
  57392=>"001001000",
  57393=>"111111111",
  57394=>"000001000",
  57395=>"000000000",
  57396=>"111111100",
  57397=>"111111111",
  57398=>"100000000",
  57399=>"000111111",
  57400=>"000000000",
  57401=>"110110011",
  57402=>"000000001",
  57403=>"000000101",
  57404=>"000001001",
  57405=>"111111111",
  57406=>"111111100",
  57407=>"000000000",
  57408=>"111111111",
  57409=>"111101111",
  57410=>"111111100",
  57411=>"000010000",
  57412=>"000111111",
  57413=>"000000000",
  57414=>"111000111",
  57415=>"111111111",
  57416=>"011011000",
  57417=>"000000000",
  57418=>"000000001",
  57419=>"100100000",
  57420=>"000000000",
  57421=>"110000011",
  57422=>"101100110",
  57423=>"000000000",
  57424=>"000000011",
  57425=>"000000000",
  57426=>"000000000",
  57427=>"000100111",
  57428=>"000000000",
  57429=>"000000000",
  57430=>"110110101",
  57431=>"011001001",
  57432=>"000000000",
  57433=>"000000000",
  57434=>"111111001",
  57435=>"001001100",
  57436=>"111111111",
  57437=>"100111111",
  57438=>"000000000",
  57439=>"000000010",
  57440=>"101111111",
  57441=>"111111111",
  57442=>"000000000",
  57443=>"111101100",
  57444=>"111101000",
  57445=>"000001011",
  57446=>"110110110",
  57447=>"000000000",
  57448=>"001001001",
  57449=>"000000000",
  57450=>"000000111",
  57451=>"111000000",
  57452=>"111111111",
  57453=>"111111111",
  57454=>"000000000",
  57455=>"110100100",
  57456=>"011011001",
  57457=>"000100111",
  57458=>"001111111",
  57459=>"011011111",
  57460=>"000000000",
  57461=>"111111111",
  57462=>"000000000",
  57463=>"000000000",
  57464=>"001111111",
  57465=>"000000000",
  57466=>"000010000",
  57467=>"000001011",
  57468=>"001001011",
  57469=>"111111001",
  57470=>"011011000",
  57471=>"000000010",
  57472=>"000000000",
  57473=>"111111111",
  57474=>"111111111",
  57475=>"111111111",
  57476=>"000000000",
  57477=>"000000100",
  57478=>"111110110",
  57479=>"001000001",
  57480=>"001111111",
  57481=>"000000000",
  57482=>"000000000",
  57483=>"000000001",
  57484=>"111111111",
  57485=>"000000000",
  57486=>"001000000",
  57487=>"010111111",
  57488=>"111101101",
  57489=>"111101000",
  57490=>"100110010",
  57491=>"111111111",
  57492=>"000000000",
  57493=>"001001000",
  57494=>"000000000",
  57495=>"000000101",
  57496=>"011001110",
  57497=>"000000000",
  57498=>"110011111",
  57499=>"000000110",
  57500=>"100100111",
  57501=>"111000000",
  57502=>"111100110",
  57503=>"010000000",
  57504=>"111111111",
  57505=>"001000000",
  57506=>"111111111",
  57507=>"111111111",
  57508=>"100110111",
  57509=>"000000100",
  57510=>"111111111",
  57511=>"100100111",
  57512=>"111111101",
  57513=>"111111111",
  57514=>"001000000",
  57515=>"010000000",
  57516=>"000000001",
  57517=>"110011010",
  57518=>"000000001",
  57519=>"001001101",
  57520=>"000110111",
  57521=>"001011000",
  57522=>"101101101",
  57523=>"111110111",
  57524=>"010011010",
  57525=>"000000000",
  57526=>"001101011",
  57527=>"000100101",
  57528=>"111000000",
  57529=>"000000000",
  57530=>"100110011",
  57531=>"100011011",
  57532=>"000000111",
  57533=>"101101101",
  57534=>"111111001",
  57535=>"000000000",
  57536=>"000000110",
  57537=>"011111000",
  57538=>"111111101",
  57539=>"111000000",
  57540=>"000000000",
  57541=>"010111111",
  57542=>"101100111",
  57543=>"000000000",
  57544=>"101111011",
  57545=>"000011011",
  57546=>"111100000",
  57547=>"000000111",
  57548=>"111111111",
  57549=>"000000000",
  57550=>"001011001",
  57551=>"000000001",
  57552=>"000010100",
  57553=>"001001111",
  57554=>"111111111",
  57555=>"000000000",
  57556=>"100100111",
  57557=>"110110111",
  57558=>"111101000",
  57559=>"110110110",
  57560=>"000000001",
  57561=>"111110000",
  57562=>"111111111",
  57563=>"101111100",
  57564=>"101111111",
  57565=>"100110110",
  57566=>"100111111",
  57567=>"000000011",
  57568=>"101111111",
  57569=>"000001111",
  57570=>"100011111",
  57571=>"111011000",
  57572=>"111110010",
  57573=>"100101001",
  57574=>"000000000",
  57575=>"110111111",
  57576=>"111111111",
  57577=>"100000000",
  57578=>"111111111",
  57579=>"000000000",
  57580=>"111111111",
  57581=>"000000000",
  57582=>"000000000",
  57583=>"111111111",
  57584=>"000101111",
  57585=>"000000000",
  57586=>"111111111",
  57587=>"000110101",
  57588=>"110111111",
  57589=>"001111111",
  57590=>"000000100",
  57591=>"111111111",
  57592=>"001111011",
  57593=>"000001001",
  57594=>"001111110",
  57595=>"111000000",
  57596=>"111110101",
  57597=>"110110111",
  57598=>"011000011",
  57599=>"010000001",
  57600=>"000000000",
  57601=>"000100100",
  57602=>"111111111",
  57603=>"000111111",
  57604=>"001001001",
  57605=>"000000111",
  57606=>"111111111",
  57607=>"100100101",
  57608=>"111111111",
  57609=>"111111101",
  57610=>"000000000",
  57611=>"100001111",
  57612=>"111001001",
  57613=>"000000111",
  57614=>"111111101",
  57615=>"011011111",
  57616=>"100111111",
  57617=>"111111000",
  57618=>"000000000",
  57619=>"000000000",
  57620=>"111001111",
  57621=>"011000110",
  57622=>"001111111",
  57623=>"111111110",
  57624=>"001101111",
  57625=>"000000000",
  57626=>"110000000",
  57627=>"000001001",
  57628=>"000000000",
  57629=>"000000000",
  57630=>"000000000",
  57631=>"111111111",
  57632=>"000000000",
  57633=>"000100101",
  57634=>"000000000",
  57635=>"000110110",
  57636=>"001000001",
  57637=>"000100000",
  57638=>"010111000",
  57639=>"000000000",
  57640=>"110010000",
  57641=>"000001000",
  57642=>"111110000",
  57643=>"000000000",
  57644=>"010011000",
  57645=>"110110000",
  57646=>"011111111",
  57647=>"101101000",
  57648=>"001000110",
  57649=>"000000000",
  57650=>"111111000",
  57651=>"010111111",
  57652=>"000000000",
  57653=>"111111001",
  57654=>"111100001",
  57655=>"111111111",
  57656=>"001000001",
  57657=>"111111111",
  57658=>"111111000",
  57659=>"111101111",
  57660=>"000010000",
  57661=>"010111000",
  57662=>"100011011",
  57663=>"111111111",
  57664=>"000100100",
  57665=>"000000000",
  57666=>"111111110",
  57667=>"111011000",
  57668=>"000001001",
  57669=>"111111111",
  57670=>"111111111",
  57671=>"111111110",
  57672=>"111111000",
  57673=>"111111111",
  57674=>"000000111",
  57675=>"000111111",
  57676=>"100111111",
  57677=>"100100111",
  57678=>"011011111",
  57679=>"111111001",
  57680=>"101111111",
  57681=>"011011111",
  57682=>"111111001",
  57683=>"000000000",
  57684=>"000000011",
  57685=>"010000000",
  57686=>"111111111",
  57687=>"111111110",
  57688=>"111111111",
  57689=>"000000111",
  57690=>"000000011",
  57691=>"010000000",
  57692=>"000100111",
  57693=>"000000010",
  57694=>"011001111",
  57695=>"000000000",
  57696=>"110100101",
  57697=>"000000000",
  57698=>"100100101",
  57699=>"100000001",
  57700=>"001011011",
  57701=>"000101111",
  57702=>"101000111",
  57703=>"111110111",
  57704=>"011011011",
  57705=>"000000000",
  57706=>"100111111",
  57707=>"111111111",
  57708=>"100000000",
  57709=>"111111000",
  57710=>"100000000",
  57711=>"000000000",
  57712=>"011000011",
  57713=>"100000000",
  57714=>"111011111",
  57715=>"110110111",
  57716=>"000100100",
  57717=>"111111111",
  57718=>"111101001",
  57719=>"101111111",
  57720=>"111111111",
  57721=>"001111111",
  57722=>"101000000",
  57723=>"100100000",
  57724=>"111111111",
  57725=>"000000000",
  57726=>"100001111",
  57727=>"111111100",
  57728=>"001011011",
  57729=>"000010000",
  57730=>"000010000",
  57731=>"000000100",
  57732=>"111111111",
  57733=>"000000000",
  57734=>"000110110",
  57735=>"011001000",
  57736=>"111111111",
  57737=>"001011110",
  57738=>"111011000",
  57739=>"000100100",
  57740=>"111111111",
  57741=>"001100100",
  57742=>"111111111",
  57743=>"010100110",
  57744=>"111111000",
  57745=>"000000000",
  57746=>"011101100",
  57747=>"001000000",
  57748=>"111111111",
  57749=>"111001001",
  57750=>"100110111",
  57751=>"011111111",
  57752=>"011111111",
  57753=>"111001011",
  57754=>"110100111",
  57755=>"111111111",
  57756=>"001011010",
  57757=>"111111111",
  57758=>"111000000",
  57759=>"000000000",
  57760=>"100000000",
  57761=>"000110111",
  57762=>"100100100",
  57763=>"111111111",
  57764=>"001000000",
  57765=>"000000101",
  57766=>"001101111",
  57767=>"101100001",
  57768=>"000000000",
  57769=>"000100100",
  57770=>"111111111",
  57771=>"000000000",
  57772=>"000000000",
  57773=>"000000000",
  57774=>"111111001",
  57775=>"110111011",
  57776=>"111111111",
  57777=>"111111001",
  57778=>"011111111",
  57779=>"010110000",
  57780=>"000000000",
  57781=>"111111110",
  57782=>"011000101",
  57783=>"000111000",
  57784=>"000100000",
  57785=>"000000000",
  57786=>"100110110",
  57787=>"000000000",
  57788=>"000000000",
  57789=>"110111111",
  57790=>"001111111",
  57791=>"000001101",
  57792=>"111111111",
  57793=>"101001000",
  57794=>"000000000",
  57795=>"111111111",
  57796=>"110100101",
  57797=>"111101101",
  57798=>"111000000",
  57799=>"111001000",
  57800=>"111111111",
  57801=>"000001111",
  57802=>"110110100",
  57803=>"001111110",
  57804=>"000010110",
  57805=>"111111111",
  57806=>"111110110",
  57807=>"111111111",
  57808=>"000100100",
  57809=>"000000000",
  57810=>"111111111",
  57811=>"101001000",
  57812=>"111111111",
  57813=>"001000000",
  57814=>"111011011",
  57815=>"111111000",
  57816=>"000000111",
  57817=>"011111000",
  57818=>"101111011",
  57819=>"111111111",
  57820=>"110111111",
  57821=>"001101111",
  57822=>"011001001",
  57823=>"011101101",
  57824=>"000101111",
  57825=>"000000111",
  57826=>"000000000",
  57827=>"011111111",
  57828=>"000000001",
  57829=>"000000000",
  57830=>"000000000",
  57831=>"000000000",
  57832=>"111111111",
  57833=>"101111111",
  57834=>"010111111",
  57835=>"111111000",
  57836=>"111100001",
  57837=>"010010111",
  57838=>"111111111",
  57839=>"011011111",
  57840=>"110101000",
  57841=>"000000000",
  57842=>"001001000",
  57843=>"001111111",
  57844=>"111111011",
  57845=>"000110000",
  57846=>"011001000",
  57847=>"110010110",
  57848=>"111111110",
  57849=>"110111011",
  57850=>"111000011",
  57851=>"000000000",
  57852=>"101001001",
  57853=>"011111110",
  57854=>"111111000",
  57855=>"000000000",
  57856=>"111101111",
  57857=>"000000000",
  57858=>"000010111",
  57859=>"000000000",
  57860=>"111111111",
  57861=>"110110010",
  57862=>"001101101",
  57863=>"111100000",
  57864=>"000000000",
  57865=>"000000000",
  57866=>"100111111",
  57867=>"000000000",
  57868=>"011111111",
  57869=>"000011111",
  57870=>"100000110",
  57871=>"010110111",
  57872=>"111001011",
  57873=>"000000000",
  57874=>"100101101",
  57875=>"111111111",
  57876=>"000000011",
  57877=>"000000110",
  57878=>"111111001",
  57879=>"011111100",
  57880=>"111111111",
  57881=>"100110111",
  57882=>"101001011",
  57883=>"011000001",
  57884=>"101101101",
  57885=>"000000001",
  57886=>"011111111",
  57887=>"000101101",
  57888=>"000000000",
  57889=>"101101001",
  57890=>"110000001",
  57891=>"111111111",
  57892=>"111111011",
  57893=>"111111110",
  57894=>"111111110",
  57895=>"000000111",
  57896=>"111111111",
  57897=>"000000000",
  57898=>"000001000",
  57899=>"000000110",
  57900=>"111111000",
  57901=>"000000000",
  57902=>"101111111",
  57903=>"000000011",
  57904=>"000000110",
  57905=>"000000111",
  57906=>"101100100",
  57907=>"110110100",
  57908=>"000110111",
  57909=>"001011011",
  57910=>"000000111",
  57911=>"011011010",
  57912=>"001011001",
  57913=>"111111111",
  57914=>"000000000",
  57915=>"111111111",
  57916=>"111000111",
  57917=>"000100111",
  57918=>"110111111",
  57919=>"000000000",
  57920=>"000000001",
  57921=>"000100110",
  57922=>"001111111",
  57923=>"111001001",
  57924=>"000010111",
  57925=>"111111111",
  57926=>"000000000",
  57927=>"000000000",
  57928=>"000010010",
  57929=>"000000000",
  57930=>"111111000",
  57931=>"000011011",
  57932=>"111111111",
  57933=>"000000000",
  57934=>"000111111",
  57935=>"111111111",
  57936=>"000001111",
  57937=>"111111111",
  57938=>"000000001",
  57939=>"000010110",
  57940=>"000000111",
  57941=>"000000000",
  57942=>"000110111",
  57943=>"101111000",
  57944=>"000000000",
  57945=>"111000000",
  57946=>"111000000",
  57947=>"000011011",
  57948=>"000000000",
  57949=>"001000000",
  57950=>"110111110",
  57951=>"000000000",
  57952=>"001000111",
  57953=>"110110111",
  57954=>"000000000",
  57955=>"000111111",
  57956=>"000100100",
  57957=>"000000001",
  57958=>"011011111",
  57959=>"000000000",
  57960=>"110110000",
  57961=>"111111111",
  57962=>"010111111",
  57963=>"000000111",
  57964=>"001011011",
  57965=>"111111111",
  57966=>"111000000",
  57967=>"000000000",
  57968=>"111110000",
  57969=>"010000111",
  57970=>"101000010",
  57971=>"000001000",
  57972=>"000111111",
  57973=>"000101111",
  57974=>"000000000",
  57975=>"000000111",
  57976=>"111000000",
  57977=>"111000001",
  57978=>"000011111",
  57979=>"000000000",
  57980=>"000000011",
  57981=>"000000000",
  57982=>"111111111",
  57983=>"000001000",
  57984=>"111111111",
  57985=>"000000000",
  57986=>"000000000",
  57987=>"000000011",
  57988=>"111111111",
  57989=>"000000100",
  57990=>"000111010",
  57991=>"010010011",
  57992=>"110111111",
  57993=>"000000100",
  57994=>"000000000",
  57995=>"100000000",
  57996=>"000000000",
  57997=>"111111111",
  57998=>"111111111",
  57999=>"000000000",
  58000=>"110110000",
  58001=>"000000010",
  58002=>"111111011",
  58003=>"000000000",
  58004=>"000001000",
  58005=>"000000000",
  58006=>"100000000",
  58007=>"010000000",
  58008=>"100011000",
  58009=>"000100000",
  58010=>"001000000",
  58011=>"110111111",
  58012=>"000000100",
  58013=>"001001000",
  58014=>"111111111",
  58015=>"100111100",
  58016=>"000000111",
  58017=>"101111111",
  58018=>"000000000",
  58019=>"111111010",
  58020=>"001001111",
  58021=>"001100110",
  58022=>"111111110",
  58023=>"000100111",
  58024=>"111111000",
  58025=>"111000100",
  58026=>"001000000",
  58027=>"111111111",
  58028=>"110111111",
  58029=>"000111101",
  58030=>"110011010",
  58031=>"000011001",
  58032=>"111111011",
  58033=>"001010000",
  58034=>"110111110",
  58035=>"111111111",
  58036=>"111111111",
  58037=>"001000001",
  58038=>"000000000",
  58039=>"100100101",
  58040=>"111010110",
  58041=>"000000000",
  58042=>"000001101",
  58043=>"111101101",
  58044=>"010001011",
  58045=>"000000011",
  58046=>"111111111",
  58047=>"101111110",
  58048=>"111111111",
  58049=>"111111111",
  58050=>"010111111",
  58051=>"111111111",
  58052=>"000000000",
  58053=>"111011000",
  58054=>"100111111",
  58055=>"001111111",
  58056=>"001001111",
  58057=>"000000000",
  58058=>"000010010",
  58059=>"000001000",
  58060=>"111000000",
  58061=>"111110000",
  58062=>"110000111",
  58063=>"000000000",
  58064=>"000000000",
  58065=>"000000010",
  58066=>"000000000",
  58067=>"000000000",
  58068=>"100100011",
  58069=>"111111111",
  58070=>"101000000",
  58071=>"000000000",
  58072=>"000000001",
  58073=>"111110100",
  58074=>"000000000",
  58075=>"111011000",
  58076=>"000000010",
  58077=>"010000000",
  58078=>"111111110",
  58079=>"000001001",
  58080=>"001000000",
  58081=>"000000010",
  58082=>"000000000",
  58083=>"000000000",
  58084=>"000000000",
  58085=>"000100100",
  58086=>"111000001",
  58087=>"000111111",
  58088=>"111111111",
  58089=>"000000101",
  58090=>"000100101",
  58091=>"010000000",
  58092=>"111111111",
  58093=>"000000000",
  58094=>"000000000",
  58095=>"100101111",
  58096=>"001000000",
  58097=>"110111100",
  58098=>"101101111",
  58099=>"001000100",
  58100=>"000000000",
  58101=>"000000000",
  58102=>"111000001",
  58103=>"111000000",
  58104=>"000000000",
  58105=>"011111001",
  58106=>"011011111",
  58107=>"111111111",
  58108=>"011011011",
  58109=>"001000000",
  58110=>"010001101",
  58111=>"011111111",
  58112=>"111010000",
  58113=>"100100000",
  58114=>"111111111",
  58115=>"111111100",
  58116=>"001001111",
  58117=>"111111000",
  58118=>"000000000",
  58119=>"111111100",
  58120=>"011111111",
  58121=>"000000000",
  58122=>"111111111",
  58123=>"000100100",
  58124=>"000000000",
  58125=>"010000000",
  58126=>"110111111",
  58127=>"111111000",
  58128=>"111001001",
  58129=>"111001000",
  58130=>"000000010",
  58131=>"000111100",
  58132=>"111000000",
  58133=>"000000001",
  58134=>"001111111",
  58135=>"000000101",
  58136=>"000011111",
  58137=>"000000001",
  58138=>"010111111",
  58139=>"010000000",
  58140=>"011111111",
  58141=>"000100110",
  58142=>"111111111",
  58143=>"100011000",
  58144=>"111111000",
  58145=>"000000010",
  58146=>"000010000",
  58147=>"000000000",
  58148=>"000000000",
  58149=>"000000000",
  58150=>"000000010",
  58151=>"000000000",
  58152=>"111111111",
  58153=>"000011111",
  58154=>"111111111",
  58155=>"111000000",
  58156=>"000000000",
  58157=>"100110110",
  58158=>"111111000",
  58159=>"000000000",
  58160=>"111111111",
  58161=>"001111111",
  58162=>"111011000",
  58163=>"111111000",
  58164=>"110000000",
  58165=>"110111110",
  58166=>"111010000",
  58167=>"000110111",
  58168=>"000000000",
  58169=>"000000101",
  58170=>"010010000",
  58171=>"111111111",
  58172=>"000000100",
  58173=>"111000000",
  58174=>"100111111",
  58175=>"111111101",
  58176=>"111100000",
  58177=>"110111111",
  58178=>"011010000",
  58179=>"000001011",
  58180=>"000000111",
  58181=>"001011111",
  58182=>"011001000",
  58183=>"101001001",
  58184=>"010110110",
  58185=>"000000111",
  58186=>"110000000",
  58187=>"111100000",
  58188=>"011000000",
  58189=>"110000000",
  58190=>"111011000",
  58191=>"111110100",
  58192=>"001111111",
  58193=>"000000111",
  58194=>"001001100",
  58195=>"010000000",
  58196=>"000000000",
  58197=>"000000001",
  58198=>"111100000",
  58199=>"110010000",
  58200=>"111000111",
  58201=>"000001111",
  58202=>"111111111",
  58203=>"000010111",
  58204=>"111000000",
  58205=>"111010000",
  58206=>"000000000",
  58207=>"000000000",
  58208=>"111111111",
  58209=>"111111111",
  58210=>"110111111",
  58211=>"101101111",
  58212=>"000000110",
  58213=>"000000001",
  58214=>"111111001",
  58215=>"000000000",
  58216=>"110100000",
  58217=>"011000000",
  58218=>"000111001",
  58219=>"101000000",
  58220=>"000000101",
  58221=>"101111000",
  58222=>"000000000",
  58223=>"111111111",
  58224=>"000000000",
  58225=>"111111110",
  58226=>"111100100",
  58227=>"000000100",
  58228=>"111111111",
  58229=>"000000000",
  58230=>"111111111",
  58231=>"000000000",
  58232=>"000000110",
  58233=>"100101111",
  58234=>"110111111",
  58235=>"111000000",
  58236=>"111111111",
  58237=>"111101001",
  58238=>"000000000",
  58239=>"001001000",
  58240=>"001001101",
  58241=>"111111111",
  58242=>"100110011",
  58243=>"111111110",
  58244=>"000000000",
  58245=>"101111111",
  58246=>"111101101",
  58247=>"000011111",
  58248=>"010010111",
  58249=>"111101101",
  58250=>"000000000",
  58251=>"111111100",
  58252=>"111101101",
  58253=>"001001011",
  58254=>"111111111",
  58255=>"110100001",
  58256=>"111111111",
  58257=>"101001001",
  58258=>"000000011",
  58259=>"011000001",
  58260=>"111111001",
  58261=>"011010000",
  58262=>"000000000",
  58263=>"001001111",
  58264=>"111111011",
  58265=>"111101111",
  58266=>"111111111",
  58267=>"000100000",
  58268=>"000000000",
  58269=>"000000100",
  58270=>"101001000",
  58271=>"000110111",
  58272=>"011111000",
  58273=>"000000011",
  58274=>"000000100",
  58275=>"111000000",
  58276=>"111110000",
  58277=>"010001111",
  58278=>"000000110",
  58279=>"000111110",
  58280=>"100111111",
  58281=>"000000000",
  58282=>"111111111",
  58283=>"111001001",
  58284=>"000000000",
  58285=>"111010010",
  58286=>"111111111",
  58287=>"000000000",
  58288=>"111000100",
  58289=>"000100100",
  58290=>"000000000",
  58291=>"011000000",
  58292=>"110111111",
  58293=>"011111111",
  58294=>"110111111",
  58295=>"000010000",
  58296=>"111111111",
  58297=>"111111111",
  58298=>"000001111",
  58299=>"001111111",
  58300=>"000000000",
  58301=>"101111111",
  58302=>"100111011",
  58303=>"000000011",
  58304=>"000000011",
  58305=>"001011110",
  58306=>"111111111",
  58307=>"111111010",
  58308=>"010111100",
  58309=>"000000111",
  58310=>"001000000",
  58311=>"000000000",
  58312=>"111111111",
  58313=>"000101111",
  58314=>"000000000",
  58315=>"000001111",
  58316=>"000000111",
  58317=>"001001011",
  58318=>"000001000",
  58319=>"110000111",
  58320=>"111100100",
  58321=>"111000000",
  58322=>"000000000",
  58323=>"000000001",
  58324=>"111111110",
  58325=>"111111001",
  58326=>"111111111",
  58327=>"000010011",
  58328=>"000111110",
  58329=>"111111111",
  58330=>"000001000",
  58331=>"000111111",
  58332=>"100100100",
  58333=>"111000000",
  58334=>"000000001",
  58335=>"001001010",
  58336=>"000000010",
  58337=>"000000000",
  58338=>"000000001",
  58339=>"111000000",
  58340=>"110010011",
  58341=>"111111111",
  58342=>"000000000",
  58343=>"011011011",
  58344=>"000000101",
  58345=>"000000111",
  58346=>"000000010",
  58347=>"000100100",
  58348=>"101000000",
  58349=>"000000100",
  58350=>"111000000",
  58351=>"000001000",
  58352=>"000000000",
  58353=>"000000110",
  58354=>"111111111",
  58355=>"001000000",
  58356=>"000000001",
  58357=>"000000000",
  58358=>"110000000",
  58359=>"000000000",
  58360=>"111101111",
  58361=>"001001111",
  58362=>"111111011",
  58363=>"110111110",
  58364=>"100111101",
  58365=>"110000000",
  58366=>"000001001",
  58367=>"101000101",
  58368=>"000000001",
  58369=>"111111111",
  58370=>"111011000",
  58371=>"111111111",
  58372=>"110110110",
  58373=>"000000000",
  58374=>"010111111",
  58375=>"011000111",
  58376=>"000110111",
  58377=>"000111111",
  58378=>"000000010",
  58379=>"010000000",
  58380=>"110111111",
  58381=>"100011000",
  58382=>"111100111",
  58383=>"110111111",
  58384=>"001111111",
  58385=>"111111111",
  58386=>"011111001",
  58387=>"000000111",
  58388=>"001000000",
  58389=>"000000000",
  58390=>"101111111",
  58391=>"000000110",
  58392=>"111000001",
  58393=>"000000000",
  58394=>"000111000",
  58395=>"100000000",
  58396=>"001000000",
  58397=>"111111111",
  58398=>"110101111",
  58399=>"000001001",
  58400=>"011010000",
  58401=>"000000000",
  58402=>"110111111",
  58403=>"101100100",
  58404=>"111111111",
  58405=>"110010010",
  58406=>"000000000",
  58407=>"000000000",
  58408=>"111111111",
  58409=>"000000000",
  58410=>"010000000",
  58411=>"111101111",
  58412=>"001001111",
  58413=>"100000000",
  58414=>"000000111",
  58415=>"000000000",
  58416=>"000000000",
  58417=>"000000011",
  58418=>"000100000",
  58419=>"101100100",
  58420=>"111111011",
  58421=>"100110110",
  58422=>"111111000",
  58423=>"000000000",
  58424=>"110111011",
  58425=>"111111111",
  58426=>"000000000",
  58427=>"111111111",
  58428=>"000000000",
  58429=>"111100100",
  58430=>"111111111",
  58431=>"111000100",
  58432=>"100100001",
  58433=>"111111111",
  58434=>"111000000",
  58435=>"000001111",
  58436=>"011001001",
  58437=>"000000100",
  58438=>"000001111",
  58439=>"000000000",
  58440=>"011000000",
  58441=>"111111111",
  58442=>"111111111",
  58443=>"111111000",
  58444=>"111011011",
  58445=>"011000000",
  58446=>"000000000",
  58447=>"111111110",
  58448=>"110111110",
  58449=>"000000000",
  58450=>"000000000",
  58451=>"001000000",
  58452=>"111011000",
  58453=>"011000000",
  58454=>"111011010",
  58455=>"111000000",
  58456=>"000000000",
  58457=>"100000001",
  58458=>"101000000",
  58459=>"000000000",
  58460=>"001000000",
  58461=>"000111111",
  58462=>"000000000",
  58463=>"110011110",
  58464=>"000000000",
  58465=>"111111111",
  58466=>"111011111",
  58467=>"000000111",
  58468=>"000000011",
  58469=>"111111110",
  58470=>"111111111",
  58471=>"000111010",
  58472=>"111111111",
  58473=>"111111111",
  58474=>"111100000",
  58475=>"111111111",
  58476=>"101101111",
  58477=>"000000000",
  58478=>"000000000",
  58479=>"000100111",
  58480=>"000000110",
  58481=>"000000000",
  58482=>"010010000",
  58483=>"000000000",
  58484=>"000000000",
  58485=>"101100100",
  58486=>"000000000",
  58487=>"011111111",
  58488=>"111000000",
  58489=>"000000000",
  58490=>"000000111",
  58491=>"000111111",
  58492=>"111101100",
  58493=>"110110000",
  58494=>"111111111",
  58495=>"001001100",
  58496=>"000000011",
  58497=>"111111111",
  58498=>"000011000",
  58499=>"001111111",
  58500=>"000000000",
  58501=>"000000011",
  58502=>"111111110",
  58503=>"111101111",
  58504=>"111111111",
  58505=>"000000001",
  58506=>"000000000",
  58507=>"111111111",
  58508=>"010111011",
  58509=>"000111001",
  58510=>"101111111",
  58511=>"000000110",
  58512=>"001000000",
  58513=>"000000000",
  58514=>"000000000",
  58515=>"111110110",
  58516=>"001111000",
  58517=>"000000000",
  58518=>"110000000",
  58519=>"000000000",
  58520=>"000000000",
  58521=>"111010000",
  58522=>"111111000",
  58523=>"001101000",
  58524=>"000000000",
  58525=>"110000110",
  58526=>"000000000",
  58527=>"000000000",
  58528=>"000111111",
  58529=>"111111000",
  58530=>"011111010",
  58531=>"100111111",
  58532=>"111111111",
  58533=>"011000000",
  58534=>"111111111",
  58535=>"011010000",
  58536=>"110101111",
  58537=>"000010010",
  58538=>"111110110",
  58539=>"001000111",
  58540=>"100000100",
  58541=>"111111111",
  58542=>"111010001",
  58543=>"111111010",
  58544=>"000000000",
  58545=>"000000000",
  58546=>"110111000",
  58547=>"110010000",
  58548=>"000000011",
  58549=>"000000000",
  58550=>"111101000",
  58551=>"000000000",
  58552=>"111110111",
  58553=>"010000000",
  58554=>"000000000",
  58555=>"111001001",
  58556=>"000010011",
  58557=>"000000000",
  58558=>"110011111",
  58559=>"000000001",
  58560=>"110100100",
  58561=>"111111111",
  58562=>"111111111",
  58563=>"000000111",
  58564=>"000111111",
  58565=>"000000000",
  58566=>"011011001",
  58567=>"011000011",
  58568=>"110010111",
  58569=>"001000001",
  58570=>"111110000",
  58571=>"111111111",
  58572=>"111111000",
  58573=>"111111100",
  58574=>"001000000",
  58575=>"110111011",
  58576=>"000000000",
  58577=>"101101001",
  58578=>"111111100",
  58579=>"000000000",
  58580=>"111111110",
  58581=>"000001001",
  58582=>"000000000",
  58583=>"100100111",
  58584=>"010000000",
  58585=>"000100110",
  58586=>"111111111",
  58587=>"000011111",
  58588=>"001000000",
  58589=>"111111111",
  58590=>"000000011",
  58591=>"000000000",
  58592=>"111111111",
  58593=>"000000111",
  58594=>"111111111",
  58595=>"000011010",
  58596=>"000000000",
  58597=>"100000010",
  58598=>"000000000",
  58599=>"000000000",
  58600=>"111111111",
  58601=>"111111011",
  58602=>"100111000",
  58603=>"001001111",
  58604=>"000000000",
  58605=>"000000000",
  58606=>"111111111",
  58607=>"000000000",
  58608=>"000111000",
  58609=>"000000011",
  58610=>"111111111",
  58611=>"011101101",
  58612=>"011111011",
  58613=>"000001001",
  58614=>"000000000",
  58615=>"000000000",
  58616=>"110110111",
  58617=>"111111111",
  58618=>"011000010",
  58619=>"000000000",
  58620=>"100100111",
  58621=>"111110110",
  58622=>"110111111",
  58623=>"100000000",
  58624=>"111111101",
  58625=>"111111011",
  58626=>"000000010",
  58627=>"010100110",
  58628=>"111001000",
  58629=>"000000000",
  58630=>"000001111",
  58631=>"011010000",
  58632=>"000000000",
  58633=>"000000000",
  58634=>"111111111",
  58635=>"100111011",
  58636=>"001001001",
  58637=>"111111111",
  58638=>"111111111",
  58639=>"111111111",
  58640=>"000000000",
  58641=>"000010111",
  58642=>"111111111",
  58643=>"000110000",
  58644=>"111111110",
  58645=>"111111111",
  58646=>"100110110",
  58647=>"000000000",
  58648=>"000000000",
  58649=>"000000000",
  58650=>"111101000",
  58651=>"000111110",
  58652=>"011011111",
  58653=>"111110110",
  58654=>"111000000",
  58655=>"111111111",
  58656=>"011100100",
  58657=>"100000110",
  58658=>"000000000",
  58659=>"111111011",
  58660=>"111110100",
  58661=>"110100000",
  58662=>"111111111",
  58663=>"000000000",
  58664=>"100100000",
  58665=>"000000001",
  58666=>"000010111",
  58667=>"111111001",
  58668=>"001001000",
  58669=>"001001001",
  58670=>"001000000",
  58671=>"111000000",
  58672=>"000000000",
  58673=>"010000000",
  58674=>"111111111",
  58675=>"100000000",
  58676=>"001000000",
  58677=>"110010011",
  58678=>"000010111",
  58679=>"111111111",
  58680=>"000000000",
  58681=>"000000111",
  58682=>"110111111",
  58683=>"000000000",
  58684=>"011000010",
  58685=>"001011011",
  58686=>"000011000",
  58687=>"111111110",
  58688=>"000000111",
  58689=>"011000100",
  58690=>"110111111",
  58691=>"111111111",
  58692=>"111011011",
  58693=>"100000000",
  58694=>"111111110",
  58695=>"000010111",
  58696=>"100000000",
  58697=>"111111000",
  58698=>"000000000",
  58699=>"010000001",
  58700=>"000000000",
  58701=>"111111000",
  58702=>"110000000",
  58703=>"110100000",
  58704=>"110110000",
  58705=>"111000111",
  58706=>"111100000",
  58707=>"111111111",
  58708=>"111111111",
  58709=>"000100111",
  58710=>"000000000",
  58711=>"110010110",
  58712=>"001000000",
  58713=>"000000000",
  58714=>"110110110",
  58715=>"000000111",
  58716=>"000011111",
  58717=>"100000000",
  58718=>"111110000",
  58719=>"111100000",
  58720=>"000011111",
  58721=>"000001111",
  58722=>"110110110",
  58723=>"111111111",
  58724=>"000000000",
  58725=>"000000111",
  58726=>"111101000",
  58727=>"000000000",
  58728=>"110111111",
  58729=>"000010010",
  58730=>"011001000",
  58731=>"000000000",
  58732=>"000000110",
  58733=>"000100000",
  58734=>"000000000",
  58735=>"011000000",
  58736=>"111000000",
  58737=>"000000000",
  58738=>"111001111",
  58739=>"000110000",
  58740=>"000000000",
  58741=>"111111111",
  58742=>"111001000",
  58743=>"111111001",
  58744=>"000000000",
  58745=>"111110100",
  58746=>"110100101",
  58747=>"111000000",
  58748=>"111101000",
  58749=>"011111011",
  58750=>"111111111",
  58751=>"001000000",
  58752=>"111101000",
  58753=>"110100000",
  58754=>"000000000",
  58755=>"111000000",
  58756=>"000000000",
  58757=>"111111111",
  58758=>"000000000",
  58759=>"111010000",
  58760=>"111100000",
  58761=>"110110110",
  58762=>"111001000",
  58763=>"111111011",
  58764=>"000000111",
  58765=>"111000011",
  58766=>"000000000",
  58767=>"011110010",
  58768=>"000001111",
  58769=>"000001111",
  58770=>"111110001",
  58771=>"100000001",
  58772=>"111111111",
  58773=>"000000000",
  58774=>"101000000",
  58775=>"000000000",
  58776=>"000111111",
  58777=>"100111110",
  58778=>"000000000",
  58779=>"000000000",
  58780=>"000000000",
  58781=>"111111110",
  58782=>"000000000",
  58783=>"000111111",
  58784=>"111111000",
  58785=>"000000000",
  58786=>"111000000",
  58787=>"111111111",
  58788=>"111111111",
  58789=>"000000000",
  58790=>"111000000",
  58791=>"111111111",
  58792=>"000000000",
  58793=>"000000000",
  58794=>"001000000",
  58795=>"111111001",
  58796=>"000110000",
  58797=>"001111111",
  58798=>"001111111",
  58799=>"111111111",
  58800=>"000000111",
  58801=>"000000010",
  58802=>"111111000",
  58803=>"000000000",
  58804=>"111111111",
  58805=>"111111111",
  58806=>"001111101",
  58807=>"000000000",
  58808=>"000001101",
  58809=>"000000000",
  58810=>"110100110",
  58811=>"111111000",
  58812=>"000000001",
  58813=>"111011000",
  58814=>"000000000",
  58815=>"001001001",
  58816=>"110111101",
  58817=>"000000000",
  58818=>"111111111",
  58819=>"000000000",
  58820=>"111111101",
  58821=>"111111110",
  58822=>"000000111",
  58823=>"000000000",
  58824=>"000000001",
  58825=>"000001000",
  58826=>"010010010",
  58827=>"000000101",
  58828=>"010010111",
  58829=>"110111011",
  58830=>"000000000",
  58831=>"111111111",
  58832=>"000000000",
  58833=>"111011011",
  58834=>"000000000",
  58835=>"000000111",
  58836=>"100111110",
  58837=>"100101111",
  58838=>"100000000",
  58839=>"011011101",
  58840=>"111110110",
  58841=>"000000000",
  58842=>"111000000",
  58843=>"000000000",
  58844=>"000010111",
  58845=>"110111000",
  58846=>"111111111",
  58847=>"011000001",
  58848=>"011001000",
  58849=>"000000111",
  58850=>"000000000",
  58851=>"111111111",
  58852=>"011001001",
  58853=>"111111111",
  58854=>"111101001",
  58855=>"111111110",
  58856=>"000010111",
  58857=>"110101100",
  58858=>"100101111",
  58859=>"000000011",
  58860=>"000000000",
  58861=>"111110110",
  58862=>"000100101",
  58863=>"111100000",
  58864=>"010010000",
  58865=>"111111111",
  58866=>"000000000",
  58867=>"110110000",
  58868=>"111111111",
  58869=>"000000000",
  58870=>"111111111",
  58871=>"111111110",
  58872=>"000000111",
  58873=>"000000000",
  58874=>"111111111",
  58875=>"000000000",
  58876=>"011011011",
  58877=>"100000001",
  58878=>"000000000",
  58879=>"000000000",
  58880=>"001011111",
  58881=>"000001001",
  58882=>"100111111",
  58883=>"101111111",
  58884=>"001111111",
  58885=>"011001100",
  58886=>"000000111",
  58887=>"111111011",
  58888=>"000000000",
  58889=>"000000000",
  58890=>"000000000",
  58891=>"011011111",
  58892=>"000110100",
  58893=>"000000000",
  58894=>"111111111",
  58895=>"111111111",
  58896=>"111111011",
  58897=>"000000001",
  58898=>"000100110",
  58899=>"111111111",
  58900=>"111000000",
  58901=>"100100111",
  58902=>"001000000",
  58903=>"001011011",
  58904=>"111111111",
  58905=>"001011011",
  58906=>"111111111",
  58907=>"111010000",
  58908=>"000000000",
  58909=>"111111110",
  58910=>"001110110",
  58911=>"111111110",
  58912=>"111001111",
  58913=>"000001111",
  58914=>"111111111",
  58915=>"111111111",
  58916=>"100101100",
  58917=>"001111111",
  58918=>"000011111",
  58919=>"000000000",
  58920=>"111111111",
  58921=>"000000000",
  58922=>"111100000",
  58923=>"111111111",
  58924=>"011111111",
  58925=>"111111111",
  58926=>"000011111",
  58927=>"110000000",
  58928=>"100001111",
  58929=>"000001001",
  58930=>"011000001",
  58931=>"111100100",
  58932=>"011001000",
  58933=>"000000011",
  58934=>"000100001",
  58935=>"011011100",
  58936=>"100111111",
  58937=>"011001111",
  58938=>"000000000",
  58939=>"110111111",
  58940=>"100000000",
  58941=>"111111110",
  58942=>"000010110",
  58943=>"111111111",
  58944=>"010011111",
  58945=>"100110111",
  58946=>"111111111",
  58947=>"111111111",
  58948=>"000011010",
  58949=>"011011000",
  58950=>"111111110",
  58951=>"111111111",
  58952=>"011011001",
  58953=>"111111111",
  58954=>"000000000",
  58955=>"111000000",
  58956=>"000000110",
  58957=>"110010111",
  58958=>"000011111",
  58959=>"000000011",
  58960=>"111111111",
  58961=>"110111011",
  58962=>"011000000",
  58963=>"000010010",
  58964=>"111111111",
  58965=>"000010000",
  58966=>"000001000",
  58967=>"110000111",
  58968=>"111111111",
  58969=>"101100000",
  58970=>"110011101",
  58971=>"111111111",
  58972=>"001001101",
  58973=>"111111111",
  58974=>"100001000",
  58975=>"111111111",
  58976=>"000000000",
  58977=>"111111111",
  58978=>"010011001",
  58979=>"111111111",
  58980=>"111110100",
  58981=>"111111111",
  58982=>"111101000",
  58983=>"000000111",
  58984=>"000000110",
  58985=>"000111111",
  58986=>"100100000",
  58987=>"000000000",
  58988=>"000001011",
  58989=>"111111111",
  58990=>"000000100",
  58991=>"010011111",
  58992=>"001011111",
  58993=>"001111111",
  58994=>"000010001",
  58995=>"000001000",
  58996=>"110100000",
  58997=>"000000000",
  58998=>"111111111",
  58999=>"111001101",
  59000=>"111001000",
  59001=>"000000000",
  59002=>"000000111",
  59003=>"111000111",
  59004=>"000000000",
  59005=>"000010000",
  59006=>"011111111",
  59007=>"000000000",
  59008=>"111111110",
  59009=>"111100111",
  59010=>"111111110",
  59011=>"011001000",
  59012=>"000000000",
  59013=>"000000101",
  59014=>"111110110",
  59015=>"000001001",
  59016=>"000000000",
  59017=>"111111100",
  59018=>"011111111",
  59019=>"011011011",
  59020=>"000000001",
  59021=>"111111111",
  59022=>"111111110",
  59023=>"000110110",
  59024=>"001000000",
  59025=>"000000000",
  59026=>"010000101",
  59027=>"001011001",
  59028=>"001101111",
  59029=>"000001000",
  59030=>"111111001",
  59031=>"000000000",
  59032=>"000001100",
  59033=>"111111010",
  59034=>"000001001",
  59035=>"000000001",
  59036=>"011111111",
  59037=>"000000000",
  59038=>"000000000",
  59039=>"000000100",
  59040=>"000111010",
  59041=>"000000111",
  59042=>"111111100",
  59043=>"111111111",
  59044=>"000000000",
  59045=>"100111001",
  59046=>"101000000",
  59047=>"000000101",
  59048=>"010000000",
  59049=>"000000010",
  59050=>"000000000",
  59051=>"000001100",
  59052=>"111111111",
  59053=>"000001000",
  59054=>"011000000",
  59055=>"111111000",
  59056=>"000000000",
  59057=>"001001001",
  59058=>"111000001",
  59059=>"000000000",
  59060=>"111111111",
  59061=>"000111100",
  59062=>"000000000",
  59063=>"001000110",
  59064=>"000001001",
  59065=>"100110110",
  59066=>"000000000",
  59067=>"111111001",
  59068=>"100100111",
  59069=>"000000001",
  59070=>"000000000",
  59071=>"111111111",
  59072=>"100100100",
  59073=>"100111101",
  59074=>"001011111",
  59075=>"000111110",
  59076=>"001011001",
  59077=>"001000000",
  59078=>"111111111",
  59079=>"111011111",
  59080=>"010101011",
  59081=>"111111111",
  59082=>"110111111",
  59083=>"110111011",
  59084=>"111111110",
  59085=>"000000000",
  59086=>"010110111",
  59087=>"000000111",
  59088=>"111111111",
  59089=>"000001111",
  59090=>"011011011",
  59091=>"111111111",
  59092=>"000010100",
  59093=>"000001011",
  59094=>"111000000",
  59095=>"000000000",
  59096=>"111111111",
  59097=>"000010010",
  59098=>"000000110",
  59099=>"111111000",
  59100=>"111111111",
  59101=>"001000001",
  59102=>"111111111",
  59103=>"111011100",
  59104=>"000000000",
  59105=>"111111111",
  59106=>"000000011",
  59107=>"111111111",
  59108=>"111100001",
  59109=>"111111111",
  59110=>"000000110",
  59111=>"000000000",
  59112=>"001100111",
  59113=>"101101101",
  59114=>"000000101",
  59115=>"001000001",
  59116=>"111111110",
  59117=>"000000000",
  59118=>"111001001",
  59119=>"000011011",
  59120=>"000000110",
  59121=>"000101100",
  59122=>"111111111",
  59123=>"000000000",
  59124=>"001011011",
  59125=>"111111111",
  59126=>"101101101",
  59127=>"111111111",
  59128=>"000000000",
  59129=>"111101000",
  59130=>"111111111",
  59131=>"100111000",
  59132=>"000000001",
  59133=>"110110000",
  59134=>"111111101",
  59135=>"000000001",
  59136=>"000000000",
  59137=>"111000000",
  59138=>"000000110",
  59139=>"111111000",
  59140=>"111111000",
  59141=>"101000000",
  59142=>"000000000",
  59143=>"101100010",
  59144=>"000000000",
  59145=>"000000000",
  59146=>"010000000",
  59147=>"100110000",
  59148=>"110100100",
  59149=>"111001000",
  59150=>"000000000",
  59151=>"110000000",
  59152=>"110000000",
  59153=>"111111101",
  59154=>"111111111",
  59155=>"111111011",
  59156=>"100010000",
  59157=>"100111111",
  59158=>"011011001",
  59159=>"111111111",
  59160=>"101111011",
  59161=>"011011111",
  59162=>"111111101",
  59163=>"111111111",
  59164=>"001001011",
  59165=>"100111111",
  59166=>"000000000",
  59167=>"000001111",
  59168=>"000100000",
  59169=>"000001000",
  59170=>"000000000",
  59171=>"111011001",
  59172=>"000000000",
  59173=>"000000000",
  59174=>"011011000",
  59175=>"000001111",
  59176=>"111110111",
  59177=>"000000011",
  59178=>"111111111",
  59179=>"000000000",
  59180=>"000000001",
  59181=>"111011000",
  59182=>"111111111",
  59183=>"111110000",
  59184=>"000000000",
  59185=>"110000000",
  59186=>"000000000",
  59187=>"101111111",
  59188=>"111110000",
  59189=>"011001111",
  59190=>"000010111",
  59191=>"011010000",
  59192=>"111111010",
  59193=>"111111000",
  59194=>"100110111",
  59195=>"000100111",
  59196=>"111111111",
  59197=>"110111101",
  59198=>"000111011",
  59199=>"011011011",
  59200=>"111111000",
  59201=>"000100110",
  59202=>"111111101",
  59203=>"111111111",
  59204=>"111000111",
  59205=>"111110110",
  59206=>"000000000",
  59207=>"000000100",
  59208=>"001001111",
  59209=>"110111010",
  59210=>"111011010",
  59211=>"111111111",
  59212=>"111111111",
  59213=>"011000000",
  59214=>"000001110",
  59215=>"001000000",
  59216=>"000010001",
  59217=>"000000000",
  59218=>"000000000",
  59219=>"111111111",
  59220=>"000000000",
  59221=>"000000000",
  59222=>"000000000",
  59223=>"111100001",
  59224=>"001001111",
  59225=>"001000011",
  59226=>"000000100",
  59227=>"111011000",
  59228=>"011111111",
  59229=>"000111001",
  59230=>"000000000",
  59231=>"011011000",
  59232=>"111111110",
  59233=>"111000100",
  59234=>"000001100",
  59235=>"101001000",
  59236=>"110111111",
  59237=>"001001001",
  59238=>"100101111",
  59239=>"001001001",
  59240=>"111111111",
  59241=>"000000000",
  59242=>"001001011",
  59243=>"111111111",
  59244=>"100000001",
  59245=>"000000111",
  59246=>"000000000",
  59247=>"000111111",
  59248=>"000000000",
  59249=>"000001011",
  59250=>"111111111",
  59251=>"000100111",
  59252=>"000000000",
  59253=>"000000000",
  59254=>"001001111",
  59255=>"000000000",
  59256=>"000000000",
  59257=>"000000000",
  59258=>"101100111",
  59259=>"000001111",
  59260=>"100111000",
  59261=>"000000000",
  59262=>"001000000",
  59263=>"100110110",
  59264=>"111111111",
  59265=>"000111111",
  59266=>"111110000",
  59267=>"111111111",
  59268=>"000000000",
  59269=>"000000110",
  59270=>"011011000",
  59271=>"000000000",
  59272=>"000000000",
  59273=>"111000011",
  59274=>"001011000",
  59275=>"100111110",
  59276=>"111111001",
  59277=>"100110100",
  59278=>"000010110",
  59279=>"000000111",
  59280=>"000000000",
  59281=>"011011111",
  59282=>"101100111",
  59283=>"001000100",
  59284=>"001000000",
  59285=>"000010010",
  59286=>"000000000",
  59287=>"000000001",
  59288=>"100111111",
  59289=>"111111111",
  59290=>"000011111",
  59291=>"111111111",
  59292=>"011000000",
  59293=>"000000001",
  59294=>"111011000",
  59295=>"111110110",
  59296=>"111111111",
  59297=>"100000000",
  59298=>"000000111",
  59299=>"000000000",
  59300=>"110000000",
  59301=>"111000110",
  59302=>"111001000",
  59303=>"011000001",
  59304=>"111111111",
  59305=>"001010000",
  59306=>"000000000",
  59307=>"000011000",
  59308=>"000000000",
  59309=>"111001000",
  59310=>"000000001",
  59311=>"100100111",
  59312=>"111011011",
  59313=>"111000000",
  59314=>"110111000",
  59315=>"111111110",
  59316=>"001000001",
  59317=>"000111001",
  59318=>"011111100",
  59319=>"111011101",
  59320=>"000100111",
  59321=>"111000000",
  59322=>"000100000",
  59323=>"111111111",
  59324=>"000000000",
  59325=>"000000000",
  59326=>"000111111",
  59327=>"011110011",
  59328=>"000000000",
  59329=>"111111111",
  59330=>"000111111",
  59331=>"000010110",
  59332=>"110110000",
  59333=>"000000000",
  59334=>"111001001",
  59335=>"100100110",
  59336=>"000000000",
  59337=>"000111110",
  59338=>"000000110",
  59339=>"000000000",
  59340=>"111011011",
  59341=>"111001111",
  59342=>"001001000",
  59343=>"000111111",
  59344=>"001111000",
  59345=>"111111110",
  59346=>"111001001",
  59347=>"111011011",
  59348=>"000100100",
  59349=>"000110100",
  59350=>"011000000",
  59351=>"000000001",
  59352=>"000000000",
  59353=>"111000000",
  59354=>"000000000",
  59355=>"000111111",
  59356=>"000001001",
  59357=>"000001011",
  59358=>"111111111",
  59359=>"001001000",
  59360=>"110110000",
  59361=>"111111111",
  59362=>"000000000",
  59363=>"000011111",
  59364=>"111100100",
  59365=>"101000001",
  59366=>"000000000",
  59367=>"111111111",
  59368=>"111111111",
  59369=>"100000000",
  59370=>"101111111",
  59371=>"111000000",
  59372=>"000000000",
  59373=>"000000101",
  59374=>"011001111",
  59375=>"000000000",
  59376=>"000010000",
  59377=>"111111111",
  59378=>"111111111",
  59379=>"111111111",
  59380=>"000111111",
  59381=>"000111111",
  59382=>"011011000",
  59383=>"110011001",
  59384=>"111111010",
  59385=>"100000111",
  59386=>"110111111",
  59387=>"000010000",
  59388=>"011111100",
  59389=>"011001111",
  59390=>"111001001",
  59391=>"010111110",
  59392=>"000000000",
  59393=>"000000110",
  59394=>"111000101",
  59395=>"000000100",
  59396=>"010111111",
  59397=>"001000010",
  59398=>"111111100",
  59399=>"000000000",
  59400=>"111111111",
  59401=>"101100100",
  59402=>"111111111",
  59403=>"000001011",
  59404=>"000000110",
  59405=>"000100000",
  59406=>"101100111",
  59407=>"000000100",
  59408=>"111111011",
  59409=>"111111101",
  59410=>"000000000",
  59411=>"111001001",
  59412=>"000000000",
  59413=>"000000000",
  59414=>"000000000",
  59415=>"111110110",
  59416=>"001011001",
  59417=>"011011011",
  59418=>"111111111",
  59419=>"001001111",
  59420=>"000000000",
  59421=>"111010000",
  59422=>"111101101",
  59423=>"111111111",
  59424=>"001010011",
  59425=>"000000000",
  59426=>"000000000",
  59427=>"000000000",
  59428=>"000000101",
  59429=>"111111111",
  59430=>"000001000",
  59431=>"100100100",
  59432=>"110100111",
  59433=>"111111111",
  59434=>"100100111",
  59435=>"111011000",
  59436=>"111111101",
  59437=>"101111100",
  59438=>"111111110",
  59439=>"101100111",
  59440=>"000000010",
  59441=>"001000000",
  59442=>"110100100",
  59443=>"111101111",
  59444=>"000100110",
  59445=>"000010110",
  59446=>"111111110",
  59447=>"011111111",
  59448=>"100111111",
  59449=>"101100000",
  59450=>"000111111",
  59451=>"010000000",
  59452=>"100000000",
  59453=>"100000001",
  59454=>"010010010",
  59455=>"000000000",
  59456=>"111111111",
  59457=>"111000000",
  59458=>"101111111",
  59459=>"111111111",
  59460=>"111111110",
  59461=>"000001001",
  59462=>"110110110",
  59463=>"111111110",
  59464=>"110110110",
  59465=>"011111111",
  59466=>"000000000",
  59467=>"000000111",
  59468=>"111110111",
  59469=>"111111101",
  59470=>"000101101",
  59471=>"111111010",
  59472=>"001000011",
  59473=>"001111011",
  59474=>"000000000",
  59475=>"000000010",
  59476=>"101111000",
  59477=>"101101000",
  59478=>"000000000",
  59479=>"000000010",
  59480=>"111011111",
  59481=>"000000000",
  59482=>"111111000",
  59483=>"111111111",
  59484=>"111001000",
  59485=>"000000000",
  59486=>"000001001",
  59487=>"011010000",
  59488=>"000001111",
  59489=>"111111111",
  59490=>"000000000",
  59491=>"000000000",
  59492=>"000000000",
  59493=>"111111111",
  59494=>"001111111",
  59495=>"111111010",
  59496=>"001111111",
  59497=>"000011000",
  59498=>"001111011",
  59499=>"000000000",
  59500=>"110000000",
  59501=>"100000101",
  59502=>"101100111",
  59503=>"011010000",
  59504=>"000100111",
  59505=>"111111111",
  59506=>"001001001",
  59507=>"010010001",
  59508=>"111111111",
  59509=>"111100101",
  59510=>"111111111",
  59511=>"111110110",
  59512=>"111111000",
  59513=>"101000000",
  59514=>"111111101",
  59515=>"001001001",
  59516=>"110111111",
  59517=>"011111111",
  59518=>"100111111",
  59519=>"000000000",
  59520=>"011111111",
  59521=>"011011111",
  59522=>"000000000",
  59523=>"000000000",
  59524=>"001001111",
  59525=>"000000001",
  59526=>"000000000",
  59527=>"111000111",
  59528=>"001000000",
  59529=>"111111011",
  59530=>"111111111",
  59531=>"110111111",
  59532=>"000000010",
  59533=>"000000000",
  59534=>"111110111",
  59535=>"000101111",
  59536=>"000000001",
  59537=>"010010000",
  59538=>"100000000",
  59539=>"101011000",
  59540=>"000000000",
  59541=>"000001101",
  59542=>"111111111",
  59543=>"000000000",
  59544=>"000000011",
  59545=>"000000011",
  59546=>"101000000",
  59547=>"000100000",
  59548=>"000000000",
  59549=>"001000000",
  59550=>"101011011",
  59551=>"110111111",
  59552=>"111111011",
  59553=>"000000000",
  59554=>"101101101",
  59555=>"000000111",
  59556=>"101000000",
  59557=>"101101111",
  59558=>"111101111",
  59559=>"001011011",
  59560=>"111111010",
  59561=>"000000100",
  59562=>"000000000",
  59563=>"001000000",
  59564=>"111111000",
  59565=>"001001001",
  59566=>"000000000",
  59567=>"001000101",
  59568=>"001111100",
  59569=>"111111111",
  59570=>"101101000",
  59571=>"111111001",
  59572=>"111100000",
  59573=>"111111011",
  59574=>"000000000",
  59575=>"110111111",
  59576=>"000010111",
  59577=>"000000000",
  59578=>"101101111",
  59579=>"001001000",
  59580=>"111000000",
  59581=>"010001000",
  59582=>"000000000",
  59583=>"011111001",
  59584=>"000000010",
  59585=>"101011111",
  59586=>"111001001",
  59587=>"000111110",
  59588=>"001001001",
  59589=>"000010011",
  59590=>"000010010",
  59591=>"000000010",
  59592=>"000000000",
  59593=>"000000000",
  59594=>"000001001",
  59595=>"000101111",
  59596=>"111101100",
  59597=>"000011111",
  59598=>"001001000",
  59599=>"000011000",
  59600=>"111111111",
  59601=>"000000010",
  59602=>"000101111",
  59603=>"100010000",
  59604=>"001000000",
  59605=>"101001000",
  59606=>"111111111",
  59607=>"011100000",
  59608=>"000111111",
  59609=>"000000000",
  59610=>"111111110",
  59611=>"111111111",
  59612=>"111000100",
  59613=>"111110111",
  59614=>"000000000",
  59615=>"010010000",
  59616=>"110010000",
  59617=>"010011011",
  59618=>"100000000",
  59619=>"100100001",
  59620=>"111101000",
  59621=>"110110100",
  59622=>"000011011",
  59623=>"000000000",
  59624=>"000000110",
  59625=>"111101111",
  59626=>"111111111",
  59627=>"111111111",
  59628=>"111111111",
  59629=>"000000111",
  59630=>"000000111",
  59631=>"000001111",
  59632=>"011111111",
  59633=>"111111111",
  59634=>"011000000",
  59635=>"000000000",
  59636=>"111101101",
  59637=>"110100001",
  59638=>"000100101",
  59639=>"010010000",
  59640=>"000000000",
  59641=>"000000000",
  59642=>"111100000",
  59643=>"010101101",
  59644=>"110111110",
  59645=>"100000000",
  59646=>"101000100",
  59647=>"111111111",
  59648=>"111111111",
  59649=>"001011001",
  59650=>"111111111",
  59651=>"111111110",
  59652=>"111011111",
  59653=>"001001001",
  59654=>"010011011",
  59655=>"111001111",
  59656=>"111111110",
  59657=>"111011111",
  59658=>"000000000",
  59659=>"111111111",
  59660=>"000000000",
  59661=>"000000000",
  59662=>"010010110",
  59663=>"000011011",
  59664=>"111011000",
  59665=>"000000000",
  59666=>"111111000",
  59667=>"011011000",
  59668=>"011001000",
  59669=>"100110111",
  59670=>"001111111",
  59671=>"000000000",
  59672=>"000000000",
  59673=>"000000001",
  59674=>"000000000",
  59675=>"111111111",
  59676=>"111111001",
  59677=>"000000000",
  59678=>"111111111",
  59679=>"111100100",
  59680=>"100100100",
  59681=>"111111010",
  59682=>"000000000",
  59683=>"111101000",
  59684=>"010110110",
  59685=>"000001111",
  59686=>"010111111",
  59687=>"000100001",
  59688=>"110100110",
  59689=>"100100000",
  59690=>"111000001",
  59691=>"111000000",
  59692=>"000000010",
  59693=>"010000000",
  59694=>"111111101",
  59695=>"000000000",
  59696=>"011111111",
  59697=>"000000000",
  59698=>"111111111",
  59699=>"111111111",
  59700=>"100000000",
  59701=>"001111100",
  59702=>"011111111",
  59703=>"000000000",
  59704=>"000000000",
  59705=>"000000001",
  59706=>"100101101",
  59707=>"011011111",
  59708=>"101111001",
  59709=>"000100110",
  59710=>"000000100",
  59711=>"000000001",
  59712=>"000000111",
  59713=>"111111111",
  59714=>"000000101",
  59715=>"000000000",
  59716=>"000001011",
  59717=>"111111111",
  59718=>"011111111",
  59719=>"111010000",
  59720=>"000101111",
  59721=>"000111111",
  59722=>"000000000",
  59723=>"010000000",
  59724=>"111100000",
  59725=>"100111111",
  59726=>"001101111",
  59727=>"000000110",
  59728=>"010000001",
  59729=>"011001000",
  59730=>"110111110",
  59731=>"111010110",
  59732=>"000111111",
  59733=>"011011001",
  59734=>"000011111",
  59735=>"111111001",
  59736=>"010110010",
  59737=>"101111111",
  59738=>"000000100",
  59739=>"111000000",
  59740=>"111000111",
  59741=>"101111111",
  59742=>"001101101",
  59743=>"110110010",
  59744=>"000001001",
  59745=>"000000000",
  59746=>"000110011",
  59747=>"000000000",
  59748=>"000010000",
  59749=>"000000000",
  59750=>"001101101",
  59751=>"000000111",
  59752=>"001011001",
  59753=>"011000100",
  59754=>"100000000",
  59755=>"011110111",
  59756=>"000110111",
  59757=>"001100000",
  59758=>"000000110",
  59759=>"000001011",
  59760=>"000000111",
  59761=>"111111111",
  59762=>"000000110",
  59763=>"111111101",
  59764=>"000000000",
  59765=>"111111111",
  59766=>"101101000",
  59767=>"001111111",
  59768=>"000000000",
  59769=>"111001001",
  59770=>"111111111",
  59771=>"111111111",
  59772=>"010110111",
  59773=>"001000000",
  59774=>"111111111",
  59775=>"000000000",
  59776=>"110110110",
  59777=>"011111110",
  59778=>"100100000",
  59779=>"111111000",
  59780=>"000000000",
  59781=>"000010111",
  59782=>"111111111",
  59783=>"000000111",
  59784=>"000101111",
  59785=>"011011110",
  59786=>"000000001",
  59787=>"011000100",
  59788=>"000000000",
  59789=>"000100111",
  59790=>"000010010",
  59791=>"101000100",
  59792=>"100110111",
  59793=>"111111100",
  59794=>"011001111",
  59795=>"000100110",
  59796=>"111111111",
  59797=>"000011001",
  59798=>"001111011",
  59799=>"011010011",
  59800=>"000100101",
  59801=>"110110111",
  59802=>"111111111",
  59803=>"000001111",
  59804=>"000001000",
  59805=>"111000000",
  59806=>"101101111",
  59807=>"111111111",
  59808=>"100000000",
  59809=>"100000001",
  59810=>"000000000",
  59811=>"000001001",
  59812=>"010010011",
  59813=>"011111111",
  59814=>"111101001",
  59815=>"111110000",
  59816=>"011111111",
  59817=>"001111111",
  59818=>"111111111",
  59819=>"111111101",
  59820=>"000000000",
  59821=>"111111101",
  59822=>"111001011",
  59823=>"101001101",
  59824=>"111001100",
  59825=>"001001101",
  59826=>"000111111",
  59827=>"111100000",
  59828=>"000110111",
  59829=>"111111111",
  59830=>"000000000",
  59831=>"111111111",
  59832=>"111111100",
  59833=>"111111001",
  59834=>"011010000",
  59835=>"110110111",
  59836=>"110000000",
  59837=>"000010011",
  59838=>"000000000",
  59839=>"001001001",
  59840=>"000000001",
  59841=>"000001111",
  59842=>"011011000",
  59843=>"110000000",
  59844=>"000001011",
  59845=>"001111110",
  59846=>"001000110",
  59847=>"011111111",
  59848=>"000000000",
  59849=>"110110111",
  59850=>"000111111",
  59851=>"000000000",
  59852=>"000000000",
  59853=>"000000000",
  59854=>"000100110",
  59855=>"111111111",
  59856=>"000001111",
  59857=>"111111111",
  59858=>"111111111",
  59859=>"000000101",
  59860=>"111110011",
  59861=>"010000000",
  59862=>"011111000",
  59863=>"000011011",
  59864=>"001001000",
  59865=>"111111111",
  59866=>"100100111",
  59867=>"111111000",
  59868=>"100100100",
  59869=>"101101111",
  59870=>"001011111",
  59871=>"000001000",
  59872=>"011111111",
  59873=>"111111011",
  59874=>"100111111",
  59875=>"100100111",
  59876=>"000100000",
  59877=>"110100111",
  59878=>"000000011",
  59879=>"111111111",
  59880=>"000000001",
  59881=>"011011000",
  59882=>"011001111",
  59883=>"000111011",
  59884=>"000010111",
  59885=>"000000000",
  59886=>"110111111",
  59887=>"111111111",
  59888=>"111111111",
  59889=>"011111110",
  59890=>"001001100",
  59891=>"001000001",
  59892=>"101001011",
  59893=>"000000000",
  59894=>"000101101",
  59895=>"011001000",
  59896=>"010000000",
  59897=>"000000000",
  59898=>"000000000",
  59899=>"000000111",
  59900=>"111100110",
  59901=>"001000110",
  59902=>"000001101",
  59903=>"001111111",
  59904=>"111111000",
  59905=>"001011000",
  59906=>"000110111",
  59907=>"011111111",
  59908=>"000111111",
  59909=>"100101000",
  59910=>"111111111",
  59911=>"101111111",
  59912=>"000001001",
  59913=>"000111010",
  59914=>"111111000",
  59915=>"111111000",
  59916=>"111111000",
  59917=>"111111011",
  59918=>"111111001",
  59919=>"111111111",
  59920=>"111111111",
  59921=>"110111111",
  59922=>"111111111",
  59923=>"000000000",
  59924=>"111111111",
  59925=>"000010111",
  59926=>"111101111",
  59927=>"100110111",
  59928=>"110111111",
  59929=>"000000001",
  59930=>"111001111",
  59931=>"111111000",
  59932=>"000000000",
  59933=>"111111111",
  59934=>"000000111",
  59935=>"000000000",
  59936=>"001011111",
  59937=>"111111111",
  59938=>"111001000",
  59939=>"111111111",
  59940=>"111111111",
  59941=>"000000000",
  59942=>"110010000",
  59943=>"001000101",
  59944=>"001111111",
  59945=>"000000011",
  59946=>"000010010",
  59947=>"101100000",
  59948=>"100111111",
  59949=>"111111111",
  59950=>"001000000",
  59951=>"111111001",
  59952=>"000011111",
  59953=>"001011111",
  59954=>"001000111",
  59955=>"111011010",
  59956=>"110010111",
  59957=>"111111111",
  59958=>"000111111",
  59959=>"000000001",
  59960=>"000000000",
  59961=>"000000111",
  59962=>"011011000",
  59963=>"110110000",
  59964=>"001000010",
  59965=>"000000000",
  59966=>"111111111",
  59967=>"111111000",
  59968=>"111000000",
  59969=>"000000011",
  59970=>"000000000",
  59971=>"000000000",
  59972=>"001001001",
  59973=>"000000000",
  59974=>"000000011",
  59975=>"111111111",
  59976=>"011001000",
  59977=>"001000000",
  59978=>"111110100",
  59979=>"001101000",
  59980=>"111000000",
  59981=>"111001011",
  59982=>"000000000",
  59983=>"000000000",
  59984=>"000000001",
  59985=>"100000111",
  59986=>"000000000",
  59987=>"110000111",
  59988=>"000000000",
  59989=>"000000000",
  59990=>"000001000",
  59991=>"100100110",
  59992=>"111111111",
  59993=>"000000000",
  59994=>"000000000",
  59995=>"000001111",
  59996=>"110111000",
  59997=>"111111100",
  59998=>"110111111",
  59999=>"111001001",
  60000=>"111100000",
  60001=>"000010111",
  60002=>"110110100",
  60003=>"111111000",
  60004=>"000000000",
  60005=>"100111100",
  60006=>"000000111",
  60007=>"000010111",
  60008=>"000000000",
  60009=>"110111111",
  60010=>"000011111",
  60011=>"011011000",
  60012=>"110110000",
  60013=>"101111100",
  60014=>"000000101",
  60015=>"111111101",
  60016=>"100000000",
  60017=>"000000110",
  60018=>"111111111",
  60019=>"010010000",
  60020=>"000000010",
  60021=>"111111111",
  60022=>"000000000",
  60023=>"000000000",
  60024=>"111111110",
  60025=>"111110000",
  60026=>"111000000",
  60027=>"000010111",
  60028=>"000111111",
  60029=>"111111111",
  60030=>"000000000",
  60031=>"001000000",
  60032=>"000000000",
  60033=>"110100001",
  60034=>"111111111",
  60035=>"111001000",
  60036=>"100000000",
  60037=>"000000000",
  60038=>"001001000",
  60039=>"111111111",
  60040=>"110000000",
  60041=>"100100100",
  60042=>"111000000",
  60043=>"111111000",
  60044=>"111111000",
  60045=>"111111111",
  60046=>"100111101",
  60047=>"001001000",
  60048=>"000000011",
  60049=>"000000000",
  60050=>"100000100",
  60051=>"111111111",
  60052=>"110111000",
  60053=>"000000000",
  60054=>"000000000",
  60055=>"000100100",
  60056=>"100000001",
  60057=>"110101100",
  60058=>"111111111",
  60059=>"000000000",
  60060=>"100111111",
  60061=>"011000000",
  60062=>"000000110",
  60063=>"000111111",
  60064=>"011011111",
  60065=>"010000000",
  60066=>"000000010",
  60067=>"111111111",
  60068=>"001001000",
  60069=>"000010000",
  60070=>"111111111",
  60071=>"110100100",
  60072=>"000110110",
  60073=>"111111111",
  60074=>"001011111",
  60075=>"000000000",
  60076=>"000110110",
  60077=>"001000000",
  60078=>"110100100",
  60079=>"011111000",
  60080=>"000000000",
  60081=>"011011111",
  60082=>"110110111",
  60083=>"000000000",
  60084=>"111011000",
  60085=>"111111111",
  60086=>"111101111",
  60087=>"110100000",
  60088=>"101101111",
  60089=>"111110100",
  60090=>"101000100",
  60091=>"101011010",
  60092=>"101111011",
  60093=>"110110111",
  60094=>"000000000",
  60095=>"000111011",
  60096=>"000111111",
  60097=>"000111111",
  60098=>"000001000",
  60099=>"000000000",
  60100=>"000001111",
  60101=>"111100110",
  60102=>"000100111",
  60103=>"100100100",
  60104=>"111111111",
  60105=>"000000111",
  60106=>"111111101",
  60107=>"101101111",
  60108=>"000000001",
  60109=>"110111111",
  60110=>"000010000",
  60111=>"111001000",
  60112=>"000000000",
  60113=>"111000000",
  60114=>"111111000",
  60115=>"000100110",
  60116=>"000000000",
  60117=>"001001110",
  60118=>"111001000",
  60119=>"000000000",
  60120=>"000000000",
  60121=>"001001000",
  60122=>"000010111",
  60123=>"000000000",
  60124=>"111011001",
  60125=>"001001000",
  60126=>"111111111",
  60127=>"100110111",
  60128=>"010000000",
  60129=>"111101000",
  60130=>"100000010",
  60131=>"000000000",
  60132=>"100100111",
  60133=>"000000011",
  60134=>"111111111",
  60135=>"111111111",
  60136=>"111111011",
  60137=>"000000000",
  60138=>"000000001",
  60139=>"000110010",
  60140=>"111111000",
  60141=>"111111001",
  60142=>"111010110",
  60143=>"111111111",
  60144=>"100000100",
  60145=>"100100000",
  60146=>"111000110",
  60147=>"011000000",
  60148=>"000000010",
  60149=>"001000000",
  60150=>"100100000",
  60151=>"000000000",
  60152=>"111111011",
  60153=>"110110111",
  60154=>"111111111",
  60155=>"000111111",
  60156=>"001000110",
  60157=>"110110110",
  60158=>"110110000",
  60159=>"001111101",
  60160=>"111000000",
  60161=>"000100100",
  60162=>"000000000",
  60163=>"000000010",
  60164=>"000010100",
  60165=>"011111111",
  60166=>"000000001",
  60167=>"011111111",
  60168=>"000111111",
  60169=>"111010000",
  60170=>"110100000",
  60171=>"001001000",
  60172=>"100000100",
  60173=>"111110111",
  60174=>"000000000",
  60175=>"111111011",
  60176=>"100100111",
  60177=>"111000000",
  60178=>"001000000",
  60179=>"000000000",
  60180=>"001011111",
  60181=>"000100111",
  60182=>"000000100",
  60183=>"111111000",
  60184=>"111111111",
  60185=>"110100000",
  60186=>"000000000",
  60187=>"111111101",
  60188=>"001000000",
  60189=>"111111010",
  60190=>"000111111",
  60191=>"111000000",
  60192=>"000000000",
  60193=>"000010000",
  60194=>"000111111",
  60195=>"011011111",
  60196=>"100000000",
  60197=>"000000011",
  60198=>"100101001",
  60199=>"000000000",
  60200=>"000001100",
  60201=>"111111111",
  60202=>"111111111",
  60203=>"111111111",
  60204=>"000000001",
  60205=>"111111110",
  60206=>"100111000",
  60207=>"100100100",
  60208=>"000000101",
  60209=>"000100111",
  60210=>"001010110",
  60211=>"000000001",
  60212=>"001001001",
  60213=>"000000100",
  60214=>"000100111",
  60215=>"111111000",
  60216=>"000000000",
  60217=>"111111111",
  60218=>"111111111",
  60219=>"100000100",
  60220=>"000000000",
  60221=>"000000000",
  60222=>"000001000",
  60223=>"000111111",
  60224=>"000000000",
  60225=>"100110000",
  60226=>"101111111",
  60227=>"010110111",
  60228=>"000000000",
  60229=>"000000000",
  60230=>"111111111",
  60231=>"111111111",
  60232=>"000100101",
  60233=>"100010000",
  60234=>"111111000",
  60235=>"110100111",
  60236=>"111101101",
  60237=>"000000000",
  60238=>"000001111",
  60239=>"000000001",
  60240=>"100100111",
  60241=>"110000010",
  60242=>"111111111",
  60243=>"000111111",
  60244=>"111101111",
  60245=>"000000011",
  60246=>"111111010",
  60247=>"010010111",
  60248=>"000000100",
  60249=>"111101000",
  60250=>"000000000",
  60251=>"111111110",
  60252=>"000000000",
  60253=>"000011000",
  60254=>"010010011",
  60255=>"111111111",
  60256=>"111111000",
  60257=>"111111111",
  60258=>"011001101",
  60259=>"000000000",
  60260=>"111111111",
  60261=>"000111111",
  60262=>"111111111",
  60263=>"001111111",
  60264=>"001001100",
  60265=>"000000000",
  60266=>"000000111",
  60267=>"001000000",
  60268=>"001011000",
  60269=>"011011000",
  60270=>"011011111",
  60271=>"011000000",
  60272=>"001101000",
  60273=>"001001000",
  60274=>"110110011",
  60275=>"111111111",
  60276=>"000000000",
  60277=>"000010010",
  60278=>"110111000",
  60279=>"111110110",
  60280=>"000000000",
  60281=>"100010011",
  60282=>"100001111",
  60283=>"000100111",
  60284=>"000000000",
  60285=>"000111111",
  60286=>"100111110",
  60287=>"100101000",
  60288=>"111111011",
  60289=>"101000000",
  60290=>"000001111",
  60291=>"000000000",
  60292=>"000010000",
  60293=>"111111110",
  60294=>"111100111",
  60295=>"111001000",
  60296=>"111111111",
  60297=>"111000000",
  60298=>"111110000",
  60299=>"011000111",
  60300=>"000000000",
  60301=>"111000000",
  60302=>"101111111",
  60303=>"100000000",
  60304=>"100111111",
  60305=>"000000000",
  60306=>"111111000",
  60307=>"000010000",
  60308=>"000000101",
  60309=>"000001011",
  60310=>"111111100",
  60311=>"001000110",
  60312=>"111001000",
  60313=>"111000000",
  60314=>"011001001",
  60315=>"111111111",
  60316=>"000000110",
  60317=>"011001111",
  60318=>"100100111",
  60319=>"110110000",
  60320=>"000100111",
  60321=>"010100110",
  60322=>"000000000",
  60323=>"011111111",
  60324=>"011111101",
  60325=>"000000000",
  60326=>"111110000",
  60327=>"111010010",
  60328=>"000001001",
  60329=>"000000000",
  60330=>"111001000",
  60331=>"111000111",
  60332=>"000000110",
  60333=>"111111110",
  60334=>"000000001",
  60335=>"000000000",
  60336=>"011111111",
  60337=>"111111111",
  60338=>"100111000",
  60339=>"010111111",
  60340=>"000000100",
  60341=>"000000111",
  60342=>"000010000",
  60343=>"010110110",
  60344=>"000000000",
  60345=>"100000000",
  60346=>"111110110",
  60347=>"100100000",
  60348=>"110100000",
  60349=>"000000101",
  60350=>"111111111",
  60351=>"100100100",
  60352=>"011010000",
  60353=>"100100110",
  60354=>"111111111",
  60355=>"000000000",
  60356=>"110111100",
  60357=>"000000001",
  60358=>"000000100",
  60359=>"001001000",
  60360=>"111111000",
  60361=>"000000011",
  60362=>"000000000",
  60363=>"110010110",
  60364=>"111111100",
  60365=>"111111111",
  60366=>"110000000",
  60367=>"110110110",
  60368=>"000000000",
  60369=>"110101000",
  60370=>"001011001",
  60371=>"000000111",
  60372=>"111111111",
  60373=>"101111110",
  60374=>"001000111",
  60375=>"110100000",
  60376=>"100010111",
  60377=>"000110110",
  60378=>"111010000",
  60379=>"100111110",
  60380=>"110111100",
  60381=>"000010000",
  60382=>"110110000",
  60383=>"000111111",
  60384=>"110010000",
  60385=>"111110101",
  60386=>"111000000",
  60387=>"000000000",
  60388=>"011011001",
  60389=>"001001000",
  60390=>"001001111",
  60391=>"000000000",
  60392=>"110111011",
  60393=>"100000000",
  60394=>"000000000",
  60395=>"001011111",
  60396=>"111111000",
  60397=>"000000000",
  60398=>"110110111",
  60399=>"110111111",
  60400=>"100001001",
  60401=>"100000111",
  60402=>"000000000",
  60403=>"111111100",
  60404=>"111111000",
  60405=>"101101111",
  60406=>"111110110",
  60407=>"001011111",
  60408=>"111111101",
  60409=>"100000001",
  60410=>"000010010",
  60411=>"000000000",
  60412=>"111111110",
  60413=>"000000100",
  60414=>"000011111",
  60415=>"101001111",
  60416=>"111100110",
  60417=>"111000100",
  60418=>"001001111",
  60419=>"000000000",
  60420=>"110111111",
  60421=>"000001001",
  60422=>"000000000",
  60423=>"111111111",
  60424=>"111111001",
  60425=>"111111111",
  60426=>"111100100",
  60427=>"111100000",
  60428=>"000000000",
  60429=>"001101111",
  60430=>"000000011",
  60431=>"110111111",
  60432=>"000000000",
  60433=>"010111011",
  60434=>"011111011",
  60435=>"001000000",
  60436=>"111111000",
  60437=>"001111111",
  60438=>"000000000",
  60439=>"100100000",
  60440=>"111101001",
  60441=>"001011111",
  60442=>"111111111",
  60443=>"000000110",
  60444=>"000000001",
  60445=>"000101000",
  60446=>"111011011",
  60447=>"001111111",
  60448=>"111000000",
  60449=>"010000000",
  60450=>"001011011",
  60451=>"000000101",
  60452=>"111111111",
  60453=>"111111111",
  60454=>"100000000",
  60455=>"111000000",
  60456=>"011111110",
  60457=>"001000000",
  60458=>"000000111",
  60459=>"000000000",
  60460=>"111001000",
  60461=>"000000000",
  60462=>"110000010",
  60463=>"111111111",
  60464=>"111100101",
  60465=>"110111000",
  60466=>"111110100",
  60467=>"000000000",
  60468=>"000000000",
  60469=>"010010010",
  60470=>"000000000",
  60471=>"111000000",
  60472=>"000000000",
  60473=>"001001001",
  60474=>"101000000",
  60475=>"111110000",
  60476=>"001001000",
  60477=>"011100000",
  60478=>"010111100",
  60479=>"111011000",
  60480=>"000000100",
  60481=>"101011000",
  60482=>"110111010",
  60483=>"101001010",
  60484=>"000000011",
  60485=>"111111110",
  60486=>"111111111",
  60487=>"111111111",
  60488=>"111100001",
  60489=>"000000111",
  60490=>"111000111",
  60491=>"110111111",
  60492=>"011000000",
  60493=>"111111111",
  60494=>"011000000",
  60495=>"111111111",
  60496=>"000000000",
  60497=>"000000000",
  60498=>"000000000",
  60499=>"011111111",
  60500=>"111001001",
  60501=>"000000000",
  60502=>"111111110",
  60503=>"110111110",
  60504=>"111011010",
  60505=>"000000000",
  60506=>"000000110",
  60507=>"011111110",
  60508=>"000000000",
  60509=>"000000000",
  60510=>"000000000",
  60511=>"000100101",
  60512=>"111101111",
  60513=>"000000000",
  60514=>"010000000",
  60515=>"111111111",
  60516=>"001011111",
  60517=>"111011001",
  60518=>"111111011",
  60519=>"000000000",
  60520=>"000000000",
  60521=>"111101111",
  60522=>"000000000",
  60523=>"110010010",
  60524=>"011011000",
  60525=>"111111111",
  60526=>"000000000",
  60527=>"000100110",
  60528=>"001001111",
  60529=>"000000110",
  60530=>"001011011",
  60531=>"000000000",
  60532=>"111111111",
  60533=>"000010111",
  60534=>"001000000",
  60535=>"000001001",
  60536=>"000000000",
  60537=>"100000000",
  60538=>"000011011",
  60539=>"000000001",
  60540=>"001001111",
  60541=>"000011010",
  60542=>"000000000",
  60543=>"000000000",
  60544=>"100111111",
  60545=>"000000000",
  60546=>"111110100",
  60547=>"100000000",
  60548=>"111100000",
  60549=>"000000000",
  60550=>"001000000",
  60551=>"111000000",
  60552=>"111011001",
  60553=>"000000101",
  60554=>"111111011",
  60555=>"000000000",
  60556=>"100000100",
  60557=>"111111010",
  60558=>"111101000",
  60559=>"011010111",
  60560=>"010000010",
  60561=>"111000001",
  60562=>"000000000",
  60563=>"101100000",
  60564=>"011000000",
  60565=>"100000111",
  60566=>"000000011",
  60567=>"110100000",
  60568=>"001000001",
  60569=>"100000000",
  60570=>"111010000",
  60571=>"101000001",
  60572=>"111111111",
  60573=>"001001111",
  60574=>"111010000",
  60575=>"000000000",
  60576=>"010111110",
  60577=>"101001101",
  60578=>"001001011",
  60579=>"110000000",
  60580=>"000110111",
  60581=>"011000111",
  60582=>"111110010",
  60583=>"011111011",
  60584=>"000000000",
  60585=>"000000000",
  60586=>"000000000",
  60587=>"111001001",
  60588=>"001111111",
  60589=>"111111001",
  60590=>"000000000",
  60591=>"100000010",
  60592=>"000000000",
  60593=>"100111111",
  60594=>"110111111",
  60595=>"100100101",
  60596=>"011010111",
  60597=>"111111111",
  60598=>"111111111",
  60599=>"111000000",
  60600=>"000000111",
  60601=>"000000000",
  60602=>"000000000",
  60603=>"111100000",
  60604=>"110010000",
  60605=>"111000000",
  60606=>"111111111",
  60607=>"000000000",
  60608=>"111111111",
  60609=>"111111111",
  60610=>"110000000",
  60611=>"000000000",
  60612=>"011000000",
  60613=>"111111111",
  60614=>"011011000",
  60615=>"110000011",
  60616=>"111000100",
  60617=>"111111111",
  60618=>"100000000",
  60619=>"110110110",
  60620=>"000000000",
  60621=>"100000001",
  60622=>"001000011",
  60623=>"000000000",
  60624=>"111000101",
  60625=>"111111010",
  60626=>"010000111",
  60627=>"000000000",
  60628=>"000000000",
  60629=>"000000000",
  60630=>"000000001",
  60631=>"000001011",
  60632=>"000110111",
  60633=>"110110100",
  60634=>"000001001",
  60635=>"000000000",
  60636=>"111101101",
  60637=>"011001010",
  60638=>"111111111",
  60639=>"001100000",
  60640=>"000000000",
  60641=>"000010000",
  60642=>"000000000",
  60643=>"001101000",
  60644=>"000000000",
  60645=>"110111111",
  60646=>"111111111",
  60647=>"111111111",
  60648=>"111110010",
  60649=>"111110100",
  60650=>"000000000",
  60651=>"101111111",
  60652=>"000110111",
  60653=>"001111111",
  60654=>"111011000",
  60655=>"110000000",
  60656=>"111111110",
  60657=>"111111011",
  60658=>"101000000",
  60659=>"000000000",
  60660=>"000000000",
  60661=>"000100000",
  60662=>"000000000",
  60663=>"111110100",
  60664=>"000000111",
  60665=>"111000001",
  60666=>"011001000",
  60667=>"111111000",
  60668=>"000011011",
  60669=>"111000000",
  60670=>"011110110",
  60671=>"000100111",
  60672=>"001000000",
  60673=>"000011011",
  60674=>"000000100",
  60675=>"000000000",
  60676=>"000110111",
  60677=>"110110010",
  60678=>"111111100",
  60679=>"000000110",
  60680=>"110111111",
  60681=>"111111111",
  60682=>"000000101",
  60683=>"000000000",
  60684=>"000000000",
  60685=>"000000000",
  60686=>"000000001",
  60687=>"100111111",
  60688=>"000001001",
  60689=>"001000001",
  60690=>"111001000",
  60691=>"000111001",
  60692=>"000000000",
  60693=>"100001110",
  60694=>"001001111",
  60695=>"111111111",
  60696=>"000000101",
  60697=>"010000111",
  60698=>"111101111",
  60699=>"111000000",
  60700=>"110110010",
  60701=>"000010011",
  60702=>"000000000",
  60703=>"111011111",
  60704=>"100111111",
  60705=>"011010110",
  60706=>"000101111",
  60707=>"111111001",
  60708=>"111111100",
  60709=>"000011111",
  60710=>"000000111",
  60711=>"001000101",
  60712=>"000000111",
  60713=>"000000000",
  60714=>"101000111",
  60715=>"100000000",
  60716=>"111111111",
  60717=>"001000011",
  60718=>"000111111",
  60719=>"000000000",
  60720=>"011011111",
  60721=>"110111000",
  60722=>"111111111",
  60723=>"111110000",
  60724=>"000000000",
  60725=>"111111111",
  60726=>"000000000",
  60727=>"001000000",
  60728=>"111110000",
  60729=>"110100110",
  60730=>"111111111",
  60731=>"111010111",
  60732=>"111111111",
  60733=>"111111110",
  60734=>"111000000",
  60735=>"111110110",
  60736=>"011000000",
  60737=>"111101111",
  60738=>"100111111",
  60739=>"000000000",
  60740=>"000010111",
  60741=>"000111111",
  60742=>"111111110",
  60743=>"000000000",
  60744=>"000000111",
  60745=>"000000111",
  60746=>"000000001",
  60747=>"001101000",
  60748=>"001001111",
  60749=>"000110000",
  60750=>"110010000",
  60751=>"100100100",
  60752=>"000000111",
  60753=>"001001101",
  60754=>"000100111",
  60755=>"000000000",
  60756=>"111111000",
  60757=>"001001001",
  60758=>"000100110",
  60759=>"000000000",
  60760=>"000001101",
  60761=>"000000001",
  60762=>"111111110",
  60763=>"110100000",
  60764=>"001001000",
  60765=>"111111111",
  60766=>"111001000",
  60767=>"000000000",
  60768=>"111101111",
  60769=>"011000000",
  60770=>"001000100",
  60771=>"100000000",
  60772=>"000111111",
  60773=>"001000000",
  60774=>"001000001",
  60775=>"110110110",
  60776=>"000001001",
  60777=>"011000110",
  60778=>"101000000",
  60779=>"111011000",
  60780=>"000000001",
  60781=>"000010100",
  60782=>"000000000",
  60783=>"111110000",
  60784=>"001100000",
  60785=>"000010110",
  60786=>"111101000",
  60787=>"111111111",
  60788=>"110110110",
  60789=>"010010000",
  60790=>"000000001",
  60791=>"000011000",
  60792=>"100000010",
  60793=>"001000000",
  60794=>"111000011",
  60795=>"000000000",
  60796=>"101101110",
  60797=>"111110110",
  60798=>"000000000",
  60799=>"000111111",
  60800=>"110110001",
  60801=>"010110011",
  60802=>"111111111",
  60803=>"000000000",
  60804=>"100000001",
  60805=>"011000000",
  60806=>"100000000",
  60807=>"000000000",
  60808=>"000000000",
  60809=>"011111111",
  60810=>"000000001",
  60811=>"000000111",
  60812=>"111111111",
  60813=>"000010011",
  60814=>"000110000",
  60815=>"000000000",
  60816=>"000000000",
  60817=>"111111111",
  60818=>"111011111",
  60819=>"111111111",
  60820=>"100111011",
  60821=>"000000000",
  60822=>"100111111",
  60823=>"111111110",
  60824=>"011111000",
  60825=>"110011011",
  60826=>"000000000",
  60827=>"000110111",
  60828=>"101101111",
  60829=>"000000000",
  60830=>"011011010",
  60831=>"000110110",
  60832=>"000000000",
  60833=>"001011011",
  60834=>"011111111",
  60835=>"000000000",
  60836=>"101100110",
  60837=>"111111001",
  60838=>"000000001",
  60839=>"000111111",
  60840=>"000000001",
  60841=>"110110000",
  60842=>"000000000",
  60843=>"011011111",
  60844=>"000000000",
  60845=>"000101001",
  60846=>"011110100",
  60847=>"110111111",
  60848=>"011111101",
  60849=>"111111111",
  60850=>"001001011",
  60851=>"000000000",
  60852=>"110111100",
  60853=>"111111100",
  60854=>"110110000",
  60855=>"000000000",
  60856=>"101111100",
  60857=>"111111111",
  60858=>"000000000",
  60859=>"000001000",
  60860=>"110100110",
  60861=>"110111110",
  60862=>"011000000",
  60863=>"000011000",
  60864=>"111111001",
  60865=>"111111111",
  60866=>"111111111",
  60867=>"110100000",
  60868=>"001001001",
  60869=>"111100110",
  60870=>"111111110",
  60871=>"001001011",
  60872=>"001000100",
  60873=>"011110000",
  60874=>"111000000",
  60875=>"000010000",
  60876=>"111011010",
  60877=>"001001000",
  60878=>"111100000",
  60879=>"111111011",
  60880=>"111011111",
  60881=>"111111011",
  60882=>"000010001",
  60883=>"000000010",
  60884=>"100000000",
  60885=>"100000000",
  60886=>"010000000",
  60887=>"001000010",
  60888=>"000001001",
  60889=>"111111000",
  60890=>"000000000",
  60891=>"111111111",
  60892=>"111111111",
  60893=>"110000110",
  60894=>"000000000",
  60895=>"000000000",
  60896=>"000000000",
  60897=>"111001111",
  60898=>"000000000",
  60899=>"001100000",
  60900=>"111001000",
  60901=>"110111111",
  60902=>"001001101",
  60903=>"111111111",
  60904=>"001000011",
  60905=>"000000010",
  60906=>"000100111",
  60907=>"111100100",
  60908=>"101001101",
  60909=>"111111101",
  60910=>"111111110",
  60911=>"010110111",
  60912=>"111111111",
  60913=>"000001011",
  60914=>"111111011",
  60915=>"010011111",
  60916=>"000011010",
  60917=>"110000101",
  60918=>"000110100",
  60919=>"011011011",
  60920=>"000110000",
  60921=>"011000000",
  60922=>"110111111",
  60923=>"000000000",
  60924=>"000000000",
  60925=>"001011011",
  60926=>"100000000",
  60927=>"000000000",
  60928=>"010111111",
  60929=>"111111111",
  60930=>"111000111",
  60931=>"111111111",
  60932=>"000100111",
  60933=>"011011000",
  60934=>"000000111",
  60935=>"110111111",
  60936=>"001000111",
  60937=>"110111111",
  60938=>"111111110",
  60939=>"110111001",
  60940=>"000100101",
  60941=>"111111111",
  60942=>"010111110",
  60943=>"000000000",
  60944=>"010110110",
  60945=>"000000111",
  60946=>"000000010",
  60947=>"110111111",
  60948=>"000000000",
  60949=>"010101100",
  60950=>"111001000",
  60951=>"000111100",
  60952=>"111111100",
  60953=>"000000000",
  60954=>"001000011",
  60955=>"011011110",
  60956=>"111111111",
  60957=>"111110000",
  60958=>"000000110",
  60959=>"100111111",
  60960=>"000000111",
  60961=>"000111111",
  60962=>"111110111",
  60963=>"000111111",
  60964=>"010000000",
  60965=>"000101111",
  60966=>"000000101",
  60967=>"111001001",
  60968=>"111001000",
  60969=>"000001011",
  60970=>"001111111",
  60971=>"000111110",
  60972=>"000000001",
  60973=>"000000000",
  60974=>"000000000",
  60975=>"111111111",
  60976=>"111101110",
  60977=>"000000000",
  60978=>"000000000",
  60979=>"101111111",
  60980=>"111111111",
  60981=>"110110110",
  60982=>"000000111",
  60983=>"000111111",
  60984=>"011000000",
  60985=>"000000000",
  60986=>"111000000",
  60987=>"000100111",
  60988=>"111100100",
  60989=>"000000000",
  60990=>"000000000",
  60991=>"111111111",
  60992=>"000000101",
  60993=>"000100000",
  60994=>"000111111",
  60995=>"111101111",
  60996=>"000000000",
  60997=>"111111111",
  60998=>"111111111",
  60999=>"111110000",
  61000=>"110111110",
  61001=>"111101101",
  61002=>"000000000",
  61003=>"110000000",
  61004=>"111001000",
  61005=>"000000111",
  61006=>"000000000",
  61007=>"000000000",
  61008=>"000001111",
  61009=>"110100000",
  61010=>"000000000",
  61011=>"111111111",
  61012=>"000000111",
  61013=>"000000101",
  61014=>"101111101",
  61015=>"111111111",
  61016=>"000000000",
  61017=>"101000000",
  61018=>"000010110",
  61019=>"000000000",
  61020=>"000000000",
  61021=>"111000000",
  61022=>"100000000",
  61023=>"000000001",
  61024=>"000000111",
  61025=>"000000000",
  61026=>"110011101",
  61027=>"000000000",
  61028=>"111000000",
  61029=>"110000000",
  61030=>"111011100",
  61031=>"000000001",
  61032=>"000000000",
  61033=>"111010000",
  61034=>"000000000",
  61035=>"000000001",
  61036=>"100001001",
  61037=>"000011111",
  61038=>"000000000",
  61039=>"111100000",
  61040=>"111011111",
  61041=>"000111111",
  61042=>"111000000",
  61043=>"000111000",
  61044=>"000100000",
  61045=>"001011111",
  61046=>"000111100",
  61047=>"000000000",
  61048=>"010000000",
  61049=>"001001000",
  61050=>"011000000",
  61051=>"000000000",
  61052=>"000000110",
  61053=>"000000000",
  61054=>"000000000",
  61055=>"111011000",
  61056=>"111111111",
  61057=>"111000000",
  61058=>"000000100",
  61059=>"111100000",
  61060=>"000101101",
  61061=>"100000011",
  61062=>"111101111",
  61063=>"111111111",
  61064=>"111111000",
  61065=>"111111111",
  61066=>"100100000",
  61067=>"111111011",
  61068=>"000000000",
  61069=>"010111000",
  61070=>"111101110",
  61071=>"111111111",
  61072=>"111000000",
  61073=>"000000111",
  61074=>"000000000",
  61075=>"111111111",
  61076=>"111111111",
  61077=>"010000001",
  61078=>"000000000",
  61079=>"111101000",
  61080=>"000000000",
  61081=>"000000000",
  61082=>"111111111",
  61083=>"000000000",
  61084=>"111000000",
  61085=>"000000000",
  61086=>"000100111",
  61087=>"111111001",
  61088=>"001001000",
  61089=>"101001111",
  61090=>"001011000",
  61091=>"101111101",
  61092=>"011001001",
  61093=>"000000000",
  61094=>"111111111",
  61095=>"000110000",
  61096=>"000001111",
  61097=>"000000000",
  61098=>"000000000",
  61099=>"111111111",
  61100=>"100100000",
  61101=>"000101111",
  61102=>"000000000",
  61103=>"000011111",
  61104=>"000011000",
  61105=>"000000001",
  61106=>"110010111",
  61107=>"100100111",
  61108=>"111111111",
  61109=>"111001000",
  61110=>"010010000",
  61111=>"101111001",
  61112=>"111011011",
  61113=>"111111111",
  61114=>"100000000",
  61115=>"111000000",
  61116=>"001001000",
  61117=>"111111100",
  61118=>"000111000",
  61119=>"110111111",
  61120=>"100000000",
  61121=>"000000111",
  61122=>"111000000",
  61123=>"111111111",
  61124=>"111111111",
  61125=>"000001111",
  61126=>"000101111",
  61127=>"000000000",
  61128=>"111111111",
  61129=>"101111111",
  61130=>"000000001",
  61131=>"111110000",
  61132=>"111101100",
  61133=>"000101000",
  61134=>"000111111",
  61135=>"000001111",
  61136=>"110010101",
  61137=>"111111111",
  61138=>"111111001",
  61139=>"000001111",
  61140=>"000000000",
  61141=>"000001011",
  61142=>"001000000",
  61143=>"111011111",
  61144=>"000000111",
  61145=>"111110100",
  61146=>"111000000",
  61147=>"111001000",
  61148=>"001001001",
  61149=>"111000000",
  61150=>"111111111",
  61151=>"001000000",
  61152=>"000000000",
  61153=>"000000000",
  61154=>"111111111",
  61155=>"001001111",
  61156=>"101100000",
  61157=>"000000000",
  61158=>"000111111",
  61159=>"111111001",
  61160=>"001101111",
  61161=>"110111111",
  61162=>"111000000",
  61163=>"000111111",
  61164=>"000000000",
  61165=>"000000001",
  61166=>"111110000",
  61167=>"111000000",
  61168=>"000101111",
  61169=>"011111111",
  61170=>"111111110",
  61171=>"101111110",
  61172=>"000111000",
  61173=>"000000000",
  61174=>"000100110",
  61175=>"111111111",
  61176=>"100110111",
  61177=>"111111111",
  61178=>"001000000",
  61179=>"111111000",
  61180=>"001111111",
  61181=>"011001001",
  61182=>"111000001",
  61183=>"111111001",
  61184=>"000000000",
  61185=>"000001001",
  61186=>"011111111",
  61187=>"110000100",
  61188=>"111001000",
  61189=>"010001111",
  61190=>"111001000",
  61191=>"001011111",
  61192=>"000001111",
  61193=>"000000000",
  61194=>"000000000",
  61195=>"101111010",
  61196=>"110111101",
  61197=>"000000000",
  61198=>"100110111",
  61199=>"000000000",
  61200=>"011111111",
  61201=>"000100110",
  61202=>"111001001",
  61203=>"001000011",
  61204=>"000000111",
  61205=>"111111111",
  61206=>"000000110",
  61207=>"111111100",
  61208=>"000000000",
  61209=>"010111111",
  61210=>"000000000",
  61211=>"110010000",
  61212=>"011111011",
  61213=>"111010000",
  61214=>"000110111",
  61215=>"111111101",
  61216=>"011000100",
  61217=>"100000001",
  61218=>"000010110",
  61219=>"111111111",
  61220=>"000000000",
  61221=>"000110111",
  61222=>"111111111",
  61223=>"110110110",
  61224=>"000000111",
  61225=>"010011000",
  61226=>"000000000",
  61227=>"111111111",
  61228=>"000111111",
  61229=>"000000000",
  61230=>"011000111",
  61231=>"110011000",
  61232=>"110111111",
  61233=>"000000111",
  61234=>"111111111",
  61235=>"101000000",
  61236=>"000000000",
  61237=>"000100111",
  61238=>"000111111",
  61239=>"001001011",
  61240=>"000000000",
  61241=>"001101111",
  61242=>"101000000",
  61243=>"000000000",
  61244=>"111111111",
  61245=>"111111111",
  61246=>"101111111",
  61247=>"111111000",
  61248=>"111111111",
  61249=>"000000000",
  61250=>"110111110",
  61251=>"111001000",
  61252=>"000111110",
  61253=>"000000000",
  61254=>"111101111",
  61255=>"100011000",
  61256=>"000000000",
  61257=>"111111111",
  61258=>"110111000",
  61259=>"101100100",
  61260=>"010000101",
  61261=>"111001010",
  61262=>"101101111",
  61263=>"111111000",
  61264=>"000111111",
  61265=>"001000000",
  61266=>"111000111",
  61267=>"001001000",
  61268=>"111001000",
  61269=>"001001001",
  61270=>"001111111",
  61271=>"000000000",
  61272=>"100111111",
  61273=>"100000000",
  61274=>"000000000",
  61275=>"100111100",
  61276=>"011000000",
  61277=>"110110000",
  61278=>"000000101",
  61279=>"110111011",
  61280=>"000000010",
  61281=>"111111111",
  61282=>"000100111",
  61283=>"000000000",
  61284=>"111111000",
  61285=>"111000000",
  61286=>"111111111",
  61287=>"000000001",
  61288=>"001001001",
  61289=>"110110100",
  61290=>"111011000",
  61291=>"111111100",
  61292=>"000000011",
  61293=>"000110110",
  61294=>"111000000",
  61295=>"101111001",
  61296=>"111111111",
  61297=>"111111111",
  61298=>"011100111",
  61299=>"000000000",
  61300=>"000110100",
  61301=>"111111110",
  61302=>"101000000",
  61303=>"000111111",
  61304=>"000000000",
  61305=>"010001000",
  61306=>"111111111",
  61307=>"000100111",
  61308=>"000000000",
  61309=>"011000000",
  61310=>"000000001",
  61311=>"111001001",
  61312=>"001001001",
  61313=>"000000100",
  61314=>"111111111",
  61315=>"000000000",
  61316=>"000000000",
  61317=>"000111100",
  61318=>"000000000",
  61319=>"111111001",
  61320=>"000000000",
  61321=>"111111110",
  61322=>"110111111",
  61323=>"000010000",
  61324=>"111111111",
  61325=>"100110110",
  61326=>"100000000",
  61327=>"000000000",
  61328=>"000000100",
  61329=>"010010000",
  61330=>"111011001",
  61331=>"111111110",
  61332=>"111111000",
  61333=>"000000010",
  61334=>"000000001",
  61335=>"011011111",
  61336=>"111111111",
  61337=>"101111111",
  61338=>"110000000",
  61339=>"111110111",
  61340=>"001001111",
  61341=>"111001111",
  61342=>"001001000",
  61343=>"111111111",
  61344=>"000100100",
  61345=>"001001000",
  61346=>"111001000",
  61347=>"000000111",
  61348=>"000000000",
  61349=>"000111111",
  61350=>"111111111",
  61351=>"111111000",
  61352=>"111001001",
  61353=>"111000000",
  61354=>"111000110",
  61355=>"000000000",
  61356=>"000000001",
  61357=>"000000000",
  61358=>"000110111",
  61359=>"000111111",
  61360=>"110000000",
  61361=>"001011000",
  61362=>"110110111",
  61363=>"111001000",
  61364=>"111111111",
  61365=>"111111111",
  61366=>"110100000",
  61367=>"111000000",
  61368=>"111000000",
  61369=>"111111000",
  61370=>"000111100",
  61371=>"111000000",
  61372=>"010000000",
  61373=>"000000000",
  61374=>"000000000",
  61375=>"000110110",
  61376=>"001000111",
  61377=>"011000000",
  61378=>"111111111",
  61379=>"110111111",
  61380=>"101111111",
  61381=>"000000000",
  61382=>"111000001",
  61383=>"000000000",
  61384=>"000000000",
  61385=>"111111111",
  61386=>"000000001",
  61387=>"000000000",
  61388=>"111111011",
  61389=>"000000111",
  61390=>"101101101",
  61391=>"000010111",
  61392=>"111000000",
  61393=>"111111111",
  61394=>"110111011",
  61395=>"111111111",
  61396=>"111000001",
  61397=>"111101000",
  61398=>"111001011",
  61399=>"110011000",
  61400=>"000000001",
  61401=>"000000000",
  61402=>"111000001",
  61403=>"111000000",
  61404=>"100111111",
  61405=>"111011111",
  61406=>"111000111",
  61407=>"000001001",
  61408=>"111010000",
  61409=>"111000000",
  61410=>"110000000",
  61411=>"111110000",
  61412=>"101111111",
  61413=>"111100010",
  61414=>"000111011",
  61415=>"110111111",
  61416=>"111111111",
  61417=>"100000110",
  61418=>"000001000",
  61419=>"111000000",
  61420=>"111000010",
  61421=>"000100111",
  61422=>"111111111",
  61423=>"000111111",
  61424=>"001000000",
  61425=>"000000111",
  61426=>"111111111",
  61427=>"111000010",
  61428=>"000000111",
  61429=>"011100000",
  61430=>"111111000",
  61431=>"110000001",
  61432=>"000000000",
  61433=>"000011111",
  61434=>"000000000",
  61435=>"111000000",
  61436=>"000000000",
  61437=>"000000000",
  61438=>"111000000",
  61439=>"000000000",
  61440=>"000000100",
  61441=>"000010010",
  61442=>"000000111",
  61443=>"111001000",
  61444=>"000000000",
  61445=>"111010010",
  61446=>"100000000",
  61447=>"111111111",
  61448=>"111111111",
  61449=>"011000000",
  61450=>"000000101",
  61451=>"000110000",
  61452=>"000000000",
  61453=>"111001001",
  61454=>"000000001",
  61455=>"011011011",
  61456=>"000000000",
  61457=>"111000000",
  61458=>"011000011",
  61459=>"000000000",
  61460=>"001001111",
  61461=>"110010110",
  61462=>"110111111",
  61463=>"011001000",
  61464=>"111111111",
  61465=>"001001011",
  61466=>"111101001",
  61467=>"110111111",
  61468=>"111101111",
  61469=>"000000000",
  61470=>"110110000",
  61471=>"000000000",
  61472=>"000000000",
  61473=>"101100000",
  61474=>"001111111",
  61475=>"100100000",
  61476=>"000000000",
  61477=>"010000000",
  61478=>"010010011",
  61479=>"000000101",
  61480=>"111111111",
  61481=>"000000000",
  61482=>"000000001",
  61483=>"000000111",
  61484=>"010010110",
  61485=>"100111111",
  61486=>"111101111",
  61487=>"000000000",
  61488=>"111111111",
  61489=>"111111101",
  61490=>"111101101",
  61491=>"101100101",
  61492=>"011111011",
  61493=>"000000000",
  61494=>"000000000",
  61495=>"001011000",
  61496=>"111111101",
  61497=>"000000000",
  61498=>"000001001",
  61499=>"000000000",
  61500=>"111001010",
  61501=>"100100101",
  61502=>"000000000",
  61503=>"000000000",
  61504=>"000000100",
  61505=>"111111111",
  61506=>"110100111",
  61507=>"000000000",
  61508=>"111111011",
  61509=>"111111110",
  61510=>"000000000",
  61511=>"101101111",
  61512=>"011011011",
  61513=>"000000111",
  61514=>"000000000",
  61515=>"101111000",
  61516=>"000000000",
  61517=>"101000000",
  61518=>"000000110",
  61519=>"000000000",
  61520=>"000000000",
  61521=>"000000000",
  61522=>"000000001",
  61523=>"010010000",
  61524=>"000000011",
  61525=>"111111111",
  61526=>"101001100",
  61527=>"001111111",
  61528=>"101000000",
  61529=>"011000111",
  61530=>"101101000",
  61531=>"111111001",
  61532=>"111111111",
  61533=>"111111111",
  61534=>"111110101",
  61535=>"111111100",
  61536=>"000000000",
  61537=>"111111111",
  61538=>"111111000",
  61539=>"111010111",
  61540=>"111001000",
  61541=>"111110111",
  61542=>"111111111",
  61543=>"111101000",
  61544=>"111111111",
  61545=>"011011111",
  61546=>"010010000",
  61547=>"110100000",
  61548=>"010000000",
  61549=>"100100000",
  61550=>"001001011",
  61551=>"111000000",
  61552=>"111111111",
  61553=>"111111001",
  61554=>"001000001",
  61555=>"001000101",
  61556=>"111111111",
  61557=>"000100101",
  61558=>"011001111",
  61559=>"000000000",
  61560=>"000000000",
  61561=>"000000000",
  61562=>"100000000",
  61563=>"000000000",
  61564=>"000000010",
  61565=>"111111001",
  61566=>"000000000",
  61567=>"000000000",
  61568=>"000000000",
  61569=>"000000000",
  61570=>"000000010",
  61571=>"001100000",
  61572=>"000000001",
  61573=>"100000000",
  61574=>"000100110",
  61575=>"000000000",
  61576=>"110011111",
  61577=>"111111111",
  61578=>"111111011",
  61579=>"111011000",
  61580=>"111101000",
  61581=>"111111000",
  61582=>"111110110",
  61583=>"101001101",
  61584=>"111111111",
  61585=>"111111111",
  61586=>"000000000",
  61587=>"111000000",
  61588=>"000000000",
  61589=>"000000000",
  61590=>"000000011",
  61591=>"000100100",
  61592=>"001111010",
  61593=>"000100111",
  61594=>"111111000",
  61595=>"000000000",
  61596=>"000010111",
  61597=>"001000001",
  61598=>"000000000",
  61599=>"000000000",
  61600=>"000011000",
  61601=>"000000001",
  61602=>"100000000",
  61603=>"100111011",
  61604=>"001001001",
  61605=>"100000000",
  61606=>"110011000",
  61607=>"000001001",
  61608=>"000000100",
  61609=>"001111111",
  61610=>"000000000",
  61611=>"010000111",
  61612=>"111111011",
  61613=>"111111110",
  61614=>"000000100",
  61615=>"001011001",
  61616=>"000000000",
  61617=>"111111000",
  61618=>"111111111",
  61619=>"111111111",
  61620=>"111111111",
  61621=>"000000110",
  61622=>"001001000",
  61623=>"000000010",
  61624=>"101101000",
  61625=>"000100111",
  61626=>"101100101",
  61627=>"001001001",
  61628=>"000111111",
  61629=>"111101101",
  61630=>"000000000",
  61631=>"000000000",
  61632=>"000000110",
  61633=>"010111000",
  61634=>"000000000",
  61635=>"000000000",
  61636=>"111111111",
  61637=>"000000000",
  61638=>"111011110",
  61639=>"000000001",
  61640=>"110010000",
  61641=>"100000000",
  61642=>"111111001",
  61643=>"100000000",
  61644=>"111111000",
  61645=>"111111111",
  61646=>"000111111",
  61647=>"000000000",
  61648=>"000000000",
  61649=>"110000001",
  61650=>"010011000",
  61651=>"111111101",
  61652=>"000000011",
  61653=>"111111110",
  61654=>"111000000",
  61655=>"001000001",
  61656=>"100111110",
  61657=>"000000001",
  61658=>"000000000",
  61659=>"000000000",
  61660=>"111010000",
  61661=>"111001001",
  61662=>"111111111",
  61663=>"000000110",
  61664=>"000000000",
  61665=>"000010000",
  61666=>"000000000",
  61667=>"000000000",
  61668=>"100000000",
  61669=>"110110000",
  61670=>"110111011",
  61671=>"110000000",
  61672=>"110111111",
  61673=>"111111111",
  61674=>"000000000",
  61675=>"110010000",
  61676=>"000010011",
  61677=>"111111111",
  61678=>"000000000",
  61679=>"000000000",
  61680=>"010110011",
  61681=>"100100111",
  61682=>"111110101",
  61683=>"001001001",
  61684=>"000000000",
  61685=>"011111001",
  61686=>"000000000",
  61687=>"000000000",
  61688=>"100000000",
  61689=>"000000000",
  61690=>"111111111",
  61691=>"000000000",
  61692=>"110110000",
  61693=>"000000001",
  61694=>"011011100",
  61695=>"001000000",
  61696=>"011011000",
  61697=>"111111111",
  61698=>"100101111",
  61699=>"000000011",
  61700=>"000111111",
  61701=>"000000000",
  61702=>"000000000",
  61703=>"000000000",
  61704=>"100111111",
  61705=>"000000111",
  61706=>"000000000",
  61707=>"111111101",
  61708=>"001000000",
  61709=>"010111111",
  61710=>"100000000",
  61711=>"000000000",
  61712=>"000000000",
  61713=>"000000011",
  61714=>"111000000",
  61715=>"000001000",
  61716=>"010011011",
  61717=>"111000000",
  61718=>"110110111",
  61719=>"111111111",
  61720=>"111111111",
  61721=>"111111011",
  61722=>"111111011",
  61723=>"110110000",
  61724=>"001111111",
  61725=>"000000100",
  61726=>"000000000",
  61727=>"000000000",
  61728=>"100100001",
  61729=>"000010111",
  61730=>"000111111",
  61731=>"001000111",
  61732=>"001000100",
  61733=>"001111011",
  61734=>"000000000",
  61735=>"011111001",
  61736=>"000000110",
  61737=>"010011011",
  61738=>"000110110",
  61739=>"111111111",
  61740=>"110111000",
  61741=>"111100110",
  61742=>"100100111",
  61743=>"100110111",
  61744=>"000000000",
  61745=>"111111111",
  61746=>"010000000",
  61747=>"100111011",
  61748=>"101110000",
  61749=>"000001111",
  61750=>"000100111",
  61751=>"111111111",
  61752=>"000000000",
  61753=>"000000000",
  61754=>"111000000",
  61755=>"111111100",
  61756=>"011111111",
  61757=>"000000111",
  61758=>"011011011",
  61759=>"000000000",
  61760=>"000010010",
  61761=>"011001000",
  61762=>"000001000",
  61763=>"001000000",
  61764=>"000010001",
  61765=>"000000000",
  61766=>"000000010",
  61767=>"111011001",
  61768=>"111010000",
  61769=>"000000111",
  61770=>"111111111",
  61771=>"111100111",
  61772=>"000000000",
  61773=>"000011111",
  61774=>"010000000",
  61775=>"110011000",
  61776=>"111001000",
  61777=>"000000000",
  61778=>"000000000",
  61779=>"000000000",
  61780=>"011000000",
  61781=>"011001001",
  61782=>"010010000",
  61783=>"000000000",
  61784=>"100100100",
  61785=>"111111111",
  61786=>"000010111",
  61787=>"001000100",
  61788=>"000000000",
  61789=>"010000000",
  61790=>"011111111",
  61791=>"111111111",
  61792=>"111111010",
  61793=>"111111110",
  61794=>"100111111",
  61795=>"001101111",
  61796=>"000000011",
  61797=>"000110000",
  61798=>"111110111",
  61799=>"000001111",
  61800=>"110000110",
  61801=>"000000000",
  61802=>"110000111",
  61803=>"011111111",
  61804=>"000010100",
  61805=>"111101111",
  61806=>"111111111",
  61807=>"001001111",
  61808=>"111111111",
  61809=>"110010000",
  61810=>"000000000",
  61811=>"111111111",
  61812=>"000000000",
  61813=>"111111111",
  61814=>"000000111",
  61815=>"010010000",
  61816=>"111001111",
  61817=>"111111111",
  61818=>"111111110",
  61819=>"111110111",
  61820=>"111111011",
  61821=>"000100000",
  61822=>"101001011",
  61823=>"000000000",
  61824=>"000000110",
  61825=>"000110111",
  61826=>"111000000",
  61827=>"000000000",
  61828=>"111111011",
  61829=>"000110111",
  61830=>"111100110",
  61831=>"000000100",
  61832=>"111110111",
  61833=>"000000000",
  61834=>"111000000",
  61835=>"111000000",
  61836=>"111111111",
  61837=>"100011000",
  61838=>"000000111",
  61839=>"000000000",
  61840=>"000000000",
  61841=>"000000000",
  61842=>"111101000",
  61843=>"011111011",
  61844=>"100000000",
  61845=>"000010000",
  61846=>"111111111",
  61847=>"000101111",
  61848=>"000000100",
  61849=>"001111111",
  61850=>"111111111",
  61851=>"110110110",
  61852=>"000010110",
  61853=>"111110100",
  61854=>"000110100",
  61855=>"000000010",
  61856=>"100100110",
  61857=>"111111110",
  61858=>"111111101",
  61859=>"000000111",
  61860=>"111101001",
  61861=>"000000000",
  61862=>"100100111",
  61863=>"000000000",
  61864=>"000000000",
  61865=>"000000010",
  61866=>"111010010",
  61867=>"000010111",
  61868=>"000000000",
  61869=>"111001000",
  61870=>"111001111",
  61871=>"101100000",
  61872=>"000000111",
  61873=>"000000000",
  61874=>"001000001",
  61875=>"000000011",
  61876=>"000000000",
  61877=>"110100101",
  61878=>"001001001",
  61879=>"001000000",
  61880=>"000000000",
  61881=>"011001000",
  61882=>"111111010",
  61883=>"111111011",
  61884=>"000000000",
  61885=>"111011111",
  61886=>"000000010",
  61887=>"011111111",
  61888=>"000000011",
  61889=>"000000000",
  61890=>"011111011",
  61891=>"011011011",
  61892=>"000001001",
  61893=>"101000001",
  61894=>"000001001",
  61895=>"111111111",
  61896=>"000000000",
  61897=>"000000110",
  61898=>"000000001",
  61899=>"111111111",
  61900=>"000011000",
  61901=>"000000000",
  61902=>"000000101",
  61903=>"111111111",
  61904=>"000110110",
  61905=>"110110100",
  61906=>"000000000",
  61907=>"111111000",
  61908=>"000000000",
  61909=>"001000000",
  61910=>"000000000",
  61911=>"000000000",
  61912=>"000000100",
  61913=>"111111000",
  61914=>"001011111",
  61915=>"111111101",
  61916=>"110111111",
  61917=>"101111111",
  61918=>"100101111",
  61919=>"001001001",
  61920=>"111111111",
  61921=>"100110111",
  61922=>"000000000",
  61923=>"000000000",
  61924=>"000010110",
  61925=>"111111000",
  61926=>"111011011",
  61927=>"101101000",
  61928=>"000000000",
  61929=>"111111111",
  61930=>"000000000",
  61931=>"000000001",
  61932=>"111111111",
  61933=>"111111001",
  61934=>"011111111",
  61935=>"111111111",
  61936=>"111100100",
  61937=>"000000000",
  61938=>"111111111",
  61939=>"000010000",
  61940=>"001001110",
  61941=>"111111100",
  61942=>"111110100",
  61943=>"001100000",
  61944=>"000000011",
  61945=>"111111111",
  61946=>"111111001",
  61947=>"000000000",
  61948=>"011001000",
  61949=>"111100101",
  61950=>"000000000",
  61951=>"111001111",
  61952=>"010010100",
  61953=>"110110010",
  61954=>"001000000",
  61955=>"100111001",
  61956=>"000000001",
  61957=>"111111110",
  61958=>"100000000",
  61959=>"000000000",
  61960=>"000000000",
  61961=>"100111111",
  61962=>"000000000",
  61963=>"000000000",
  61964=>"000001011",
  61965=>"111000000",
  61966=>"000000100",
  61967=>"001100111",
  61968=>"000000000",
  61969=>"100100100",
  61970=>"000000000",
  61971=>"001000110",
  61972=>"111111111",
  61973=>"111111111",
  61974=>"110110111",
  61975=>"000000000",
  61976=>"010010111",
  61977=>"101111011",
  61978=>"111111111",
  61979=>"111000000",
  61980=>"100000000",
  61981=>"000000001",
  61982=>"110100100",
  61983=>"111111110",
  61984=>"000001001",
  61985=>"110000000",
  61986=>"011111111",
  61987=>"000100110",
  61988=>"000100000",
  61989=>"111111011",
  61990=>"000000000",
  61991=>"000000000",
  61992=>"110111001",
  61993=>"001001111",
  61994=>"111111111",
  61995=>"100000000",
  61996=>"001001100",
  61997=>"000000001",
  61998=>"110111111",
  61999=>"111111111",
  62000=>"100011001",
  62001=>"001001011",
  62002=>"010010011",
  62003=>"110000000",
  62004=>"000000000",
  62005=>"000011011",
  62006=>"101000001",
  62007=>"000110101",
  62008=>"000000101",
  62009=>"101001111",
  62010=>"111111111",
  62011=>"000000000",
  62012=>"111100101",
  62013=>"100000100",
  62014=>"111111111",
  62015=>"100000000",
  62016=>"000000100",
  62017=>"000011010",
  62018=>"000000000",
  62019=>"111111111",
  62020=>"010010011",
  62021=>"110110111",
  62022=>"001000000",
  62023=>"001000000",
  62024=>"000110111",
  62025=>"111111101",
  62026=>"000000000",
  62027=>"000110111",
  62028=>"110101111",
  62029=>"100100000",
  62030=>"111010011",
  62031=>"100111111",
  62032=>"100000100",
  62033=>"001000011",
  62034=>"111111111",
  62035=>"000000011",
  62036=>"000000000",
  62037=>"101000000",
  62038=>"011011000",
  62039=>"000000000",
  62040=>"000000000",
  62041=>"000000100",
  62042=>"111111100",
  62043=>"110011011",
  62044=>"111101000",
  62045=>"000101000",
  62046=>"110000110",
  62047=>"111110100",
  62048=>"000101100",
  62049=>"000000000",
  62050=>"000011111",
  62051=>"011000011",
  62052=>"000000001",
  62053=>"000111111",
  62054=>"011000001",
  62055=>"000000000",
  62056=>"010111111",
  62057=>"111111111",
  62058=>"011111111",
  62059=>"000000000",
  62060=>"110110011",
  62061=>"000000000",
  62062=>"000000000",
  62063=>"111011111",
  62064=>"000110110",
  62065=>"100000000",
  62066=>"001000111",
  62067=>"011000000",
  62068=>"111111111",
  62069=>"111111001",
  62070=>"000000111",
  62071=>"000000000",
  62072=>"000000000",
  62073=>"111111000",
  62074=>"111001000",
  62075=>"111000000",
  62076=>"000011111",
  62077=>"111111001",
  62078=>"111111111",
  62079=>"000000000",
  62080=>"000000000",
  62081=>"001000000",
  62082=>"111111111",
  62083=>"111000000",
  62084=>"000101111",
  62085=>"001001111",
  62086=>"111111111",
  62087=>"100000000",
  62088=>"111111001",
  62089=>"000000001",
  62090=>"111111111",
  62091=>"001101000",
  62092=>"000000000",
  62093=>"000000000",
  62094=>"101000110",
  62095=>"000111010",
  62096=>"000000000",
  62097=>"111111000",
  62098=>"000000000",
  62099=>"111111100",
  62100=>"101111111",
  62101=>"000100111",
  62102=>"011110000",
  62103=>"001000000",
  62104=>"001000000",
  62105=>"111111111",
  62106=>"111111100",
  62107=>"000000000",
  62108=>"001001111",
  62109=>"110110100",
  62110=>"000000000",
  62111=>"000111111",
  62112=>"111111111",
  62113=>"000000000",
  62114=>"000000001",
  62115=>"101111111",
  62116=>"100011011",
  62117=>"001000000",
  62118=>"001000000",
  62119=>"110111111",
  62120=>"111111111",
  62121=>"000100111",
  62122=>"111111000",
  62123=>"111111111",
  62124=>"111111111",
  62125=>"110111111",
  62126=>"001011111",
  62127=>"001001101",
  62128=>"000111111",
  62129=>"110110110",
  62130=>"000101000",
  62131=>"011000000",
  62132=>"000000000",
  62133=>"100111111",
  62134=>"100111111",
  62135=>"001101001",
  62136=>"100110111",
  62137=>"000000000",
  62138=>"110111001",
  62139=>"101001001",
  62140=>"011011011",
  62141=>"000101001",
  62142=>"111111011",
  62143=>"000111111",
  62144=>"011111111",
  62145=>"101000001",
  62146=>"111111100",
  62147=>"011111000",
  62148=>"011011111",
  62149=>"111001011",
  62150=>"000001111",
  62151=>"000000111",
  62152=>"000000111",
  62153=>"111000101",
  62154=>"111001011",
  62155=>"000100111",
  62156=>"000011111",
  62157=>"000111111",
  62158=>"000000000",
  62159=>"100000000",
  62160=>"111110101",
  62161=>"001111111",
  62162=>"011001011",
  62163=>"000000000",
  62164=>"000000011",
  62165=>"000000001",
  62166=>"000000010",
  62167=>"010010001",
  62168=>"111111111",
  62169=>"011011001",
  62170=>"111000000",
  62171=>"001011111",
  62172=>"000000001",
  62173=>"110111111",
  62174=>"111011001",
  62175=>"111101101",
  62176=>"000000000",
  62177=>"000000011",
  62178=>"111111111",
  62179=>"111101100",
  62180=>"111001001",
  62181=>"000000110",
  62182=>"101000000",
  62183=>"001111111",
  62184=>"000000000",
  62185=>"111111111",
  62186=>"000100101",
  62187=>"001000001",
  62188=>"111111111",
  62189=>"111111100",
  62190=>"100000111",
  62191=>"111110000",
  62192=>"111011010",
  62193=>"000000000",
  62194=>"010111111",
  62195=>"001001001",
  62196=>"000000000",
  62197=>"001001000",
  62198=>"100001001",
  62199=>"011111011",
  62200=>"000000000",
  62201=>"000100111",
  62202=>"111111011",
  62203=>"000111111",
  62204=>"110111001",
  62205=>"001111001",
  62206=>"100000000",
  62207=>"111111111",
  62208=>"000001001",
  62209=>"110110110",
  62210=>"101101000",
  62211=>"111101111",
  62212=>"000000000",
  62213=>"000100111",
  62214=>"111110111",
  62215=>"100110110",
  62216=>"100000100",
  62217=>"000000000",
  62218=>"001001001",
  62219=>"000000001",
  62220=>"000000000",
  62221=>"000000000",
  62222=>"000000000",
  62223=>"000000001",
  62224=>"000001000",
  62225=>"101101001",
  62226=>"000000000",
  62227=>"000111111",
  62228=>"001001000",
  62229=>"101000000",
  62230=>"000000100",
  62231=>"111101011",
  62232=>"111001001",
  62233=>"000000000",
  62234=>"000000000",
  62235=>"101001111",
  62236=>"010011000",
  62237=>"000000000",
  62238=>"010110110",
  62239=>"111000000",
  62240=>"000010110",
  62241=>"110111111",
  62242=>"000000001",
  62243=>"000000000",
  62244=>"100110110",
  62245=>"111111111",
  62246=>"111111111",
  62247=>"111000111",
  62248=>"000000010",
  62249=>"000001101",
  62250=>"000000000",
  62251=>"000000000",
  62252=>"111010011",
  62253=>"101110111",
  62254=>"111000000",
  62255=>"001000000",
  62256=>"000000000",
  62257=>"100000001",
  62258=>"000000000",
  62259=>"000111011",
  62260=>"111111111",
  62261=>"111111111",
  62262=>"100111000",
  62263=>"111111110",
  62264=>"001011000",
  62265=>"000000100",
  62266=>"100110111",
  62267=>"111110000",
  62268=>"100111111",
  62269=>"001001111",
  62270=>"110110100",
  62271=>"110010000",
  62272=>"000000000",
  62273=>"111000000",
  62274=>"000001011",
  62275=>"010010010",
  62276=>"001000000",
  62277=>"001001001",
  62278=>"111111111",
  62279=>"000000100",
  62280=>"000000000",
  62281=>"111111000",
  62282=>"100000001",
  62283=>"110110100",
  62284=>"111111111",
  62285=>"011011111",
  62286=>"101100100",
  62287=>"000011011",
  62288=>"111111111",
  62289=>"000100110",
  62290=>"111111111",
  62291=>"100000000",
  62292=>"000100101",
  62293=>"011000011",
  62294=>"111111111",
  62295=>"111000101",
  62296=>"111111111",
  62297=>"011011001",
  62298=>"011000101",
  62299=>"111000000",
  62300=>"011001011",
  62301=>"111111111",
  62302=>"000000001",
  62303=>"011011111",
  62304=>"011011001",
  62305=>"111111101",
  62306=>"100000000",
  62307=>"001000000",
  62308=>"000001011",
  62309=>"000000001",
  62310=>"000000000",
  62311=>"111111111",
  62312=>"111111101",
  62313=>"000000000",
  62314=>"101110110",
  62315=>"110110000",
  62316=>"100101111",
  62317=>"110110000",
  62318=>"000000000",
  62319=>"111111111",
  62320=>"100000000",
  62321=>"000000100",
  62322=>"000000000",
  62323=>"100100100",
  62324=>"111111111",
  62325=>"110111111",
  62326=>"111000110",
  62327=>"100000010",
  62328=>"000000111",
  62329=>"111111111",
  62330=>"100100111",
  62331=>"100001001",
  62332=>"000000000",
  62333=>"111111111",
  62334=>"111010010",
  62335=>"000000010",
  62336=>"100001001",
  62337=>"000000000",
  62338=>"011110110",
  62339=>"111111111",
  62340=>"000000111",
  62341=>"010011011",
  62342=>"000110111",
  62343=>"000011111",
  62344=>"111111111",
  62345=>"001011111",
  62346=>"001001000",
  62347=>"001001000",
  62348=>"111111111",
  62349=>"000000101",
  62350=>"000000000",
  62351=>"111111000",
  62352=>"000000000",
  62353=>"000001000",
  62354=>"010011111",
  62355=>"110101001",
  62356=>"001111011",
  62357=>"000111111",
  62358=>"000000000",
  62359=>"010011011",
  62360=>"100001000",
  62361=>"111110110",
  62362=>"111111111",
  62363=>"111111111",
  62364=>"000000000",
  62365=>"000100100",
  62366=>"100001001",
  62367=>"011111000",
  62368=>"001001111",
  62369=>"101100111",
  62370=>"001011000",
  62371=>"000000000",
  62372=>"000000001",
  62373=>"000000111",
  62374=>"111111101",
  62375=>"111000000",
  62376=>"000001111",
  62377=>"110110000",
  62378=>"001001001",
  62379=>"000011011",
  62380=>"111111111",
  62381=>"000000000",
  62382=>"100000100",
  62383=>"111111111",
  62384=>"000000111",
  62385=>"000000111",
  62386=>"110101111",
  62387=>"111101001",
  62388=>"000101111",
  62389=>"000000000",
  62390=>"111111111",
  62391=>"000000011",
  62392=>"000111011",
  62393=>"000111111",
  62394=>"111111001",
  62395=>"111000000",
  62396=>"001001001",
  62397=>"000000010",
  62398=>"000000000",
  62399=>"001101101",
  62400=>"111111111",
  62401=>"110100100",
  62402=>"111111011",
  62403=>"111111100",
  62404=>"000000000",
  62405=>"011001001",
  62406=>"100110111",
  62407=>"011111111",
  62408=>"101101111",
  62409=>"100111111",
  62410=>"001000000",
  62411=>"101001011",
  62412=>"001001000",
  62413=>"110010000",
  62414=>"111111010",
  62415=>"111111111",
  62416=>"000000001",
  62417=>"000001000",
  62418=>"000101001",
  62419=>"011001100",
  62420=>"111110110",
  62421=>"111000110",
  62422=>"000000001",
  62423=>"100111111",
  62424=>"001000000",
  62425=>"111110100",
  62426=>"000000111",
  62427=>"001001000",
  62428=>"001000000",
  62429=>"101110000",
  62430=>"000000100",
  62431=>"101001011",
  62432=>"010111111",
  62433=>"110111111",
  62434=>"111100111",
  62435=>"000110111",
  62436=>"000000111",
  62437=>"001001001",
  62438=>"000000000",
  62439=>"111111111",
  62440=>"111111111",
  62441=>"111111000",
  62442=>"100000100",
  62443=>"010110111",
  62444=>"000000110",
  62445=>"111111000",
  62446=>"000000100",
  62447=>"111111011",
  62448=>"110111111",
  62449=>"000111111",
  62450=>"000000000",
  62451=>"000000000",
  62452=>"101000000",
  62453=>"001111111",
  62454=>"111111111",
  62455=>"101111111",
  62456=>"011001001",
  62457=>"000000000",
  62458=>"000000100",
  62459=>"011000000",
  62460=>"000000000",
  62461=>"111011011",
  62462=>"001001011",
  62463=>"000000000",
  62464=>"010010011",
  62465=>"000000010",
  62466=>"101111111",
  62467=>"011111011",
  62468=>"001011001",
  62469=>"110110000",
  62470=>"000000000",
  62471=>"111111111",
  62472=>"000000000",
  62473=>"111000000",
  62474=>"110111111",
  62475=>"111110111",
  62476=>"100101011",
  62477=>"001000000",
  62478=>"000000000",
  62479=>"111111111",
  62480=>"000000000",
  62481=>"111111111",
  62482=>"011111110",
  62483=>"001000101",
  62484=>"010010010",
  62485=>"101101000",
  62486=>"000000001",
  62487=>"011001011",
  62488=>"000010000",
  62489=>"001001000",
  62490=>"000000000",
  62491=>"000000000",
  62492=>"000000000",
  62493=>"000000001",
  62494=>"000011110",
  62495=>"011111111",
  62496=>"110000000",
  62497=>"111111111",
  62498=>"001000111",
  62499=>"111000000",
  62500=>"100110000",
  62501=>"101000000",
  62502=>"010111111",
  62503=>"011101000",
  62504=>"011011011",
  62505=>"000000000",
  62506=>"111111111",
  62507=>"111111111",
  62508=>"111111101",
  62509=>"111111001",
  62510=>"001111110",
  62511=>"000010010",
  62512=>"001011110",
  62513=>"000000000",
  62514=>"010000001",
  62515=>"011010000",
  62516=>"110100110",
  62517=>"011011011",
  62518=>"110111110",
  62519=>"000110110",
  62520=>"000000000",
  62521=>"000001111",
  62522=>"000000000",
  62523=>"101100100",
  62524=>"000000000",
  62525=>"111001100",
  62526=>"110110111",
  62527=>"111000100",
  62528=>"100101111",
  62529=>"101000000",
  62530=>"000000000",
  62531=>"010000000",
  62532=>"000000000",
  62533=>"110000001",
  62534=>"000000000",
  62535=>"000000100",
  62536=>"000011011",
  62537=>"000001101",
  62538=>"111111111",
  62539=>"000001000",
  62540=>"111111111",
  62541=>"000101111",
  62542=>"000000000",
  62543=>"000000110",
  62544=>"111111011",
  62545=>"000000110",
  62546=>"100000000",
  62547=>"000100101",
  62548=>"000000000",
  62549=>"011001001",
  62550=>"000100000",
  62551=>"000000101",
  62552=>"000000000",
  62553=>"111111111",
  62554=>"111111011",
  62555=>"011011111",
  62556=>"111111000",
  62557=>"111110111",
  62558=>"111001011",
  62559=>"111111101",
  62560=>"000000000",
  62561=>"000000000",
  62562=>"000000101",
  62563=>"111111110",
  62564=>"101001000",
  62565=>"111111111",
  62566=>"000000000",
  62567=>"000000000",
  62568=>"000000000",
  62569=>"100100000",
  62570=>"011111111",
  62571=>"101101111",
  62572=>"000000000",
  62573=>"101000000",
  62574=>"110000000",
  62575=>"111000000",
  62576=>"000000011",
  62577=>"000100111",
  62578=>"111000000",
  62579=>"000000000",
  62580=>"111000111",
  62581=>"110111111",
  62582=>"111101110",
  62583=>"001000111",
  62584=>"011111101",
  62585=>"111111111",
  62586=>"000000000",
  62587=>"010000000",
  62588=>"101000001",
  62589=>"000000000",
  62590=>"000000000",
  62591=>"000000000",
  62592=>"001001000",
  62593=>"011111111",
  62594=>"000000000",
  62595=>"110110110",
  62596=>"111111111",
  62597=>"111101111",
  62598=>"000000000",
  62599=>"000000000",
  62600=>"111111011",
  62601=>"100000000",
  62602=>"101111000",
  62603=>"000000000",
  62604=>"111111111",
  62605=>"111111100",
  62606=>"111111001",
  62607=>"111000001",
  62608=>"111111011",
  62609=>"111111110",
  62610=>"000000111",
  62611=>"100100000",
  62612=>"010111011",
  62613=>"000101000",
  62614=>"000100101",
  62615=>"000000000",
  62616=>"011011000",
  62617=>"000010111",
  62618=>"000000000",
  62619=>"000000000",
  62620=>"000000110",
  62621=>"001000000",
  62622=>"111111111",
  62623=>"100000000",
  62624=>"111111000",
  62625=>"001000000",
  62626=>"000000000",
  62627=>"000000000",
  62628=>"000000000",
  62629=>"111111111",
  62630=>"010111010",
  62631=>"111110000",
  62632=>"011000111",
  62633=>"011111111",
  62634=>"111111111",
  62635=>"000000000",
  62636=>"000000000",
  62637=>"111110110",
  62638=>"101001101",
  62639=>"000010010",
  62640=>"010111000",
  62641=>"111110000",
  62642=>"110111111",
  62643=>"111011000",
  62644=>"000001110",
  62645=>"000000110",
  62646=>"000000111",
  62647=>"111101101",
  62648=>"000000001",
  62649=>"000000000",
  62650=>"000000000",
  62651=>"010000010",
  62652=>"101000001",
  62653=>"011000000",
  62654=>"000000000",
  62655=>"000000111",
  62656=>"100000100",
  62657=>"000111111",
  62658=>"110100101",
  62659=>"001001000",
  62660=>"100111111",
  62661=>"110111111",
  62662=>"000000000",
  62663=>"110000000",
  62664=>"111111000",
  62665=>"000000000",
  62666=>"000000000",
  62667=>"111111111",
  62668=>"000000001",
  62669=>"111111111",
  62670=>"111111001",
  62671=>"000000000",
  62672=>"111111111",
  62673=>"001011011",
  62674=>"000000000",
  62675=>"000000000",
  62676=>"000000000",
  62677=>"100000001",
  62678=>"111001000",
  62679=>"111110110",
  62680=>"110110111",
  62681=>"001001111",
  62682=>"000011000",
  62683=>"001000000",
  62684=>"111111111",
  62685=>"000000000",
  62686=>"111111111",
  62687=>"000000100",
  62688=>"111111111",
  62689=>"000000101",
  62690=>"111111111",
  62691=>"111101101",
  62692=>"000000111",
  62693=>"100110110",
  62694=>"000000000",
  62695=>"000111011",
  62696=>"001000000",
  62697=>"011001110",
  62698=>"001000000",
  62699=>"000000000",
  62700=>"011000100",
  62701=>"000000001",
  62702=>"000011110",
  62703=>"000001111",
  62704=>"111101001",
  62705=>"000110110",
  62706=>"111111101",
  62707=>"000000000",
  62708=>"011011000",
  62709=>"100100100",
  62710=>"000000000",
  62711=>"000000000",
  62712=>"000000001",
  62713=>"111110110",
  62714=>"000000000",
  62715=>"000000000",
  62716=>"110110110",
  62717=>"000000111",
  62718=>"111011011",
  62719=>"111111111",
  62720=>"000000000",
  62721=>"111000000",
  62722=>"000000000",
  62723=>"000111111",
  62724=>"111011000",
  62725=>"001000100",
  62726=>"111111111",
  62727=>"000100111",
  62728=>"000100000",
  62729=>"111111111",
  62730=>"111000000",
  62731=>"100100000",
  62732=>"001111111",
  62733=>"100110111",
  62734=>"001011110",
  62735=>"000100110",
  62736=>"000011111",
  62737=>"000000000",
  62738=>"101101111",
  62739=>"001011000",
  62740=>"000000000",
  62741=>"111111001",
  62742=>"011000000",
  62743=>"111001000",
  62744=>"111111111",
  62745=>"000000000",
  62746=>"000110111",
  62747=>"001000000",
  62748=>"000000100",
  62749=>"001000001",
  62750=>"001111111",
  62751=>"000111111",
  62752=>"011011011",
  62753=>"001011000",
  62754=>"000000000",
  62755=>"011011111",
  62756=>"111111111",
  62757=>"000000000",
  62758=>"000000000",
  62759=>"000000111",
  62760=>"001111011",
  62761=>"100000000",
  62762=>"000100110",
  62763=>"000111111",
  62764=>"000000001",
  62765=>"111000101",
  62766=>"000000111",
  62767=>"111111011",
  62768=>"000000011",
  62769=>"010000000",
  62770=>"111111011",
  62771=>"111111111",
  62772=>"111011011",
  62773=>"000000000",
  62774=>"000100100",
  62775=>"000000000",
  62776=>"000000000",
  62777=>"111101101",
  62778=>"000000111",
  62779=>"000011111",
  62780=>"111111001",
  62781=>"000111111",
  62782=>"000000010",
  62783=>"111000001",
  62784=>"000000010",
  62785=>"111111111",
  62786=>"111111110",
  62787=>"000000000",
  62788=>"111000001",
  62789=>"011001001",
  62790=>"111000100",
  62791=>"000000000",
  62792=>"111111111",
  62793=>"000000011",
  62794=>"001000111",
  62795=>"010110111",
  62796=>"000011000",
  62797=>"000101111",
  62798=>"000011111",
  62799=>"111000000",
  62800=>"100000000",
  62801=>"000010101",
  62802=>"000000111",
  62803=>"111100111",
  62804=>"000000111",
  62805=>"000011000",
  62806=>"011010011",
  62807=>"111111111",
  62808=>"000000000",
  62809=>"111111111",
  62810=>"011010000",
  62811=>"111111100",
  62812=>"000000000",
  62813=>"000000000",
  62814=>"001000010",
  62815=>"111111111",
  62816=>"010111111",
  62817=>"111111010",
  62818=>"100001001",
  62819=>"000000000",
  62820=>"000000000",
  62821=>"000000111",
  62822=>"000000010",
  62823=>"110011011",
  62824=>"110111111",
  62825=>"111001000",
  62826=>"000000000",
  62827=>"000000001",
  62828=>"100110000",
  62829=>"000011010",
  62830=>"111111100",
  62831=>"000000110",
  62832=>"111110111",
  62833=>"000010000",
  62834=>"000010000",
  62835=>"000100110",
  62836=>"000000000",
  62837=>"000100101",
  62838=>"011111000",
  62839=>"111111111",
  62840=>"000001111",
  62841=>"111111111",
  62842=>"100000000",
  62843=>"000010000",
  62844=>"000000000",
  62845=>"111111110",
  62846=>"011111000",
  62847=>"001000000",
  62848=>"011111111",
  62849=>"111111111",
  62850=>"011110110",
  62851=>"111111111",
  62852=>"110000001",
  62853=>"001101000",
  62854=>"111111111",
  62855=>"000000000",
  62856=>"000000000",
  62857=>"111011111",
  62858=>"110111111",
  62859=>"001000000",
  62860=>"101001000",
  62861=>"001001111",
  62862=>"001000000",
  62863=>"100100000",
  62864=>"001011011",
  62865=>"111111111",
  62866=>"011011000",
  62867=>"111111000",
  62868=>"111101000",
  62869=>"000000001",
  62870=>"111111111",
  62871=>"010110110",
  62872=>"000110110",
  62873=>"010000011",
  62874=>"111110000",
  62875=>"000000001",
  62876=>"110000000",
  62877=>"000000110",
  62878=>"000000000",
  62879=>"000000000",
  62880=>"001101111",
  62881=>"011011011",
  62882=>"110111111",
  62883=>"111111111",
  62884=>"111001001",
  62885=>"111111111",
  62886=>"010010000",
  62887=>"110101111",
  62888=>"001110110",
  62889=>"110111111",
  62890=>"000000000",
  62891=>"000000000",
  62892=>"000000001",
  62893=>"000000011",
  62894=>"111000001",
  62895=>"111111001",
  62896=>"000000111",
  62897=>"000000000",
  62898=>"111001001",
  62899=>"111111111",
  62900=>"000000000",
  62901=>"111000000",
  62902=>"111000000",
  62903=>"111111001",
  62904=>"000010000",
  62905=>"000000111",
  62906=>"000000100",
  62907=>"011100100",
  62908=>"000100100",
  62909=>"111001001",
  62910=>"011000011",
  62911=>"111111111",
  62912=>"111100000",
  62913=>"000000000",
  62914=>"000011000",
  62915=>"000000011",
  62916=>"111101101",
  62917=>"100000001",
  62918=>"110110111",
  62919=>"111001000",
  62920=>"000000000",
  62921=>"000000000",
  62922=>"000000000",
  62923=>"110111111",
  62924=>"000000000",
  62925=>"110110100",
  62926=>"000000000",
  62927=>"001111000",
  62928=>"011000000",
  62929=>"111111111",
  62930=>"111111110",
  62931=>"111111011",
  62932=>"000000110",
  62933=>"000001111",
  62934=>"000000101",
  62935=>"101001111",
  62936=>"111111110",
  62937=>"001001111",
  62938=>"000000000",
  62939=>"000000001",
  62940=>"000101101",
  62941=>"000000111",
  62942=>"100000111",
  62943=>"001001001",
  62944=>"000000000",
  62945=>"111110110",
  62946=>"000000000",
  62947=>"111110111",
  62948=>"000111111",
  62949=>"111110100",
  62950=>"111111110",
  62951=>"000000111",
  62952=>"001000000",
  62953=>"111111111",
  62954=>"001000000",
  62955=>"111111000",
  62956=>"101000000",
  62957=>"111111011",
  62958=>"000111111",
  62959=>"000010111",
  62960=>"000000000",
  62961=>"000000000",
  62962=>"000000000",
  62963=>"110111110",
  62964=>"100000000",
  62965=>"000010011",
  62966=>"111011111",
  62967=>"011111110",
  62968=>"000000000",
  62969=>"100100100",
  62970=>"000000000",
  62971=>"000111100",
  62972=>"000111001",
  62973=>"111111111",
  62974=>"000011011",
  62975=>"100111110",
  62976=>"000000000",
  62977=>"101000001",
  62978=>"001000001",
  62979=>"111111111",
  62980=>"110110110",
  62981=>"000000000",
  62982=>"001001111",
  62983=>"110111111",
  62984=>"111111110",
  62985=>"011011111",
  62986=>"101000111",
  62987=>"000000001",
  62988=>"000000000",
  62989=>"000000110",
  62990=>"011011000",
  62991=>"001111000",
  62992=>"010001001",
  62993=>"000000001",
  62994=>"000000000",
  62995=>"000110011",
  62996=>"000111000",
  62997=>"011000110",
  62998=>"111110110",
  62999=>"000110110",
  63000=>"000000000",
  63001=>"111101111",
  63002=>"111000000",
  63003=>"000000000",
  63004=>"111111000",
  63005=>"001000010",
  63006=>"111111110",
  63007=>"100000001",
  63008=>"000000000",
  63009=>"000001000",
  63010=>"111111011",
  63011=>"111111111",
  63012=>"100100111",
  63013=>"111110100",
  63014=>"111111111",
  63015=>"100000000",
  63016=>"100101001",
  63017=>"100000000",
  63018=>"000000000",
  63019=>"000010010",
  63020=>"111111111",
  63021=>"011111111",
  63022=>"001001000",
  63023=>"111111111",
  63024=>"000000000",
  63025=>"111111111",
  63026=>"100111111",
  63027=>"000001111",
  63028=>"101101101",
  63029=>"111001000",
  63030=>"000000000",
  63031=>"100001000",
  63032=>"111111111",
  63033=>"000010111",
  63034=>"000000000",
  63035=>"000111111",
  63036=>"101001011",
  63037=>"000010110",
  63038=>"001000000",
  63039=>"000000000",
  63040=>"011001000",
  63041=>"000000000",
  63042=>"010011000",
  63043=>"010110111",
  63044=>"111111011",
  63045=>"000000000",
  63046=>"011000000",
  63047=>"111111111",
  63048=>"111111000",
  63049=>"000000100",
  63050=>"000000001",
  63051=>"111101000",
  63052=>"111111111",
  63053=>"100000000",
  63054=>"000111111",
  63055=>"000000000",
  63056=>"000111111",
  63057=>"111000100",
  63058=>"111111001",
  63059=>"000000000",
  63060=>"001000101",
  63061=>"110111000",
  63062=>"111111111",
  63063=>"001000100",
  63064=>"001000110",
  63065=>"110000101",
  63066=>"111111111",
  63067=>"000001000",
  63068=>"111111111",
  63069=>"111011111",
  63070=>"000000000",
  63071=>"110110000",
  63072=>"001111010",
  63073=>"000100000",
  63074=>"000000000",
  63075=>"000000001",
  63076=>"111011111",
  63077=>"000001001",
  63078=>"100110011",
  63079=>"111011111",
  63080=>"100110000",
  63081=>"000000101",
  63082=>"000000100",
  63083=>"110100000",
  63084=>"000000000",
  63085=>"000000000",
  63086=>"000000000",
  63087=>"000000011",
  63088=>"000000000",
  63089=>"111111111",
  63090=>"100100110",
  63091=>"000011001",
  63092=>"010010111",
  63093=>"000000000",
  63094=>"111111111",
  63095=>"000111111",
  63096=>"000100100",
  63097=>"111111111",
  63098=>"011000000",
  63099=>"000000000",
  63100=>"100000000",
  63101=>"000000000",
  63102=>"000100111",
  63103=>"000000000",
  63104=>"000000001",
  63105=>"000111111",
  63106=>"000001000",
  63107=>"000000000",
  63108=>"111111111",
  63109=>"000000101",
  63110=>"100100000",
  63111=>"100011011",
  63112=>"111000000",
  63113=>"111111111",
  63114=>"000011011",
  63115=>"111010000",
  63116=>"111111111",
  63117=>"111000000",
  63118=>"111111111",
  63119=>"000000000",
  63120=>"000000000",
  63121=>"111101101",
  63122=>"111111111",
  63123=>"111001001",
  63124=>"001001001",
  63125=>"110011111",
  63126=>"000101101",
  63127=>"111110111",
  63128=>"000000000",
  63129=>"111100101",
  63130=>"111010000",
  63131=>"111111111",
  63132=>"000000000",
  63133=>"110100100",
  63134=>"000000001",
  63135=>"000000000",
  63136=>"000000100",
  63137=>"000111111",
  63138=>"000000000",
  63139=>"111110100",
  63140=>"111111111",
  63141=>"010110111",
  63142=>"111001101",
  63143=>"000010010",
  63144=>"000000000",
  63145=>"000111111",
  63146=>"000000000",
  63147=>"000000001",
  63148=>"010001011",
  63149=>"110110110",
  63150=>"000000101",
  63151=>"000011000",
  63152=>"000100000",
  63153=>"111111111",
  63154=>"111111010",
  63155=>"111100100",
  63156=>"111110000",
  63157=>"111000000",
  63158=>"000001111",
  63159=>"110111000",
  63160=>"111111111",
  63161=>"111001001",
  63162=>"111011011",
  63163=>"110110100",
  63164=>"001001000",
  63165=>"000000000",
  63166=>"000000111",
  63167=>"001001101",
  63168=>"000100111",
  63169=>"111000010",
  63170=>"101000000",
  63171=>"001111001",
  63172=>"000111111",
  63173=>"001111111",
  63174=>"000110111",
  63175=>"001001111",
  63176=>"000000111",
  63177=>"001001011",
  63178=>"000000000",
  63179=>"111111111",
  63180=>"000100111",
  63181=>"000000001",
  63182=>"010010000",
  63183=>"000000011",
  63184=>"010010000",
  63185=>"101000100",
  63186=>"110111111",
  63187=>"101000000",
  63188=>"100110010",
  63189=>"111111000",
  63190=>"000000000",
  63191=>"000000000",
  63192=>"100100111",
  63193=>"111111100",
  63194=>"000000000",
  63195=>"000111111",
  63196=>"110110000",
  63197=>"000001000",
  63198=>"110101111",
  63199=>"000110111",
  63200=>"100111111",
  63201=>"111001000",
  63202=>"000110111",
  63203=>"000010000",
  63204=>"111111110",
  63205=>"011111101",
  63206=>"111111111",
  63207=>"111111111",
  63208=>"111000000",
  63209=>"111101101",
  63210=>"000000001",
  63211=>"111111111",
  63212=>"000000001",
  63213=>"000111111",
  63214=>"000000111",
  63215=>"111100011",
  63216=>"000000000",
  63217=>"110110111",
  63218=>"001100100",
  63219=>"000000000",
  63220=>"011111111",
  63221=>"111000000",
  63222=>"000100000",
  63223=>"000000000",
  63224=>"110111111",
  63225=>"011001001",
  63226=>"111111111",
  63227=>"001001111",
  63228=>"111111111",
  63229=>"111111000",
  63230=>"010110111",
  63231=>"010010111",
  63232=>"000000000",
  63233=>"110110011",
  63234=>"111110111",
  63235=>"000000001",
  63236=>"000100101",
  63237=>"001001001",
  63238=>"000100111",
  63239=>"111101001",
  63240=>"000111111",
  63241=>"000101111",
  63242=>"111111100",
  63243=>"000000000",
  63244=>"111001101",
  63245=>"001000000",
  63246=>"000100000",
  63247=>"000001001",
  63248=>"111111000",
  63249=>"000111111",
  63250=>"101000000",
  63251=>"000010011",
  63252=>"000000000",
  63253=>"000000000",
  63254=>"100000111",
  63255=>"101101000",
  63256=>"111111111",
  63257=>"001011011",
  63258=>"111111100",
  63259=>"010110000",
  63260=>"011011011",
  63261=>"000000000",
  63262=>"000000000",
  63263=>"011111111",
  63264=>"010010011",
  63265=>"000000001",
  63266=>"111000000",
  63267=>"000000000",
  63268=>"001011001",
  63269=>"000000001",
  63270=>"000011111",
  63271=>"000111000",
  63272=>"111011000",
  63273=>"010111111",
  63274=>"111111011",
  63275=>"111111111",
  63276=>"000000110",
  63277=>"000000000",
  63278=>"100000000",
  63279=>"001001111",
  63280=>"000000000",
  63281=>"000000100",
  63282=>"100110111",
  63283=>"010010010",
  63284=>"000000001",
  63285=>"111100100",
  63286=>"000000011",
  63287=>"001011000",
  63288=>"000101100",
  63289=>"111000000",
  63290=>"010010010",
  63291=>"000000000",
  63292=>"010011111",
  63293=>"011111111",
  63294=>"111011001",
  63295=>"000000000",
  63296=>"101101111",
  63297=>"111111111",
  63298=>"000000000",
  63299=>"000000000",
  63300=>"111111110",
  63301=>"110111111",
  63302=>"000000011",
  63303=>"111111001",
  63304=>"001011111",
  63305=>"000000111",
  63306=>"000000000",
  63307=>"000000000",
  63308=>"111111111",
  63309=>"111101000",
  63310=>"111111111",
  63311=>"101001000",
  63312=>"011011111",
  63313=>"010011001",
  63314=>"000000011",
  63315=>"000000000",
  63316=>"000000000",
  63317=>"011011011",
  63318=>"111011111",
  63319=>"000000000",
  63320=>"111111111",
  63321=>"000000110",
  63322=>"111111000",
  63323=>"000111111",
  63324=>"000000000",
  63325=>"000001000",
  63326=>"111111100",
  63327=>"111111000",
  63328=>"111111111",
  63329=>"000010000",
  63330=>"100100100",
  63331=>"111111111",
  63332=>"111111100",
  63333=>"000000000",
  63334=>"111000000",
  63335=>"111111111",
  63336=>"100100000",
  63337=>"100111000",
  63338=>"000000000",
  63339=>"011011111",
  63340=>"000001011",
  63341=>"000000111",
  63342=>"000000000",
  63343=>"000000000",
  63344=>"000000000",
  63345=>"010000010",
  63346=>"000111111",
  63347=>"011111011",
  63348=>"000110110",
  63349=>"000000000",
  63350=>"100100110",
  63351=>"000000000",
  63352=>"000000111",
  63353=>"111111111",
  63354=>"000001111",
  63355=>"000011011",
  63356=>"011010000",
  63357=>"111111111",
  63358=>"000000000",
  63359=>"000101111",
  63360=>"100100001",
  63361=>"111011101",
  63362=>"000000000",
  63363=>"110111111",
  63364=>"010001011",
  63365=>"110001100",
  63366=>"000100000",
  63367=>"001110111",
  63368=>"111111101",
  63369=>"000010111",
  63370=>"101000011",
  63371=>"100101100",
  63372=>"100111111",
  63373=>"110111000",
  63374=>"111100000",
  63375=>"000001000",
  63376=>"000000000",
  63377=>"000000000",
  63378=>"000101001",
  63379=>"001000001",
  63380=>"111111000",
  63381=>"000000000",
  63382=>"001000000",
  63383=>"000000010",
  63384=>"000000000",
  63385=>"010111011",
  63386=>"000000001",
  63387=>"100000000",
  63388=>"000000000",
  63389=>"011000001",
  63390=>"101101111",
  63391=>"000000000",
  63392=>"000000000",
  63393=>"001011000",
  63394=>"000000000",
  63395=>"011011000",
  63396=>"110110111",
  63397=>"000111111",
  63398=>"100000000",
  63399=>"000011111",
  63400=>"111111111",
  63401=>"110011011",
  63402=>"000000000",
  63403=>"101101111",
  63404=>"000000000",
  63405=>"000000000",
  63406=>"000000000",
  63407=>"011111111",
  63408=>"111110000",
  63409=>"111111111",
  63410=>"100101111",
  63411=>"000000000",
  63412=>"101111101",
  63413=>"111110000",
  63414=>"100111111",
  63415=>"110110000",
  63416=>"100110000",
  63417=>"111111011",
  63418=>"000000011",
  63419=>"000000010",
  63420=>"011111001",
  63421=>"111111110",
  63422=>"111111101",
  63423=>"100100000",
  63424=>"111111011",
  63425=>"000000111",
  63426=>"001000000",
  63427=>"000000000",
  63428=>"111111111",
  63429=>"000000100",
  63430=>"000000011",
  63431=>"001001101",
  63432=>"000000000",
  63433=>"001011011",
  63434=>"000000000",
  63435=>"011001000",
  63436=>"000000000",
  63437=>"001111011",
  63438=>"100000001",
  63439=>"111111111",
  63440=>"101100100",
  63441=>"000000000",
  63442=>"111000000",
  63443=>"000001111",
  63444=>"111111011",
  63445=>"111111111",
  63446=>"111011010",
  63447=>"000011110",
  63448=>"100110100",
  63449=>"000100100",
  63450=>"111010000",
  63451=>"000000000",
  63452=>"000000000",
  63453=>"000001111",
  63454=>"000000000",
  63455=>"110000000",
  63456=>"111111111",
  63457=>"111011010",
  63458=>"001000000",
  63459=>"101111111",
  63460=>"111111000",
  63461=>"110000000",
  63462=>"000000100",
  63463=>"010000000",
  63464=>"100100101",
  63465=>"000000000",
  63466=>"111010000",
  63467=>"000000000",
  63468=>"011111101",
  63469=>"001000001",
  63470=>"111100111",
  63471=>"000111111",
  63472=>"111001011",
  63473=>"111110100",
  63474=>"101110111",
  63475=>"000000000",
  63476=>"111111111",
  63477=>"000000000",
  63478=>"000101001",
  63479=>"000000000",
  63480=>"111111111",
  63481=>"001001001",
  63482=>"010010000",
  63483=>"000000101",
  63484=>"111011000",
  63485=>"000000000",
  63486=>"000011110",
  63487=>"000000111",
  63488=>"111011111",
  63489=>"000111111",
  63490=>"111111111",
  63491=>"000000000",
  63492=>"100000111",
  63493=>"000000000",
  63494=>"011111110",
  63495=>"101111111",
  63496=>"111001101",
  63497=>"100000000",
  63498=>"010000000",
  63499=>"111111111",
  63500=>"000001001",
  63501=>"111100000",
  63502=>"000001011",
  63503=>"000000000",
  63504=>"111111000",
  63505=>"000000000",
  63506=>"000000001",
  63507=>"000000010",
  63508=>"000000100",
  63509=>"111001000",
  63510=>"111111101",
  63511=>"100001011",
  63512=>"000000001",
  63513=>"111111111",
  63514=>"000101111",
  63515=>"100100000",
  63516=>"110111011",
  63517=>"100000000",
  63518=>"110111111",
  63519=>"110100111",
  63520=>"000000000",
  63521=>"111111111",
  63522=>"111000001",
  63523=>"111001001",
  63524=>"111111111",
  63525=>"000110110",
  63526=>"001000001",
  63527=>"000000001",
  63528=>"110000000",
  63529=>"111100000",
  63530=>"000011111",
  63531=>"000111111",
  63532=>"001000000",
  63533=>"000000111",
  63534=>"011010111",
  63535=>"111100000",
  63536=>"001001001",
  63537=>"000000000",
  63538=>"010000000",
  63539=>"000100111",
  63540=>"111111111",
  63541=>"000000010",
  63542=>"011111111",
  63543=>"011001000",
  63544=>"001001000",
  63545=>"000000011",
  63546=>"000000000",
  63547=>"111111000",
  63548=>"111111111",
  63549=>"111011000",
  63550=>"011111111",
  63551=>"001001000",
  63552=>"111010010",
  63553=>"000010010",
  63554=>"000000001",
  63555=>"001001111",
  63556=>"011001000",
  63557=>"100101111",
  63558=>"111000111",
  63559=>"111111111",
  63560=>"111111011",
  63561=>"111100000",
  63562=>"111111111",
  63563=>"110110111",
  63564=>"111111000",
  63565=>"110010111",
  63566=>"001010010",
  63567=>"000011000",
  63568=>"111111101",
  63569=>"111111011",
  63570=>"000101111",
  63571=>"010011001",
  63572=>"000000000",
  63573=>"000000000",
  63574=>"001000000",
  63575=>"000001001",
  63576=>"110111011",
  63577=>"101101111",
  63578=>"100100100",
  63579=>"000000000",
  63580=>"000100000",
  63581=>"101101101",
  63582=>"001111111",
  63583=>"111011000",
  63584=>"000011111",
  63585=>"001001000",
  63586=>"111101001",
  63587=>"010000100",
  63588=>"000011010",
  63589=>"110000000",
  63590=>"001000000",
  63591=>"000100111",
  63592=>"111111110",
  63593=>"111101000",
  63594=>"011111111",
  63595=>"111100000",
  63596=>"111111011",
  63597=>"111111111",
  63598=>"111111111",
  63599=>"001111111",
  63600=>"000000000",
  63601=>"111111000",
  63602=>"111011011",
  63603=>"111011011",
  63604=>"000000000",
  63605=>"000000000",
  63606=>"000000000",
  63607=>"000001111",
  63608=>"100100000",
  63609=>"101001100",
  63610=>"000000000",
  63611=>"000010000",
  63612=>"111111010",
  63613=>"000110000",
  63614=>"011011011",
  63615=>"111111111",
  63616=>"000100111",
  63617=>"111000000",
  63618=>"111111111",
  63619=>"000000011",
  63620=>"100100100",
  63621=>"111111111",
  63622=>"111000111",
  63623=>"000001000",
  63624=>"111111111",
  63625=>"011011001",
  63626=>"011010111",
  63627=>"110100110",
  63628=>"000111111",
  63629=>"000001101",
  63630=>"000000000",
  63631=>"000000000",
  63632=>"111111111",
  63633=>"000000000",
  63634=>"101001001",
  63635=>"000000000",
  63636=>"000010110",
  63637=>"000000111",
  63638=>"111111111",
  63639=>"111111111",
  63640=>"000101000",
  63641=>"111100101",
  63642=>"000001111",
  63643=>"111111011",
  63644=>"111111111",
  63645=>"000000000",
  63646=>"111100100",
  63647=>"000000111",
  63648=>"000000000",
  63649=>"111111110",
  63650=>"110000101",
  63651=>"000000000",
  63652=>"110110000",
  63653=>"101111111",
  63654=>"001000000",
  63655=>"011111110",
  63656=>"111111101",
  63657=>"000000000",
  63658=>"111111111",
  63659=>"110000000",
  63660=>"111111111",
  63661=>"001001011",
  63662=>"001011001",
  63663=>"000000110",
  63664=>"000111111",
  63665=>"110111111",
  63666=>"011111011",
  63667=>"111111100",
  63668=>"000100000",
  63669=>"111000000",
  63670=>"000001001",
  63671=>"000000100",
  63672=>"111111011",
  63673=>"111111111",
  63674=>"000000000",
  63675=>"000000000",
  63676=>"111111111",
  63677=>"110111000",
  63678=>"111111111",
  63679=>"100000000",
  63680=>"000000000",
  63681=>"000000011",
  63682=>"011111111",
  63683=>"001000000",
  63684=>"111101111",
  63685=>"111111100",
  63686=>"000000000",
  63687=>"000100000",
  63688=>"001001111",
  63689=>"111111111",
  63690=>"111011001",
  63691=>"111110111",
  63692=>"000011111",
  63693=>"111000001",
  63694=>"111111000",
  63695=>"101111001",
  63696=>"101101100",
  63697=>"001000000",
  63698=>"011111111",
  63699=>"110111111",
  63700=>"110000000",
  63701=>"001000100",
  63702=>"000000101",
  63703=>"000001001",
  63704=>"101000100",
  63705=>"110111111",
  63706=>"000000000",
  63707=>"000100101",
  63708=>"111111101",
  63709=>"000000000",
  63710=>"000001001",
  63711=>"111111111",
  63712=>"011000000",
  63713=>"000000000",
  63714=>"111111111",
  63715=>"111111111",
  63716=>"101111111",
  63717=>"100110000",
  63718=>"001000000",
  63719=>"000000000",
  63720=>"000000000",
  63721=>"101001001",
  63722=>"000000000",
  63723=>"111111100",
  63724=>"000000010",
  63725=>"000000100",
  63726=>"110000111",
  63727=>"111111111",
  63728=>"001000000",
  63729=>"111000000",
  63730=>"111111111",
  63731=>"111111000",
  63732=>"100100111",
  63733=>"111111000",
  63734=>"110010000",
  63735=>"111111111",
  63736=>"111101111",
  63737=>"011000000",
  63738=>"111111000",
  63739=>"111011000",
  63740=>"001111111",
  63741=>"110101001",
  63742=>"001000000",
  63743=>"000100100",
  63744=>"000000001",
  63745=>"001011111",
  63746=>"111111111",
  63747=>"111101000",
  63748=>"100111000",
  63749=>"000010010",
  63750=>"111111000",
  63751=>"011001111",
  63752=>"111111001",
  63753=>"000000000",
  63754=>"100100000",
  63755=>"111111011",
  63756=>"001001011",
  63757=>"111111111",
  63758=>"000001111",
  63759=>"110111111",
  63760=>"111000000",
  63761=>"001001111",
  63762=>"000000000",
  63763=>"111001101",
  63764=>"001001001",
  63765=>"000000000",
  63766=>"111011001",
  63767=>"100000000",
  63768=>"110110000",
  63769=>"111111111",
  63770=>"000000001",
  63771=>"001000111",
  63772=>"111111110",
  63773=>"111001000",
  63774=>"111101101",
  63775=>"101000010",
  63776=>"111111001",
  63777=>"100100000",
  63778=>"100100101",
  63779=>"011000000",
  63780=>"000000000",
  63781=>"000000001",
  63782=>"100111111",
  63783=>"011011010",
  63784=>"111111111",
  63785=>"000000000",
  63786=>"000100001",
  63787=>"111111111",
  63788=>"001111111",
  63789=>"000000000",
  63790=>"000000000",
  63791=>"001000101",
  63792=>"110110111",
  63793=>"111100111",
  63794=>"001111110",
  63795=>"000000000",
  63796=>"100100000",
  63797=>"000011011",
  63798=>"111111101",
  63799=>"100000000",
  63800=>"010011000",
  63801=>"101000000",
  63802=>"111000000",
  63803=>"110111001",
  63804=>"000000100",
  63805=>"100100100",
  63806=>"000000000",
  63807=>"001000000",
  63808=>"000000111",
  63809=>"111110000",
  63810=>"000000001",
  63811=>"000000000",
  63812=>"001001000",
  63813=>"000000111",
  63814=>"000000000",
  63815=>"000001001",
  63816=>"101000000",
  63817=>"000000100",
  63818=>"001111111",
  63819=>"111111111",
  63820=>"001001000",
  63821=>"000001111",
  63822=>"001111111",
  63823=>"110111111",
  63824=>"100100100",
  63825=>"000000000",
  63826=>"000100111",
  63827=>"100000111",
  63828=>"000000000",
  63829=>"001000000",
  63830=>"111111111",
  63831=>"111111010",
  63832=>"111110111",
  63833=>"100000000",
  63834=>"100111010",
  63835=>"000000000",
  63836=>"100100000",
  63837=>"000000001",
  63838=>"001111111",
  63839=>"100000011",
  63840=>"100000000",
  63841=>"100001001",
  63842=>"111000001",
  63843=>"101111111",
  63844=>"111111111",
  63845=>"001000000",
  63846=>"100000000",
  63847=>"111111001",
  63848=>"111111101",
  63849=>"111101101",
  63850=>"000000000",
  63851=>"111010000",
  63852=>"010011011",
  63853=>"110000000",
  63854=>"000000000",
  63855=>"111111111",
  63856=>"101000000",
  63857=>"001011000",
  63858=>"111000000",
  63859=>"011010000",
  63860=>"000000000",
  63861=>"111111111",
  63862=>"010000000",
  63863=>"000000000",
  63864=>"000000000",
  63865=>"111001000",
  63866=>"000000000",
  63867=>"001000000",
  63868=>"111110000",
  63869=>"000000001",
  63870=>"001000001",
  63871=>"000000000",
  63872=>"111001011",
  63873=>"001001000",
  63874=>"001100110",
  63875=>"011011110",
  63876=>"000000111",
  63877=>"011000000",
  63878=>"111000000",
  63879=>"101000000",
  63880=>"000001111",
  63881=>"100110100",
  63882=>"111111111",
  63883=>"111111111",
  63884=>"000000000",
  63885=>"111011000",
  63886=>"010111111",
  63887=>"000000001",
  63888=>"110000001",
  63889=>"111111111",
  63890=>"100100111",
  63891=>"000000001",
  63892=>"000111111",
  63893=>"000000000",
  63894=>"111111111",
  63895=>"110000000",
  63896=>"000001001",
  63897=>"111111011",
  63898=>"111111111",
  63899=>"000001111",
  63900=>"111101100",
  63901=>"111111000",
  63902=>"111111111",
  63903=>"000000000",
  63904=>"101101000",
  63905=>"111011011",
  63906=>"110011001",
  63907=>"111100000",
  63908=>"000000000",
  63909=>"011000011",
  63910=>"000000000",
  63911=>"100000000",
  63912=>"110000000",
  63913=>"111101111",
  63914=>"000000000",
  63915=>"000000000",
  63916=>"100110111",
  63917=>"000000000",
  63918=>"111100000",
  63919=>"111111111",
  63920=>"111011011",
  63921=>"111111110",
  63922=>"111110111",
  63923=>"011011101",
  63924=>"111111010",
  63925=>"000000000",
  63926=>"001111111",
  63927=>"111111111",
  63928=>"111111111",
  63929=>"111101000",
  63930=>"101100000",
  63931=>"000100100",
  63932=>"111111111",
  63933=>"100111111",
  63934=>"111111111",
  63935=>"111011000",
  63936=>"111111111",
  63937=>"000000000",
  63938=>"111111111",
  63939=>"111001001",
  63940=>"001000001",
  63941=>"011000000",
  63942=>"000000101",
  63943=>"111111101",
  63944=>"000101101",
  63945=>"001000001",
  63946=>"101111111",
  63947=>"111110000",
  63948=>"000000010",
  63949=>"111110111",
  63950=>"111101001",
  63951=>"111001111",
  63952=>"001111111",
  63953=>"000000000",
  63954=>"001111011",
  63955=>"111111111",
  63956=>"111111111",
  63957=>"110100011",
  63958=>"000000000",
  63959=>"010110110",
  63960=>"110011000",
  63961=>"111111111",
  63962=>"000010000",
  63963=>"001000001",
  63964=>"000000000",
  63965=>"110110000",
  63966=>"000000000",
  63967=>"000100111",
  63968=>"001111111",
  63969=>"001001100",
  63970=>"100110111",
  63971=>"000111011",
  63972=>"111111010",
  63973=>"000000000",
  63974=>"000010111",
  63975=>"101100000",
  63976=>"010000000",
  63977=>"100000000",
  63978=>"000000000",
  63979=>"000000111",
  63980=>"000111111",
  63981=>"000000000",
  63982=>"000111111",
  63983=>"111101101",
  63984=>"111111011",
  63985=>"111111111",
  63986=>"111111010",
  63987=>"111111111",
  63988=>"111011000",
  63989=>"111111111",
  63990=>"101111111",
  63991=>"001001111",
  63992=>"111111100",
  63993=>"111100000",
  63994=>"001001001",
  63995=>"111001111",
  63996=>"111000000",
  63997=>"001011000",
  63998=>"111011011",
  63999=>"000000000",
  64000=>"011011111",
  64001=>"000000000",
  64002=>"000111011",
  64003=>"111110011",
  64004=>"100000000",
  64005=>"111101101",
  64006=>"001001101",
  64007=>"011011000",
  64008=>"100110110",
  64009=>"000000100",
  64010=>"100111111",
  64011=>"000011111",
  64012=>"000000000",
  64013=>"111111111",
  64014=>"111111111",
  64015=>"000000000",
  64016=>"111000101",
  64017=>"000000111",
  64018=>"000011000",
  64019=>"111110110",
  64020=>"111100101",
  64021=>"111111111",
  64022=>"111111111",
  64023=>"000000000",
  64024=>"001001011",
  64025=>"000001001",
  64026=>"111111010",
  64027=>"000100111",
  64028=>"111111000",
  64029=>"111011001",
  64030=>"011000000",
  64031=>"000000011",
  64032=>"111111110",
  64033=>"000100110",
  64034=>"111111001",
  64035=>"011111111",
  64036=>"100000111",
  64037=>"111111111",
  64038=>"000000000",
  64039=>"000000000",
  64040=>"100000001",
  64041=>"111111111",
  64042=>"000000000",
  64043=>"100100101",
  64044=>"000000000",
  64045=>"110111011",
  64046=>"111111111",
  64047=>"111111001",
  64048=>"111111111",
  64049=>"111111000",
  64050=>"100100001",
  64051=>"100100111",
  64052=>"101100100",
  64053=>"010010111",
  64054=>"000000000",
  64055=>"000111111",
  64056=>"110111111",
  64057=>"000000000",
  64058=>"101101000",
  64059=>"100111111",
  64060=>"011000111",
  64061=>"000000111",
  64062=>"000000111",
  64063=>"111111111",
  64064=>"111011100",
  64065=>"011111111",
  64066=>"000000000",
  64067=>"100100000",
  64068=>"011011111",
  64069=>"011111011",
  64070=>"000000000",
  64071=>"000000000",
  64072=>"110000000",
  64073=>"001001001",
  64074=>"111101111",
  64075=>"000000000",
  64076=>"000011011",
  64077=>"111111110",
  64078=>"101000000",
  64079=>"000100111",
  64080=>"000011111",
  64081=>"111111111",
  64082=>"110110111",
  64083=>"001011111",
  64084=>"111111111",
  64085=>"000111111",
  64086=>"000000110",
  64087=>"000000000",
  64088=>"111000000",
  64089=>"111100111",
  64090=>"000000000",
  64091=>"001001001",
  64092=>"000000000",
  64093=>"001001000",
  64094=>"001001001",
  64095=>"111111110",
  64096=>"111101011",
  64097=>"111111011",
  64098=>"110010100",
  64099=>"111000000",
  64100=>"011110110",
  64101=>"101111101",
  64102=>"011000000",
  64103=>"000101111",
  64104=>"101100000",
  64105=>"111111111",
  64106=>"000000000",
  64107=>"000000000",
  64108=>"011111100",
  64109=>"000000000",
  64110=>"111111000",
  64111=>"001000101",
  64112=>"111111011",
  64113=>"111111111",
  64114=>"000110110",
  64115=>"000010011",
  64116=>"111110110",
  64117=>"000000000",
  64118=>"111111000",
  64119=>"111111111",
  64120=>"011000001",
  64121=>"110111111",
  64122=>"000000000",
  64123=>"111000000",
  64124=>"111110110",
  64125=>"001000000",
  64126=>"000000000",
  64127=>"111111010",
  64128=>"000000000",
  64129=>"000000111",
  64130=>"111111101",
  64131=>"110011000",
  64132=>"001001100",
  64133=>"111001111",
  64134=>"001000111",
  64135=>"111111111",
  64136=>"000000000",
  64137=>"111111111",
  64138=>"000001001",
  64139=>"111111111",
  64140=>"000000000",
  64141=>"101111111",
  64142=>"111011001",
  64143=>"000000000",
  64144=>"000000000",
  64145=>"000000000",
  64146=>"111100100",
  64147=>"000000000",
  64148=>"111111111",
  64149=>"000001000",
  64150=>"111111111",
  64151=>"000000000",
  64152=>"111100100",
  64153=>"000010111",
  64154=>"000000111",
  64155=>"111111100",
  64156=>"110110111",
  64157=>"000101001",
  64158=>"000000000",
  64159=>"000000010",
  64160=>"111100100",
  64161=>"000010000",
  64162=>"011110000",
  64163=>"101101100",
  64164=>"000000000",
  64165=>"111001101",
  64166=>"111111000",
  64167=>"101000000",
  64168=>"000000100",
  64169=>"001000000",
  64170=>"000000000",
  64171=>"111111111",
  64172=>"000000000",
  64173=>"001000100",
  64174=>"000000001",
  64175=>"000100100",
  64176=>"111111111",
  64177=>"000000000",
  64178=>"000111010",
  64179=>"111111100",
  64180=>"011010111",
  64181=>"111111111",
  64182=>"000000000",
  64183=>"010000000",
  64184=>"001001110",
  64185=>"100100000",
  64186=>"111110110",
  64187=>"010000100",
  64188=>"111111111",
  64189=>"111111111",
  64190=>"111111111",
  64191=>"111111110",
  64192=>"000000011",
  64193=>"111111000",
  64194=>"000000011",
  64195=>"000000000",
  64196=>"000100111",
  64197=>"000000000",
  64198=>"011111000",
  64199=>"000100100",
  64200=>"001001011",
  64201=>"111111111",
  64202=>"000001001",
  64203=>"111100000",
  64204=>"000000000",
  64205=>"000000111",
  64206=>"000000001",
  64207=>"000000001",
  64208=>"100111001",
  64209=>"111111101",
  64210=>"101001000",
  64211=>"101000111",
  64212=>"001001011",
  64213=>"000010110",
  64214=>"110110110",
  64215=>"111000101",
  64216=>"000000000",
  64217=>"111011111",
  64218=>"000000110",
  64219=>"000110011",
  64220=>"111000000",
  64221=>"111111111",
  64222=>"000010000",
  64223=>"000111111",
  64224=>"000111111",
  64225=>"110111111",
  64226=>"000000000",
  64227=>"100110111",
  64228=>"111111010",
  64229=>"100100110",
  64230=>"111111111",
  64231=>"111111111",
  64232=>"111111111",
  64233=>"000000000",
  64234=>"111111000",
  64235=>"000000000",
  64236=>"000110000",
  64237=>"000000110",
  64238=>"000001111",
  64239=>"000000001",
  64240=>"011011111",
  64241=>"000000000",
  64242=>"110000000",
  64243=>"100100100",
  64244=>"000000100",
  64245=>"111111001",
  64246=>"111111111",
  64247=>"111111111",
  64248=>"000000000",
  64249=>"111100000",
  64250=>"111000111",
  64251=>"000000000",
  64252=>"110110000",
  64253=>"111011011",
  64254=>"000000100",
  64255=>"100110111",
  64256=>"100100111",
  64257=>"001000000",
  64258=>"111111011",
  64259=>"111111111",
  64260=>"011111111",
  64261=>"111111000",
  64262=>"000001100",
  64263=>"000000001",
  64264=>"000000000",
  64265=>"000000000",
  64266=>"111111111",
  64267=>"101111111",
  64268=>"000000110",
  64269=>"000010010",
  64270=>"011000111",
  64271=>"111111111",
  64272=>"000000000",
  64273=>"000000001",
  64274=>"111111000",
  64275=>"011111111",
  64276=>"000000011",
  64277=>"000000000",
  64278=>"100100000",
  64279=>"101101101",
  64280=>"000000011",
  64281=>"111111111",
  64282=>"000000000",
  64283=>"000100111",
  64284=>"000000110",
  64285=>"111111111",
  64286=>"111111111",
  64287=>"111101000",
  64288=>"100100000",
  64289=>"000000001",
  64290=>"111111111",
  64291=>"001001001",
  64292=>"000000000",
  64293=>"100100111",
  64294=>"000100100",
  64295=>"101111000",
  64296=>"001000000",
  64297=>"011111111",
  64298=>"000000000",
  64299=>"100000111",
  64300=>"000000000",
  64301=>"000000000",
  64302=>"111111111",
  64303=>"001000000",
  64304=>"111111111",
  64305=>"011001001",
  64306=>"111111101",
  64307=>"111000000",
  64308=>"111111111",
  64309=>"000100111",
  64310=>"111010000",
  64311=>"111111111",
  64312=>"000000000",
  64313=>"000000000",
  64314=>"001111110",
  64315=>"100110100",
  64316=>"001000111",
  64317=>"000000000",
  64318=>"000111111",
  64319=>"011001001",
  64320=>"010111111",
  64321=>"000000000",
  64322=>"111111100",
  64323=>"000000010",
  64324=>"000000000",
  64325=>"111111111",
  64326=>"000011010",
  64327=>"000000000",
  64328=>"111111111",
  64329=>"001000000",
  64330=>"011100100",
  64331=>"111111111",
  64332=>"111111011",
  64333=>"001000111",
  64334=>"011001001",
  64335=>"110111101",
  64336=>"000000110",
  64337=>"111100111",
  64338=>"111000000",
  64339=>"011001000",
  64340=>"111011000",
  64341=>"001011011",
  64342=>"111111111",
  64343=>"001000000",
  64344=>"111111000",
  64345=>"111111111",
  64346=>"111111111",
  64347=>"111101000",
  64348=>"000100111",
  64349=>"111111011",
  64350=>"111111000",
  64351=>"000000000",
  64352=>"111000000",
  64353=>"111111111",
  64354=>"000000001",
  64355=>"000011011",
  64356=>"000000110",
  64357=>"111111111",
  64358=>"000000000",
  64359=>"111000111",
  64360=>"011001000",
  64361=>"110110011",
  64362=>"011111011",
  64363=>"101111111",
  64364=>"001001001",
  64365=>"111100111",
  64366=>"000000000",
  64367=>"001000010",
  64368=>"111111100",
  64369=>"111000111",
  64370=>"011100101",
  64371=>"111111111",
  64372=>"111100100",
  64373=>"011001001",
  64374=>"111110000",
  64375=>"101111110",
  64376=>"000000000",
  64377=>"000100000",
  64378=>"011011111",
  64379=>"000000000",
  64380=>"111111111",
  64381=>"111110111",
  64382=>"101000000",
  64383=>"000000110",
  64384=>"000000111",
  64385=>"111011111",
  64386=>"100000000",
  64387=>"110000110",
  64388=>"111111011",
  64389=>"100000111",
  64390=>"100000000",
  64391=>"000000000",
  64392=>"111111010",
  64393=>"111111101",
  64394=>"111111111",
  64395=>"000101101",
  64396=>"000000111",
  64397=>"111110110",
  64398=>"011111111",
  64399=>"100000000",
  64400=>"101000000",
  64401=>"101001001",
  64402=>"111111011",
  64403=>"000000011",
  64404=>"110111111",
  64405=>"000000011",
  64406=>"110111111",
  64407=>"000000000",
  64408=>"111111111",
  64409=>"111011111",
  64410=>"111111011",
  64411=>"000000000",
  64412=>"000000100",
  64413=>"000000000",
  64414=>"111000000",
  64415=>"111111110",
  64416=>"011011111",
  64417=>"011000001",
  64418=>"111100111",
  64419=>"000000000",
  64420=>"111111111",
  64421=>"111111000",
  64422=>"111111011",
  64423=>"000010111",
  64424=>"001000000",
  64425=>"110110110",
  64426=>"000111111",
  64427=>"000000000",
  64428=>"000000000",
  64429=>"000000000",
  64430=>"000000000",
  64431=>"010000001",
  64432=>"001111111",
  64433=>"110111010",
  64434=>"110000000",
  64435=>"001100000",
  64436=>"111001111",
  64437=>"111011111",
  64438=>"111111111",
  64439=>"000000000",
  64440=>"111111111",
  64441=>"000100100",
  64442=>"000000100",
  64443=>"011111111",
  64444=>"000000000",
  64445=>"000000000",
  64446=>"100100100",
  64447=>"011000000",
  64448=>"100111011",
  64449=>"111010000",
  64450=>"001000000",
  64451=>"001111111",
  64452=>"000000000",
  64453=>"000010111",
  64454=>"000000000",
  64455=>"000000000",
  64456=>"111000000",
  64457=>"100111000",
  64458=>"001000000",
  64459=>"011111111",
  64460=>"111111111",
  64461=>"001001001",
  64462=>"111111000",
  64463=>"110111111",
  64464=>"111011011",
  64465=>"000000000",
  64466=>"111011111",
  64467=>"011011011",
  64468=>"100000001",
  64469=>"000110010",
  64470=>"111101100",
  64471=>"000000010",
  64472=>"000000000",
  64473=>"111011000",
  64474=>"000010000",
  64475=>"111001000",
  64476=>"000000011",
  64477=>"000000101",
  64478=>"000000000",
  64479=>"001000011",
  64480=>"100110111",
  64481=>"000000000",
  64482=>"010110110",
  64483=>"000111101",
  64484=>"000111111",
  64485=>"111111111",
  64486=>"111110111",
  64487=>"111111111",
  64488=>"000000111",
  64489=>"000000000",
  64490=>"111010000",
  64491=>"000000000",
  64492=>"111100011",
  64493=>"101101001",
  64494=>"111001011",
  64495=>"000001111",
  64496=>"000000000",
  64497=>"001001111",
  64498=>"111111111",
  64499=>"000111001",
  64500=>"100100000",
  64501=>"011111111",
  64502=>"111101111",
  64503=>"000000001",
  64504=>"001001111",
  64505=>"000000100",
  64506=>"110000000",
  64507=>"000000000",
  64508=>"001011011",
  64509=>"111111101",
  64510=>"000000001",
  64511=>"111001111",
  64512=>"001000000",
  64513=>"110110010",
  64514=>"010110111",
  64515=>"000000000",
  64516=>"100110111",
  64517=>"011011011",
  64518=>"100000001",
  64519=>"111111111",
  64520=>"011111000",
  64521=>"111111111",
  64522=>"000000000",
  64523=>"000000000",
  64524=>"000000110",
  64525=>"100000011",
  64526=>"011111111",
  64527=>"111001001",
  64528=>"001001000",
  64529=>"100110111",
  64530=>"100100101",
  64531=>"000000100",
  64532=>"000000000",
  64533=>"000100111",
  64534=>"010000011",
  64535=>"100100000",
  64536=>"000000000",
  64537=>"000000011",
  64538=>"111000000",
  64539=>"011001001",
  64540=>"000001110",
  64541=>"111101111",
  64542=>"110110111",
  64543=>"111111111",
  64544=>"110110110",
  64545=>"000001000",
  64546=>"001001001",
  64547=>"111010000",
  64548=>"000000000",
  64549=>"000000110",
  64550=>"111111111",
  64551=>"000000100",
  64552=>"111111111",
  64553=>"000110000",
  64554=>"100000000",
  64555=>"111111111",
  64556=>"101011010",
  64557=>"001001011",
  64558=>"000100111",
  64559=>"011011111",
  64560=>"011011111",
  64561=>"000000000",
  64562=>"000000000",
  64563=>"000000000",
  64564=>"001001011",
  64565=>"000000000",
  64566=>"111001001",
  64567=>"000011011",
  64568=>"000000000",
  64569=>"000000000",
  64570=>"111111111",
  64571=>"010110000",
  64572=>"000111001",
  64573=>"011001001",
  64574=>"111110111",
  64575=>"000000001",
  64576=>"011001111",
  64577=>"000110000",
  64578=>"111111111",
  64579=>"000000111",
  64580=>"001001001",
  64581=>"111101011",
  64582=>"111011001",
  64583=>"111111111",
  64584=>"011010000",
  64585=>"000000000",
  64586=>"000000110",
  64587=>"001011001",
  64588=>"001000111",
  64589=>"110110110",
  64590=>"111000000",
  64591=>"001001001",
  64592=>"000000000",
  64593=>"000000011",
  64594=>"111111111",
  64595=>"001001111",
  64596=>"100100111",
  64597=>"100100111",
  64598=>"001000000",
  64599=>"111111111",
  64600=>"111111111",
  64601=>"000000000",
  64602=>"111011001",
  64603=>"011111011",
  64604=>"110110011",
  64605=>"111111111",
  64606=>"111111111",
  64607=>"111111110",
  64608=>"111000000",
  64609=>"001010000",
  64610=>"010111111",
  64611=>"111111111",
  64612=>"001001011",
  64613=>"110111111",
  64614=>"010000010",
  64615=>"111111111",
  64616=>"111101111",
  64617=>"001100111",
  64618=>"100000000",
  64619=>"000000000",
  64620=>"111101001",
  64621=>"101111111",
  64622=>"110111111",
  64623=>"100110100",
  64624=>"111111110",
  64625=>"101111011",
  64626=>"111111111",
  64627=>"110110110",
  64628=>"000000000",
  64629=>"110111100",
  64630=>"000000000",
  64631=>"100000001",
  64632=>"000000000",
  64633=>"010000000",
  64634=>"111110101",
  64635=>"000000110",
  64636=>"000100110",
  64637=>"000001011",
  64638=>"111000000",
  64639=>"111111111",
  64640=>"000000000",
  64641=>"000000001",
  64642=>"111111111",
  64643=>"011010000",
  64644=>"000011011",
  64645=>"000000000",
  64646=>"000010111",
  64647=>"011001111",
  64648=>"000000011",
  64649=>"111111111",
  64650=>"000110100",
  64651=>"000000001",
  64652=>"111111111",
  64653=>"111111111",
  64654=>"001000000",
  64655=>"101001101",
  64656=>"111111111",
  64657=>"110000000",
  64658=>"111000011",
  64659=>"000000000",
  64660=>"011010000",
  64661=>"111111111",
  64662=>"111111111",
  64663=>"001001000",
  64664=>"000000011",
  64665=>"101000011",
  64666=>"111111111",
  64667=>"011011011",
  64668=>"001011000",
  64669=>"110111001",
  64670=>"000000000",
  64671=>"010000000",
  64672=>"101000000",
  64673=>"110101101",
  64674=>"011000001",
  64675=>"010111011",
  64676=>"111100000",
  64677=>"000100110",
  64678=>"000101111",
  64679=>"001001001",
  64680=>"000000011",
  64681=>"111000101",
  64682=>"111111111",
  64683=>"100100110",
  64684=>"111111111",
  64685=>"000000000",
  64686=>"011000000",
  64687=>"111000000",
  64688=>"111111111",
  64689=>"001111010",
  64690=>"000000000",
  64691=>"010001001",
  64692=>"000000100",
  64693=>"011111100",
  64694=>"111111111",
  64695=>"111000000",
  64696=>"111001011",
  64697=>"001000101",
  64698=>"001110110",
  64699=>"000000011",
  64700=>"111111111",
  64701=>"111111111",
  64702=>"000000000",
  64703=>"000000000",
  64704=>"111111111",
  64705=>"110111011",
  64706=>"111111111",
  64707=>"000000000",
  64708=>"011001010",
  64709=>"000000000",
  64710=>"001011000",
  64711=>"011111010",
  64712=>"100111111",
  64713=>"011000101",
  64714=>"111111011",
  64715=>"111111111",
  64716=>"011011111",
  64717=>"000001111",
  64718=>"111011011",
  64719=>"111101110",
  64720=>"000000111",
  64721=>"000010011",
  64722=>"101100111",
  64723=>"000000000",
  64724=>"111101111",
  64725=>"100000000",
  64726=>"111011000",
  64727=>"000000001",
  64728=>"001000001",
  64729=>"100001111",
  64730=>"111011000",
  64731=>"011111001",
  64732=>"111011110",
  64733=>"011111111",
  64734=>"111001111",
  64735=>"000000000",
  64736=>"000010011",
  64737=>"000000000",
  64738=>"111111111",
  64739=>"111111011",
  64740=>"110110110",
  64741=>"100110100",
  64742=>"110111110",
  64743=>"001011001",
  64744=>"011111111",
  64745=>"000111111",
  64746=>"000100111",
  64747=>"100000001",
  64748=>"111111111",
  64749=>"111001001",
  64750=>"111111111",
  64751=>"000010111",
  64752=>"110110110",
  64753=>"111001110",
  64754=>"000000011",
  64755=>"000000000",
  64756=>"111011011",
  64757=>"110101111",
  64758=>"000000000",
  64759=>"111011000",
  64760=>"100000000",
  64761=>"111111111",
  64762=>"001000011",
  64763=>"000000010",
  64764=>"100010000",
  64765=>"000000001",
  64766=>"111111000",
  64767=>"111111111",
  64768=>"001000000",
  64769=>"000000000",
  64770=>"000000000",
  64771=>"000000001",
  64772=>"111111111",
  64773=>"100100111",
  64774=>"111011111",
  64775=>"000000001",
  64776=>"111110010",
  64777=>"111110110",
  64778=>"000001111",
  64779=>"100111111",
  64780=>"110110110",
  64781=>"011101101",
  64782=>"000000000",
  64783=>"000000001",
  64784=>"111111110",
  64785=>"100111111",
  64786=>"100100100",
  64787=>"000100100",
  64788=>"111111111",
  64789=>"111111110",
  64790=>"000000000",
  64791=>"110100111",
  64792=>"001101111",
  64793=>"111111111",
  64794=>"111111000",
  64795=>"000000000",
  64796=>"000000000",
  64797=>"101101111",
  64798=>"110110011",
  64799=>"111110111",
  64800=>"000100100",
  64801=>"110111010",
  64802=>"111111111",
  64803=>"111100111",
  64804=>"000000000",
  64805=>"010010111",
  64806=>"000001011",
  64807=>"111111111",
  64808=>"001011000",
  64809=>"011111111",
  64810=>"111111111",
  64811=>"011110110",
  64812=>"111111000",
  64813=>"000001001",
  64814=>"111111111",
  64815=>"000000000",
  64816=>"111111110",
  64817=>"111111001",
  64818=>"000000111",
  64819=>"000100111",
  64820=>"111011111",
  64821=>"000000000",
  64822=>"001011111",
  64823=>"000010010",
  64824=>"111011011",
  64825=>"000000000",
  64826=>"110110110",
  64827=>"000111001",
  64828=>"100000000",
  64829=>"001001111",
  64830=>"000100100",
  64831=>"000000000",
  64832=>"001000000",
  64833=>"000000000",
  64834=>"000000000",
  64835=>"111011011",
  64836=>"000000000",
  64837=>"111001001",
  64838=>"101101100",
  64839=>"110011011",
  64840=>"110000000",
  64841=>"110110111",
  64842=>"110111111",
  64843=>"111011001",
  64844=>"111111111",
  64845=>"000000100",
  64846=>"111111110",
  64847=>"100100111",
  64848=>"011011110",
  64849=>"000000110",
  64850=>"110110110",
  64851=>"000000000",
  64852=>"000000000",
  64853=>"100100101",
  64854=>"000000111",
  64855=>"011000001",
  64856=>"000000000",
  64857=>"111111111",
  64858=>"111000000",
  64859=>"000000011",
  64860=>"110111111",
  64861=>"100100111",
  64862=>"100100001",
  64863=>"001001111",
  64864=>"001101110",
  64865=>"111101111",
  64866=>"111111010",
  64867=>"000000011",
  64868=>"000001001",
  64869=>"011000000",
  64870=>"100110110",
  64871=>"010001001",
  64872=>"000000010",
  64873=>"001011001",
  64874=>"100100100",
  64875=>"000010000",
  64876=>"110110100",
  64877=>"111111111",
  64878=>"010011010",
  64879=>"000110100",
  64880=>"111110000",
  64881=>"111111110",
  64882=>"001101001",
  64883=>"111101101",
  64884=>"100100100",
  64885=>"000000000",
  64886=>"111111011",
  64887=>"110000010",
  64888=>"111111110",
  64889=>"110000000",
  64890=>"110000010",
  64891=>"000000000",
  64892=>"000000000",
  64893=>"111000000",
  64894=>"111101111",
  64895=>"000000101",
  64896=>"000001111",
  64897=>"111011011",
  64898=>"111101100",
  64899=>"100110110",
  64900=>"000000110",
  64901=>"000000000",
  64902=>"110111111",
  64903=>"111110111",
  64904=>"110101000",
  64905=>"000000001",
  64906=>"010011011",
  64907=>"000000000",
  64908=>"111111111",
  64909=>"000000000",
  64910=>"011011011",
  64911=>"000000000",
  64912=>"010011000",
  64913=>"001001001",
  64914=>"000000000",
  64915=>"000000000",
  64916=>"000000011",
  64917=>"000000000",
  64918=>"111110000",
  64919=>"000001001",
  64920=>"000111111",
  64921=>"000000001",
  64922=>"001001111",
  64923=>"000101000",
  64924=>"010010010",
  64925=>"001001001",
  64926=>"000000011",
  64927=>"000000000",
  64928=>"111100101",
  64929=>"111111111",
  64930=>"011000000",
  64931=>"111111111",
  64932=>"011111111",
  64933=>"001111011",
  64934=>"100000000",
  64935=>"111011111",
  64936=>"111011001",
  64937=>"110110111",
  64938=>"011011001",
  64939=>"000010010",
  64940=>"110000000",
  64941=>"000000110",
  64942=>"110010010",
  64943=>"111111111",
  64944=>"000010000",
  64945=>"000000000",
  64946=>"110111111",
  64947=>"101000000",
  64948=>"011011001",
  64949=>"111000100",
  64950=>"000000000",
  64951=>"100000010",
  64952=>"000111111",
  64953=>"001001000",
  64954=>"111111111",
  64955=>"000000001",
  64956=>"010000000",
  64957=>"000000010",
  64958=>"010000011",
  64959=>"000000000",
  64960=>"000010000",
  64961=>"010110111",
  64962=>"000000010",
  64963=>"111111111",
  64964=>"000000111",
  64965=>"000000100",
  64966=>"000000000",
  64967=>"000000001",
  64968=>"110000000",
  64969=>"111010000",
  64970=>"001110111",
  64971=>"111111111",
  64972=>"011010000",
  64973=>"001001111",
  64974=>"000001011",
  64975=>"111110111",
  64976=>"010000000",
  64977=>"000001111",
  64978=>"100111111",
  64979=>"100100100",
  64980=>"000000000",
  64981=>"110110011",
  64982=>"010110110",
  64983=>"101000100",
  64984=>"011111010",
  64985=>"111111111",
  64986=>"000110110",
  64987=>"010000000",
  64988=>"111111111",
  64989=>"111011111",
  64990=>"111111111",
  64991=>"000100000",
  64992=>"011001111",
  64993=>"010111111",
  64994=>"111111001",
  64995=>"011111110",
  64996=>"111110110",
  64997=>"111111111",
  64998=>"100100110",
  64999=>"111111000",
  65000=>"000001111",
  65001=>"001111000",
  65002=>"000000000",
  65003=>"000000001",
  65004=>"110101111",
  65005=>"111111111",
  65006=>"001000000",
  65007=>"000000111",
  65008=>"101101111",
  65009=>"100111111",
  65010=>"011010000",
  65011=>"011011011",
  65012=>"111001001",
  65013=>"100100110",
  65014=>"000000000",
  65015=>"111001001",
  65016=>"110111011",
  65017=>"111111011",
  65018=>"100110110",
  65019=>"111000000",
  65020=>"000000000",
  65021=>"010110111",
  65022=>"000011011",
  65023=>"000010011",
  65024=>"111111111",
  65025=>"100100001",
  65026=>"000000000",
  65027=>"111111111",
  65028=>"100111111",
  65029=>"000000000",
  65030=>"000000000",
  65031=>"100000000",
  65032=>"000010000",
  65033=>"000000000",
  65034=>"111111111",
  65035=>"000000100",
  65036=>"000000000",
  65037=>"100000000",
  65038=>"110111111",
  65039=>"111111111",
  65040=>"010000000",
  65041=>"000100111",
  65042=>"000000000",
  65043=>"000000000",
  65044=>"000000111",
  65045=>"000000000",
  65046=>"000000000",
  65047=>"000000001",
  65048=>"100110111",
  65049=>"000000010",
  65050=>"111000000",
  65051=>"000110001",
  65052=>"000000000",
  65053=>"000000000",
  65054=>"000000000",
  65055=>"011111111",
  65056=>"111110100",
  65057=>"111111111",
  65058=>"111011111",
  65059=>"110111111",
  65060=>"000000000",
  65061=>"011111111",
  65062=>"111111000",
  65063=>"000000000",
  65064=>"111011111",
  65065=>"111111111",
  65066=>"000000000",
  65067=>"111000000",
  65068=>"111111111",
  65069=>"110000111",
  65070=>"111001000",
  65071=>"011111111",
  65072=>"000000001",
  65073=>"000000000",
  65074=>"000000001",
  65075=>"000000000",
  65076=>"100111100",
  65077=>"111111111",
  65078=>"001000111",
  65079=>"000000000",
  65080=>"000000110",
  65081=>"000000000",
  65082=>"000000000",
  65083=>"010110110",
  65084=>"111101000",
  65085=>"000000000",
  65086=>"000000000",
  65087=>"111111111",
  65088=>"000000100",
  65089=>"000111111",
  65090=>"100100100",
  65091=>"000000000",
  65092=>"111111111",
  65093=>"111111111",
  65094=>"000000000",
  65095=>"000000001",
  65096=>"111111011",
  65097=>"111111111",
  65098=>"111111111",
  65099=>"111111111",
  65100=>"000000000",
  65101=>"000100111",
  65102=>"001000101",
  65103=>"001000000",
  65104=>"000000000",
  65105=>"001001000",
  65106=>"111111111",
  65107=>"011001100",
  65108=>"100111111",
  65109=>"000000101",
  65110=>"100000000",
  65111=>"111111111",
  65112=>"000000111",
  65113=>"111100100",
  65114=>"000100101",
  65115=>"000000000",
  65116=>"111100000",
  65117=>"111110000",
  65118=>"000011001",
  65119=>"110111111",
  65120=>"111111111",
  65121=>"000000000",
  65122=>"000000000",
  65123=>"110111111",
  65124=>"111111111",
  65125=>"000001010",
  65126=>"000000000",
  65127=>"000100101",
  65128=>"000011011",
  65129=>"111001000",
  65130=>"000000000",
  65131=>"001000000",
  65132=>"000000000",
  65133=>"111111110",
  65134=>"111111111",
  65135=>"110111111",
  65136=>"000111111",
  65137=>"001011111",
  65138=>"111111100",
  65139=>"010000000",
  65140=>"000000000",
  65141=>"111111111",
  65142=>"110100110",
  65143=>"101001111",
  65144=>"011111111",
  65145=>"110111111",
  65146=>"010000000",
  65147=>"011101011",
  65148=>"100100110",
  65149=>"111111000",
  65150=>"000000000",
  65151=>"011001000",
  65152=>"011111111",
  65153=>"001000000",
  65154=>"111110110",
  65155=>"000000000",
  65156=>"100100111",
  65157=>"111101111",
  65158=>"111111111",
  65159=>"000000000",
  65160=>"000000000",
  65161=>"111111111",
  65162=>"110011111",
  65163=>"010110100",
  65164=>"011000111",
  65165=>"111111111",
  65166=>"111111111",
  65167=>"111011000",
  65168=>"000000000",
  65169=>"111111111",
  65170=>"100100000",
  65171=>"000000000",
  65172=>"000100000",
  65173=>"000111111",
  65174=>"111111111",
  65175=>"000000111",
  65176=>"100101111",
  65177=>"111001111",
  65178=>"111011111",
  65179=>"000111110",
  65180=>"011000011",
  65181=>"100001101",
  65182=>"111111111",
  65183=>"000111011",
  65184=>"000000000",
  65185=>"100000000",
  65186=>"010011111",
  65187=>"011000111",
  65188=>"100000101",
  65189=>"111111111",
  65190=>"000000011",
  65191=>"000000000",
  65192=>"111111111",
  65193=>"000000000",
  65194=>"111111111",
  65195=>"001011011",
  65196=>"000000000",
  65197=>"000000000",
  65198=>"000000000",
  65199=>"100101001",
  65200=>"111111011",
  65201=>"111111111",
  65202=>"111111111",
  65203=>"001000000",
  65204=>"110111000",
  65205=>"111111011",
  65206=>"001011011",
  65207=>"000000000",
  65208=>"111111111",
  65209=>"111001000",
  65210=>"001001111",
  65211=>"011111011",
  65212=>"100110000",
  65213=>"111111111",
  65214=>"000000000",
  65215=>"000000000",
  65216=>"000000000",
  65217=>"000000000",
  65218=>"000000000",
  65219=>"000000000",
  65220=>"111111111",
  65221=>"000000000",
  65222=>"111111110",
  65223=>"111111111",
  65224=>"000000000",
  65225=>"111111000",
  65226=>"111111111",
  65227=>"110111111",
  65228=>"000001011",
  65229=>"000111111",
  65230=>"000000000",
  65231=>"000000000",
  65232=>"000000000",
  65233=>"000000000",
  65234=>"000000000",
  65235=>"000000000",
  65236=>"111111111",
  65237=>"110100100",
  65238=>"111110111",
  65239=>"101001101",
  65240=>"000000000",
  65241=>"000010111",
  65242=>"001000000",
  65243=>"000111111",
  65244=>"000000000",
  65245=>"000000000",
  65246=>"000000000",
  65247=>"000000000",
  65248=>"011011111",
  65249=>"001101111",
  65250=>"111111111",
  65251=>"111111111",
  65252=>"000000000",
  65253=>"110110000",
  65254=>"111111111",
  65255=>"111000000",
  65256=>"111111110",
  65257=>"111111111",
  65258=>"000000001",
  65259=>"000000100",
  65260=>"000000000",
  65261=>"001001111",
  65262=>"000000000",
  65263=>"000000100",
  65264=>"000000000",
  65265=>"000000000",
  65266=>"001111111",
  65267=>"001001000",
  65268=>"000000000",
  65269=>"111011011",
  65270=>"001011111",
  65271=>"111111111",
  65272=>"111000000",
  65273=>"000000000",
  65274=>"000000000",
  65275=>"010000000",
  65276=>"000000000",
  65277=>"000111110",
  65278=>"000110010",
  65279=>"000010111",
  65280=>"111001000",
  65281=>"000000000",
  65282=>"000000000",
  65283=>"111011001",
  65284=>"111111111",
  65285=>"011011111",
  65286=>"111111111",
  65287=>"000000111",
  65288=>"111011110",
  65289=>"100110000",
  65290=>"000000011",
  65291=>"000000000",
  65292=>"100000000",
  65293=>"000001000",
  65294=>"111111111",
  65295=>"111111111",
  65296=>"111100111",
  65297=>"111111111",
  65298=>"000000111",
  65299=>"000000000",
  65300=>"000000010",
  65301=>"111111111",
  65302=>"000000000",
  65303=>"000000000",
  65304=>"000000000",
  65305=>"010110010",
  65306=>"000110000",
  65307=>"010010001",
  65308=>"111011111",
  65309=>"111000000",
  65310=>"111011111",
  65311=>"111111111",
  65312=>"111111011",
  65313=>"100111111",
  65314=>"000000000",
  65315=>"111111111",
  65316=>"101000000",
  65317=>"111111111",
  65318=>"000000101",
  65319=>"011000111",
  65320=>"000000000",
  65321=>"000000000",
  65322=>"111000011",
  65323=>"111110000",
  65324=>"011111111",
  65325=>"000000100",
  65326=>"001000111",
  65327=>"000000001",
  65328=>"000000000",
  65329=>"000000000",
  65330=>"000000000",
  65331=>"000000000",
  65332=>"111111111",
  65333=>"111101001",
  65334=>"111111001",
  65335=>"111111111",
  65336=>"000011000",
  65337=>"111111111",
  65338=>"001001000",
  65339=>"000000000",
  65340=>"000000000",
  65341=>"000000110",
  65342=>"111000110",
  65343=>"011011011",
  65344=>"111111000",
  65345=>"100000000",
  65346=>"111011111",
  65347=>"010000010",
  65348=>"000001111",
  65349=>"111011111",
  65350=>"111111111",
  65351=>"111000000",
  65352=>"000000000",
  65353=>"000000000",
  65354=>"101111111",
  65355=>"000000000",
  65356=>"000000011",
  65357=>"111001011",
  65358=>"000000000",
  65359=>"001011111",
  65360=>"000000000",
  65361=>"000000111",
  65362=>"001000000",
  65363=>"111111111",
  65364=>"000100100",
  65365=>"011011011",
  65366=>"111111111",
  65367=>"111000000",
  65368=>"110000111",
  65369=>"000010000",
  65370=>"000000000",
  65371=>"000100110",
  65372=>"011000000",
  65373=>"000000000",
  65374=>"000000000",
  65375=>"111111111",
  65376=>"000010010",
  65377=>"011001001",
  65378=>"000000000",
  65379=>"111111111",
  65380=>"110110111",
  65381=>"111000000",
  65382=>"111111111",
  65383=>"000000001",
  65384=>"000000000",
  65385=>"111111111",
  65386=>"000000000",
  65387=>"110111111",
  65388=>"000000000",
  65389=>"111001001",
  65390=>"000000000",
  65391=>"000000000",
  65392=>"010000001",
  65393=>"010011011",
  65394=>"000000000",
  65395=>"000000111",
  65396=>"001001000",
  65397=>"000000000",
  65398=>"000000000",
  65399=>"111111111",
  65400=>"111111111",
  65401=>"111011000",
  65402=>"000000000",
  65403=>"101100000",
  65404=>"111000000",
  65405=>"000111011",
  65406=>"000110100",
  65407=>"000100111",
  65408=>"110111111",
  65409=>"111111111",
  65410=>"111111111",
  65411=>"111111111",
  65412=>"011111111",
  65413=>"000000111",
  65414=>"000000000",
  65415=>"000101111",
  65416=>"000101111",
  65417=>"011011000",
  65418=>"010011001",
  65419=>"110111010",
  65420=>"111111111",
  65421=>"000000110",
  65422=>"001001011",
  65423=>"000000011",
  65424=>"000000000",
  65425=>"000000000",
  65426=>"111111111",
  65427=>"000000000",
  65428=>"111111010",
  65429=>"000010000",
  65430=>"000000000",
  65431=>"000000000",
  65432=>"011011100",
  65433=>"111000000",
  65434=>"111111111",
  65435=>"000000010",
  65436=>"111111111",
  65437=>"000000000",
  65438=>"111111011",
  65439=>"000000000",
  65440=>"011100000",
  65441=>"000000000",
  65442=>"010000010",
  65443=>"111111111",
  65444=>"000000000",
  65445=>"000000011",
  65446=>"000000000",
  65447=>"000000000",
  65448=>"000000000",
  65449=>"000000000",
  65450=>"011000000",
  65451=>"000100111",
  65452=>"000000111",
  65453=>"001001000",
  65454=>"000111111",
  65455=>"111110110",
  65456=>"100000000",
  65457=>"111111111",
  65458=>"111111111",
  65459=>"001000110",
  65460=>"000000000",
  65461=>"111111001",
  65462=>"110111111",
  65463=>"111111110",
  65464=>"000000000",
  65465=>"110100000",
  65466=>"110000000",
  65467=>"000000010",
  65468=>"000000000",
  65469=>"000000000",
  65470=>"000101111",
  65471=>"000000000",
  65472=>"111111111",
  65473=>"000000110",
  65474=>"111111111",
  65475=>"000000000",
  65476=>"011111111",
  65477=>"001001001",
  65478=>"111111111",
  65479=>"001001001",
  65480=>"101000100",
  65481=>"011110100",
  65482=>"000000111",
  65483=>"110111111",
  65484=>"000100100",
  65485=>"110111110",
  65486=>"000000000",
  65487=>"000111111",
  65488=>"000001111",
  65489=>"000000001",
  65490=>"111111111",
  65491=>"111111111",
  65492=>"110111110",
  65493=>"000000000",
  65494=>"001111111",
  65495=>"001000001",
  65496=>"000000000",
  65497=>"000001111",
  65498=>"111111111",
  65499=>"111111111",
  65500=>"111111111",
  65501=>"101111111",
  65502=>"111111111",
  65503=>"001110000",
  65504=>"000000000",
  65505=>"111110110",
  65506=>"000000000",
  65507=>"111111001",
  65508=>"000000011",
  65509=>"111111111",
  65510=>"000000011",
  65511=>"111111111",
  65512=>"111111111",
  65513=>"111111011",
  65514=>"000100101",
  65515=>"111111111",
  65516=>"111111111",
  65517=>"000000000",
  65518=>"001000000",
  65519=>"000000011",
  65520=>"000000100",
  65521=>"110011011",
  65522=>"111000111",
  65523=>"110000000",
  65524=>"000111111",
  65525=>"010111011",
  65526=>"000000000",
  65527=>"110100000",
  65528=>"001111111",
  65529=>"000000000",
  65530=>"111111111",
  65531=>"000000000",
  65532=>"000011011",
  65533=>"111111111",
  65534=>"010001000",
  65535=>"000000000");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;