LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L8_13_WROM IS
  PORT (
    weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    address : IN unsigned(weightsbitsAddress(8)-1 DOWNTO 0));
END L8_13_WROM;

ARCHITECTURE RTL OF L8_13_WROM IS

  TYPE ROM_mem IS ARRAY (0 TO 65535) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

  CONSTANT ROM_content : ROM_mem := (0=>"100001110",
  1=>"110011110",
  2=>"100000010",
  3=>"000010000",
  4=>"000001001",
  5=>"111011110",
  6=>"111110100",
  7=>"110011111",
  8=>"111000101",
  9=>"010000010",
  10=>"010011100",
  11=>"010101011",
  12=>"100000110",
  13=>"110001000",
  14=>"001101011",
  15=>"100100000",
  16=>"001011101",
  17=>"010110010",
  18=>"101101111",
  19=>"110110100",
  20=>"010001001",
  21=>"101001101",
  22=>"101001101",
  23=>"111100001",
  24=>"001010101",
  25=>"110000011",
  26=>"101000001",
  27=>"110110110",
  28=>"010110001",
  29=>"101000110",
  30=>"010010101",
  31=>"111001110",
  32=>"001110110",
  33=>"001111010",
  34=>"000000100",
  35=>"100000101",
  36=>"110011111",
  37=>"010100100",
  38=>"001011100",
  39=>"010111011",
  40=>"110000010",
  41=>"010110000",
  42=>"000010110",
  43=>"010011000",
  44=>"001110010",
  45=>"001100001",
  46=>"100100100",
  47=>"110101000",
  48=>"100100100",
  49=>"001000111",
  50=>"110111100",
  51=>"100000001",
  52=>"010111111",
  53=>"001101110",
  54=>"110111011",
  55=>"000000101",
  56=>"001001010",
  57=>"110101110",
  58=>"010000011",
  59=>"101010100",
  60=>"100001001",
  61=>"110010001",
  62=>"111010001",
  63=>"000101101",
  64=>"101001000",
  65=>"101110000",
  66=>"010001011",
  67=>"110000000",
  68=>"100010110",
  69=>"111110100",
  70=>"100110010",
  71=>"111010000",
  72=>"011100011",
  73=>"011101111",
  74=>"100011011",
  75=>"000010000",
  76=>"010100111",
  77=>"011101100",
  78=>"110011100",
  79=>"011111111",
  80=>"000001100",
  81=>"000110000",
  82=>"100001011",
  83=>"001101100",
  84=>"101111011",
  85=>"010010100",
  86=>"010011111",
  87=>"000010101",
  88=>"100010010",
  89=>"010100111",
  90=>"101001001",
  91=>"011001111",
  92=>"010000110",
  93=>"111100000",
  94=>"010010001",
  95=>"100000100",
  96=>"110011101",
  97=>"000001111",
  98=>"010010000",
  99=>"111010010",
  100=>"010011000",
  101=>"001011011",
  102=>"111101011",
  103=>"010100000",
  104=>"110101100",
  105=>"111010011",
  106=>"010100000",
  107=>"100110010",
  108=>"101000001",
  109=>"010010010",
  110=>"001011110",
  111=>"011010110",
  112=>"110101011",
  113=>"010100010",
  114=>"111011001",
  115=>"000000010",
  116=>"110111000",
  117=>"001101011",
  118=>"011101000",
  119=>"011110101",
  120=>"111101111",
  121=>"000110110",
  122=>"111111010",
  123=>"110001100",
  124=>"111100000",
  125=>"010100000",
  126=>"011011100",
  127=>"110100100",
  128=>"011000111",
  129=>"010011000",
  130=>"101100000",
  131=>"011101011",
  132=>"100110100",
  133=>"100001101",
  134=>"101011000",
  135=>"111010101",
  136=>"001000101",
  137=>"101010001",
  138=>"010000111",
  139=>"100111111",
  140=>"011101111",
  141=>"101100011",
  142=>"100001111",
  143=>"000100000",
  144=>"110000001",
  145=>"110000101",
  146=>"010100111",
  147=>"011101111",
  148=>"101111111",
  149=>"011101011",
  150=>"011010101",
  151=>"111011101",
  152=>"011001111",
  153=>"111000010",
  154=>"110111010",
  155=>"010110110",
  156=>"110001100",
  157=>"000111110",
  158=>"000001101",
  159=>"011000111",
  160=>"001110111",
  161=>"100010101",
  162=>"010100000",
  163=>"100100000",
  164=>"100011000",
  165=>"100010110",
  166=>"111011000",
  167=>"111001011",
  168=>"111110110",
  169=>"000000011",
  170=>"000101001",
  171=>"011101101",
  172=>"001000000",
  173=>"000010010",
  174=>"011000100",
  175=>"010000111",
  176=>"110000000",
  177=>"111001101",
  178=>"111011111",
  179=>"010100010",
  180=>"001011001",
  181=>"000101001",
  182=>"101110011",
  183=>"000110000",
  184=>"011111111",
  185=>"110101010",
  186=>"110001110",
  187=>"001101000",
  188=>"100111010",
  189=>"110000000",
  190=>"011111111",
  191=>"010010110",
  192=>"101001100",
  193=>"010110001",
  194=>"000101111",
  195=>"110010111",
  196=>"001000101",
  197=>"100101001",
  198=>"010110011",
  199=>"100011000",
  200=>"000110111",
  201=>"101110000",
  202=>"101010001",
  203=>"100110100",
  204=>"101101010",
  205=>"101011101",
  206=>"000110001",
  207=>"000110100",
  208=>"110110111",
  209=>"011011011",
  210=>"110100100",
  211=>"000010111",
  212=>"001011110",
  213=>"110111100",
  214=>"110111001",
  215=>"100100001",
  216=>"101100101",
  217=>"110001001",
  218=>"010000000",
  219=>"101111010",
  220=>"100100101",
  221=>"010000111",
  222=>"111110101",
  223=>"110011101",
  224=>"000011000",
  225=>"111010101",
  226=>"001000101",
  227=>"000110110",
  228=>"101110011",
  229=>"010000101",
  230=>"011111111",
  231=>"011111001",
  232=>"111000010",
  233=>"111011111",
  234=>"101111010",
  235=>"010100001",
  236=>"110100100",
  237=>"100101110",
  238=>"011011101",
  239=>"010010000",
  240=>"110011011",
  241=>"110000010",
  242=>"110111111",
  243=>"010000011",
  244=>"101110001",
  245=>"000011000",
  246=>"111011001",
  247=>"100000010",
  248=>"110001010",
  249=>"011100111",
  250=>"010101011",
  251=>"010100010",
  252=>"000101010",
  253=>"000000001",
  254=>"110100001",
  255=>"011001010",
  256=>"001010111",
  257=>"000010001",
  258=>"111101001",
  259=>"100000110",
  260=>"010100100",
  261=>"011000010",
  262=>"000010100",
  263=>"101001001",
  264=>"001011111",
  265=>"111011001",
  266=>"001011010",
  267=>"110101101",
  268=>"001011000",
  269=>"101111111",
  270=>"100100110",
  271=>"101001101",
  272=>"011100000",
  273=>"111110100",
  274=>"011111010",
  275=>"011111100",
  276=>"100000110",
  277=>"011011000",
  278=>"110011010",
  279=>"101100000",
  280=>"000101111",
  281=>"111101110",
  282=>"101100010",
  283=>"101011011",
  284=>"000111110",
  285=>"000110000",
  286=>"100110011",
  287=>"000001111",
  288=>"110101110",
  289=>"010000100",
  290=>"000000100",
  291=>"010110100",
  292=>"001111111",
  293=>"011110111",
  294=>"001001100",
  295=>"101110101",
  296=>"001111100",
  297=>"010110111",
  298=>"100000011",
  299=>"000000001",
  300=>"110011010",
  301=>"110101111",
  302=>"010111100",
  303=>"011001011",
  304=>"101000110",
  305=>"011110011",
  306=>"000111010",
  307=>"110010001",
  308=>"000110001",
  309=>"111011101",
  310=>"010011001",
  311=>"001100010",
  312=>"000011101",
  313=>"100011001",
  314=>"011111010",
  315=>"010011100",
  316=>"111001101",
  317=>"111010110",
  318=>"111000111",
  319=>"001010100",
  320=>"110000111",
  321=>"011000011",
  322=>"100011000",
  323=>"111110011",
  324=>"010011100",
  325=>"111101010",
  326=>"110000110",
  327=>"011100001",
  328=>"011110011",
  329=>"111100000",
  330=>"110110110",
  331=>"000100011",
  332=>"010110111",
  333=>"010011001",
  334=>"110100011",
  335=>"011001110",
  336=>"111001001",
  337=>"010101010",
  338=>"001000101",
  339=>"001111111",
  340=>"101000010",
  341=>"010000000",
  342=>"100000101",
  343=>"011111110",
  344=>"101101010",
  345=>"010101101",
  346=>"101111000",
  347=>"001011010",
  348=>"000011100",
  349=>"001100111",
  350=>"000110100",
  351=>"100100011",
  352=>"100011101",
  353=>"100111000",
  354=>"100110011",
  355=>"010111011",
  356=>"110110000",
  357=>"101001011",
  358=>"011000011",
  359=>"011000101",
  360=>"101100100",
  361=>"111111011",
  362=>"001011100",
  363=>"010100100",
  364=>"101000000",
  365=>"100111011",
  366=>"011000011",
  367=>"101100001",
  368=>"101000111",
  369=>"101001010",
  370=>"000011001",
  371=>"011100111",
  372=>"111101111",
  373=>"110110110",
  374=>"110010011",
  375=>"110001111",
  376=>"100001000",
  377=>"110000110",
  378=>"111010010",
  379=>"010000010",
  380=>"001100011",
  381=>"000010011",
  382=>"001110111",
  383=>"111101110",
  384=>"011101001",
  385=>"000101110",
  386=>"101111011",
  387=>"100010100",
  388=>"101001101",
  389=>"010010100",
  390=>"101100001",
  391=>"101010101",
  392=>"100000101",
  393=>"100111000",
  394=>"110001001",
  395=>"001110100",
  396=>"010100000",
  397=>"011001001",
  398=>"110111011",
  399=>"111110011",
  400=>"100001110",
  401=>"110001101",
  402=>"001001011",
  403=>"010010011",
  404=>"000000010",
  405=>"000011101",
  406=>"101111010",
  407=>"111110001",
  408=>"010001100",
  409=>"000011010",
  410=>"111111101",
  411=>"000111000",
  412=>"110100010",
  413=>"111001000",
  414=>"110101110",
  415=>"110010100",
  416=>"011010011",
  417=>"001111001",
  418=>"111101010",
  419=>"011101110",
  420=>"101110001",
  421=>"101101100",
  422=>"001111111",
  423=>"101100110",
  424=>"111111100",
  425=>"000001101",
  426=>"000001011",
  427=>"010111011",
  428=>"000110101",
  429=>"111111000",
  430=>"000110000",
  431=>"001001110",
  432=>"110101000",
  433=>"000011100",
  434=>"011010101",
  435=>"101111010",
  436=>"100001000",
  437=>"111010001",
  438=>"000010010",
  439=>"111111001",
  440=>"111011111",
  441=>"101111110",
  442=>"001111011",
  443=>"010001101",
  444=>"101011000",
  445=>"000000001",
  446=>"001110111",
  447=>"010000010",
  448=>"000010101",
  449=>"111110010",
  450=>"111001110",
  451=>"001100111",
  452=>"001001011",
  453=>"011000011",
  454=>"111110111",
  455=>"100101001",
  456=>"010100011",
  457=>"101100001",
  458=>"110110000",
  459=>"111111010",
  460=>"000110100",
  461=>"111100101",
  462=>"010001001",
  463=>"001001101",
  464=>"111001111",
  465=>"010000011",
  466=>"011100110",
  467=>"001101111",
  468=>"111011011",
  469=>"100100000",
  470=>"110001101",
  471=>"110001010",
  472=>"101111110",
  473=>"101001000",
  474=>"000110101",
  475=>"100100010",
  476=>"001000010",
  477=>"111000001",
  478=>"000000000",
  479=>"110111110",
  480=>"001000101",
  481=>"100101011",
  482=>"001100101",
  483=>"011011011",
  484=>"111010111",
  485=>"100111100",
  486=>"100010111",
  487=>"100011000",
  488=>"101000111",
  489=>"100001010",
  490=>"110000110",
  491=>"100001001",
  492=>"001000100",
  493=>"110100010",
  494=>"111011010",
  495=>"001001110",
  496=>"011110011",
  497=>"001100000",
  498=>"000000000",
  499=>"010010110",
  500=>"011101011",
  501=>"100110011",
  502=>"011010001",
  503=>"000100110",
  504=>"111101110",
  505=>"111000011",
  506=>"000000110",
  507=>"100010010",
  508=>"000100000",
  509=>"110101111",
  510=>"100000010",
  511=>"110000100",
  512=>"000101011",
  513=>"000000111",
  514=>"010110000",
  515=>"100000000",
  516=>"000111100",
  517=>"111010110",
  518=>"011001111",
  519=>"101010110",
  520=>"000110111",
  521=>"101100011",
  522=>"011100100",
  523=>"101010010",
  524=>"110000000",
  525=>"010011111",
  526=>"000000001",
  527=>"011011101",
  528=>"001110110",
  529=>"011111010",
  530=>"010000101",
  531=>"110100110",
  532=>"101000100",
  533=>"100110000",
  534=>"101011101",
  535=>"111111110",
  536=>"011010010",
  537=>"100110100",
  538=>"001101101",
  539=>"010110100",
  540=>"001001111",
  541=>"001110011",
  542=>"011000000",
  543=>"101101011",
  544=>"001010011",
  545=>"101011111",
  546=>"010100001",
  547=>"010001011",
  548=>"100010111",
  549=>"110100100",
  550=>"010110000",
  551=>"001111100",
  552=>"010001000",
  553=>"011100000",
  554=>"111011111",
  555=>"111011001",
  556=>"000010010",
  557=>"010110011",
  558=>"010010111",
  559=>"000011000",
  560=>"001111110",
  561=>"001010110",
  562=>"001010011",
  563=>"001010000",
  564=>"101011110",
  565=>"011010001",
  566=>"011111101",
  567=>"101101000",
  568=>"000001001",
  569=>"001011100",
  570=>"110110000",
  571=>"000110111",
  572=>"101100111",
  573=>"000010110",
  574=>"001111000",
  575=>"001101110",
  576=>"101010101",
  577=>"011110011",
  578=>"010100000",
  579=>"010001110",
  580=>"100110110",
  581=>"110100110",
  582=>"111110011",
  583=>"000001111",
  584=>"010100110",
  585=>"000010101",
  586=>"011011101",
  587=>"101000111",
  588=>"101010011",
  589=>"110101010",
  590=>"100100010",
  591=>"000100000",
  592=>"110001100",
  593=>"101001010",
  594=>"101010110",
  595=>"001010011",
  596=>"001000100",
  597=>"111110100",
  598=>"111000101",
  599=>"111001010",
  600=>"110010001",
  601=>"001111110",
  602=>"110100010",
  603=>"001011101",
  604=>"100111010",
  605=>"001101111",
  606=>"001000001",
  607=>"111101011",
  608=>"100101011",
  609=>"000101000",
  610=>"000000000",
  611=>"010101010",
  612=>"101101000",
  613=>"000110001",
  614=>"100011101",
  615=>"111111101",
  616=>"011000110",
  617=>"100001100",
  618=>"000011000",
  619=>"111110101",
  620=>"100111000",
  621=>"101011010",
  622=>"101010010",
  623=>"100100110",
  624=>"011011000",
  625=>"000100000",
  626=>"111101101",
  627=>"011011101",
  628=>"111010010",
  629=>"001010001",
  630=>"001000010",
  631=>"111100010",
  632=>"001111001",
  633=>"110101100",
  634=>"111110001",
  635=>"100111110",
  636=>"110011110",
  637=>"101100101",
  638=>"111001101",
  639=>"011101101",
  640=>"111011110",
  641=>"100100101",
  642=>"011110110",
  643=>"000001001",
  644=>"000000010",
  645=>"011110000",
  646=>"000011011",
  647=>"000100110",
  648=>"010011011",
  649=>"000000011",
  650=>"001101010",
  651=>"011110000",
  652=>"100101100",
  653=>"010010110",
  654=>"110101001",
  655=>"101101010",
  656=>"011011100",
  657=>"000110111",
  658=>"111111011",
  659=>"011010000",
  660=>"100000110",
  661=>"010100001",
  662=>"000000100",
  663=>"011011100",
  664=>"001100011",
  665=>"100010111",
  666=>"010010010",
  667=>"010000010",
  668=>"100000111",
  669=>"101110010",
  670=>"110101001",
  671=>"101011000",
  672=>"111111100",
  673=>"011011010",
  674=>"010011110",
  675=>"101101100",
  676=>"011010100",
  677=>"101111111",
  678=>"001110010",
  679=>"000010000",
  680=>"010100011",
  681=>"110111011",
  682=>"100101110",
  683=>"111100101",
  684=>"010111011",
  685=>"110110100",
  686=>"011001100",
  687=>"010101001",
  688=>"100100001",
  689=>"101100111",
  690=>"111111011",
  691=>"011010100",
  692=>"101110010",
  693=>"010101111",
  694=>"110000001",
  695=>"000000000",
  696=>"100101011",
  697=>"011111001",
  698=>"001000010",
  699=>"101011111",
  700=>"011100010",
  701=>"001111110",
  702=>"100000011",
  703=>"110110110",
  704=>"100010001",
  705=>"101110010",
  706=>"101000010",
  707=>"100101110",
  708=>"011011011",
  709=>"010000101",
  710=>"000111011",
  711=>"111110101",
  712=>"101100111",
  713=>"011110011",
  714=>"111000110",
  715=>"000001010",
  716=>"111110001",
  717=>"011001111",
  718=>"011111100",
  719=>"011110000",
  720=>"000011110",
  721=>"011100001",
  722=>"100110101",
  723=>"001010100",
  724=>"110101111",
  725=>"110111010",
  726=>"010101111",
  727=>"001001001",
  728=>"010100000",
  729=>"101100000",
  730=>"010111110",
  731=>"100001100",
  732=>"100001100",
  733=>"000111011",
  734=>"101111001",
  735=>"110010110",
  736=>"000101110",
  737=>"100011011",
  738=>"110111111",
  739=>"010100110",
  740=>"110000111",
  741=>"101110111",
  742=>"111010100",
  743=>"000000111",
  744=>"110111001",
  745=>"000011101",
  746=>"101010110",
  747=>"110001100",
  748=>"000111001",
  749=>"110000011",
  750=>"101110111",
  751=>"111110010",
  752=>"010110001",
  753=>"110000011",
  754=>"111000000",
  755=>"010011111",
  756=>"111000110",
  757=>"100111100",
  758=>"010111011",
  759=>"001101010",
  760=>"001101101",
  761=>"111110001",
  762=>"010011110",
  763=>"011100100",
  764=>"000010100",
  765=>"010001100",
  766=>"001111010",
  767=>"000010001",
  768=>"111010011",
  769=>"000110100",
  770=>"011001000",
  771=>"100100001",
  772=>"111110101",
  773=>"010001010",
  774=>"101111101",
  775=>"110111000",
  776=>"001001110",
  777=>"111111010",
  778=>"111111100",
  779=>"111101101",
  780=>"010001111",
  781=>"111110011",
  782=>"111011111",
  783=>"001011000",
  784=>"101111001",
  785=>"110011001",
  786=>"111000000",
  787=>"010011000",
  788=>"011101001",
  789=>"001111110",
  790=>"101110001",
  791=>"100100100",
  792=>"110000000",
  793=>"110110111",
  794=>"110111000",
  795=>"000111011",
  796=>"110010110",
  797=>"101101100",
  798=>"101100101",
  799=>"111001101",
  800=>"010011101",
  801=>"100100101",
  802=>"101111101",
  803=>"110001101",
  804=>"101011010",
  805=>"110110100",
  806=>"000000000",
  807=>"000111111",
  808=>"000001110",
  809=>"111110110",
  810=>"010111001",
  811=>"010110000",
  812=>"100101110",
  813=>"100011111",
  814=>"000000000",
  815=>"100001000",
  816=>"011011011",
  817=>"000011100",
  818=>"111111100",
  819=>"110111001",
  820=>"010011000",
  821=>"011101011",
  822=>"010001011",
  823=>"001000010",
  824=>"010100110",
  825=>"000000011",
  826=>"001111010",
  827=>"001101110",
  828=>"100000001",
  829=>"100111000",
  830=>"101011001",
  831=>"000101100",
  832=>"101101110",
  833=>"110111000",
  834=>"111110001",
  835=>"110010101",
  836=>"100011101",
  837=>"010101100",
  838=>"101000000",
  839=>"011101000",
  840=>"011110111",
  841=>"001110010",
  842=>"011000100",
  843=>"101001000",
  844=>"011011011",
  845=>"011000001",
  846=>"001100010",
  847=>"110001010",
  848=>"010110000",
  849=>"111111111",
  850=>"100100101",
  851=>"001000111",
  852=>"010001001",
  853=>"110010101",
  854=>"010101010",
  855=>"010011101",
  856=>"111111011",
  857=>"010010101",
  858=>"111110100",
  859=>"000011111",
  860=>"110010111",
  861=>"100110001",
  862=>"000001111",
  863=>"001001000",
  864=>"111111101",
  865=>"110100001",
  866=>"100101101",
  867=>"110011001",
  868=>"100001101",
  869=>"000001011",
  870=>"001001001",
  871=>"011101010",
  872=>"100100010",
  873=>"100101001",
  874=>"011110111",
  875=>"111110011",
  876=>"100010001",
  877=>"000111011",
  878=>"000110110",
  879=>"111001101",
  880=>"000101000",
  881=>"011111010",
  882=>"100111010",
  883=>"011010100",
  884=>"000001100",
  885=>"010100011",
  886=>"011100111",
  887=>"111101010",
  888=>"010101100",
  889=>"101100011",
  890=>"100110001",
  891=>"011000100",
  892=>"111101100",
  893=>"010110110",
  894=>"011010101",
  895=>"011011100",
  896=>"101001101",
  897=>"110001101",
  898=>"010100111",
  899=>"110100111",
  900=>"011010010",
  901=>"000000101",
  902=>"100011111",
  903=>"100010101",
  904=>"010101000",
  905=>"111111001",
  906=>"111001111",
  907=>"111000110",
  908=>"101001110",
  909=>"110010101",
  910=>"111000110",
  911=>"010100001",
  912=>"100010010",
  913=>"111000111",
  914=>"100000001",
  915=>"100000001",
  916=>"101010111",
  917=>"010111010",
  918=>"100011110",
  919=>"011011011",
  920=>"000000001",
  921=>"010010100",
  922=>"111101000",
  923=>"000101000",
  924=>"111001100",
  925=>"100001110",
  926=>"100110010",
  927=>"100000000",
  928=>"111010110",
  929=>"110101101",
  930=>"111100010",
  931=>"111111000",
  932=>"100000000",
  933=>"010001110",
  934=>"001111101",
  935=>"000100101",
  936=>"011100000",
  937=>"100110001",
  938=>"010101011",
  939=>"110111010",
  940=>"010101100",
  941=>"010110010",
  942=>"110101101",
  943=>"110101100",
  944=>"000100001",
  945=>"101001000",
  946=>"000010100",
  947=>"101111111",
  948=>"011000000",
  949=>"111011100",
  950=>"101011111",
  951=>"011100111",
  952=>"110110011",
  953=>"100000000",
  954=>"111010011",
  955=>"100001110",
  956=>"110010000",
  957=>"001001111",
  958=>"111101111",
  959=>"101010000",
  960=>"100111011",
  961=>"000001000",
  962=>"111100001",
  963=>"111101010",
  964=>"101000111",
  965=>"101111010",
  966=>"001010110",
  967=>"101111111",
  968=>"000011100",
  969=>"000111011",
  970=>"000100010",
  971=>"111001101",
  972=>"011010001",
  973=>"100000110",
  974=>"000011000",
  975=>"000110111",
  976=>"000001111",
  977=>"101100000",
  978=>"000001100",
  979=>"110001100",
  980=>"011000001",
  981=>"111110100",
  982=>"011111011",
  983=>"111101100",
  984=>"111100011",
  985=>"110000001",
  986=>"001000110",
  987=>"111101101",
  988=>"111110110",
  989=>"011101101",
  990=>"101010111",
  991=>"111011110",
  992=>"101000110",
  993=>"000001011",
  994=>"111101000",
  995=>"110110100",
  996=>"011000001",
  997=>"111110010",
  998=>"110000000",
  999=>"000001010",
  1000=>"110110011",
  1001=>"111111011",
  1002=>"100111110",
  1003=>"100101011",
  1004=>"000110011",
  1005=>"111101010",
  1006=>"010000011",
  1007=>"010001001",
  1008=>"011010111",
  1009=>"010010010",
  1010=>"100000100",
  1011=>"010000101",
  1012=>"010111101",
  1013=>"011001000",
  1014=>"001110001",
  1015=>"001001011",
  1016=>"001100000",
  1017=>"101000101",
  1018=>"100010010",
  1019=>"101111000",
  1020=>"000100101",
  1021=>"111110101",
  1022=>"110100001",
  1023=>"101110110",
  1024=>"100000010",
  1025=>"010101001",
  1026=>"110001001",
  1027=>"110011101",
  1028=>"101000001",
  1029=>"111110101",
  1030=>"000001111",
  1031=>"011111010",
  1032=>"111111110",
  1033=>"100110100",
  1034=>"111001101",
  1035=>"111001011",
  1036=>"110010000",
  1037=>"110101111",
  1038=>"000001101",
  1039=>"101100101",
  1040=>"111100001",
  1041=>"011000010",
  1042=>"011010101",
  1043=>"010101000",
  1044=>"000111110",
  1045=>"101101101",
  1046=>"101101100",
  1047=>"100010101",
  1048=>"001000001",
  1049=>"101000011",
  1050=>"111010100",
  1051=>"011000101",
  1052=>"000010101",
  1053=>"001101100",
  1054=>"000000000",
  1055=>"001110000",
  1056=>"110111010",
  1057=>"011110101",
  1058=>"000111010",
  1059=>"001001000",
  1060=>"100101101",
  1061=>"111111001",
  1062=>"110111111",
  1063=>"001111001",
  1064=>"010110100",
  1065=>"000110000",
  1066=>"111101110",
  1067=>"001110110",
  1068=>"101100001",
  1069=>"000100011",
  1070=>"101011101",
  1071=>"110010101",
  1072=>"001100010",
  1073=>"000110011",
  1074=>"111111100",
  1075=>"001000100",
  1076=>"011111111",
  1077=>"110100100",
  1078=>"100100111",
  1079=>"001011101",
  1080=>"000011110",
  1081=>"100001000",
  1082=>"011100011",
  1083=>"010011101",
  1084=>"110100000",
  1085=>"010010001",
  1086=>"010001001",
  1087=>"101111101",
  1088=>"011010100",
  1089=>"001000101",
  1090=>"010000001",
  1091=>"100001011",
  1092=>"101010001",
  1093=>"110101111",
  1094=>"100111111",
  1095=>"100010010",
  1096=>"011010001",
  1097=>"111001100",
  1098=>"000000100",
  1099=>"000111011",
  1100=>"011011110",
  1101=>"100101010",
  1102=>"110101110",
  1103=>"110001001",
  1104=>"000010110",
  1105=>"111111011",
  1106=>"000100011",
  1107=>"101110111",
  1108=>"100101110",
  1109=>"111100001",
  1110=>"011010101",
  1111=>"000010000",
  1112=>"110001111",
  1113=>"100111010",
  1114=>"010110000",
  1115=>"111110111",
  1116=>"100011111",
  1117=>"001011110",
  1118=>"101111101",
  1119=>"000111000",
  1120=>"101000111",
  1121=>"001101100",
  1122=>"010001010",
  1123=>"000011000",
  1124=>"110100001",
  1125=>"001011111",
  1126=>"001110010",
  1127=>"000001111",
  1128=>"100000000",
  1129=>"000010011",
  1130=>"010111000",
  1131=>"010010001",
  1132=>"110011001",
  1133=>"100110101",
  1134=>"110010101",
  1135=>"100100011",
  1136=>"111111110",
  1137=>"101100010",
  1138=>"010011011",
  1139=>"110011000",
  1140=>"100101110",
  1141=>"101011101",
  1142=>"010101100",
  1143=>"111101011",
  1144=>"101001100",
  1145=>"101011010",
  1146=>"111010101",
  1147=>"101101100",
  1148=>"010111011",
  1149=>"100101000",
  1150=>"110010001",
  1151=>"111111001",
  1152=>"100001000",
  1153=>"110111001",
  1154=>"000001101",
  1155=>"100010011",
  1156=>"000010011",
  1157=>"110100110",
  1158=>"010011000",
  1159=>"110100010",
  1160=>"111111100",
  1161=>"000111011",
  1162=>"010011000",
  1163=>"100111101",
  1164=>"100000111",
  1165=>"000100111",
  1166=>"010111001",
  1167=>"101000101",
  1168=>"001010011",
  1169=>"000010010",
  1170=>"010011101",
  1171=>"101000011",
  1172=>"111011000",
  1173=>"010000001",
  1174=>"100110000",
  1175=>"000111001",
  1176=>"110001000",
  1177=>"010010000",
  1178=>"110111111",
  1179=>"011001111",
  1180=>"010100001",
  1181=>"100001010",
  1182=>"010100111",
  1183=>"100000100",
  1184=>"100101000",
  1185=>"011111101",
  1186=>"010100110",
  1187=>"101000000",
  1188=>"100111100",
  1189=>"101101101",
  1190=>"010111000",
  1191=>"000111010",
  1192=>"101101111",
  1193=>"101101011",
  1194=>"001110001",
  1195=>"011100001",
  1196=>"100100101",
  1197=>"101110101",
  1198=>"000011000",
  1199=>"000111111",
  1200=>"001110001",
  1201=>"011000011",
  1202=>"001001111",
  1203=>"000110110",
  1204=>"101101101",
  1205=>"101111000",
  1206=>"100011101",
  1207=>"000010100",
  1208=>"000011010",
  1209=>"001101101",
  1210=>"110010100",
  1211=>"001011101",
  1212=>"010011001",
  1213=>"000000011",
  1214=>"100110001",
  1215=>"010111011",
  1216=>"011000000",
  1217=>"011000001",
  1218=>"010001111",
  1219=>"111110110",
  1220=>"111000101",
  1221=>"100010000",
  1222=>"010110011",
  1223=>"100000101",
  1224=>"011110100",
  1225=>"110000111",
  1226=>"111010110",
  1227=>"010110010",
  1228=>"111110010",
  1229=>"011101010",
  1230=>"000011101",
  1231=>"111010100",
  1232=>"110111110",
  1233=>"011010100",
  1234=>"011011110",
  1235=>"011100111",
  1236=>"100100111",
  1237=>"101000110",
  1238=>"010101011",
  1239=>"111001100",
  1240=>"010111110",
  1241=>"001110010",
  1242=>"110101111",
  1243=>"000001001",
  1244=>"111100010",
  1245=>"001001010",
  1246=>"001010000",
  1247=>"001111010",
  1248=>"100000010",
  1249=>"100001100",
  1250=>"011011011",
  1251=>"000011110",
  1252=>"110001111",
  1253=>"010100000",
  1254=>"100011100",
  1255=>"011000101",
  1256=>"011000001",
  1257=>"101100101",
  1258=>"101101110",
  1259=>"100110111",
  1260=>"101000110",
  1261=>"011100100",
  1262=>"010011110",
  1263=>"000110010",
  1264=>"111111010",
  1265=>"011101010",
  1266=>"000011110",
  1267=>"000110010",
  1268=>"101101101",
  1269=>"100001101",
  1270=>"011010111",
  1271=>"011001000",
  1272=>"110101111",
  1273=>"101101011",
  1274=>"000000110",
  1275=>"111000010",
  1276=>"000100110",
  1277=>"000011110",
  1278=>"110111010",
  1279=>"110111000",
  1280=>"101010001",
  1281=>"001111101",
  1282=>"110111111",
  1283=>"000110100",
  1284=>"101101011",
  1285=>"000010100",
  1286=>"100010001",
  1287=>"000000111",
  1288=>"010010011",
  1289=>"100001100",
  1290=>"010011111",
  1291=>"000011011",
  1292=>"001000101",
  1293=>"000110111",
  1294=>"110001110",
  1295=>"000100110",
  1296=>"011100011",
  1297=>"001111000",
  1298=>"111000011",
  1299=>"101100100",
  1300=>"001000111",
  1301=>"011001011",
  1302=>"011101010",
  1303=>"100110111",
  1304=>"111010101",
  1305=>"000110010",
  1306=>"000000000",
  1307=>"111000010",
  1308=>"101100101",
  1309=>"101011000",
  1310=>"101111101",
  1311=>"000011101",
  1312=>"001010001",
  1313=>"000010000",
  1314=>"100100011",
  1315=>"111101011",
  1316=>"011110001",
  1317=>"010011001",
  1318=>"010111110",
  1319=>"011001101",
  1320=>"000110101",
  1321=>"000011000",
  1322=>"111001000",
  1323=>"000101000",
  1324=>"010000001",
  1325=>"010001010",
  1326=>"010011010",
  1327=>"010100000",
  1328=>"111110101",
  1329=>"101111001",
  1330=>"010010000",
  1331=>"001011111",
  1332=>"001110010",
  1333=>"100001001",
  1334=>"000010111",
  1335=>"110010100",
  1336=>"001010110",
  1337=>"101011110",
  1338=>"010101111",
  1339=>"110111100",
  1340=>"001101100",
  1341=>"110011110",
  1342=>"110001110",
  1343=>"101010100",
  1344=>"001110101",
  1345=>"111100110",
  1346=>"100000100",
  1347=>"111101101",
  1348=>"001101110",
  1349=>"111111010",
  1350=>"001000001",
  1351=>"000100101",
  1352=>"011000000",
  1353=>"001010101",
  1354=>"100001001",
  1355=>"001001101",
  1356=>"101100110",
  1357=>"110101010",
  1358=>"111101100",
  1359=>"000110100",
  1360=>"011011110",
  1361=>"011110001",
  1362=>"011010111",
  1363=>"010000001",
  1364=>"110000011",
  1365=>"000101111",
  1366=>"101100100",
  1367=>"101101001",
  1368=>"000000011",
  1369=>"000110101",
  1370=>"001100010",
  1371=>"001101000",
  1372=>"110111110",
  1373=>"000100111",
  1374=>"101001000",
  1375=>"010000011",
  1376=>"010001101",
  1377=>"011100111",
  1378=>"101100000",
  1379=>"000100000",
  1380=>"110011010",
  1381=>"010010111",
  1382=>"111011001",
  1383=>"110101111",
  1384=>"111000100",
  1385=>"000000001",
  1386=>"110100101",
  1387=>"010010001",
  1388=>"001001000",
  1389=>"000000000",
  1390=>"000000010",
  1391=>"010111101",
  1392=>"000010110",
  1393=>"000011111",
  1394=>"001000000",
  1395=>"010001000",
  1396=>"110110101",
  1397=>"101001010",
  1398=>"000110111",
  1399=>"110000010",
  1400=>"010010101",
  1401=>"100111100",
  1402=>"001111001",
  1403=>"101011000",
  1404=>"101011000",
  1405=>"001001001",
  1406=>"101100011",
  1407=>"000110010",
  1408=>"000001000",
  1409=>"111000010",
  1410=>"010011010",
  1411=>"111111001",
  1412=>"100011100",
  1413=>"010111111",
  1414=>"001111000",
  1415=>"100100010",
  1416=>"110010001",
  1417=>"101111111",
  1418=>"001000010",
  1419=>"100001101",
  1420=>"101110011",
  1421=>"001100001",
  1422=>"110011011",
  1423=>"010110100",
  1424=>"001110001",
  1425=>"000000001",
  1426=>"001000001",
  1427=>"111111110",
  1428=>"101100111",
  1429=>"000000100",
  1430=>"010000000",
  1431=>"000100000",
  1432=>"010010010",
  1433=>"010000011",
  1434=>"100010001",
  1435=>"110100001",
  1436=>"011110111",
  1437=>"110101100",
  1438=>"000011010",
  1439=>"110110110",
  1440=>"010010000",
  1441=>"001101000",
  1442=>"111100110",
  1443=>"001000001",
  1444=>"011011110",
  1445=>"110001100",
  1446=>"011110001",
  1447=>"100101111",
  1448=>"101000011",
  1449=>"111111000",
  1450=>"001000001",
  1451=>"010100111",
  1452=>"110110001",
  1453=>"110011010",
  1454=>"100000101",
  1455=>"110001110",
  1456=>"110111001",
  1457=>"101001000",
  1458=>"010001010",
  1459=>"110010001",
  1460=>"110001110",
  1461=>"101010011",
  1462=>"001110101",
  1463=>"110100101",
  1464=>"101101001",
  1465=>"000010000",
  1466=>"000111000",
  1467=>"110101001",
  1468=>"111000000",
  1469=>"111001011",
  1470=>"000010001",
  1471=>"111010011",
  1472=>"101101000",
  1473=>"010110101",
  1474=>"000101100",
  1475=>"110001000",
  1476=>"000110110",
  1477=>"110000100",
  1478=>"100011110",
  1479=>"100000000",
  1480=>"011110100",
  1481=>"001000100",
  1482=>"100110000",
  1483=>"000010001",
  1484=>"100110001",
  1485=>"010100010",
  1486=>"111001011",
  1487=>"111110100",
  1488=>"110100111",
  1489=>"000000001",
  1490=>"110000011",
  1491=>"110111011",
  1492=>"001000111",
  1493=>"010110101",
  1494=>"111100101",
  1495=>"101011010",
  1496=>"110100001",
  1497=>"000001110",
  1498=>"011101110",
  1499=>"010101110",
  1500=>"010100001",
  1501=>"111000010",
  1502=>"100011000",
  1503=>"011011101",
  1504=>"000001110",
  1505=>"111010011",
  1506=>"010001011",
  1507=>"000100111",
  1508=>"101100111",
  1509=>"001100000",
  1510=>"110111110",
  1511=>"110000001",
  1512=>"001101100",
  1513=>"100001110",
  1514=>"000101101",
  1515=>"010110100",
  1516=>"001000100",
  1517=>"101010001",
  1518=>"100101101",
  1519=>"010100010",
  1520=>"011110100",
  1521=>"111001100",
  1522=>"011111001",
  1523=>"011110000",
  1524=>"110101000",
  1525=>"010100011",
  1526=>"100100011",
  1527=>"100010010",
  1528=>"001010000",
  1529=>"101001111",
  1530=>"011110000",
  1531=>"011110001",
  1532=>"000001110",
  1533=>"001001000",
  1534=>"100111001",
  1535=>"000101001",
  1536=>"011000011",
  1537=>"111101000",
  1538=>"110101111",
  1539=>"110110001",
  1540=>"000101011",
  1541=>"000010111",
  1542=>"100011100",
  1543=>"100001001",
  1544=>"110110000",
  1545=>"110011101",
  1546=>"010101000",
  1547=>"110110111",
  1548=>"111011110",
  1549=>"000011011",
  1550=>"101000100",
  1551=>"101001001",
  1552=>"010001101",
  1553=>"001100101",
  1554=>"111111101",
  1555=>"111010101",
  1556=>"011000010",
  1557=>"001010000",
  1558=>"011010110",
  1559=>"101010110",
  1560=>"010000100",
  1561=>"111101010",
  1562=>"101010111",
  1563=>"111111100",
  1564=>"011111000",
  1565=>"011011010",
  1566=>"110010011",
  1567=>"000010001",
  1568=>"100110011",
  1569=>"101000010",
  1570=>"010011001",
  1571=>"001010110",
  1572=>"100011011",
  1573=>"001100000",
  1574=>"011101011",
  1575=>"101110000",
  1576=>"110100000",
  1577=>"111011010",
  1578=>"111001011",
  1579=>"000001001",
  1580=>"000101101",
  1581=>"010111001",
  1582=>"011110000",
  1583=>"100111101",
  1584=>"100011000",
  1585=>"010010010",
  1586=>"011111100",
  1587=>"111100101",
  1588=>"000011111",
  1589=>"110000000",
  1590=>"011111100",
  1591=>"011111001",
  1592=>"100010100",
  1593=>"010001100",
  1594=>"100100001",
  1595=>"000100110",
  1596=>"000000111",
  1597=>"001010010",
  1598=>"100001011",
  1599=>"110011101",
  1600=>"111011011",
  1601=>"000100100",
  1602=>"101010000",
  1603=>"101100011",
  1604=>"001110001",
  1605=>"100010110",
  1606=>"010011000",
  1607=>"001010011",
  1608=>"111001100",
  1609=>"100110001",
  1610=>"100010000",
  1611=>"010100111",
  1612=>"100010010",
  1613=>"010010010",
  1614=>"000001100",
  1615=>"011010010",
  1616=>"001011101",
  1617=>"101101110",
  1618=>"110000101",
  1619=>"101101111",
  1620=>"100011000",
  1621=>"000001101",
  1622=>"000100100",
  1623=>"010111100",
  1624=>"111111110",
  1625=>"111111111",
  1626=>"101001000",
  1627=>"111111010",
  1628=>"000011100",
  1629=>"001100000",
  1630=>"010110000",
  1631=>"001100011",
  1632=>"101011110",
  1633=>"000100001",
  1634=>"110101110",
  1635=>"101000001",
  1636=>"000010100",
  1637=>"111110110",
  1638=>"000000000",
  1639=>"110111000",
  1640=>"000110010",
  1641=>"010001011",
  1642=>"000101011",
  1643=>"011001001",
  1644=>"000010111",
  1645=>"101111111",
  1646=>"111101110",
  1647=>"110001010",
  1648=>"010011001",
  1649=>"001000001",
  1650=>"000010101",
  1651=>"000101011",
  1652=>"100010111",
  1653=>"000000110",
  1654=>"010101000",
  1655=>"011000001",
  1656=>"111100011",
  1657=>"101111111",
  1658=>"000110111",
  1659=>"101011011",
  1660=>"011000101",
  1661=>"001011010",
  1662=>"101001100",
  1663=>"000000011",
  1664=>"001100010",
  1665=>"100111101",
  1666=>"110000111",
  1667=>"000011100",
  1668=>"110010111",
  1669=>"111001001",
  1670=>"111010101",
  1671=>"111101101",
  1672=>"111110110",
  1673=>"000011100",
  1674=>"001010101",
  1675=>"000100011",
  1676=>"000111110",
  1677=>"111011110",
  1678=>"011110100",
  1679=>"110000110",
  1680=>"010101011",
  1681=>"001100110",
  1682=>"111100011",
  1683=>"000101111",
  1684=>"010000011",
  1685=>"101100001",
  1686=>"101111000",
  1687=>"010010100",
  1688=>"011101111",
  1689=>"111111001",
  1690=>"000000100",
  1691=>"100101111",
  1692=>"111101110",
  1693=>"011110100",
  1694=>"011011111",
  1695=>"101111011",
  1696=>"001010110",
  1697=>"000111110",
  1698=>"010011111",
  1699=>"101101001",
  1700=>"100101010",
  1701=>"010101001",
  1702=>"001011000",
  1703=>"000001000",
  1704=>"000011001",
  1705=>"010000001",
  1706=>"010011010",
  1707=>"000011001",
  1708=>"001001010",
  1709=>"101100101",
  1710=>"111100001",
  1711=>"100000001",
  1712=>"011001110",
  1713=>"011010100",
  1714=>"001001110",
  1715=>"000000011",
  1716=>"010010111",
  1717=>"100001111",
  1718=>"111101001",
  1719=>"000110011",
  1720=>"101100101",
  1721=>"100010000",
  1722=>"111111111",
  1723=>"110110000",
  1724=>"101010111",
  1725=>"110111011",
  1726=>"001101001",
  1727=>"100101101",
  1728=>"100101111",
  1729=>"000111100",
  1730=>"110000111",
  1731=>"001100110",
  1732=>"100111100",
  1733=>"000110101",
  1734=>"010101101",
  1735=>"100011000",
  1736=>"111001001",
  1737=>"001111001",
  1738=>"011011100",
  1739=>"000000011",
  1740=>"100000001",
  1741=>"101011010",
  1742=>"001111000",
  1743=>"001001010",
  1744=>"110001000",
  1745=>"110010111",
  1746=>"110010101",
  1747=>"000001010",
  1748=>"111010110",
  1749=>"011010010",
  1750=>"011010101",
  1751=>"111111111",
  1752=>"111101000",
  1753=>"000001011",
  1754=>"111011100",
  1755=>"001000000",
  1756=>"111110101",
  1757=>"000010111",
  1758=>"110101001",
  1759=>"111101100",
  1760=>"111001001",
  1761=>"000010000",
  1762=>"011100101",
  1763=>"010111010",
  1764=>"000111000",
  1765=>"010110010",
  1766=>"000000100",
  1767=>"010110100",
  1768=>"010101101",
  1769=>"010011100",
  1770=>"000010000",
  1771=>"111111101",
  1772=>"001001010",
  1773=>"001011001",
  1774=>"001100111",
  1775=>"010100111",
  1776=>"100001011",
  1777=>"010100100",
  1778=>"100100000",
  1779=>"111011111",
  1780=>"001100110",
  1781=>"111010001",
  1782=>"110101110",
  1783=>"000000101",
  1784=>"110011010",
  1785=>"011110110",
  1786=>"101011010",
  1787=>"101000010",
  1788=>"011011011",
  1789=>"010000010",
  1790=>"101100011",
  1791=>"101011100",
  1792=>"100000001",
  1793=>"000001000",
  1794=>"111010111",
  1795=>"011101011",
  1796=>"000110000",
  1797=>"001001010",
  1798=>"010100111",
  1799=>"101001001",
  1800=>"101100111",
  1801=>"000111100",
  1802=>"111001100",
  1803=>"100010111",
  1804=>"010111001",
  1805=>"000011000",
  1806=>"000001011",
  1807=>"111100101",
  1808=>"100000000",
  1809=>"001001110",
  1810=>"000010100",
  1811=>"100100001",
  1812=>"111110011",
  1813=>"000110000",
  1814=>"011011010",
  1815=>"010101000",
  1816=>"100001111",
  1817=>"001011101",
  1818=>"111111101",
  1819=>"111010010",
  1820=>"000100100",
  1821=>"111010100",
  1822=>"001011010",
  1823=>"001101000",
  1824=>"000010101",
  1825=>"000101011",
  1826=>"010111000",
  1827=>"000011010",
  1828=>"110101110",
  1829=>"001111000",
  1830=>"010011110",
  1831=>"110001111",
  1832=>"000011010",
  1833=>"111010100",
  1834=>"000010110",
  1835=>"110111001",
  1836=>"111011110",
  1837=>"001011101",
  1838=>"001110000",
  1839=>"001100000",
  1840=>"100000010",
  1841=>"110110000",
  1842=>"000100001",
  1843=>"010111100",
  1844=>"100100010",
  1845=>"110101000",
  1846=>"100010100",
  1847=>"000011000",
  1848=>"110001100",
  1849=>"000001010",
  1850=>"111111001",
  1851=>"110001000",
  1852=>"010101100",
  1853=>"010101001",
  1854=>"001100101",
  1855=>"100100010",
  1856=>"001111110",
  1857=>"100001001",
  1858=>"101110011",
  1859=>"100011011",
  1860=>"100110101",
  1861=>"101000000",
  1862=>"111000100",
  1863=>"000110010",
  1864=>"110101110",
  1865=>"110111111",
  1866=>"001000000",
  1867=>"011010101",
  1868=>"100110011",
  1869=>"100100001",
  1870=>"100100001",
  1871=>"100010110",
  1872=>"100000110",
  1873=>"001011101",
  1874=>"110111110",
  1875=>"001100111",
  1876=>"000011010",
  1877=>"111111110",
  1878=>"011000000",
  1879=>"001010001",
  1880=>"101000010",
  1881=>"010100111",
  1882=>"110000101",
  1883=>"011111110",
  1884=>"101010111",
  1885=>"000111100",
  1886=>"000101110",
  1887=>"000110110",
  1888=>"000100000",
  1889=>"101101001",
  1890=>"000001000",
  1891=>"000001100",
  1892=>"100001100",
  1893=>"001011100",
  1894=>"111110100",
  1895=>"101110010",
  1896=>"000010010",
  1897=>"111000011",
  1898=>"000100000",
  1899=>"010111000",
  1900=>"000101110",
  1901=>"111100010",
  1902=>"111100111",
  1903=>"010001111",
  1904=>"010000000",
  1905=>"111001110",
  1906=>"111111101",
  1907=>"011000001",
  1908=>"000101100",
  1909=>"100100110",
  1910=>"100100110",
  1911=>"001010000",
  1912=>"010101000",
  1913=>"100101110",
  1914=>"000110011",
  1915=>"101000111",
  1916=>"101010100",
  1917=>"011000010",
  1918=>"100101000",
  1919=>"111011001",
  1920=>"111100110",
  1921=>"000001101",
  1922=>"010111110",
  1923=>"001000001",
  1924=>"010000000",
  1925=>"101010000",
  1926=>"000111110",
  1927=>"000100000",
  1928=>"101111000",
  1929=>"101011100",
  1930=>"000001000",
  1931=>"110000000",
  1932=>"011100010",
  1933=>"001101100",
  1934=>"100100000",
  1935=>"111010101",
  1936=>"011011101",
  1937=>"101111101",
  1938=>"000101111",
  1939=>"001000011",
  1940=>"010010111",
  1941=>"010111111",
  1942=>"100000100",
  1943=>"101101110",
  1944=>"101000000",
  1945=>"011001010",
  1946=>"101101100",
  1947=>"001000000",
  1948=>"111100001",
  1949=>"000001001",
  1950=>"011011000",
  1951=>"100000110",
  1952=>"011010000",
  1953=>"001110110",
  1954=>"101100001",
  1955=>"000100001",
  1956=>"000000001",
  1957=>"101110000",
  1958=>"111011010",
  1959=>"000010010",
  1960=>"111110110",
  1961=>"111010100",
  1962=>"111000001",
  1963=>"111110000",
  1964=>"101111100",
  1965=>"110111110",
  1966=>"101110010",
  1967=>"110010010",
  1968=>"100110010",
  1969=>"001000111",
  1970=>"010011111",
  1971=>"010010101",
  1972=>"001011111",
  1973=>"100110100",
  1974=>"111011101",
  1975=>"110011010",
  1976=>"111010000",
  1977=>"100111000",
  1978=>"111101110",
  1979=>"010000001",
  1980=>"000010000",
  1981=>"011100000",
  1982=>"101010111",
  1983=>"111000111",
  1984=>"000111011",
  1985=>"011011010",
  1986=>"101111000",
  1987=>"000000010",
  1988=>"001100111",
  1989=>"011111011",
  1990=>"111101010",
  1991=>"100010111",
  1992=>"000101010",
  1993=>"111001000",
  1994=>"011010011",
  1995=>"010110001",
  1996=>"110011010",
  1997=>"001000000",
  1998=>"011000001",
  1999=>"100101000",
  2000=>"110111101",
  2001=>"000101101",
  2002=>"110110100",
  2003=>"101000111",
  2004=>"100011101",
  2005=>"000000011",
  2006=>"110101000",
  2007=>"101101011",
  2008=>"100111011",
  2009=>"000010011",
  2010=>"000011111",
  2011=>"111001001",
  2012=>"111111111",
  2013=>"101100101",
  2014=>"100101000",
  2015=>"001100011",
  2016=>"001111101",
  2017=>"111010000",
  2018=>"111101011",
  2019=>"100111101",
  2020=>"011000010",
  2021=>"011001101",
  2022=>"000011100",
  2023=>"000111100",
  2024=>"000010010",
  2025=>"011001111",
  2026=>"000010000",
  2027=>"110101110",
  2028=>"010100101",
  2029=>"010101111",
  2030=>"000111111",
  2031=>"111101011",
  2032=>"101011100",
  2033=>"011011000",
  2034=>"000011011",
  2035=>"101001000",
  2036=>"101011010",
  2037=>"101000100",
  2038=>"111111100",
  2039=>"111000110",
  2040=>"010110101",
  2041=>"101111110",
  2042=>"100100100",
  2043=>"011001001",
  2044=>"110010110",
  2045=>"001010110",
  2046=>"010110011",
  2047=>"101111110",
  2048=>"010001011",
  2049=>"101110000",
  2050=>"110000100",
  2051=>"100011011",
  2052=>"110101101",
  2053=>"111101101",
  2054=>"100110010",
  2055=>"111101000",
  2056=>"110001011",
  2057=>"001000001",
  2058=>"101010110",
  2059=>"010110100",
  2060=>"110010000",
  2061=>"110101000",
  2062=>"100110001",
  2063=>"000111100",
  2064=>"000111100",
  2065=>"111101011",
  2066=>"001100000",
  2067=>"111111010",
  2068=>"000011110",
  2069=>"100000001",
  2070=>"101110010",
  2071=>"110101000",
  2072=>"000001111",
  2073=>"101011101",
  2074=>"010100100",
  2075=>"111100011",
  2076=>"110000110",
  2077=>"101110001",
  2078=>"000101110",
  2079=>"111011011",
  2080=>"111111011",
  2081=>"001011000",
  2082=>"000010100",
  2083=>"000000111",
  2084=>"101101110",
  2085=>"111111101",
  2086=>"101010000",
  2087=>"010110111",
  2088=>"100010110",
  2089=>"001001110",
  2090=>"000100100",
  2091=>"011101011",
  2092=>"011000101",
  2093=>"000100011",
  2094=>"011111010",
  2095=>"100011010",
  2096=>"110001100",
  2097=>"100111111",
  2098=>"000001100",
  2099=>"110111111",
  2100=>"100101111",
  2101=>"100010110",
  2102=>"001110100",
  2103=>"100110010",
  2104=>"101100011",
  2105=>"001011101",
  2106=>"011010011",
  2107=>"010001011",
  2108=>"111000101",
  2109=>"010000101",
  2110=>"010110001",
  2111=>"010101010",
  2112=>"000110100",
  2113=>"010101111",
  2114=>"001101011",
  2115=>"000011011",
  2116=>"110111011",
  2117=>"011111001",
  2118=>"011011010",
  2119=>"110101001",
  2120=>"110111000",
  2121=>"001100100",
  2122=>"010011001",
  2123=>"010101000",
  2124=>"100000100",
  2125=>"010110100",
  2126=>"111110011",
  2127=>"111011110",
  2128=>"010000011",
  2129=>"100101101",
  2130=>"101101000",
  2131=>"011100011",
  2132=>"010000000",
  2133=>"011101000",
  2134=>"100010111",
  2135=>"010011111",
  2136=>"111110111",
  2137=>"101101000",
  2138=>"101011010",
  2139=>"001101100",
  2140=>"011000010",
  2141=>"010000100",
  2142=>"110010110",
  2143=>"011111100",
  2144=>"101110001",
  2145=>"101011000",
  2146=>"110001011",
  2147=>"111100011",
  2148=>"100011010",
  2149=>"100010001",
  2150=>"101000000",
  2151=>"010010010",
  2152=>"111111110",
  2153=>"011110001",
  2154=>"101011010",
  2155=>"110000111",
  2156=>"001110110",
  2157=>"100111110",
  2158=>"001100110",
  2159=>"010101011",
  2160=>"000111111",
  2161=>"010001010",
  2162=>"111010010",
  2163=>"100110111",
  2164=>"011111001",
  2165=>"010000101",
  2166=>"001100001",
  2167=>"011100101",
  2168=>"010111001",
  2169=>"000001000",
  2170=>"000000101",
  2171=>"110111111",
  2172=>"111110100",
  2173=>"100101000",
  2174=>"101011011",
  2175=>"001100110",
  2176=>"110011101",
  2177=>"111101000",
  2178=>"110011111",
  2179=>"001101110",
  2180=>"001001101",
  2181=>"110101101",
  2182=>"101110001",
  2183=>"011100110",
  2184=>"011011011",
  2185=>"000000011",
  2186=>"101001110",
  2187=>"111010111",
  2188=>"011000000",
  2189=>"111101000",
  2190=>"000001100",
  2191=>"011011111",
  2192=>"100111110",
  2193=>"111111000",
  2194=>"100001101",
  2195=>"101111011",
  2196=>"010001001",
  2197=>"101011100",
  2198=>"011011111",
  2199=>"100010100",
  2200=>"111011001",
  2201=>"010000100",
  2202=>"000001100",
  2203=>"001000111",
  2204=>"110001000",
  2205=>"010100110",
  2206=>"110011101",
  2207=>"010110110",
  2208=>"111110000",
  2209=>"100011111",
  2210=>"011111110",
  2211=>"110001101",
  2212=>"010100110",
  2213=>"110111011",
  2214=>"111110111",
  2215=>"101000101",
  2216=>"111010000",
  2217=>"101110010",
  2218=>"011010101",
  2219=>"011111111",
  2220=>"010011001",
  2221=>"101110110",
  2222=>"100100001",
  2223=>"011011001",
  2224=>"100011011",
  2225=>"111000000",
  2226=>"010010001",
  2227=>"101000101",
  2228=>"111101111",
  2229=>"111000001",
  2230=>"101000010",
  2231=>"000011110",
  2232=>"110010110",
  2233=>"001000010",
  2234=>"110000010",
  2235=>"000001010",
  2236=>"000101011",
  2237=>"001110111",
  2238=>"001000000",
  2239=>"110101011",
  2240=>"000010000",
  2241=>"100100010",
  2242=>"011111111",
  2243=>"000100001",
  2244=>"110111111",
  2245=>"011010110",
  2246=>"000110110",
  2247=>"001111010",
  2248=>"111010000",
  2249=>"001100110",
  2250=>"101000001",
  2251=>"110100011",
  2252=>"101100110",
  2253=>"000001010",
  2254=>"011011100",
  2255=>"111100101",
  2256=>"100111000",
  2257=>"100010101",
  2258=>"010001000",
  2259=>"101110011",
  2260=>"011110110",
  2261=>"000010001",
  2262=>"010100001",
  2263=>"011110001",
  2264=>"100111111",
  2265=>"000100011",
  2266=>"011001110",
  2267=>"001110011",
  2268=>"011111000",
  2269=>"011111101",
  2270=>"001001001",
  2271=>"101100001",
  2272=>"010111101",
  2273=>"010000000",
  2274=>"000011100",
  2275=>"111011101",
  2276=>"110101111",
  2277=>"011111000",
  2278=>"111101010",
  2279=>"010110110",
  2280=>"110001101",
  2281=>"001001001",
  2282=>"111011010",
  2283=>"010001111",
  2284=>"001010000",
  2285=>"100101101",
  2286=>"001000111",
  2287=>"000000010",
  2288=>"000111110",
  2289=>"101101010",
  2290=>"101010001",
  2291=>"001011101",
  2292=>"100111001",
  2293=>"011100110",
  2294=>"001101110",
  2295=>"001001000",
  2296=>"001100101",
  2297=>"001100101",
  2298=>"010000110",
  2299=>"001101101",
  2300=>"011010110",
  2301=>"010110111",
  2302=>"111101000",
  2303=>"111100100",
  2304=>"101100010",
  2305=>"110001110",
  2306=>"110011011",
  2307=>"010000000",
  2308=>"111101101",
  2309=>"101111100",
  2310=>"100111111",
  2311=>"100000001",
  2312=>"110010000",
  2313=>"110010001",
  2314=>"101000000",
  2315=>"101111011",
  2316=>"000000101",
  2317=>"000000110",
  2318=>"001101101",
  2319=>"001000000",
  2320=>"010000101",
  2321=>"110000111",
  2322=>"110010111",
  2323=>"100010010",
  2324=>"101100111",
  2325=>"010001001",
  2326=>"000001100",
  2327=>"110101111",
  2328=>"111001000",
  2329=>"000110100",
  2330=>"010010100",
  2331=>"010010010",
  2332=>"000011100",
  2333=>"010000011",
  2334=>"010110010",
  2335=>"111110001",
  2336=>"101101110",
  2337=>"100101101",
  2338=>"000011001",
  2339=>"110111001",
  2340=>"101110010",
  2341=>"011111001",
  2342=>"000011000",
  2343=>"111111101",
  2344=>"100001001",
  2345=>"111101111",
  2346=>"010100000",
  2347=>"001101110",
  2348=>"101000110",
  2349=>"111000010",
  2350=>"111011111",
  2351=>"000001100",
  2352=>"000011000",
  2353=>"011100010",
  2354=>"111000101",
  2355=>"110101011",
  2356=>"011011000",
  2357=>"011100000",
  2358=>"001110011",
  2359=>"010111111",
  2360=>"010000000",
  2361=>"101001110",
  2362=>"001101110",
  2363=>"100011000",
  2364=>"000000010",
  2365=>"000110100",
  2366=>"010000000",
  2367=>"111100011",
  2368=>"100101111",
  2369=>"001001000",
  2370=>"111001010",
  2371=>"011000001",
  2372=>"011110111",
  2373=>"001000000",
  2374=>"101111100",
  2375=>"000111011",
  2376=>"000101111",
  2377=>"111111110",
  2378=>"111111101",
  2379=>"000001011",
  2380=>"011101100",
  2381=>"000111000",
  2382=>"011000000",
  2383=>"110101010",
  2384=>"010000111",
  2385=>"100101010",
  2386=>"101001101",
  2387=>"001110010",
  2388=>"110101110",
  2389=>"101100100",
  2390=>"001010100",
  2391=>"001000110",
  2392=>"000000001",
  2393=>"110000111",
  2394=>"000001001",
  2395=>"111000011",
  2396=>"001111011",
  2397=>"010011001",
  2398=>"010111110",
  2399=>"001101001",
  2400=>"111111111",
  2401=>"001000001",
  2402=>"111110010",
  2403=>"011110100",
  2404=>"001000000",
  2405=>"010010000",
  2406=>"101011010",
  2407=>"000000010",
  2408=>"001100010",
  2409=>"011000001",
  2410=>"111111100",
  2411=>"010010001",
  2412=>"110111000",
  2413=>"001110011",
  2414=>"001110100",
  2415=>"001110000",
  2416=>"110011101",
  2417=>"010101000",
  2418=>"110111111",
  2419=>"011010111",
  2420=>"110010110",
  2421=>"001010110",
  2422=>"111010110",
  2423=>"011101011",
  2424=>"000010001",
  2425=>"100111011",
  2426=>"111110111",
  2427=>"011101011",
  2428=>"101011101",
  2429=>"100010001",
  2430=>"001000101",
  2431=>"111001011",
  2432=>"011101110",
  2433=>"011101000",
  2434=>"101100011",
  2435=>"011010111",
  2436=>"000001001",
  2437=>"010011110",
  2438=>"001101111",
  2439=>"000101110",
  2440=>"101101111",
  2441=>"110110111",
  2442=>"010001101",
  2443=>"111100100",
  2444=>"110111000",
  2445=>"001000011",
  2446=>"100110111",
  2447=>"111001000",
  2448=>"100010110",
  2449=>"111100110",
  2450=>"100001100",
  2451=>"111111000",
  2452=>"100010100",
  2453=>"111001010",
  2454=>"011001000",
  2455=>"101001100",
  2456=>"100010101",
  2457=>"011000101",
  2458=>"011110001",
  2459=>"110001100",
  2460=>"011000100",
  2461=>"010001011",
  2462=>"101110100",
  2463=>"110001100",
  2464=>"001100100",
  2465=>"110000010",
  2466=>"110100011",
  2467=>"001001100",
  2468=>"011011100",
  2469=>"110011111",
  2470=>"111010010",
  2471=>"111011100",
  2472=>"111111110",
  2473=>"101011001",
  2474=>"001000000",
  2475=>"100011110",
  2476=>"110100110",
  2477=>"011101010",
  2478=>"000011110",
  2479=>"110001011",
  2480=>"110110000",
  2481=>"000010001",
  2482=>"011011111",
  2483=>"010101001",
  2484=>"100100000",
  2485=>"011111000",
  2486=>"100001010",
  2487=>"011101100",
  2488=>"111100110",
  2489=>"011110100",
  2490=>"101001101",
  2491=>"110101101",
  2492=>"110010110",
  2493=>"000011011",
  2494=>"110101000",
  2495=>"110110011",
  2496=>"100110100",
  2497=>"100101110",
  2498=>"010011000",
  2499=>"011110101",
  2500=>"001111011",
  2501=>"111101011",
  2502=>"100000101",
  2503=>"000010000",
  2504=>"001001001",
  2505=>"000101101",
  2506=>"101101110",
  2507=>"100011101",
  2508=>"000110001",
  2509=>"101111010",
  2510=>"101101100",
  2511=>"010001000",
  2512=>"101001101",
  2513=>"110000000",
  2514=>"111011000",
  2515=>"000100001",
  2516=>"001100011",
  2517=>"101010000",
  2518=>"100110000",
  2519=>"101000000",
  2520=>"100110010",
  2521=>"110011110",
  2522=>"010010001",
  2523=>"001001111",
  2524=>"000000010",
  2525=>"010110111",
  2526=>"011100010",
  2527=>"000101010",
  2528=>"001100101",
  2529=>"100101001",
  2530=>"111011001",
  2531=>"000001100",
  2532=>"000010111",
  2533=>"111000101",
  2534=>"111001101",
  2535=>"000111111",
  2536=>"010101110",
  2537=>"101111000",
  2538=>"101111101",
  2539=>"010000000",
  2540=>"001000001",
  2541=>"000000111",
  2542=>"111011111",
  2543=>"110011000",
  2544=>"011000000",
  2545=>"100110001",
  2546=>"000001000",
  2547=>"101001111",
  2548=>"111000001",
  2549=>"010010010",
  2550=>"011110101",
  2551=>"011111100",
  2552=>"100001100",
  2553=>"000101001",
  2554=>"011111101",
  2555=>"010100000",
  2556=>"101000000",
  2557=>"001010111",
  2558=>"110000111",
  2559=>"010100001",
  2560=>"000101011",
  2561=>"010000111",
  2562=>"110111100",
  2563=>"001001000",
  2564=>"101010101",
  2565=>"110000011",
  2566=>"010011100",
  2567=>"100001000",
  2568=>"101010111",
  2569=>"110100100",
  2570=>"000111001",
  2571=>"100011001",
  2572=>"011011100",
  2573=>"110001001",
  2574=>"001011100",
  2575=>"011100101",
  2576=>"110110010",
  2577=>"101001111",
  2578=>"100001111",
  2579=>"100101011",
  2580=>"010001011",
  2581=>"101011001",
  2582=>"001011001",
  2583=>"000010101",
  2584=>"001101000",
  2585=>"011000010",
  2586=>"001010111",
  2587=>"000000000",
  2588=>"001101001",
  2589=>"110111011",
  2590=>"111001001",
  2591=>"111110101",
  2592=>"011010001",
  2593=>"011100111",
  2594=>"001110111",
  2595=>"000010111",
  2596=>"000000101",
  2597=>"010111011",
  2598=>"111111011",
  2599=>"000010111",
  2600=>"111011111",
  2601=>"010111001",
  2602=>"100011000",
  2603=>"010001111",
  2604=>"100010111",
  2605=>"000101000",
  2606=>"101010110",
  2607=>"010100010",
  2608=>"001000101",
  2609=>"101000010",
  2610=>"111101100",
  2611=>"001111100",
  2612=>"001111110",
  2613=>"111111000",
  2614=>"001110110",
  2615=>"101101010",
  2616=>"000100001",
  2617=>"110101000",
  2618=>"110000101",
  2619=>"111100011",
  2620=>"011111111",
  2621=>"111101001",
  2622=>"101010011",
  2623=>"110011100",
  2624=>"000011111",
  2625=>"110011010",
  2626=>"101011011",
  2627=>"010110100",
  2628=>"111111110",
  2629=>"111010011",
  2630=>"000000000",
  2631=>"110101111",
  2632=>"000100111",
  2633=>"111111110",
  2634=>"001011010",
  2635=>"011100101",
  2636=>"110011110",
  2637=>"011010000",
  2638=>"001001000",
  2639=>"110001110",
  2640=>"010001011",
  2641=>"011010001",
  2642=>"001011010",
  2643=>"100011001",
  2644=>"000100110",
  2645=>"100000000",
  2646=>"100100110",
  2647=>"110110010",
  2648=>"111110111",
  2649=>"101100101",
  2650=>"000010101",
  2651=>"001010000",
  2652=>"010001000",
  2653=>"011101000",
  2654=>"001000100",
  2655=>"110111100",
  2656=>"100010100",
  2657=>"010011011",
  2658=>"010001110",
  2659=>"110110111",
  2660=>"000001100",
  2661=>"101100111",
  2662=>"111101010",
  2663=>"011010110",
  2664=>"111111110",
  2665=>"101110011",
  2666=>"010010101",
  2667=>"011000000",
  2668=>"111011011",
  2669=>"100000101",
  2670=>"101101000",
  2671=>"011011110",
  2672=>"111101000",
  2673=>"010110111",
  2674=>"110011101",
  2675=>"011000001",
  2676=>"000010111",
  2677=>"011101101",
  2678=>"100010001",
  2679=>"111000111",
  2680=>"111010101",
  2681=>"101000001",
  2682=>"110101010",
  2683=>"001010100",
  2684=>"110010001",
  2685=>"101010000",
  2686=>"011100100",
  2687=>"000000011",
  2688=>"100010000",
  2689=>"010100100",
  2690=>"111110010",
  2691=>"001001000",
  2692=>"111001110",
  2693=>"011000001",
  2694=>"011101011",
  2695=>"100000000",
  2696=>"001000111",
  2697=>"110101010",
  2698=>"001011110",
  2699=>"110011101",
  2700=>"100100110",
  2701=>"111111110",
  2702=>"101101101",
  2703=>"001000010",
  2704=>"010111010",
  2705=>"100011101",
  2706=>"100001011",
  2707=>"001101101",
  2708=>"100001001",
  2709=>"011111011",
  2710=>"100100100",
  2711=>"111011111",
  2712=>"000100001",
  2713=>"101001011",
  2714=>"011001110",
  2715=>"110100110",
  2716=>"000011111",
  2717=>"001000001",
  2718=>"000011100",
  2719=>"111000010",
  2720=>"011110101",
  2721=>"001100111",
  2722=>"110100101",
  2723=>"111110110",
  2724=>"110011011",
  2725=>"111110101",
  2726=>"101101010",
  2727=>"000000010",
  2728=>"001010101",
  2729=>"000111111",
  2730=>"111000111",
  2731=>"001000001",
  2732=>"100100000",
  2733=>"111000011",
  2734=>"000010000",
  2735=>"001001010",
  2736=>"010000001",
  2737=>"100011101",
  2738=>"111111010",
  2739=>"111101010",
  2740=>"010000010",
  2741=>"000101010",
  2742=>"000011010",
  2743=>"101001010",
  2744=>"111100111",
  2745=>"101001001",
  2746=>"011011011",
  2747=>"100100110",
  2748=>"111100100",
  2749=>"111110011",
  2750=>"011010000",
  2751=>"011110111",
  2752=>"100101010",
  2753=>"100010001",
  2754=>"001111100",
  2755=>"010000001",
  2756=>"000000100",
  2757=>"111001000",
  2758=>"101000111",
  2759=>"111000110",
  2760=>"111111111",
  2761=>"100000111",
  2762=>"011111000",
  2763=>"111100001",
  2764=>"011101101",
  2765=>"001001111",
  2766=>"011001011",
  2767=>"100001110",
  2768=>"011111100",
  2769=>"111101010",
  2770=>"110100111",
  2771=>"111000100",
  2772=>"111011101",
  2773=>"111000001",
  2774=>"101100000",
  2775=>"001010010",
  2776=>"110111100",
  2777=>"011101011",
  2778=>"001101001",
  2779=>"111011101",
  2780=>"011010000",
  2781=>"100110010",
  2782=>"000010001",
  2783=>"100111000",
  2784=>"000001111",
  2785=>"011100100",
  2786=>"100101010",
  2787=>"101111011",
  2788=>"001001101",
  2789=>"010010100",
  2790=>"011101101",
  2791=>"011010111",
  2792=>"100001011",
  2793=>"100011101",
  2794=>"011101111",
  2795=>"000101110",
  2796=>"110010011",
  2797=>"110010010",
  2798=>"110011101",
  2799=>"000110111",
  2800=>"011011010",
  2801=>"001101100",
  2802=>"010001100",
  2803=>"110100001",
  2804=>"101111101",
  2805=>"010100000",
  2806=>"010110110",
  2807=>"100110011",
  2808=>"010001010",
  2809=>"000100001",
  2810=>"011011101",
  2811=>"010010010",
  2812=>"100010011",
  2813=>"101011100",
  2814=>"111010010",
  2815=>"100011000",
  2816=>"001100000",
  2817=>"000101111",
  2818=>"111101101",
  2819=>"001100000",
  2820=>"111000010",
  2821=>"000011111",
  2822=>"111101110",
  2823=>"111010010",
  2824=>"010110110",
  2825=>"011011101",
  2826=>"110111000",
  2827=>"101011010",
  2828=>"110001101",
  2829=>"011111010",
  2830=>"011000011",
  2831=>"001110110",
  2832=>"111000011",
  2833=>"110010101",
  2834=>"010010000",
  2835=>"100101011",
  2836=>"111000100",
  2837=>"110010000",
  2838=>"101111110",
  2839=>"001010101",
  2840=>"001011000",
  2841=>"000100010",
  2842=>"000101010",
  2843=>"111101011",
  2844=>"111000000",
  2845=>"110111001",
  2846=>"000100010",
  2847=>"011111000",
  2848=>"111111001",
  2849=>"101111011",
  2850=>"110010010",
  2851=>"111010011",
  2852=>"011010101",
  2853=>"010000010",
  2854=>"111111010",
  2855=>"001110010",
  2856=>"110010111",
  2857=>"100111110",
  2858=>"111111100",
  2859=>"011000110",
  2860=>"101000100",
  2861=>"000000010",
  2862=>"011111000",
  2863=>"111000100",
  2864=>"000001110",
  2865=>"000101001",
  2866=>"111111111",
  2867=>"010100110",
  2868=>"111011011",
  2869=>"001111100",
  2870=>"111101110",
  2871=>"011110010",
  2872=>"101100110",
  2873=>"000001000",
  2874=>"110101110",
  2875=>"110010000",
  2876=>"010011000",
  2877=>"100100100",
  2878=>"111111011",
  2879=>"001000100",
  2880=>"101010000",
  2881=>"100110111",
  2882=>"101001100",
  2883=>"011001011",
  2884=>"000101010",
  2885=>"010000001",
  2886=>"100001100",
  2887=>"101000001",
  2888=>"011110000",
  2889=>"101101100",
  2890=>"000110111",
  2891=>"000101001",
  2892=>"101110001",
  2893=>"000010000",
  2894=>"110100111",
  2895=>"100010010",
  2896=>"101001000",
  2897=>"111111101",
  2898=>"001011001",
  2899=>"101110001",
  2900=>"001101100",
  2901=>"100000010",
  2902=>"000011110",
  2903=>"000011110",
  2904=>"000000111",
  2905=>"011111111",
  2906=>"110101100",
  2907=>"110101011",
  2908=>"000011101",
  2909=>"100000001",
  2910=>"101011011",
  2911=>"111101101",
  2912=>"111110001",
  2913=>"101110100",
  2914=>"001101001",
  2915=>"011111101",
  2916=>"100010000",
  2917=>"001000001",
  2918=>"100110010",
  2919=>"000111110",
  2920=>"000100110",
  2921=>"010011110",
  2922=>"011010111",
  2923=>"111011010",
  2924=>"001101100",
  2925=>"011001001",
  2926=>"000111100",
  2927=>"000011011",
  2928=>"101011111",
  2929=>"001001001",
  2930=>"101010000",
  2931=>"101100001",
  2932=>"001011011",
  2933=>"100011110",
  2934=>"111110000",
  2935=>"111011000",
  2936=>"010000011",
  2937=>"100000110",
  2938=>"101011001",
  2939=>"011010011",
  2940=>"000011111",
  2941=>"011101001",
  2942=>"001101001",
  2943=>"011001111",
  2944=>"000010100",
  2945=>"110010000",
  2946=>"010000110",
  2947=>"111000001",
  2948=>"100001010",
  2949=>"000000110",
  2950=>"111101001",
  2951=>"110100100",
  2952=>"100010101",
  2953=>"111000111",
  2954=>"000101010",
  2955=>"110111111",
  2956=>"000000000",
  2957=>"111110000",
  2958=>"011001100",
  2959=>"111101000",
  2960=>"010111100",
  2961=>"111011101",
  2962=>"111000011",
  2963=>"001011100",
  2964=>"101000001",
  2965=>"101111001",
  2966=>"011101111",
  2967=>"011110100",
  2968=>"110111100",
  2969=>"001010100",
  2970=>"000101111",
  2971=>"111010111",
  2972=>"000000010",
  2973=>"101011010",
  2974=>"010110011",
  2975=>"000001110",
  2976=>"111110010",
  2977=>"011111101",
  2978=>"010001101",
  2979=>"001110000",
  2980=>"111111000",
  2981=>"100110011",
  2982=>"101100010",
  2983=>"100101111",
  2984=>"100001010",
  2985=>"110000101",
  2986=>"011000110",
  2987=>"001000110",
  2988=>"011101101",
  2989=>"101000000",
  2990=>"000011011",
  2991=>"000011000",
  2992=>"000000000",
  2993=>"111111010",
  2994=>"110001101",
  2995=>"100110011",
  2996=>"000111100",
  2997=>"000101010",
  2998=>"010111110",
  2999=>"111110011",
  3000=>"000011111",
  3001=>"111101111",
  3002=>"110101011",
  3003=>"101101110",
  3004=>"110000110",
  3005=>"111000101",
  3006=>"111100010",
  3007=>"000011010",
  3008=>"111111101",
  3009=>"101100010",
  3010=>"000100010",
  3011=>"000110001",
  3012=>"111010010",
  3013=>"000011011",
  3014=>"011111111",
  3015=>"101111101",
  3016=>"100010011",
  3017=>"110110101",
  3018=>"101001111",
  3019=>"111101100",
  3020=>"001011111",
  3021=>"101110010",
  3022=>"010111101",
  3023=>"011100011",
  3024=>"110010011",
  3025=>"000101000",
  3026=>"110110001",
  3027=>"101111111",
  3028=>"111001001",
  3029=>"110001111",
  3030=>"101010010",
  3031=>"111111100",
  3032=>"010011010",
  3033=>"001101110",
  3034=>"000011001",
  3035=>"001011111",
  3036=>"100111001",
  3037=>"000111001",
  3038=>"011110101",
  3039=>"111001000",
  3040=>"101011111",
  3041=>"100001010",
  3042=>"011100101",
  3043=>"001000110",
  3044=>"111111001",
  3045=>"001101101",
  3046=>"001010111",
  3047=>"000001010",
  3048=>"001101111",
  3049=>"010010010",
  3050=>"011010001",
  3051=>"101001110",
  3052=>"101110010",
  3053=>"110111111",
  3054=>"000000001",
  3055=>"010111010",
  3056=>"110100100",
  3057=>"100111111",
  3058=>"010000111",
  3059=>"110010011",
  3060=>"010111000",
  3061=>"110110111",
  3062=>"100100001",
  3063=>"011010011",
  3064=>"100010010",
  3065=>"100000100",
  3066=>"001001101",
  3067=>"110110010",
  3068=>"001010100",
  3069=>"001101101",
  3070=>"010111101",
  3071=>"110111000",
  3072=>"101111110",
  3073=>"011010001",
  3074=>"011101011",
  3075=>"100010010",
  3076=>"100001000",
  3077=>"111010011",
  3078=>"010110111",
  3079=>"100000011",
  3080=>"011101000",
  3081=>"001100101",
  3082=>"011010111",
  3083=>"001111100",
  3084=>"011000011",
  3085=>"111001100",
  3086=>"000101100",
  3087=>"010110001",
  3088=>"000010110",
  3089=>"010100111",
  3090=>"011000111",
  3091=>"101010111",
  3092=>"101011000",
  3093=>"101010110",
  3094=>"100100101",
  3095=>"110010001",
  3096=>"101011100",
  3097=>"011010101",
  3098=>"001111111",
  3099=>"111001111",
  3100=>"110111101",
  3101=>"000000100",
  3102=>"011110101",
  3103=>"100010010",
  3104=>"011011000",
  3105=>"111101100",
  3106=>"010100010",
  3107=>"100111001",
  3108=>"001000001",
  3109=>"010101000",
  3110=>"110100111",
  3111=>"100001101",
  3112=>"010000000",
  3113=>"110111110",
  3114=>"111001000",
  3115=>"001000011",
  3116=>"111100011",
  3117=>"010011010",
  3118=>"000000101",
  3119=>"010000110",
  3120=>"010111100",
  3121=>"000001110",
  3122=>"000010111",
  3123=>"110000010",
  3124=>"000110100",
  3125=>"110001000",
  3126=>"010111010",
  3127=>"000000111",
  3128=>"000101111",
  3129=>"000110111",
  3130=>"111101100",
  3131=>"010000111",
  3132=>"111011000",
  3133=>"101001011",
  3134=>"100010000",
  3135=>"001001111",
  3136=>"000111100",
  3137=>"000101011",
  3138=>"011101100",
  3139=>"011101111",
  3140=>"110101001",
  3141=>"100011101",
  3142=>"010010000",
  3143=>"000111110",
  3144=>"010111110",
  3145=>"110001101",
  3146=>"100001101",
  3147=>"000100001",
  3148=>"101000000",
  3149=>"101100111",
  3150=>"000110010",
  3151=>"011001001",
  3152=>"100000011",
  3153=>"000010110",
  3154=>"111000111",
  3155=>"110000010",
  3156=>"110111011",
  3157=>"001100101",
  3158=>"000000111",
  3159=>"010010001",
  3160=>"010110001",
  3161=>"101000110",
  3162=>"101011000",
  3163=>"111111000",
  3164=>"110001010",
  3165=>"010100110",
  3166=>"000011111",
  3167=>"010111010",
  3168=>"101101111",
  3169=>"000011110",
  3170=>"110000011",
  3171=>"011101001",
  3172=>"100001110",
  3173=>"010111110",
  3174=>"001011010",
  3175=>"011100111",
  3176=>"101101111",
  3177=>"111101101",
  3178=>"010111000",
  3179=>"101010001",
  3180=>"111100001",
  3181=>"010101010",
  3182=>"100011100",
  3183=>"010100011",
  3184=>"001110110",
  3185=>"010000110",
  3186=>"011110110",
  3187=>"110111000",
  3188=>"111001111",
  3189=>"001000110",
  3190=>"010111100",
  3191=>"110100110",
  3192=>"100101100",
  3193=>"101111000",
  3194=>"011000001",
  3195=>"100111010",
  3196=>"111100101",
  3197=>"001111011",
  3198=>"101010100",
  3199=>"001000010",
  3200=>"001100000",
  3201=>"000000000",
  3202=>"101100010",
  3203=>"111010011",
  3204=>"001100000",
  3205=>"101101010",
  3206=>"000000010",
  3207=>"101001000",
  3208=>"101010100",
  3209=>"100011000",
  3210=>"010000011",
  3211=>"001111110",
  3212=>"011010110",
  3213=>"000010001",
  3214=>"001111100",
  3215=>"000101000",
  3216=>"111111010",
  3217=>"001011111",
  3218=>"001111110",
  3219=>"011000000",
  3220=>"000111010",
  3221=>"011110011",
  3222=>"000010101",
  3223=>"011000111",
  3224=>"000000111",
  3225=>"110100001",
  3226=>"010010111",
  3227=>"100000100",
  3228=>"100110010",
  3229=>"011111110",
  3230=>"001111001",
  3231=>"101000011",
  3232=>"001001010",
  3233=>"100011111",
  3234=>"111110110",
  3235=>"110011001",
  3236=>"010101111",
  3237=>"010101100",
  3238=>"111100010",
  3239=>"101010010",
  3240=>"010001100",
  3241=>"010011010",
  3242=>"010100001",
  3243=>"011100101",
  3244=>"000010100",
  3245=>"100110100",
  3246=>"000111000",
  3247=>"000010000",
  3248=>"100011001",
  3249=>"100000100",
  3250=>"011010100",
  3251=>"100100010",
  3252=>"101011001",
  3253=>"001010100",
  3254=>"110111001",
  3255=>"101111101",
  3256=>"010011001",
  3257=>"111110101",
  3258=>"000010110",
  3259=>"001100010",
  3260=>"011101101",
  3261=>"011101011",
  3262=>"010100001",
  3263=>"000010100",
  3264=>"100000101",
  3265=>"101001111",
  3266=>"101011101",
  3267=>"100010100",
  3268=>"101111000",
  3269=>"001010001",
  3270=>"011010111",
  3271=>"010100001",
  3272=>"100100100",
  3273=>"100010000",
  3274=>"010011100",
  3275=>"101111111",
  3276=>"000110101",
  3277=>"110101111",
  3278=>"100011101",
  3279=>"010000000",
  3280=>"111100111",
  3281=>"110111110",
  3282=>"000100110",
  3283=>"101000110",
  3284=>"010001000",
  3285=>"111100011",
  3286=>"000000011",
  3287=>"000110001",
  3288=>"101001011",
  3289=>"010111100",
  3290=>"011100000",
  3291=>"000101000",
  3292=>"001011101",
  3293=>"100111101",
  3294=>"111010000",
  3295=>"001111110",
  3296=>"000011000",
  3297=>"101100101",
  3298=>"111111010",
  3299=>"100010110",
  3300=>"110010100",
  3301=>"110000000",
  3302=>"001010101",
  3303=>"011011010",
  3304=>"100000100",
  3305=>"000011101",
  3306=>"111010001",
  3307=>"111110010",
  3308=>"000100011",
  3309=>"100001111",
  3310=>"000010101",
  3311=>"100011000",
  3312=>"110101011",
  3313=>"011010000",
  3314=>"101001101",
  3315=>"111001011",
  3316=>"110000001",
  3317=>"010000000",
  3318=>"000000000",
  3319=>"100010000",
  3320=>"011011000",
  3321=>"010111001",
  3322=>"011111101",
  3323=>"100001010",
  3324=>"011000001",
  3325=>"010111110",
  3326=>"111011011",
  3327=>"011011101",
  3328=>"010001011",
  3329=>"000010101",
  3330=>"100100100",
  3331=>"001101001",
  3332=>"011111111",
  3333=>"110000100",
  3334=>"000100101",
  3335=>"011110011",
  3336=>"001010011",
  3337=>"001010010",
  3338=>"101010000",
  3339=>"010000001",
  3340=>"000001011",
  3341=>"001111100",
  3342=>"010000100",
  3343=>"100000010",
  3344=>"001111001",
  3345=>"011111001",
  3346=>"010000100",
  3347=>"110000101",
  3348=>"001111111",
  3349=>"111001011",
  3350=>"100000001",
  3351=>"111100100",
  3352=>"001111111",
  3353=>"001001100",
  3354=>"011100101",
  3355=>"101010111",
  3356=>"111110000",
  3357=>"001000000",
  3358=>"011101000",
  3359=>"001001011",
  3360=>"000000001",
  3361=>"001000111",
  3362=>"001100010",
  3363=>"010000011",
  3364=>"110000001",
  3365=>"101110010",
  3366=>"001111111",
  3367=>"101001101",
  3368=>"010100010",
  3369=>"110100110",
  3370=>"110101001",
  3371=>"110110010",
  3372=>"100111111",
  3373=>"000100010",
  3374=>"110010000",
  3375=>"111000000",
  3376=>"111000010",
  3377=>"011011111",
  3378=>"011110000",
  3379=>"111001011",
  3380=>"000100111",
  3381=>"111110101",
  3382=>"000111101",
  3383=>"011000010",
  3384=>"110110111",
  3385=>"101110000",
  3386=>"101110111",
  3387=>"000110011",
  3388=>"010010011",
  3389=>"010110011",
  3390=>"000110000",
  3391=>"001010000",
  3392=>"111101111",
  3393=>"010001001",
  3394=>"111000101",
  3395=>"010010000",
  3396=>"001101010",
  3397=>"010111110",
  3398=>"100000111",
  3399=>"010001011",
  3400=>"100100000",
  3401=>"011010001",
  3402=>"101001110",
  3403=>"010000111",
  3404=>"010011011",
  3405=>"101011100",
  3406=>"001101010",
  3407=>"101111111",
  3408=>"110001111",
  3409=>"010100011",
  3410=>"100011000",
  3411=>"101111110",
  3412=>"100011000",
  3413=>"010110001",
  3414=>"000000001",
  3415=>"001011001",
  3416=>"010010010",
  3417=>"110101111",
  3418=>"010110000",
  3419=>"010011100",
  3420=>"110000110",
  3421=>"011011011",
  3422=>"101101111",
  3423=>"101001000",
  3424=>"010101111",
  3425=>"011101100",
  3426=>"001100110",
  3427=>"101101001",
  3428=>"001101000",
  3429=>"101011111",
  3430=>"011001000",
  3431=>"100101000",
  3432=>"101101000",
  3433=>"010011001",
  3434=>"001011010",
  3435=>"000011110",
  3436=>"010011000",
  3437=>"010111001",
  3438=>"110100010",
  3439=>"001000100",
  3440=>"100001101",
  3441=>"101011111",
  3442=>"111001110",
  3443=>"001001110",
  3444=>"001101101",
  3445=>"110110100",
  3446=>"111110100",
  3447=>"010110111",
  3448=>"000010000",
  3449=>"100010110",
  3450=>"000110001",
  3451=>"001110010",
  3452=>"000001110",
  3453=>"101100111",
  3454=>"000011110",
  3455=>"100011001",
  3456=>"010001110",
  3457=>"010011110",
  3458=>"111010010",
  3459=>"100101011",
  3460=>"001011111",
  3461=>"101000101",
  3462=>"011001100",
  3463=>"010010001",
  3464=>"010000010",
  3465=>"111110101",
  3466=>"010101100",
  3467=>"101101110",
  3468=>"101011111",
  3469=>"001011001",
  3470=>"110000101",
  3471=>"110110110",
  3472=>"011010010",
  3473=>"001010000",
  3474=>"010000011",
  3475=>"111100100",
  3476=>"101010111",
  3477=>"011001110",
  3478=>"110101000",
  3479=>"110101110",
  3480=>"001010111",
  3481=>"000110101",
  3482=>"001000101",
  3483=>"010001110",
  3484=>"001011001",
  3485=>"000000110",
  3486=>"010010101",
  3487=>"011001000",
  3488=>"110100001",
  3489=>"111100000",
  3490=>"010000111",
  3491=>"111010011",
  3492=>"111001100",
  3493=>"010000000",
  3494=>"100011101",
  3495=>"000000000",
  3496=>"100001000",
  3497=>"100011010",
  3498=>"000001101",
  3499=>"000000000",
  3500=>"110010110",
  3501=>"001000011",
  3502=>"000100111",
  3503=>"011010011",
  3504=>"111111110",
  3505=>"100000100",
  3506=>"001101111",
  3507=>"011010111",
  3508=>"100011000",
  3509=>"110110111",
  3510=>"000000101",
  3511=>"100111111",
  3512=>"010010110",
  3513=>"101111110",
  3514=>"100111100",
  3515=>"111111101",
  3516=>"100110101",
  3517=>"000101010",
  3518=>"110100101",
  3519=>"110110111",
  3520=>"001110000",
  3521=>"110101010",
  3522=>"000010111",
  3523=>"000011000",
  3524=>"000101011",
  3525=>"101000010",
  3526=>"101100010",
  3527=>"100111100",
  3528=>"101101100",
  3529=>"000001010",
  3530=>"111100011",
  3531=>"111011111",
  3532=>"100110110",
  3533=>"100110110",
  3534=>"010000011",
  3535=>"110001110",
  3536=>"110010010",
  3537=>"000110001",
  3538=>"011001110",
  3539=>"111011111",
  3540=>"100011111",
  3541=>"000011111",
  3542=>"000000100",
  3543=>"111101000",
  3544=>"010101001",
  3545=>"110101101",
  3546=>"001100010",
  3547=>"000101001",
  3548=>"100011111",
  3549=>"000100100",
  3550=>"000101111",
  3551=>"000000010",
  3552=>"001000001",
  3553=>"101001111",
  3554=>"011101110",
  3555=>"001011010",
  3556=>"001001010",
  3557=>"100001100",
  3558=>"101101011",
  3559=>"010001000",
  3560=>"101000010",
  3561=>"001001110",
  3562=>"100001101",
  3563=>"100100001",
  3564=>"000010000",
  3565=>"110110000",
  3566=>"101101111",
  3567=>"101100000",
  3568=>"010000001",
  3569=>"000101101",
  3570=>"011010110",
  3571=>"110111101",
  3572=>"111100001",
  3573=>"101101110",
  3574=>"001110110",
  3575=>"111001001",
  3576=>"100000100",
  3577=>"111111100",
  3578=>"000101000",
  3579=>"100110011",
  3580=>"011101101",
  3581=>"010000000",
  3582=>"001000111",
  3583=>"101101110",
  3584=>"000110110",
  3585=>"001101001",
  3586=>"001001010",
  3587=>"110111010",
  3588=>"000010000",
  3589=>"011101101",
  3590=>"111100001",
  3591=>"100001010",
  3592=>"101001100",
  3593=>"111110011",
  3594=>"001000101",
  3595=>"001001110",
  3596=>"110000111",
  3597=>"100110100",
  3598=>"111100101",
  3599=>"110110001",
  3600=>"011011110",
  3601=>"000110110",
  3602=>"100100100",
  3603=>"000000110",
  3604=>"000111111",
  3605=>"100001010",
  3606=>"110001100",
  3607=>"101000100",
  3608=>"010111011",
  3609=>"001001101",
  3610=>"010111111",
  3611=>"101111101",
  3612=>"011000001",
  3613=>"111111111",
  3614=>"000011010",
  3615=>"110001001",
  3616=>"101001011",
  3617=>"110001100",
  3618=>"000001011",
  3619=>"010011111",
  3620=>"111011101",
  3621=>"010101101",
  3622=>"111101101",
  3623=>"011101110",
  3624=>"011000011",
  3625=>"110101011",
  3626=>"110110010",
  3627=>"101010110",
  3628=>"111010111",
  3629=>"000001111",
  3630=>"100011100",
  3631=>"101100110",
  3632=>"000100000",
  3633=>"010010010",
  3634=>"100101110",
  3635=>"010110111",
  3636=>"000011100",
  3637=>"011010000",
  3638=>"000101111",
  3639=>"111111100",
  3640=>"110110101",
  3641=>"111001010",
  3642=>"000001100",
  3643=>"000010110",
  3644=>"110101111",
  3645=>"011100100",
  3646=>"111110010",
  3647=>"111100101",
  3648=>"110100110",
  3649=>"110000001",
  3650=>"111111010",
  3651=>"000001001",
  3652=>"001010101",
  3653=>"111100110",
  3654=>"001111110",
  3655=>"101111101",
  3656=>"101001011",
  3657=>"100111100",
  3658=>"000000001",
  3659=>"110100110",
  3660=>"100111110",
  3661=>"000010111",
  3662=>"101010101",
  3663=>"111001001",
  3664=>"110111011",
  3665=>"101011001",
  3666=>"000001110",
  3667=>"110000111",
  3668=>"011011100",
  3669=>"100000101",
  3670=>"100100010",
  3671=>"101101011",
  3672=>"111101101",
  3673=>"010101001",
  3674=>"111111000",
  3675=>"001000111",
  3676=>"001101101",
  3677=>"101010101",
  3678=>"000010011",
  3679=>"100100011",
  3680=>"010100110",
  3681=>"001000000",
  3682=>"100001111",
  3683=>"001001000",
  3684=>"011110111",
  3685=>"111100100",
  3686=>"111011000",
  3687=>"100111101",
  3688=>"010001101",
  3689=>"110011111",
  3690=>"000110111",
  3691=>"001000001",
  3692=>"001001001",
  3693=>"010101111",
  3694=>"110001101",
  3695=>"100110010",
  3696=>"000110000",
  3697=>"110000100",
  3698=>"111010101",
  3699=>"111000111",
  3700=>"101010100",
  3701=>"110101110",
  3702=>"101010011",
  3703=>"001001101",
  3704=>"011100100",
  3705=>"110000110",
  3706=>"000101101",
  3707=>"001000101",
  3708=>"001100011",
  3709=>"111111011",
  3710=>"100010011",
  3711=>"110110010",
  3712=>"101011010",
  3713=>"110101001",
  3714=>"111010100",
  3715=>"001000011",
  3716=>"100000101",
  3717=>"001110001",
  3718=>"010011000",
  3719=>"111001111",
  3720=>"100110111",
  3721=>"001011001",
  3722=>"111111011",
  3723=>"101000010",
  3724=>"101110000",
  3725=>"001011001",
  3726=>"101000010",
  3727=>"011111101",
  3728=>"110100001",
  3729=>"100111001",
  3730=>"011101111",
  3731=>"101101111",
  3732=>"000001001",
  3733=>"111000011",
  3734=>"101010000",
  3735=>"100001001",
  3736=>"101010110",
  3737=>"010011111",
  3738=>"111110000",
  3739=>"100001000",
  3740=>"101010010",
  3741=>"101001101",
  3742=>"101100010",
  3743=>"100011010",
  3744=>"001110100",
  3745=>"110001111",
  3746=>"111111000",
  3747=>"101010011",
  3748=>"010110010",
  3749=>"010111001",
  3750=>"110000010",
  3751=>"000000111",
  3752=>"111111111",
  3753=>"111111111",
  3754=>"100001100",
  3755=>"010000101",
  3756=>"100100110",
  3757=>"000100010",
  3758=>"101111000",
  3759=>"010001000",
  3760=>"100001000",
  3761=>"101010100",
  3762=>"100111001",
  3763=>"111001100",
  3764=>"110110110",
  3765=>"110101001",
  3766=>"101110001",
  3767=>"000110011",
  3768=>"000000110",
  3769=>"111011010",
  3770=>"101011111",
  3771=>"010101011",
  3772=>"001101011",
  3773=>"010111101",
  3774=>"000101011",
  3775=>"100111001",
  3776=>"100010111",
  3777=>"101010110",
  3778=>"010000111",
  3779=>"001010111",
  3780=>"101000011",
  3781=>"000110111",
  3782=>"011101101",
  3783=>"110100011",
  3784=>"000010101",
  3785=>"111100110",
  3786=>"011011001",
  3787=>"111011100",
  3788=>"110110000",
  3789=>"111000101",
  3790=>"110101111",
  3791=>"100000110",
  3792=>"001111001",
  3793=>"000011001",
  3794=>"101010111",
  3795=>"001101001",
  3796=>"001100101",
  3797=>"011001100",
  3798=>"000111010",
  3799=>"110010111",
  3800=>"000010000",
  3801=>"111001011",
  3802=>"111011001",
  3803=>"101010100",
  3804=>"100010010",
  3805=>"101101000",
  3806=>"101101111",
  3807=>"111110001",
  3808=>"001000000",
  3809=>"100001100",
  3810=>"111001000",
  3811=>"000011010",
  3812=>"000001000",
  3813=>"101011001",
  3814=>"110000111",
  3815=>"011001101",
  3816=>"100000000",
  3817=>"100010101",
  3818=>"111101001",
  3819=>"001110111",
  3820=>"111101001",
  3821=>"111101101",
  3822=>"110011000",
  3823=>"111101101",
  3824=>"011000101",
  3825=>"011100011",
  3826=>"110101100",
  3827=>"111101001",
  3828=>"110011110",
  3829=>"011001001",
  3830=>"010001111",
  3831=>"010000000",
  3832=>"001110111",
  3833=>"100000000",
  3834=>"011001010",
  3835=>"101110110",
  3836=>"010010010",
  3837=>"011100101",
  3838=>"001100101",
  3839=>"011011011",
  3840=>"000100000",
  3841=>"110001011",
  3842=>"000011010",
  3843=>"010000110",
  3844=>"100000011",
  3845=>"011000001",
  3846=>"110000111",
  3847=>"100100010",
  3848=>"010000010",
  3849=>"010111001",
  3850=>"000111001",
  3851=>"010100111",
  3852=>"110110110",
  3853=>"001011100",
  3854=>"010011101",
  3855=>"101110110",
  3856=>"010000100",
  3857=>"010110100",
  3858=>"111011001",
  3859=>"001100101",
  3860=>"001110100",
  3861=>"000110000",
  3862=>"001011100",
  3863=>"001000101",
  3864=>"010100100",
  3865=>"010001100",
  3866=>"111100101",
  3867=>"110110100",
  3868=>"001001111",
  3869=>"111001101",
  3870=>"111000110",
  3871=>"111011110",
  3872=>"111100111",
  3873=>"101100001",
  3874=>"001101000",
  3875=>"110100000",
  3876=>"010010001",
  3877=>"111001110",
  3878=>"100000000",
  3879=>"010011011",
  3880=>"110101000",
  3881=>"111011111",
  3882=>"110001001",
  3883=>"000001000",
  3884=>"011010001",
  3885=>"110110110",
  3886=>"000011100",
  3887=>"110111001",
  3888=>"001001110",
  3889=>"100001011",
  3890=>"001000110",
  3891=>"000011110",
  3892=>"110101111",
  3893=>"010100101",
  3894=>"010000100",
  3895=>"100011010",
  3896=>"111110110",
  3897=>"011111001",
  3898=>"100100110",
  3899=>"100111010",
  3900=>"100000101",
  3901=>"111101100",
  3902=>"010100110",
  3903=>"001111010",
  3904=>"011000111",
  3905=>"101100001",
  3906=>"011011100",
  3907=>"010010110",
  3908=>"010101100",
  3909=>"000010111",
  3910=>"100011111",
  3911=>"111001001",
  3912=>"011100101",
  3913=>"100110110",
  3914=>"100101101",
  3915=>"011101111",
  3916=>"100000111",
  3917=>"111010010",
  3918=>"000000000",
  3919=>"110110111",
  3920=>"111110001",
  3921=>"000111011",
  3922=>"011101111",
  3923=>"001001011",
  3924=>"001001110",
  3925=>"011000001",
  3926=>"101010000",
  3927=>"000011001",
  3928=>"010100011",
  3929=>"000000111",
  3930=>"001101000",
  3931=>"100010111",
  3932=>"001001000",
  3933=>"000101000",
  3934=>"111000001",
  3935=>"000111010",
  3936=>"110011001",
  3937=>"110001111",
  3938=>"100111001",
  3939=>"001001100",
  3940=>"101100101",
  3941=>"001101010",
  3942=>"100000100",
  3943=>"110100011",
  3944=>"110111001",
  3945=>"111001100",
  3946=>"001010010",
  3947=>"100010001",
  3948=>"101100001",
  3949=>"110100000",
  3950=>"100110100",
  3951=>"011100100",
  3952=>"001101111",
  3953=>"000010110",
  3954=>"011110001",
  3955=>"101100010",
  3956=>"010000010",
  3957=>"110001111",
  3958=>"101100110",
  3959=>"010101100",
  3960=>"000101100",
  3961=>"100000011",
  3962=>"010101100",
  3963=>"100111101",
  3964=>"110000011",
  3965=>"001000001",
  3966=>"011011000",
  3967=>"100100001",
  3968=>"101011110",
  3969=>"010001000",
  3970=>"011011000",
  3971=>"010001100",
  3972=>"000000011",
  3973=>"001101000",
  3974=>"010001000",
  3975=>"110110100",
  3976=>"010110110",
  3977=>"011000000",
  3978=>"011110111",
  3979=>"001100100",
  3980=>"000010100",
  3981=>"011101000",
  3982=>"111001100",
  3983=>"110001101",
  3984=>"101011000",
  3985=>"110010010",
  3986=>"000000100",
  3987=>"100011010",
  3988=>"101111101",
  3989=>"101011110",
  3990=>"101010100",
  3991=>"000100101",
  3992=>"100111011",
  3993=>"000011011",
  3994=>"111100101",
  3995=>"011100001",
  3996=>"000010100",
  3997=>"010101000",
  3998=>"100001000",
  3999=>"101011111",
  4000=>"101000011",
  4001=>"001000110",
  4002=>"010010101",
  4003=>"110000000",
  4004=>"101001011",
  4005=>"101101110",
  4006=>"110101110",
  4007=>"011111011",
  4008=>"000011111",
  4009=>"000010001",
  4010=>"011010011",
  4011=>"111000000",
  4012=>"101101100",
  4013=>"001101110",
  4014=>"111111110",
  4015=>"000000111",
  4016=>"010000000",
  4017=>"101000011",
  4018=>"111010000",
  4019=>"110011110",
  4020=>"101000100",
  4021=>"100000001",
  4022=>"011110110",
  4023=>"000100010",
  4024=>"111101011",
  4025=>"000011100",
  4026=>"010101110",
  4027=>"101010111",
  4028=>"011011111",
  4029=>"111100001",
  4030=>"100100101",
  4031=>"001010100",
  4032=>"000001101",
  4033=>"000011011",
  4034=>"111100001",
  4035=>"011100101",
  4036=>"001001111",
  4037=>"111000000",
  4038=>"001110101",
  4039=>"111100111",
  4040=>"110000101",
  4041=>"011100001",
  4042=>"111001000",
  4043=>"011101011",
  4044=>"000011001",
  4045=>"011100101",
  4046=>"101011110",
  4047=>"001010001",
  4048=>"100101101",
  4049=>"001010010",
  4050=>"011000001",
  4051=>"001100100",
  4052=>"111101111",
  4053=>"101101110",
  4054=>"110011010",
  4055=>"110111101",
  4056=>"010000001",
  4057=>"110110001",
  4058=>"000100010",
  4059=>"011110000",
  4060=>"101000110",
  4061=>"101110000",
  4062=>"000001101",
  4063=>"110001110",
  4064=>"010110011",
  4065=>"000000011",
  4066=>"010000011",
  4067=>"000010001",
  4068=>"111111100",
  4069=>"010011001",
  4070=>"000111011",
  4071=>"000011001",
  4072=>"000001101",
  4073=>"010000110",
  4074=>"000000111",
  4075=>"100011100",
  4076=>"001100111",
  4077=>"001101010",
  4078=>"101111010",
  4079=>"101111100",
  4080=>"101111110",
  4081=>"111110001",
  4082=>"011110101",
  4083=>"011010001",
  4084=>"100110100",
  4085=>"011110111",
  4086=>"111101111",
  4087=>"011011111",
  4088=>"000001111",
  4089=>"100010000",
  4090=>"110001111",
  4091=>"100111110",
  4092=>"101001101",
  4093=>"100001010",
  4094=>"111100001",
  4095=>"110001111",
  4096=>"011000011",
  4097=>"001010110",
  4098=>"110010111",
  4099=>"011110101",
  4100=>"100101010",
  4101=>"000100011",
  4102=>"111000110",
  4103=>"100100011",
  4104=>"111010010",
  4105=>"100001010",
  4106=>"010011110",
  4107=>"101100010",
  4108=>"101011000",
  4109=>"000111101",
  4110=>"100100101",
  4111=>"000001001",
  4112=>"010101110",
  4113=>"111101100",
  4114=>"010111001",
  4115=>"111101101",
  4116=>"001010011",
  4117=>"100000001",
  4118=>"010100111",
  4119=>"001011101",
  4120=>"000001001",
  4121=>"110111010",
  4122=>"001111110",
  4123=>"101100110",
  4124=>"001011010",
  4125=>"111101100",
  4126=>"011110000",
  4127=>"010100000",
  4128=>"101001010",
  4129=>"011100011",
  4130=>"001101001",
  4131=>"000000110",
  4132=>"111100000",
  4133=>"110000001",
  4134=>"001000011",
  4135=>"001000101",
  4136=>"110000100",
  4137=>"111100101",
  4138=>"000011110",
  4139=>"000100101",
  4140=>"100010010",
  4141=>"010011011",
  4142=>"011010010",
  4143=>"001101011",
  4144=>"011000100",
  4145=>"011111001",
  4146=>"001000001",
  4147=>"000010110",
  4148=>"000000000",
  4149=>"110011100",
  4150=>"001100010",
  4151=>"001100111",
  4152=>"011000000",
  4153=>"001111110",
  4154=>"011100011",
  4155=>"000111010",
  4156=>"101110001",
  4157=>"000000000",
  4158=>"110000000",
  4159=>"110100100",
  4160=>"111111111",
  4161=>"001010101",
  4162=>"011000100",
  4163=>"001010100",
  4164=>"011011001",
  4165=>"111101110",
  4166=>"111011000",
  4167=>"111100010",
  4168=>"101011011",
  4169=>"101100111",
  4170=>"011001010",
  4171=>"000100100",
  4172=>"111111001",
  4173=>"000000011",
  4174=>"011001101",
  4175=>"110000011",
  4176=>"000010011",
  4177=>"100101001",
  4178=>"110111010",
  4179=>"010110001",
  4180=>"111000010",
  4181=>"101010000",
  4182=>"111010010",
  4183=>"111010011",
  4184=>"001101000",
  4185=>"111110110",
  4186=>"101010110",
  4187=>"001101000",
  4188=>"011101010",
  4189=>"110100010",
  4190=>"110010111",
  4191=>"101010101",
  4192=>"101000101",
  4193=>"011010010",
  4194=>"000000111",
  4195=>"001100101",
  4196=>"111010110",
  4197=>"001010111",
  4198=>"010101101",
  4199=>"011100100",
  4200=>"000111010",
  4201=>"100010000",
  4202=>"011111111",
  4203=>"000011100",
  4204=>"010011100",
  4205=>"111011011",
  4206=>"000001110",
  4207=>"001001000",
  4208=>"001110000",
  4209=>"000110101",
  4210=>"110101110",
  4211=>"111101111",
  4212=>"000010000",
  4213=>"100110010",
  4214=>"110011110",
  4215=>"101110000",
  4216=>"110111111",
  4217=>"110101011",
  4218=>"100000101",
  4219=>"000101101",
  4220=>"001010111",
  4221=>"010111010",
  4222=>"011010000",
  4223=>"101111001",
  4224=>"111011110",
  4225=>"111010100",
  4226=>"101001110",
  4227=>"010000011",
  4228=>"111000100",
  4229=>"010111001",
  4230=>"110000110",
  4231=>"110101001",
  4232=>"010100111",
  4233=>"100000001",
  4234=>"001110011",
  4235=>"110100101",
  4236=>"101100000",
  4237=>"001001001",
  4238=>"011000011",
  4239=>"111010111",
  4240=>"110000001",
  4241=>"010011111",
  4242=>"101111100",
  4243=>"100011001",
  4244=>"101100000",
  4245=>"101011001",
  4246=>"000110101",
  4247=>"111010011",
  4248=>"010000000",
  4249=>"011100100",
  4250=>"010101111",
  4251=>"010101110",
  4252=>"110010100",
  4253=>"100100001",
  4254=>"000101010",
  4255=>"110110011",
  4256=>"111101001",
  4257=>"010110110",
  4258=>"110100001",
  4259=>"010001111",
  4260=>"010001011",
  4261=>"110111000",
  4262=>"011111011",
  4263=>"111110110",
  4264=>"110001001",
  4265=>"000000010",
  4266=>"010101000",
  4267=>"101010010",
  4268=>"000111100",
  4269=>"110111100",
  4270=>"001101000",
  4271=>"100000101",
  4272=>"010011000",
  4273=>"110001111",
  4274=>"000110101",
  4275=>"111101101",
  4276=>"001101000",
  4277=>"100100110",
  4278=>"000001000",
  4279=>"100011001",
  4280=>"100101101",
  4281=>"101010011",
  4282=>"010010111",
  4283=>"100111100",
  4284=>"010011000",
  4285=>"010010001",
  4286=>"010000101",
  4287=>"001110011",
  4288=>"101000000",
  4289=>"111000101",
  4290=>"100111011",
  4291=>"110100011",
  4292=>"111100010",
  4293=>"101100101",
  4294=>"100011110",
  4295=>"010101010",
  4296=>"101000011",
  4297=>"001000101",
  4298=>"010110010",
  4299=>"100010100",
  4300=>"001001111",
  4301=>"101111001",
  4302=>"000101111",
  4303=>"001111110",
  4304=>"010001000",
  4305=>"011000001",
  4306=>"011101011",
  4307=>"001000101",
  4308=>"010100001",
  4309=>"111111011",
  4310=>"011110111",
  4311=>"001110001",
  4312=>"111010110",
  4313=>"001111110",
  4314=>"100001100",
  4315=>"011101101",
  4316=>"000101001",
  4317=>"110011110",
  4318=>"010110011",
  4319=>"111001010",
  4320=>"000100001",
  4321=>"110111111",
  4322=>"100011001",
  4323=>"011111111",
  4324=>"110011111",
  4325=>"001111010",
  4326=>"101100011",
  4327=>"101000010",
  4328=>"011001101",
  4329=>"000101010",
  4330=>"011010101",
  4331=>"011000001",
  4332=>"001101001",
  4333=>"011001000",
  4334=>"111110001",
  4335=>"111000101",
  4336=>"111001110",
  4337=>"101101111",
  4338=>"111001001",
  4339=>"010101110",
  4340=>"111101011",
  4341=>"101000001",
  4342=>"001011000",
  4343=>"011010101",
  4344=>"100111001",
  4345=>"011110101",
  4346=>"000100001",
  4347=>"101001011",
  4348=>"111001111",
  4349=>"011111100",
  4350=>"111100000",
  4351=>"101000001",
  4352=>"101000100",
  4353=>"101011110",
  4354=>"010001101",
  4355=>"110000101",
  4356=>"101101001",
  4357=>"000001100",
  4358=>"101110111",
  4359=>"000101001",
  4360=>"100011100",
  4361=>"100111010",
  4362=>"110111111",
  4363=>"010111001",
  4364=>"100010110",
  4365=>"101001010",
  4366=>"101111001",
  4367=>"010110110",
  4368=>"011001000",
  4369=>"111000101",
  4370=>"110011001",
  4371=>"100101111",
  4372=>"100111010",
  4373=>"010110111",
  4374=>"100000111",
  4375=>"001101111",
  4376=>"000000001",
  4377=>"001101001",
  4378=>"001010001",
  4379=>"101011000",
  4380=>"101101001",
  4381=>"000010100",
  4382=>"000001110",
  4383=>"001011100",
  4384=>"110111110",
  4385=>"000011100",
  4386=>"011100111",
  4387=>"100111011",
  4388=>"101110110",
  4389=>"000110011",
  4390=>"100111110",
  4391=>"011000101",
  4392=>"110100010",
  4393=>"001100011",
  4394=>"110000101",
  4395=>"001101001",
  4396=>"100111011",
  4397=>"011010010",
  4398=>"110110010",
  4399=>"011001100",
  4400=>"010011101",
  4401=>"010111101",
  4402=>"001100011",
  4403=>"110111100",
  4404=>"101001001",
  4405=>"000010101",
  4406=>"011000010",
  4407=>"110100111",
  4408=>"010101000",
  4409=>"011001011",
  4410=>"011011101",
  4411=>"011110010",
  4412=>"110001101",
  4413=>"110010001",
  4414=>"100001101",
  4415=>"100001101",
  4416=>"110111111",
  4417=>"101111101",
  4418=>"110010110",
  4419=>"010100001",
  4420=>"111111001",
  4421=>"001011010",
  4422=>"100101001",
  4423=>"111100010",
  4424=>"001001111",
  4425=>"000110011",
  4426=>"011110000",
  4427=>"010101010",
  4428=>"011101110",
  4429=>"000101011",
  4430=>"011001000",
  4431=>"011010001",
  4432=>"001011101",
  4433=>"001111111",
  4434=>"000101010",
  4435=>"111010111",
  4436=>"100101000",
  4437=>"110111110",
  4438=>"011111110",
  4439=>"101101100",
  4440=>"001101011",
  4441=>"000001000",
  4442=>"111011001",
  4443=>"000111011",
  4444=>"001001100",
  4445=>"111110100",
  4446=>"000111100",
  4447=>"110110010",
  4448=>"101011100",
  4449=>"000001101",
  4450=>"001110110",
  4451=>"100000110",
  4452=>"000111011",
  4453=>"000110100",
  4454=>"101110110",
  4455=>"011100110",
  4456=>"101100100",
  4457=>"001011011",
  4458=>"111110110",
  4459=>"010001000",
  4460=>"111111000",
  4461=>"001000110",
  4462=>"001000111",
  4463=>"010001111",
  4464=>"010111110",
  4465=>"111010001",
  4466=>"110101100",
  4467=>"011001000",
  4468=>"100001110",
  4469=>"110000101",
  4470=>"011001000",
  4471=>"010001001",
  4472=>"001000111",
  4473=>"001100111",
  4474=>"000001010",
  4475=>"011011100",
  4476=>"011111110",
  4477=>"000011101",
  4478=>"011010000",
  4479=>"110010010",
  4480=>"111111111",
  4481=>"110111101",
  4482=>"000001001",
  4483=>"111100010",
  4484=>"010011101",
  4485=>"101100100",
  4486=>"010000111",
  4487=>"010010101",
  4488=>"010011001",
  4489=>"011100000",
  4490=>"100010111",
  4491=>"101110111",
  4492=>"001100000",
  4493=>"010111101",
  4494=>"110000110",
  4495=>"010000111",
  4496=>"100000001",
  4497=>"011111110",
  4498=>"111101001",
  4499=>"001010000",
  4500=>"000000111",
  4501=>"001000101",
  4502=>"000000010",
  4503=>"100111111",
  4504=>"111000010",
  4505=>"101011100",
  4506=>"000110011",
  4507=>"001000111",
  4508=>"101010010",
  4509=>"000001110",
  4510=>"000001101",
  4511=>"010110000",
  4512=>"111111101",
  4513=>"100000000",
  4514=>"111001111",
  4515=>"100001010",
  4516=>"111001011",
  4517=>"100111000",
  4518=>"010000001",
  4519=>"011000001",
  4520=>"101111101",
  4521=>"111110101",
  4522=>"010000110",
  4523=>"010011001",
  4524=>"100110011",
  4525=>"110000111",
  4526=>"100110101",
  4527=>"000000000",
  4528=>"100011101",
  4529=>"110111100",
  4530=>"010000110",
  4531=>"001111101",
  4532=>"011110001",
  4533=>"111101000",
  4534=>"101000111",
  4535=>"000100111",
  4536=>"111100010",
  4537=>"001100101",
  4538=>"111101110",
  4539=>"101100111",
  4540=>"100011000",
  4541=>"010110000",
  4542=>"000001010",
  4543=>"001100011",
  4544=>"010000101",
  4545=>"110000101",
  4546=>"001010011",
  4547=>"100000111",
  4548=>"111010010",
  4549=>"001110001",
  4550=>"001111000",
  4551=>"001100010",
  4552=>"000100100",
  4553=>"100111001",
  4554=>"110110111",
  4555=>"001100101",
  4556=>"000110000",
  4557=>"110010011",
  4558=>"011100111",
  4559=>"011000001",
  4560=>"101110010",
  4561=>"000001001",
  4562=>"011100101",
  4563=>"101100010",
  4564=>"100111110",
  4565=>"111001111",
  4566=>"000100000",
  4567=>"001001110",
  4568=>"010110010",
  4569=>"110011110",
  4570=>"100101111",
  4571=>"111001110",
  4572=>"111111011",
  4573=>"100000001",
  4574=>"010101011",
  4575=>"100110111",
  4576=>"010111111",
  4577=>"001101110",
  4578=>"001101011",
  4579=>"011000010",
  4580=>"011000110",
  4581=>"010101001",
  4582=>"001110010",
  4583=>"100100100",
  4584=>"101010000",
  4585=>"011111011",
  4586=>"010011110",
  4587=>"101100010",
  4588=>"001100011",
  4589=>"001110010",
  4590=>"111001011",
  4591=>"010000101",
  4592=>"111110001",
  4593=>"011010111",
  4594=>"011001101",
  4595=>"000001100",
  4596=>"001110110",
  4597=>"000110100",
  4598=>"001001001",
  4599=>"011111011",
  4600=>"000011011",
  4601=>"100110010",
  4602=>"001101110",
  4603=>"101100011",
  4604=>"000101110",
  4605=>"100000001",
  4606=>"100111110",
  4607=>"110011111",
  4608=>"010011011",
  4609=>"100000011",
  4610=>"110101101",
  4611=>"010101011",
  4612=>"100101111",
  4613=>"010111111",
  4614=>"110010110",
  4615=>"110011101",
  4616=>"001001010",
  4617=>"111110000",
  4618=>"011010111",
  4619=>"001101010",
  4620=>"101011010",
  4621=>"000100110",
  4622=>"001100101",
  4623=>"111101111",
  4624=>"011101101",
  4625=>"011000001",
  4626=>"011010111",
  4627=>"101011101",
  4628=>"000000010",
  4629=>"010101111",
  4630=>"000001111",
  4631=>"111000101",
  4632=>"000100101",
  4633=>"100001100",
  4634=>"101010001",
  4635=>"011000110",
  4636=>"010100111",
  4637=>"111110110",
  4638=>"100011000",
  4639=>"110111011",
  4640=>"000000001",
  4641=>"011010001",
  4642=>"001100010",
  4643=>"011000110",
  4644=>"010110101",
  4645=>"100001001",
  4646=>"110010101",
  4647=>"010001111",
  4648=>"010100011",
  4649=>"101000101",
  4650=>"001001011",
  4651=>"011000101",
  4652=>"011000000",
  4653=>"101100001",
  4654=>"010001011",
  4655=>"100001000",
  4656=>"111011100",
  4657=>"011111001",
  4658=>"101001000",
  4659=>"001011101",
  4660=>"111100110",
  4661=>"111010001",
  4662=>"010000110",
  4663=>"111001001",
  4664=>"110110000",
  4665=>"010000010",
  4666=>"110011101",
  4667=>"000111011",
  4668=>"011011101",
  4669=>"011110010",
  4670=>"110101111",
  4671=>"110100001",
  4672=>"001000111",
  4673=>"101111011",
  4674=>"010110000",
  4675=>"111011010",
  4676=>"110000001",
  4677=>"101010100",
  4678=>"010000111",
  4679=>"011000011",
  4680=>"011010010",
  4681=>"011110000",
  4682=>"010011111",
  4683=>"000110111",
  4684=>"111100101",
  4685=>"100001000",
  4686=>"101101110",
  4687=>"101111010",
  4688=>"010000111",
  4689=>"011110000",
  4690=>"100101110",
  4691=>"110110001",
  4692=>"010011110",
  4693=>"000000100",
  4694=>"100001111",
  4695=>"101011010",
  4696=>"010111110",
  4697=>"000101111",
  4698=>"001001010",
  4699=>"100001010",
  4700=>"010011110",
  4701=>"111101111",
  4702=>"011011010",
  4703=>"101000000",
  4704=>"000011011",
  4705=>"000010001",
  4706=>"000011001",
  4707=>"101000010",
  4708=>"111010110",
  4709=>"000011111",
  4710=>"001111110",
  4711=>"110011011",
  4712=>"101111011",
  4713=>"110010100",
  4714=>"100110111",
  4715=>"110000100",
  4716=>"100011010",
  4717=>"101001011",
  4718=>"011101011",
  4719=>"111100011",
  4720=>"101010100",
  4721=>"100011010",
  4722=>"111100111",
  4723=>"111011011",
  4724=>"111010100",
  4725=>"101111111",
  4726=>"101110100",
  4727=>"010000011",
  4728=>"101110110",
  4729=>"001101011",
  4730=>"001000111",
  4731=>"110100100",
  4732=>"111010101",
  4733=>"110001111",
  4734=>"110010101",
  4735=>"101010000",
  4736=>"010100000",
  4737=>"000111100",
  4738=>"111011111",
  4739=>"001000101",
  4740=>"100011001",
  4741=>"011010001",
  4742=>"101101110",
  4743=>"100101010",
  4744=>"111011001",
  4745=>"000001101",
  4746=>"010011101",
  4747=>"100001111",
  4748=>"111000111",
  4749=>"100111000",
  4750=>"111100011",
  4751=>"111001011",
  4752=>"010000010",
  4753=>"010111100",
  4754=>"101100011",
  4755=>"101100000",
  4756=>"101101010",
  4757=>"001100010",
  4758=>"101111010",
  4759=>"010000011",
  4760=>"011101010",
  4761=>"001101011",
  4762=>"000001011",
  4763=>"100000111",
  4764=>"110111001",
  4765=>"011111001",
  4766=>"100001100",
  4767=>"111001101",
  4768=>"010100000",
  4769=>"000111010",
  4770=>"101000111",
  4771=>"101000100",
  4772=>"111001101",
  4773=>"011110011",
  4774=>"111001100",
  4775=>"000001000",
  4776=>"010101110",
  4777=>"100010010",
  4778=>"011000010",
  4779=>"100000100",
  4780=>"010000111",
  4781=>"011000001",
  4782=>"001000100",
  4783=>"110100001",
  4784=>"011011111",
  4785=>"000000111",
  4786=>"001011111",
  4787=>"110100001",
  4788=>"101111110",
  4789=>"011101101",
  4790=>"011000001",
  4791=>"100000100",
  4792=>"110001011",
  4793=>"010110101",
  4794=>"011000011",
  4795=>"101101111",
  4796=>"111110110",
  4797=>"100111110",
  4798=>"111000000",
  4799=>"000101011",
  4800=>"110111100",
  4801=>"110011111",
  4802=>"000101000",
  4803=>"100001111",
  4804=>"111011011",
  4805=>"001110110",
  4806=>"110111101",
  4807=>"001111110",
  4808=>"011110110",
  4809=>"101001010",
  4810=>"001010111",
  4811=>"011011011",
  4812=>"000001001",
  4813=>"010111011",
  4814=>"010000111",
  4815=>"011000011",
  4816=>"110011111",
  4817=>"011100010",
  4818=>"010001100",
  4819=>"011001011",
  4820=>"000110011",
  4821=>"110000010",
  4822=>"001010011",
  4823=>"111101101",
  4824=>"010100000",
  4825=>"001100011",
  4826=>"111111000",
  4827=>"001100000",
  4828=>"001111110",
  4829=>"011110000",
  4830=>"011111111",
  4831=>"111100011",
  4832=>"110000000",
  4833=>"110110011",
  4834=>"001000011",
  4835=>"010011110",
  4836=>"110100000",
  4837=>"011000101",
  4838=>"000011111",
  4839=>"000000111",
  4840=>"101111111",
  4841=>"001100001",
  4842=>"011111000",
  4843=>"010100101",
  4844=>"011111110",
  4845=>"110110010",
  4846=>"110010010",
  4847=>"000000101",
  4848=>"101001110",
  4849=>"010111011",
  4850=>"010110111",
  4851=>"011001001",
  4852=>"000110001",
  4853=>"001111100",
  4854=>"001001001",
  4855=>"000001110",
  4856=>"100111111",
  4857=>"011010100",
  4858=>"001010010",
  4859=>"000001100",
  4860=>"110010000",
  4861=>"010100101",
  4862=>"111000000",
  4863=>"001100110",
  4864=>"010000001",
  4865=>"110111101",
  4866=>"110001011",
  4867=>"110001011",
  4868=>"000101101",
  4869=>"101100001",
  4870=>"111111010",
  4871=>"101101100",
  4872=>"101111101",
  4873=>"111011110",
  4874=>"111010011",
  4875=>"110110000",
  4876=>"001001000",
  4877=>"000010001",
  4878=>"000000001",
  4879=>"110110010",
  4880=>"110011110",
  4881=>"111110111",
  4882=>"011100100",
  4883=>"010101110",
  4884=>"001011110",
  4885=>"110010111",
  4886=>"011111100",
  4887=>"111101100",
  4888=>"100110000",
  4889=>"101000000",
  4890=>"000000000",
  4891=>"011011111",
  4892=>"011011101",
  4893=>"011010100",
  4894=>"010010000",
  4895=>"101101000",
  4896=>"000101111",
  4897=>"110011000",
  4898=>"101100010",
  4899=>"011001100",
  4900=>"111011010",
  4901=>"001101111",
  4902=>"111000111",
  4903=>"011001010",
  4904=>"100011011",
  4905=>"101100001",
  4906=>"101000011",
  4907=>"110011000",
  4908=>"000001010",
  4909=>"111011111",
  4910=>"010110010",
  4911=>"000101111",
  4912=>"111110001",
  4913=>"110100001",
  4914=>"001101010",
  4915=>"111100011",
  4916=>"100101000",
  4917=>"000010101",
  4918=>"111100100",
  4919=>"100101111",
  4920=>"111100011",
  4921=>"010001110",
  4922=>"000010111",
  4923=>"000000010",
  4924=>"110001110",
  4925=>"111111111",
  4926=>"010101011",
  4927=>"101011110",
  4928=>"001100011",
  4929=>"011111110",
  4930=>"101110111",
  4931=>"010010111",
  4932=>"011100110",
  4933=>"001011010",
  4934=>"000001101",
  4935=>"111111111",
  4936=>"100011101",
  4937=>"111111001",
  4938=>"111110001",
  4939=>"101000001",
  4940=>"101000111",
  4941=>"110011110",
  4942=>"110011010",
  4943=>"011010100",
  4944=>"101101100",
  4945=>"101101000",
  4946=>"010101001",
  4947=>"001110110",
  4948=>"010100100",
  4949=>"001111101",
  4950=>"110000010",
  4951=>"101111101",
  4952=>"011100101",
  4953=>"110011100",
  4954=>"101111111",
  4955=>"111110011",
  4956=>"111101100",
  4957=>"100111111",
  4958=>"110011111",
  4959=>"001011111",
  4960=>"101100001",
  4961=>"010110010",
  4962=>"011001101",
  4963=>"000111111",
  4964=>"100001100",
  4965=>"100101101",
  4966=>"000000000",
  4967=>"011101110",
  4968=>"110001001",
  4969=>"110111110",
  4970=>"000000001",
  4971=>"000001000",
  4972=>"000100000",
  4973=>"100001000",
  4974=>"000111010",
  4975=>"000100101",
  4976=>"111011110",
  4977=>"000001101",
  4978=>"110001010",
  4979=>"011001010",
  4980=>"101100011",
  4981=>"000101010",
  4982=>"001111011",
  4983=>"110010111",
  4984=>"110001110",
  4985=>"001001011",
  4986=>"000110111",
  4987=>"010110101",
  4988=>"010100111",
  4989=>"010100110",
  4990=>"010110011",
  4991=>"001111001",
  4992=>"110011101",
  4993=>"001111101",
  4994=>"110010011",
  4995=>"001110100",
  4996=>"101100011",
  4997=>"101000010",
  4998=>"100000010",
  4999=>"011001110",
  5000=>"111010000",
  5001=>"110011001",
  5002=>"110010011",
  5003=>"011011000",
  5004=>"111010001",
  5005=>"111000110",
  5006=>"000101100",
  5007=>"111000100",
  5008=>"010111010",
  5009=>"010010010",
  5010=>"000000000",
  5011=>"100110101",
  5012=>"001100100",
  5013=>"011010100",
  5014=>"001010101",
  5015=>"110000010",
  5016=>"111111101",
  5017=>"001000010",
  5018=>"001000010",
  5019=>"110001001",
  5020=>"000100111",
  5021=>"011000110",
  5022=>"000001111",
  5023=>"011011010",
  5024=>"101100111",
  5025=>"000001011",
  5026=>"001101110",
  5027=>"001110011",
  5028=>"100001111",
  5029=>"001101100",
  5030=>"010110101",
  5031=>"110101111",
  5032=>"001011100",
  5033=>"101001000",
  5034=>"111110100",
  5035=>"001010111",
  5036=>"110010111",
  5037=>"001111011",
  5038=>"010111100",
  5039=>"000011001",
  5040=>"010101101",
  5041=>"110111000",
  5042=>"011101101",
  5043=>"101000101",
  5044=>"100001001",
  5045=>"001111011",
  5046=>"101010101",
  5047=>"000010111",
  5048=>"010110100",
  5049=>"001000010",
  5050=>"100011100",
  5051=>"100010010",
  5052=>"111010011",
  5053=>"110100110",
  5054=>"000101110",
  5055=>"000001010",
  5056=>"011101110",
  5057=>"010000011",
  5058=>"010110101",
  5059=>"100111100",
  5060=>"111001101",
  5061=>"111010110",
  5062=>"011101001",
  5063=>"011001011",
  5064=>"101101111",
  5065=>"000011100",
  5066=>"110110100",
  5067=>"001100100",
  5068=>"011010001",
  5069=>"010000101",
  5070=>"111000010",
  5071=>"000110011",
  5072=>"110011100",
  5073=>"101101001",
  5074=>"100011011",
  5075=>"010001000",
  5076=>"001000010",
  5077=>"100001101",
  5078=>"000010101",
  5079=>"101010000",
  5080=>"000000111",
  5081=>"011000100",
  5082=>"000110000",
  5083=>"000110111",
  5084=>"010100010",
  5085=>"100100100",
  5086=>"010101000",
  5087=>"010101010",
  5088=>"111101100",
  5089=>"001001001",
  5090=>"100000000",
  5091=>"000011110",
  5092=>"010100111",
  5093=>"011011010",
  5094=>"101110110",
  5095=>"000000000",
  5096=>"111000000",
  5097=>"010101010",
  5098=>"001110101",
  5099=>"111011101",
  5100=>"011111101",
  5101=>"000000001",
  5102=>"100011110",
  5103=>"001110101",
  5104=>"001010101",
  5105=>"110110110",
  5106=>"011000001",
  5107=>"000010010",
  5108=>"010010011",
  5109=>"111101111",
  5110=>"111101000",
  5111=>"100100110",
  5112=>"011100101",
  5113=>"110110000",
  5114=>"010000111",
  5115=>"110110010",
  5116=>"100100110",
  5117=>"011000000",
  5118=>"110111001",
  5119=>"000101011",
  5120=>"010000011",
  5121=>"001011011",
  5122=>"010000110",
  5123=>"010101000",
  5124=>"010111100",
  5125=>"010001001",
  5126=>"111110110",
  5127=>"101000000",
  5128=>"111001001",
  5129=>"110101111",
  5130=>"110001001",
  5131=>"111100101",
  5132=>"010100100",
  5133=>"100001001",
  5134=>"010001001",
  5135=>"110111110",
  5136=>"110001010",
  5137=>"011010011",
  5138=>"100101011",
  5139=>"100000111",
  5140=>"110110111",
  5141=>"110011111",
  5142=>"111111010",
  5143=>"001100000",
  5144=>"011011001",
  5145=>"000010111",
  5146=>"110111110",
  5147=>"011100000",
  5148=>"010011000",
  5149=>"110001100",
  5150=>"010000110",
  5151=>"001010110",
  5152=>"000000010",
  5153=>"100010100",
  5154=>"001001010",
  5155=>"100001000",
  5156=>"101100011",
  5157=>"011010110",
  5158=>"111000111",
  5159=>"001011010",
  5160=>"011110110",
  5161=>"110110111",
  5162=>"100010100",
  5163=>"101000100",
  5164=>"100001011",
  5165=>"110101010",
  5166=>"010111010",
  5167=>"110111111",
  5168=>"000110001",
  5169=>"100000110",
  5170=>"011000101",
  5171=>"001011110",
  5172=>"111000110",
  5173=>"010011000",
  5174=>"011010011",
  5175=>"101111100",
  5176=>"110001000",
  5177=>"000110100",
  5178=>"101100010",
  5179=>"100100010",
  5180=>"101110000",
  5181=>"010001001",
  5182=>"101111000",
  5183=>"011011100",
  5184=>"010010001",
  5185=>"101100000",
  5186=>"001011010",
  5187=>"111010100",
  5188=>"011110101",
  5189=>"001000101",
  5190=>"111011011",
  5191=>"110111110",
  5192=>"101001010",
  5193=>"001010001",
  5194=>"101000100",
  5195=>"111110001",
  5196=>"100100010",
  5197=>"110111100",
  5198=>"111000100",
  5199=>"110001010",
  5200=>"100110111",
  5201=>"001001000",
  5202=>"111110000",
  5203=>"101000010",
  5204=>"011000010",
  5205=>"011101011",
  5206=>"000101100",
  5207=>"100101111",
  5208=>"011110000",
  5209=>"110000011",
  5210=>"011101010",
  5211=>"001010110",
  5212=>"111011011",
  5213=>"100010010",
  5214=>"100111110",
  5215=>"001100100",
  5216=>"001000101",
  5217=>"111001000",
  5218=>"110000101",
  5219=>"011010001",
  5220=>"010010110",
  5221=>"111000001",
  5222=>"111011101",
  5223=>"010100100",
  5224=>"000110001",
  5225=>"100101001",
  5226=>"101000110",
  5227=>"010010000",
  5228=>"110111101",
  5229=>"111010000",
  5230=>"110011000",
  5231=>"111101010",
  5232=>"100000010",
  5233=>"101110100",
  5234=>"110101011",
  5235=>"101010111",
  5236=>"001100000",
  5237=>"100001011",
  5238=>"001011101",
  5239=>"010000011",
  5240=>"010001101",
  5241=>"000001010",
  5242=>"011111101",
  5243=>"000110001",
  5244=>"110100011",
  5245=>"110011011",
  5246=>"000000111",
  5247=>"011110000",
  5248=>"010000100",
  5249=>"101111100",
  5250=>"101101101",
  5251=>"100010101",
  5252=>"111101101",
  5253=>"000000001",
  5254=>"011101010",
  5255=>"001000101",
  5256=>"111111101",
  5257=>"101010001",
  5258=>"110001100",
  5259=>"010011001",
  5260=>"001000011",
  5261=>"110110000",
  5262=>"010000111",
  5263=>"001110101",
  5264=>"101101111",
  5265=>"011001110",
  5266=>"111100100",
  5267=>"010111110",
  5268=>"111101111",
  5269=>"100010100",
  5270=>"110000101",
  5271=>"110110100",
  5272=>"000110001",
  5273=>"010001011",
  5274=>"111111000",
  5275=>"010101111",
  5276=>"011000001",
  5277=>"111111001",
  5278=>"100110000",
  5279=>"110010100",
  5280=>"000010101",
  5281=>"010000100",
  5282=>"001100111",
  5283=>"101010110",
  5284=>"100111110",
  5285=>"000110001",
  5286=>"000001000",
  5287=>"100110110",
  5288=>"111101010",
  5289=>"101010010",
  5290=>"101011001",
  5291=>"101110011",
  5292=>"000111110",
  5293=>"110011001",
  5294=>"000001101",
  5295=>"010111010",
  5296=>"000000111",
  5297=>"011010111",
  5298=>"111010110",
  5299=>"001100011",
  5300=>"000011011",
  5301=>"011011111",
  5302=>"010001010",
  5303=>"011100001",
  5304=>"000100100",
  5305=>"010100001",
  5306=>"100110110",
  5307=>"011110010",
  5308=>"000110100",
  5309=>"011101001",
  5310=>"000100010",
  5311=>"011000111",
  5312=>"010011110",
  5313=>"110101001",
  5314=>"101111101",
  5315=>"011000100",
  5316=>"011101000",
  5317=>"100100100",
  5318=>"010000100",
  5319=>"011000010",
  5320=>"111011010",
  5321=>"100101000",
  5322=>"100100110",
  5323=>"111011111",
  5324=>"110100100",
  5325=>"110111001",
  5326=>"001100100",
  5327=>"001011010",
  5328=>"110001000",
  5329=>"111110010",
  5330=>"000010010",
  5331=>"000111100",
  5332=>"111110100",
  5333=>"111110000",
  5334=>"100000100",
  5335=>"111100001",
  5336=>"100010100",
  5337=>"010010110",
  5338=>"100001100",
  5339=>"110111111",
  5340=>"000010001",
  5341=>"111110111",
  5342=>"101001110",
  5343=>"111010110",
  5344=>"100110001",
  5345=>"011110100",
  5346=>"001111000",
  5347=>"110010000",
  5348=>"110100011",
  5349=>"101111101",
  5350=>"011111110",
  5351=>"011111011",
  5352=>"010001010",
  5353=>"001110101",
  5354=>"010000100",
  5355=>"000111001",
  5356=>"111010001",
  5357=>"011000101",
  5358=>"000001101",
  5359=>"001010101",
  5360=>"100110000",
  5361=>"111011000",
  5362=>"010101000",
  5363=>"101000111",
  5364=>"111011100",
  5365=>"010110100",
  5366=>"011110000",
  5367=>"110000111",
  5368=>"001110010",
  5369=>"101011000",
  5370=>"010100101",
  5371=>"000011110",
  5372=>"000000010",
  5373=>"000000111",
  5374=>"101010000",
  5375=>"011111111",
  5376=>"000000111",
  5377=>"111101001",
  5378=>"111111000",
  5379=>"000100001",
  5380=>"110011100",
  5381=>"011011100",
  5382=>"011101011",
  5383=>"110101011",
  5384=>"000111001",
  5385=>"111001110",
  5386=>"110100100",
  5387=>"100000010",
  5388=>"010110110",
  5389=>"000101000",
  5390=>"010100101",
  5391=>"001010110",
  5392=>"101000110",
  5393=>"000100101",
  5394=>"001001110",
  5395=>"111110010",
  5396=>"010100111",
  5397=>"111110000",
  5398=>"110010001",
  5399=>"000000100",
  5400=>"110010010",
  5401=>"000110001",
  5402=>"001100010",
  5403=>"101010000",
  5404=>"101111101",
  5405=>"000000001",
  5406=>"010101111",
  5407=>"001010011",
  5408=>"001010101",
  5409=>"111100010",
  5410=>"110011000",
  5411=>"010001110",
  5412=>"001010010",
  5413=>"010111011",
  5414=>"101001001",
  5415=>"001111011",
  5416=>"000001100",
  5417=>"000000000",
  5418=>"111010001",
  5419=>"101011000",
  5420=>"100010010",
  5421=>"001011000",
  5422=>"001000111",
  5423=>"001111001",
  5424=>"011001001",
  5425=>"110001001",
  5426=>"000010101",
  5427=>"101110010",
  5428=>"001110101",
  5429=>"111100111",
  5430=>"000101010",
  5431=>"100000000",
  5432=>"000001001",
  5433=>"010010110",
  5434=>"010101011",
  5435=>"000100101",
  5436=>"100000110",
  5437=>"001110101",
  5438=>"100010010",
  5439=>"100000001",
  5440=>"110100010",
  5441=>"110101010",
  5442=>"010011110",
  5443=>"000010101",
  5444=>"010011101",
  5445=>"001111000",
  5446=>"001100001",
  5447=>"110010001",
  5448=>"011000001",
  5449=>"100000110",
  5450=>"101111001",
  5451=>"001100001",
  5452=>"110111011",
  5453=>"111111110",
  5454=>"010011110",
  5455=>"111011011",
  5456=>"110110011",
  5457=>"101010011",
  5458=>"011010101",
  5459=>"110111010",
  5460=>"101001100",
  5461=>"110111101",
  5462=>"111000001",
  5463=>"000011001",
  5464=>"000111110",
  5465=>"000100011",
  5466=>"101100111",
  5467=>"110000000",
  5468=>"000100011",
  5469=>"001011110",
  5470=>"001011001",
  5471=>"110110101",
  5472=>"011000100",
  5473=>"011010010",
  5474=>"110000100",
  5475=>"000000001",
  5476=>"001001000",
  5477=>"001000011",
  5478=>"001001001",
  5479=>"010101011",
  5480=>"000011001",
  5481=>"101000010",
  5482=>"111101111",
  5483=>"101001010",
  5484=>"000110101",
  5485=>"101001111",
  5486=>"000000100",
  5487=>"011100111",
  5488=>"000101111",
  5489=>"101011101",
  5490=>"110100110",
  5491=>"100101101",
  5492=>"100011010",
  5493=>"011001101",
  5494=>"101000001",
  5495=>"001010111",
  5496=>"010100011",
  5497=>"010011011",
  5498=>"001101100",
  5499=>"110000001",
  5500=>"011000101",
  5501=>"000011010",
  5502=>"111111101",
  5503=>"101001010",
  5504=>"011110001",
  5505=>"100100001",
  5506=>"100100111",
  5507=>"111101011",
  5508=>"011011001",
  5509=>"110011101",
  5510=>"111101111",
  5511=>"000010001",
  5512=>"100011100",
  5513=>"111110101",
  5514=>"010110000",
  5515=>"110101110",
  5516=>"110000001",
  5517=>"011001111",
  5518=>"101110100",
  5519=>"000001101",
  5520=>"010110100",
  5521=>"000010101",
  5522=>"010100101",
  5523=>"110011011",
  5524=>"001110111",
  5525=>"110100100",
  5526=>"111010111",
  5527=>"110001010",
  5528=>"010000001",
  5529=>"110100001",
  5530=>"110001101",
  5531=>"001100001",
  5532=>"011101000",
  5533=>"000000011",
  5534=>"011011100",
  5535=>"011100111",
  5536=>"100111001",
  5537=>"001000010",
  5538=>"000000000",
  5539=>"100000100",
  5540=>"010001000",
  5541=>"000000010",
  5542=>"100010000",
  5543=>"101010000",
  5544=>"001010111",
  5545=>"101111110",
  5546=>"100101111",
  5547=>"110011110",
  5548=>"010111000",
  5549=>"010010000",
  5550=>"100000101",
  5551=>"001100111",
  5552=>"011001011",
  5553=>"000100100",
  5554=>"101101010",
  5555=>"110011110",
  5556=>"010010100",
  5557=>"101001111",
  5558=>"101111011",
  5559=>"111011000",
  5560=>"111101011",
  5561=>"111111010",
  5562=>"100101111",
  5563=>"000011011",
  5564=>"110110001",
  5565=>"010001100",
  5566=>"100010100",
  5567=>"100001110",
  5568=>"001100000",
  5569=>"110000011",
  5570=>"110000001",
  5571=>"000101001",
  5572=>"110001110",
  5573=>"100111101",
  5574=>"000101010",
  5575=>"000001000",
  5576=>"100000010",
  5577=>"100001101",
  5578=>"000011100",
  5579=>"100010110",
  5580=>"111011001",
  5581=>"110100010",
  5582=>"100011000",
  5583=>"110110110",
  5584=>"010010000",
  5585=>"001101001",
  5586=>"000001110",
  5587=>"011011001",
  5588=>"001100101",
  5589=>"001000010",
  5590=>"010010000",
  5591=>"010101111",
  5592=>"001110101",
  5593=>"111111101",
  5594=>"001010000",
  5595=>"000000000",
  5596=>"010011001",
  5597=>"011100101",
  5598=>"011101000",
  5599=>"101110101",
  5600=>"111011111",
  5601=>"101111011",
  5602=>"010100010",
  5603=>"111010110",
  5604=>"101000100",
  5605=>"001010011",
  5606=>"111100001",
  5607=>"100101001",
  5608=>"101000000",
  5609=>"011101101",
  5610=>"100100011",
  5611=>"100100101",
  5612=>"100101010",
  5613=>"100010000",
  5614=>"110001000",
  5615=>"100100101",
  5616=>"111111111",
  5617=>"100011001",
  5618=>"010011000",
  5619=>"100100001",
  5620=>"001101011",
  5621=>"101111100",
  5622=>"000001110",
  5623=>"000111110",
  5624=>"010000001",
  5625=>"110010101",
  5626=>"001100001",
  5627=>"110000000",
  5628=>"101100110",
  5629=>"000101011",
  5630=>"110001101",
  5631=>"110000000",
  5632=>"000111000",
  5633=>"110100111",
  5634=>"000001100",
  5635=>"111001011",
  5636=>"011111100",
  5637=>"001000111",
  5638=>"100100010",
  5639=>"000100111",
  5640=>"011011101",
  5641=>"001001110",
  5642=>"101010010",
  5643=>"000001010",
  5644=>"010011100",
  5645=>"110101110",
  5646=>"001100001",
  5647=>"001000100",
  5648=>"000110011",
  5649=>"100000000",
  5650=>"100001110",
  5651=>"011100000",
  5652=>"001000010",
  5653=>"100111111",
  5654=>"111100011",
  5655=>"111100101",
  5656=>"100000001",
  5657=>"001111111",
  5658=>"001110111",
  5659=>"001000100",
  5660=>"001001001",
  5661=>"010110111",
  5662=>"011011001",
  5663=>"000011111",
  5664=>"101000101",
  5665=>"110100000",
  5666=>"100111010",
  5667=>"110010000",
  5668=>"111000001",
  5669=>"001000111",
  5670=>"101010000",
  5671=>"110011100",
  5672=>"000100110",
  5673=>"110101100",
  5674=>"001010001",
  5675=>"101110110",
  5676=>"000101000",
  5677=>"001001110",
  5678=>"010110100",
  5679=>"000011100",
  5680=>"100000101",
  5681=>"111011010",
  5682=>"111110100",
  5683=>"101110100",
  5684=>"010110100",
  5685=>"010110001",
  5686=>"100101001",
  5687=>"001001100",
  5688=>"110011000",
  5689=>"010010101",
  5690=>"001010100",
  5691=>"010011101",
  5692=>"101011000",
  5693=>"000010011",
  5694=>"010000011",
  5695=>"000101100",
  5696=>"111101111",
  5697=>"110100100",
  5698=>"101100100",
  5699=>"001111111",
  5700=>"111000110",
  5701=>"111000110",
  5702=>"011100100",
  5703=>"110111001",
  5704=>"110011011",
  5705=>"011110101",
  5706=>"111001000",
  5707=>"111001111",
  5708=>"000000000",
  5709=>"110101001",
  5710=>"001000011",
  5711=>"110101110",
  5712=>"011010111",
  5713=>"100001010",
  5714=>"110111001",
  5715=>"000100001",
  5716=>"101011110",
  5717=>"011101100",
  5718=>"101001111",
  5719=>"100110010",
  5720=>"100000111",
  5721=>"011000110",
  5722=>"000000110",
  5723=>"101000010",
  5724=>"000010001",
  5725=>"010101100",
  5726=>"011110111",
  5727=>"111111111",
  5728=>"111101011",
  5729=>"110101110",
  5730=>"100110011",
  5731=>"000001010",
  5732=>"101111111",
  5733=>"111010010",
  5734=>"011100101",
  5735=>"101101101",
  5736=>"010010011",
  5737=>"000001100",
  5738=>"001111010",
  5739=>"100010100",
  5740=>"101001010",
  5741=>"011011001",
  5742=>"111101011",
  5743=>"101101100",
  5744=>"111000101",
  5745=>"010101000",
  5746=>"011101000",
  5747=>"010100000",
  5748=>"101101100",
  5749=>"110111110",
  5750=>"101110001",
  5751=>"010000111",
  5752=>"110011111",
  5753=>"101011011",
  5754=>"101010101",
  5755=>"011111010",
  5756=>"000000100",
  5757=>"111011000",
  5758=>"001010100",
  5759=>"000111110",
  5760=>"000000000",
  5761=>"000111111",
  5762=>"110001110",
  5763=>"100100100",
  5764=>"011010111",
  5765=>"001100000",
  5766=>"110000011",
  5767=>"110001001",
  5768=>"010111011",
  5769=>"101001001",
  5770=>"011110100",
  5771=>"101111100",
  5772=>"000000101",
  5773=>"000100101",
  5774=>"000011000",
  5775=>"101011111",
  5776=>"000111110",
  5777=>"000101001",
  5778=>"101000011",
  5779=>"101010101",
  5780=>"001001100",
  5781=>"100001011",
  5782=>"001001000",
  5783=>"011101011",
  5784=>"000000001",
  5785=>"011011101",
  5786=>"000100000",
  5787=>"110111110",
  5788=>"011010111",
  5789=>"001000100",
  5790=>"011100101",
  5791=>"111000101",
  5792=>"110111110",
  5793=>"110111100",
  5794=>"100000000",
  5795=>"011011001",
  5796=>"111011100",
  5797=>"101111001",
  5798=>"000001001",
  5799=>"110111010",
  5800=>"010000111",
  5801=>"111111111",
  5802=>"111001001",
  5803=>"001110100",
  5804=>"100011001",
  5805=>"110001010",
  5806=>"010011111",
  5807=>"001011000",
  5808=>"000100111",
  5809=>"111100000",
  5810=>"100000100",
  5811=>"000110101",
  5812=>"100101010",
  5813=>"111111001",
  5814=>"111100000",
  5815=>"111011011",
  5816=>"001111000",
  5817=>"100010011",
  5818=>"101011100",
  5819=>"100010001",
  5820=>"101010110",
  5821=>"000000000",
  5822=>"110000011",
  5823=>"000010001",
  5824=>"001100110",
  5825=>"010010011",
  5826=>"000010010",
  5827=>"111100110",
  5828=>"111010100",
  5829=>"100011100",
  5830=>"000100010",
  5831=>"110010010",
  5832=>"000110001",
  5833=>"101000001",
  5834=>"011110011",
  5835=>"010000000",
  5836=>"101101101",
  5837=>"100010001",
  5838=>"011111111",
  5839=>"010011101",
  5840=>"011111000",
  5841=>"000111001",
  5842=>"100111001",
  5843=>"111001000",
  5844=>"101101110",
  5845=>"001000001",
  5846=>"001111101",
  5847=>"101101111",
  5848=>"011100100",
  5849=>"111110101",
  5850=>"000110011",
  5851=>"000010000",
  5852=>"000001010",
  5853=>"000111000",
  5854=>"010000110",
  5855=>"111011010",
  5856=>"011010111",
  5857=>"100000011",
  5858=>"100000101",
  5859=>"111110100",
  5860=>"000000000",
  5861=>"111110110",
  5862=>"011100000",
  5863=>"101011111",
  5864=>"000001011",
  5865=>"000100101",
  5866=>"011010111",
  5867=>"110111101",
  5868=>"010001100",
  5869=>"010110101",
  5870=>"101010100",
  5871=>"100010100",
  5872=>"000101011",
  5873=>"001001111",
  5874=>"010001011",
  5875=>"101110110",
  5876=>"100010011",
  5877=>"011010111",
  5878=>"000011001",
  5879=>"010001010",
  5880=>"110010101",
  5881=>"011001101",
  5882=>"000001010",
  5883=>"000111101",
  5884=>"101101001",
  5885=>"000011000",
  5886=>"011101000",
  5887=>"101001101",
  5888=>"011011011",
  5889=>"000011011",
  5890=>"111100010",
  5891=>"001110100",
  5892=>"010011001",
  5893=>"000000111",
  5894=>"000001101",
  5895=>"001010110",
  5896=>"000001101",
  5897=>"110101010",
  5898=>"110111001",
  5899=>"100001111",
  5900=>"000000111",
  5901=>"010011100",
  5902=>"011111100",
  5903=>"010000000",
  5904=>"010100011",
  5905=>"100101000",
  5906=>"011100111",
  5907=>"110001100",
  5908=>"111100111",
  5909=>"100011100",
  5910=>"011010001",
  5911=>"000010011",
  5912=>"001000111",
  5913=>"110110010",
  5914=>"100100100",
  5915=>"010001001",
  5916=>"000000001",
  5917=>"101101010",
  5918=>"010110101",
  5919=>"000010111",
  5920=>"000000011",
  5921=>"011101110",
  5922=>"010011101",
  5923=>"011110000",
  5924=>"111001011",
  5925=>"011011001",
  5926=>"111111110",
  5927=>"011100111",
  5928=>"011010010",
  5929=>"010001100",
  5930=>"100101000",
  5931=>"011101110",
  5932=>"111101101",
  5933=>"100010011",
  5934=>"001000101",
  5935=>"100111110",
  5936=>"100001001",
  5937=>"011100101",
  5938=>"110000100",
  5939=>"101110001",
  5940=>"101111010",
  5941=>"110101010",
  5942=>"111001110",
  5943=>"001100111",
  5944=>"100101110",
  5945=>"001110111",
  5946=>"010011111",
  5947=>"101110100",
  5948=>"110110110",
  5949=>"011101001",
  5950=>"110100000",
  5951=>"100110011",
  5952=>"010010010",
  5953=>"110010000",
  5954=>"000000110",
  5955=>"110101110",
  5956=>"111010111",
  5957=>"110010010",
  5958=>"101000101",
  5959=>"011100011",
  5960=>"101110100",
  5961=>"010111011",
  5962=>"111111100",
  5963=>"010101100",
  5964=>"001000011",
  5965=>"111110111",
  5966=>"000100011",
  5967=>"111011010",
  5968=>"000010111",
  5969=>"101111000",
  5970=>"001000100",
  5971=>"100010000",
  5972=>"011010011",
  5973=>"011000001",
  5974=>"001110010",
  5975=>"000110010",
  5976=>"111101101",
  5977=>"000110100",
  5978=>"011010110",
  5979=>"001011111",
  5980=>"000000001",
  5981=>"000001011",
  5982=>"010011011",
  5983=>"000010010",
  5984=>"001001010",
  5985=>"011000110",
  5986=>"001000010",
  5987=>"110000011",
  5988=>"010000011",
  5989=>"111101100",
  5990=>"010000011",
  5991=>"110011000",
  5992=>"001000000",
  5993=>"111010000",
  5994=>"110001111",
  5995=>"010100011",
  5996=>"101111011",
  5997=>"110011010",
  5998=>"000000010",
  5999=>"111100000",
  6000=>"010100100",
  6001=>"110101001",
  6002=>"000100011",
  6003=>"101101000",
  6004=>"000010110",
  6005=>"011000010",
  6006=>"100000000",
  6007=>"000011111",
  6008=>"000001101",
  6009=>"011000111",
  6010=>"001000101",
  6011=>"000100111",
  6012=>"001101110",
  6013=>"001111100",
  6014=>"110101001",
  6015=>"100010001",
  6016=>"101100111",
  6017=>"110111001",
  6018=>"010100111",
  6019=>"010010110",
  6020=>"000001010",
  6021=>"100101000",
  6022=>"000001011",
  6023=>"100001011",
  6024=>"011110101",
  6025=>"101001000",
  6026=>"011100001",
  6027=>"011000011",
  6028=>"010000011",
  6029=>"010011010",
  6030=>"001001011",
  6031=>"011001011",
  6032=>"111010001",
  6033=>"101111101",
  6034=>"101000011",
  6035=>"111101010",
  6036=>"000010110",
  6037=>"001000101",
  6038=>"111011001",
  6039=>"101000111",
  6040=>"001110010",
  6041=>"010010001",
  6042=>"111111010",
  6043=>"000011111",
  6044=>"011100110",
  6045=>"010101111",
  6046=>"011100001",
  6047=>"000001100",
  6048=>"111100000",
  6049=>"110100000",
  6050=>"001010110",
  6051=>"000100000",
  6052=>"000100010",
  6053=>"111010000",
  6054=>"011101001",
  6055=>"110011110",
  6056=>"101010100",
  6057=>"100101100",
  6058=>"110010111",
  6059=>"101101111",
  6060=>"100101000",
  6061=>"000001111",
  6062=>"111100000",
  6063=>"010110011",
  6064=>"010110001",
  6065=>"111100110",
  6066=>"000000000",
  6067=>"101101100",
  6068=>"001000111",
  6069=>"110011101",
  6070=>"111011100",
  6071=>"101000010",
  6072=>"110011101",
  6073=>"111111110",
  6074=>"111001010",
  6075=>"010111101",
  6076=>"101001000",
  6077=>"101000111",
  6078=>"010110101",
  6079=>"101011101",
  6080=>"010011010",
  6081=>"100111111",
  6082=>"001111111",
  6083=>"110001111",
  6084=>"000110111",
  6085=>"001001100",
  6086=>"100110100",
  6087=>"111101001",
  6088=>"000001010",
  6089=>"011110100",
  6090=>"000000010",
  6091=>"001101000",
  6092=>"010101111",
  6093=>"111100000",
  6094=>"000100001",
  6095=>"000111100",
  6096=>"011111111",
  6097=>"011101000",
  6098=>"010110100",
  6099=>"100100101",
  6100=>"110010000",
  6101=>"100000010",
  6102=>"111111110",
  6103=>"101010101",
  6104=>"100001101",
  6105=>"101101000",
  6106=>"110001000",
  6107=>"101111001",
  6108=>"110000111",
  6109=>"011010101",
  6110=>"111100010",
  6111=>"010001111",
  6112=>"111111000",
  6113=>"100010010",
  6114=>"001100101",
  6115=>"010001101",
  6116=>"001110010",
  6117=>"000010000",
  6118=>"101100010",
  6119=>"110110111",
  6120=>"110001111",
  6121=>"110010001",
  6122=>"100001011",
  6123=>"000101111",
  6124=>"101000011",
  6125=>"100011001",
  6126=>"001000000",
  6127=>"001010100",
  6128=>"101111001",
  6129=>"111110001",
  6130=>"111001001",
  6131=>"011010000",
  6132=>"110101011",
  6133=>"001000101",
  6134=>"001101010",
  6135=>"011000111",
  6136=>"001111011",
  6137=>"101110001",
  6138=>"000011000",
  6139=>"110010100",
  6140=>"111110111",
  6141=>"110001000",
  6142=>"011100111",
  6143=>"000110100",
  6144=>"111100111",
  6145=>"101011101",
  6146=>"000101011",
  6147=>"100100001",
  6148=>"001111111",
  6149=>"011010111",
  6150=>"000110010",
  6151=>"000110000",
  6152=>"100001010",
  6153=>"000100011",
  6154=>"011010111",
  6155=>"000110111",
  6156=>"010110111",
  6157=>"000010101",
  6158=>"011100010",
  6159=>"011001001",
  6160=>"100101001",
  6161=>"001001111",
  6162=>"001000101",
  6163=>"111110000",
  6164=>"011111011",
  6165=>"111111110",
  6166=>"011000101",
  6167=>"000000000",
  6168=>"111000011",
  6169=>"000001100",
  6170=>"101101110",
  6171=>"010010001",
  6172=>"000001111",
  6173=>"100001110",
  6174=>"011101000",
  6175=>"111010100",
  6176=>"001010010",
  6177=>"110101110",
  6178=>"100000100",
  6179=>"100000000",
  6180=>"111100000",
  6181=>"010001111",
  6182=>"110111100",
  6183=>"001011010",
  6184=>"111010101",
  6185=>"100100011",
  6186=>"011010101",
  6187=>"101101000",
  6188=>"100100000",
  6189=>"000101011",
  6190=>"111000010",
  6191=>"101100011",
  6192=>"011100111",
  6193=>"110010100",
  6194=>"100000001",
  6195=>"010000110",
  6196=>"111001101",
  6197=>"110010000",
  6198=>"001010010",
  6199=>"110011101",
  6200=>"111111110",
  6201=>"011111011",
  6202=>"101101101",
  6203=>"001001000",
  6204=>"110110111",
  6205=>"100110100",
  6206=>"101110100",
  6207=>"101011000",
  6208=>"000000011",
  6209=>"101101001",
  6210=>"110111010",
  6211=>"100011111",
  6212=>"100110110",
  6213=>"100010011",
  6214=>"100000110",
  6215=>"100100001",
  6216=>"000001110",
  6217=>"110110010",
  6218=>"101100010",
  6219=>"011001111",
  6220=>"001100111",
  6221=>"010001001",
  6222=>"100010110",
  6223=>"010000001",
  6224=>"010000001",
  6225=>"110100100",
  6226=>"001110111",
  6227=>"111001101",
  6228=>"100001010",
  6229=>"010110100",
  6230=>"111011001",
  6231=>"010010011",
  6232=>"001000100",
  6233=>"001000011",
  6234=>"001011000",
  6235=>"100110001",
  6236=>"111000101",
  6237=>"011101101",
  6238=>"011110100",
  6239=>"000110011",
  6240=>"101111001",
  6241=>"000011000",
  6242=>"000010101",
  6243=>"000011000",
  6244=>"011100001",
  6245=>"000011100",
  6246=>"011111001",
  6247=>"100010010",
  6248=>"011011101",
  6249=>"001101110",
  6250=>"010010101",
  6251=>"110100100",
  6252=>"010100000",
  6253=>"010001001",
  6254=>"000011111",
  6255=>"000000111",
  6256=>"101100110",
  6257=>"110000110",
  6258=>"001011010",
  6259=>"101111111",
  6260=>"000100110",
  6261=>"001010001",
  6262=>"000011110",
  6263=>"101110111",
  6264=>"000011001",
  6265=>"111010110",
  6266=>"110101110",
  6267=>"010111001",
  6268=>"001110100",
  6269=>"111100011",
  6270=>"111100100",
  6271=>"110001101",
  6272=>"101111001",
  6273=>"111101010",
  6274=>"010001010",
  6275=>"001011100",
  6276=>"001010110",
  6277=>"010010001",
  6278=>"111001101",
  6279=>"100100110",
  6280=>"001010100",
  6281=>"101100001",
  6282=>"010001101",
  6283=>"101001101",
  6284=>"001100010",
  6285=>"111010001",
  6286=>"011101000",
  6287=>"000111101",
  6288=>"000101101",
  6289=>"011111111",
  6290=>"111110011",
  6291=>"110111011",
  6292=>"111000101",
  6293=>"000110110",
  6294=>"101100110",
  6295=>"010001000",
  6296=>"000000100",
  6297=>"011011010",
  6298=>"111101101",
  6299=>"110100010",
  6300=>"000010010",
  6301=>"000001111",
  6302=>"100001100",
  6303=>"101000111",
  6304=>"111110011",
  6305=>"110101110",
  6306=>"100110010",
  6307=>"010010111",
  6308=>"011111001",
  6309=>"001001001",
  6310=>"111010110",
  6311=>"110011000",
  6312=>"101100000",
  6313=>"010000111",
  6314=>"001010100",
  6315=>"110000011",
  6316=>"000011110",
  6317=>"011000010",
  6318=>"000111100",
  6319=>"000001010",
  6320=>"011100110",
  6321=>"110101011",
  6322=>"011011000",
  6323=>"010000110",
  6324=>"100001101",
  6325=>"001101111",
  6326=>"001101101",
  6327=>"001010000",
  6328=>"110111001",
  6329=>"100000111",
  6330=>"111000100",
  6331=>"010111100",
  6332=>"000000100",
  6333=>"101111011",
  6334=>"110101000",
  6335=>"111011100",
  6336=>"101110001",
  6337=>"011101011",
  6338=>"110010001",
  6339=>"010100000",
  6340=>"111111011",
  6341=>"110110010",
  6342=>"000011110",
  6343=>"000011010",
  6344=>"111110011",
  6345=>"111101001",
  6346=>"111011100",
  6347=>"001111011",
  6348=>"101111011",
  6349=>"111111011",
  6350=>"100111111",
  6351=>"000100110",
  6352=>"011011000",
  6353=>"000100111",
  6354=>"001010111",
  6355=>"011100100",
  6356=>"010011000",
  6357=>"101110101",
  6358=>"111000110",
  6359=>"001000111",
  6360=>"100100100",
  6361=>"111111011",
  6362=>"001011010",
  6363=>"010001101",
  6364=>"010111000",
  6365=>"101110001",
  6366=>"001000010",
  6367=>"000010001",
  6368=>"011010000",
  6369=>"100111000",
  6370=>"111111000",
  6371=>"100011010",
  6372=>"001111000",
  6373=>"010101001",
  6374=>"010100101",
  6375=>"111101111",
  6376=>"000000101",
  6377=>"000110100",
  6378=>"010001111",
  6379=>"101111010",
  6380=>"110101110",
  6381=>"011110110",
  6382=>"010111011",
  6383=>"001110111",
  6384=>"000100000",
  6385=>"010111011",
  6386=>"001111001",
  6387=>"110001010",
  6388=>"110010011",
  6389=>"000011110",
  6390=>"000000101",
  6391=>"010101011",
  6392=>"001101111",
  6393=>"000111001",
  6394=>"110001111",
  6395=>"000010001",
  6396=>"001101001",
  6397=>"101101101",
  6398=>"000010101",
  6399=>"101100000",
  6400=>"000011001",
  6401=>"110110101",
  6402=>"011111110",
  6403=>"000000000",
  6404=>"011100111",
  6405=>"100011011",
  6406=>"000000001",
  6407=>"010011111",
  6408=>"011100111",
  6409=>"110110100",
  6410=>"001011100",
  6411=>"011000110",
  6412=>"011001011",
  6413=>"111000111",
  6414=>"000101000",
  6415=>"110101100",
  6416=>"011111011",
  6417=>"000010111",
  6418=>"010010001",
  6419=>"011010011",
  6420=>"110111001",
  6421=>"010010101",
  6422=>"111110110",
  6423=>"100011101",
  6424=>"011111001",
  6425=>"001101110",
  6426=>"000000101",
  6427=>"010001101",
  6428=>"000000011",
  6429=>"111111011",
  6430=>"011001001",
  6431=>"001011101",
  6432=>"101010000",
  6433=>"001011011",
  6434=>"000010010",
  6435=>"100101100",
  6436=>"111100000",
  6437=>"000001010",
  6438=>"100010010",
  6439=>"101011100",
  6440=>"111111000",
  6441=>"111000000",
  6442=>"101000011",
  6443=>"011101011",
  6444=>"011111110",
  6445=>"010011000",
  6446=>"110101111",
  6447=>"011101010",
  6448=>"001011101",
  6449=>"100000010",
  6450=>"011011110",
  6451=>"001101110",
  6452=>"110101111",
  6453=>"101110111",
  6454=>"010100001",
  6455=>"011110111",
  6456=>"001000001",
  6457=>"001010110",
  6458=>"011110101",
  6459=>"111101111",
  6460=>"110000000",
  6461=>"111011011",
  6462=>"101110101",
  6463=>"111111011",
  6464=>"110001010",
  6465=>"110000010",
  6466=>"101100000",
  6467=>"001100101",
  6468=>"111010001",
  6469=>"101100000",
  6470=>"111010110",
  6471=>"011101100",
  6472=>"000000010",
  6473=>"000110010",
  6474=>"111110110",
  6475=>"001110110",
  6476=>"001011101",
  6477=>"111011110",
  6478=>"101011100",
  6479=>"011000010",
  6480=>"000000000",
  6481=>"001100101",
  6482=>"101001110",
  6483=>"101111111",
  6484=>"010000000",
  6485=>"011010011",
  6486=>"111110100",
  6487=>"001100011",
  6488=>"000001010",
  6489=>"010010010",
  6490=>"000000101",
  6491=>"000001010",
  6492=>"011101001",
  6493=>"111111000",
  6494=>"101100011",
  6495=>"000010010",
  6496=>"000110011",
  6497=>"100100011",
  6498=>"100001110",
  6499=>"010101011",
  6500=>"011001000",
  6501=>"011101010",
  6502=>"011011101",
  6503=>"001011000",
  6504=>"000010011",
  6505=>"100001010",
  6506=>"101111101",
  6507=>"010011110",
  6508=>"110011100",
  6509=>"100001011",
  6510=>"101001010",
  6511=>"100000111",
  6512=>"001000100",
  6513=>"001010000",
  6514=>"011100110",
  6515=>"101111101",
  6516=>"101011011",
  6517=>"011110101",
  6518=>"101101001",
  6519=>"010010010",
  6520=>"000001111",
  6521=>"010101001",
  6522=>"111111110",
  6523=>"111101111",
  6524=>"101100010",
  6525=>"111110111",
  6526=>"011100011",
  6527=>"110010010",
  6528=>"010010101",
  6529=>"101100010",
  6530=>"110011011",
  6531=>"011100110",
  6532=>"101111010",
  6533=>"010101111",
  6534=>"111101011",
  6535=>"010100100",
  6536=>"101111110",
  6537=>"101001111",
  6538=>"111100111",
  6539=>"011100000",
  6540=>"101100100",
  6541=>"001111111",
  6542=>"100110100",
  6543=>"010101111",
  6544=>"010010010",
  6545=>"110011000",
  6546=>"011101101",
  6547=>"011010110",
  6548=>"110001010",
  6549=>"110001001",
  6550=>"011001111",
  6551=>"000011100",
  6552=>"011111111",
  6553=>"010101000",
  6554=>"011111101",
  6555=>"001110010",
  6556=>"100100100",
  6557=>"110110100",
  6558=>"000101101",
  6559=>"101111111",
  6560=>"100100001",
  6561=>"010110111",
  6562=>"101010000",
  6563=>"001000010",
  6564=>"001010100",
  6565=>"000101111",
  6566=>"111110110",
  6567=>"110011100",
  6568=>"001101101",
  6569=>"110010100",
  6570=>"011010110",
  6571=>"100011001",
  6572=>"101100000",
  6573=>"001101110",
  6574=>"010011110",
  6575=>"111010000",
  6576=>"110001111",
  6577=>"110110010",
  6578=>"111001110",
  6579=>"011010110",
  6580=>"010001000",
  6581=>"100110100",
  6582=>"000100001",
  6583=>"101011011",
  6584=>"101010011",
  6585=>"000110000",
  6586=>"111001100",
  6587=>"010110110",
  6588=>"101110110",
  6589=>"011000001",
  6590=>"111011111",
  6591=>"110101100",
  6592=>"100001000",
  6593=>"111111111",
  6594=>"101000100",
  6595=>"001111101",
  6596=>"111110111",
  6597=>"011010111",
  6598=>"101011101",
  6599=>"110111000",
  6600=>"010101100",
  6601=>"100011110",
  6602=>"010001010",
  6603=>"111000001",
  6604=>"011100111",
  6605=>"001011101",
  6606=>"001101101",
  6607=>"101111100",
  6608=>"110001011",
  6609=>"101110000",
  6610=>"000111100",
  6611=>"111110011",
  6612=>"110111101",
  6613=>"110010110",
  6614=>"001010100",
  6615=>"011111100",
  6616=>"010001010",
  6617=>"111110010",
  6618=>"011010111",
  6619=>"100111000",
  6620=>"010001000",
  6621=>"011011110",
  6622=>"010000000",
  6623=>"100001110",
  6624=>"010000111",
  6625=>"101011010",
  6626=>"110111000",
  6627=>"010001100",
  6628=>"100111100",
  6629=>"000001101",
  6630=>"111111101",
  6631=>"100100010",
  6632=>"001010100",
  6633=>"110011000",
  6634=>"101011101",
  6635=>"011110100",
  6636=>"010001111",
  6637=>"010110111",
  6638=>"010011100",
  6639=>"001000001",
  6640=>"100000001",
  6641=>"110100011",
  6642=>"000010111",
  6643=>"010110101",
  6644=>"110010111",
  6645=>"101110011",
  6646=>"111111100",
  6647=>"001000001",
  6648=>"000101100",
  6649=>"110100111",
  6650=>"011111011",
  6651=>"011000110",
  6652=>"000101010",
  6653=>"001000111",
  6654=>"011111011",
  6655=>"101000011",
  6656=>"000000010",
  6657=>"000010101",
  6658=>"011010110",
  6659=>"000000111",
  6660=>"100101110",
  6661=>"011001110",
  6662=>"101111110",
  6663=>"100000011",
  6664=>"010100000",
  6665=>"110001100",
  6666=>"010010001",
  6667=>"001000101",
  6668=>"111011110",
  6669=>"100000000",
  6670=>"011000100",
  6671=>"000001010",
  6672=>"100001110",
  6673=>"001001001",
  6674=>"100111011",
  6675=>"001111100",
  6676=>"110010101",
  6677=>"000001010",
  6678=>"010101110",
  6679=>"010001111",
  6680=>"101110010",
  6681=>"101001001",
  6682=>"111100011",
  6683=>"010101101",
  6684=>"110111111",
  6685=>"001111011",
  6686=>"100100000",
  6687=>"001111111",
  6688=>"100110001",
  6689=>"000100001",
  6690=>"000000000",
  6691=>"011101111",
  6692=>"001100100",
  6693=>"111011110",
  6694=>"000001100",
  6695=>"110100011",
  6696=>"010100111",
  6697=>"101010011",
  6698=>"011111111",
  6699=>"101110000",
  6700=>"010011110",
  6701=>"101000001",
  6702=>"111111110",
  6703=>"010010110",
  6704=>"111101111",
  6705=>"111111101",
  6706=>"010101010",
  6707=>"000011001",
  6708=>"010110111",
  6709=>"111101010",
  6710=>"111000101",
  6711=>"110011000",
  6712=>"111001001",
  6713=>"001000110",
  6714=>"001100100",
  6715=>"010100010",
  6716=>"000101011",
  6717=>"000011000",
  6718=>"001011110",
  6719=>"101000111",
  6720=>"100011100",
  6721=>"101000010",
  6722=>"111111110",
  6723=>"110000100",
  6724=>"110110101",
  6725=>"011001101",
  6726=>"111011000",
  6727=>"101111011",
  6728=>"110110111",
  6729=>"011101001",
  6730=>"010100000",
  6731=>"100101110",
  6732=>"011011001",
  6733=>"110111011",
  6734=>"111100110",
  6735=>"000111110",
  6736=>"011010010",
  6737=>"011001101",
  6738=>"011110001",
  6739=>"100000110",
  6740=>"001000001",
  6741=>"001001100",
  6742=>"111111000",
  6743=>"101100110",
  6744=>"000011010",
  6745=>"101011000",
  6746=>"100010011",
  6747=>"001111010",
  6748=>"100011100",
  6749=>"000000010",
  6750=>"010000110",
  6751=>"010100000",
  6752=>"101101010",
  6753=>"000000000",
  6754=>"001111010",
  6755=>"001111010",
  6756=>"111101001",
  6757=>"100111101",
  6758=>"001111001",
  6759=>"101001100",
  6760=>"000001010",
  6761=>"011001111",
  6762=>"011010111",
  6763=>"101110000",
  6764=>"100011111",
  6765=>"000000001",
  6766=>"000011111",
  6767=>"001010001",
  6768=>"011010110",
  6769=>"010101011",
  6770=>"011101111",
  6771=>"100000010",
  6772=>"000101101",
  6773=>"110011100",
  6774=>"010100011",
  6775=>"101010001",
  6776=>"010111100",
  6777=>"011100101",
  6778=>"011101101",
  6779=>"100000100",
  6780=>"010100010",
  6781=>"111010010",
  6782=>"100101110",
  6783=>"100110001",
  6784=>"001100010",
  6785=>"011110110",
  6786=>"111110101",
  6787=>"000001000",
  6788=>"011101001",
  6789=>"000111111",
  6790=>"101000110",
  6791=>"001111001",
  6792=>"000011000",
  6793=>"000101110",
  6794=>"100000110",
  6795=>"010001000",
  6796=>"101010100",
  6797=>"101010110",
  6798=>"110101001",
  6799=>"111000110",
  6800=>"100000000",
  6801=>"110111111",
  6802=>"100011000",
  6803=>"111011101",
  6804=>"100010001",
  6805=>"001001111",
  6806=>"111101111",
  6807=>"001000011",
  6808=>"000011101",
  6809=>"110010111",
  6810=>"111011110",
  6811=>"101110010",
  6812=>"010010110",
  6813=>"011100110",
  6814=>"110100101",
  6815=>"001011100",
  6816=>"010010110",
  6817=>"100110011",
  6818=>"010011011",
  6819=>"010011111",
  6820=>"101000000",
  6821=>"101110111",
  6822=>"101000001",
  6823=>"000010000",
  6824=>"001000011",
  6825=>"110000110",
  6826=>"001111111",
  6827=>"111010000",
  6828=>"001000001",
  6829=>"000100111",
  6830=>"000000000",
  6831=>"001101011",
  6832=>"101010101",
  6833=>"100110100",
  6834=>"111001110",
  6835=>"100110101",
  6836=>"111010001",
  6837=>"010110000",
  6838=>"101001001",
  6839=>"110011000",
  6840=>"010000111",
  6841=>"110111100",
  6842=>"000010010",
  6843=>"000101101",
  6844=>"100111011",
  6845=>"100011000",
  6846=>"000001100",
  6847=>"000001110",
  6848=>"010110010",
  6849=>"100101000",
  6850=>"011001101",
  6851=>"111101111",
  6852=>"000011000",
  6853=>"100110110",
  6854=>"110110110",
  6855=>"001101101",
  6856=>"001100001",
  6857=>"011010110",
  6858=>"111111101",
  6859=>"010101110",
  6860=>"110110100",
  6861=>"111101100",
  6862=>"011000001",
  6863=>"010000001",
  6864=>"010101001",
  6865=>"011011111",
  6866=>"001101100",
  6867=>"010100011",
  6868=>"100001011",
  6869=>"011011111",
  6870=>"110100110",
  6871=>"010100111",
  6872=>"100011111",
  6873=>"010101110",
  6874=>"111110101",
  6875=>"000111000",
  6876=>"000111010",
  6877=>"110111110",
  6878=>"110001100",
  6879=>"101011100",
  6880=>"000100101",
  6881=>"000000010",
  6882=>"011101010",
  6883=>"011101111",
  6884=>"010100001",
  6885=>"110011110",
  6886=>"000001011",
  6887=>"101110000",
  6888=>"111001001",
  6889=>"000000011",
  6890=>"111100001",
  6891=>"100000100",
  6892=>"111001110",
  6893=>"000101110",
  6894=>"101101000",
  6895=>"000110101",
  6896=>"101011000",
  6897=>"000010111",
  6898=>"000101001",
  6899=>"000010111",
  6900=>"100100110",
  6901=>"000110111",
  6902=>"110010111",
  6903=>"011001000",
  6904=>"000000000",
  6905=>"111000010",
  6906=>"011011011",
  6907=>"001011100",
  6908=>"100000110",
  6909=>"110111111",
  6910=>"000101100",
  6911=>"110101011",
  6912=>"000000011",
  6913=>"001101001",
  6914=>"100111111",
  6915=>"011001111",
  6916=>"001110101",
  6917=>"000011010",
  6918=>"000110011",
  6919=>"110110010",
  6920=>"100101101",
  6921=>"000111100",
  6922=>"010001101",
  6923=>"000000111",
  6924=>"111011110",
  6925=>"000011110",
  6926=>"100001110",
  6927=>"001100100",
  6928=>"011010101",
  6929=>"100110001",
  6930=>"101100000",
  6931=>"111100000",
  6932=>"111001001",
  6933=>"000001100",
  6934=>"110010110",
  6935=>"011111010",
  6936=>"000000001",
  6937=>"000001100",
  6938=>"101011101",
  6939=>"010110011",
  6940=>"100100111",
  6941=>"111000101",
  6942=>"101010100",
  6943=>"001001010",
  6944=>"100001001",
  6945=>"000010000",
  6946=>"101011111",
  6947=>"101010010",
  6948=>"100000110",
  6949=>"010000000",
  6950=>"001100111",
  6951=>"011000100",
  6952=>"111111011",
  6953=>"100101110",
  6954=>"101110001",
  6955=>"011000100",
  6956=>"010100001",
  6957=>"100101111",
  6958=>"101000000",
  6959=>"111000111",
  6960=>"000001001",
  6961=>"010100010",
  6962=>"001000111",
  6963=>"011110011",
  6964=>"101000111",
  6965=>"001001100",
  6966=>"000110101",
  6967=>"100110000",
  6968=>"110110001",
  6969=>"000000101",
  6970=>"101111101",
  6971=>"110000010",
  6972=>"100001010",
  6973=>"110101110",
  6974=>"011000011",
  6975=>"011011110",
  6976=>"000010100",
  6977=>"010101000",
  6978=>"111001100",
  6979=>"000000110",
  6980=>"111111110",
  6981=>"010110010",
  6982=>"011101100",
  6983=>"110101101",
  6984=>"010010111",
  6985=>"001110001",
  6986=>"001101101",
  6987=>"010001001",
  6988=>"100010101",
  6989=>"000110111",
  6990=>"100111100",
  6991=>"111111111",
  6992=>"110110101",
  6993=>"000100111",
  6994=>"110111010",
  6995=>"001110010",
  6996=>"100001000",
  6997=>"001000010",
  6998=>"000000000",
  6999=>"110001010",
  7000=>"011010101",
  7001=>"110011000",
  7002=>"010010111",
  7003=>"000000011",
  7004=>"101110000",
  7005=>"011011100",
  7006=>"011111000",
  7007=>"000000000",
  7008=>"110011011",
  7009=>"101100100",
  7010=>"010110101",
  7011=>"001000111",
  7012=>"110010001",
  7013=>"100110101",
  7014=>"000110111",
  7015=>"110110001",
  7016=>"100010011",
  7017=>"011010001",
  7018=>"111010001",
  7019=>"000000000",
  7020=>"010001000",
  7021=>"001110000",
  7022=>"110100101",
  7023=>"010001000",
  7024=>"111000101",
  7025=>"011111001",
  7026=>"110111101",
  7027=>"000100100",
  7028=>"100110110",
  7029=>"011111100",
  7030=>"111100110",
  7031=>"111010110",
  7032=>"101001010",
  7033=>"111010100",
  7034=>"010011011",
  7035=>"000110000",
  7036=>"000110001",
  7037=>"111101100",
  7038=>"111100100",
  7039=>"110001101",
  7040=>"001101101",
  7041=>"000111100",
  7042=>"011011001",
  7043=>"011111111",
  7044=>"101001110",
  7045=>"011101011",
  7046=>"010011011",
  7047=>"100010000",
  7048=>"100011011",
  7049=>"001110110",
  7050=>"101111001",
  7051=>"100010000",
  7052=>"000000000",
  7053=>"100010000",
  7054=>"100011011",
  7055=>"000000101",
  7056=>"101111111",
  7057=>"110000010",
  7058=>"101000001",
  7059=>"011111001",
  7060=>"001011011",
  7061=>"000001110",
  7062=>"100101101",
  7063=>"010010010",
  7064=>"110111001",
  7065=>"110011010",
  7066=>"000000111",
  7067=>"111011111",
  7068=>"001010100",
  7069=>"000000011",
  7070=>"000000000",
  7071=>"011011101",
  7072=>"001010001",
  7073=>"101011011",
  7074=>"010111111",
  7075=>"001110101",
  7076=>"010110000",
  7077=>"011001001",
  7078=>"110111111",
  7079=>"111111110",
  7080=>"000001011",
  7081=>"110011101",
  7082=>"110000001",
  7083=>"011011110",
  7084=>"101100001",
  7085=>"000011100",
  7086=>"110110101",
  7087=>"111101001",
  7088=>"000011011",
  7089=>"010101011",
  7090=>"011001011",
  7091=>"110000110",
  7092=>"100011011",
  7093=>"001101101",
  7094=>"001001011",
  7095=>"111001010",
  7096=>"111111110",
  7097=>"000011101",
  7098=>"101101010",
  7099=>"111111010",
  7100=>"011010011",
  7101=>"011000000",
  7102=>"111100100",
  7103=>"111110110",
  7104=>"111100110",
  7105=>"111011011",
  7106=>"100000001",
  7107=>"001110011",
  7108=>"111101110",
  7109=>"011110100",
  7110=>"001001001",
  7111=>"010100001",
  7112=>"110111011",
  7113=>"011110000",
  7114=>"001101001",
  7115=>"100010011",
  7116=>"011010110",
  7117=>"001001010",
  7118=>"110100110",
  7119=>"110111001",
  7120=>"110100001",
  7121=>"011001100",
  7122=>"001000110",
  7123=>"000101011",
  7124=>"100001010",
  7125=>"111000110",
  7126=>"110011111",
  7127=>"010111000",
  7128=>"100100011",
  7129=>"110001001",
  7130=>"101110000",
  7131=>"111011000",
  7132=>"110001101",
  7133=>"000010100",
  7134=>"001100101",
  7135=>"000001000",
  7136=>"000001100",
  7137=>"111101111",
  7138=>"100011110",
  7139=>"100110100",
  7140=>"100111000",
  7141=>"011110001",
  7142=>"001011111",
  7143=>"010010100",
  7144=>"001101000",
  7145=>"011010010",
  7146=>"001110101",
  7147=>"011000011",
  7148=>"101011010",
  7149=>"001010000",
  7150=>"000001001",
  7151=>"101001010",
  7152=>"010000011",
  7153=>"110111010",
  7154=>"100110011",
  7155=>"010000110",
  7156=>"000000001",
  7157=>"100011011",
  7158=>"110100011",
  7159=>"000111110",
  7160=>"010110010",
  7161=>"101001111",
  7162=>"010101000",
  7163=>"011001011",
  7164=>"111101001",
  7165=>"011110011",
  7166=>"100011001",
  7167=>"111100000",
  7168=>"010110010",
  7169=>"011010000",
  7170=>"000010101",
  7171=>"010111111",
  7172=>"100100110",
  7173=>"000001001",
  7174=>"100111100",
  7175=>"110001010",
  7176=>"101111010",
  7177=>"100001010",
  7178=>"010110001",
  7179=>"001110111",
  7180=>"101101000",
  7181=>"011001111",
  7182=>"011001100",
  7183=>"110110100",
  7184=>"101101111",
  7185=>"000010011",
  7186=>"110101010",
  7187=>"010101000",
  7188=>"111001010",
  7189=>"110101100",
  7190=>"100111000",
  7191=>"000000001",
  7192=>"000110001",
  7193=>"111101100",
  7194=>"101100010",
  7195=>"010001000",
  7196=>"101010111",
  7197=>"110001000",
  7198=>"101110110",
  7199=>"011101011",
  7200=>"010101010",
  7201=>"000000010",
  7202=>"000111001",
  7203=>"000110100",
  7204=>"010011100",
  7205=>"001000000",
  7206=>"010111001",
  7207=>"000110101",
  7208=>"100100111",
  7209=>"010011111",
  7210=>"100010110",
  7211=>"100000001",
  7212=>"110000101",
  7213=>"111111101",
  7214=>"110000011",
  7215=>"001101111",
  7216=>"100110101",
  7217=>"011011011",
  7218=>"101000000",
  7219=>"010010000",
  7220=>"010000001",
  7221=>"011000011",
  7222=>"001101110",
  7223=>"011001110",
  7224=>"111100111",
  7225=>"110101111",
  7226=>"000110101",
  7227=>"111100000",
  7228=>"000011011",
  7229=>"111110011",
  7230=>"001011111",
  7231=>"010110110",
  7232=>"100101011",
  7233=>"101001011",
  7234=>"010010000",
  7235=>"001010000",
  7236=>"010101011",
  7237=>"010100011",
  7238=>"110110001",
  7239=>"110100010",
  7240=>"001001101",
  7241=>"101010010",
  7242=>"110000100",
  7243=>"100010011",
  7244=>"001011001",
  7245=>"100110011",
  7246=>"111110011",
  7247=>"000001111",
  7248=>"101001111",
  7249=>"000110111",
  7250=>"111101010",
  7251=>"001111101",
  7252=>"101010110",
  7253=>"111011000",
  7254=>"011010111",
  7255=>"001010011",
  7256=>"100100111",
  7257=>"111111101",
  7258=>"010101111",
  7259=>"000011110",
  7260=>"111111111",
  7261=>"111110111",
  7262=>"111101001",
  7263=>"110111100",
  7264=>"000100011",
  7265=>"011101100",
  7266=>"010001010",
  7267=>"000101010",
  7268=>"000001101",
  7269=>"001001101",
  7270=>"100101000",
  7271=>"001111110",
  7272=>"100011001",
  7273=>"100000101",
  7274=>"100111101",
  7275=>"111101111",
  7276=>"101110011",
  7277=>"111001010",
  7278=>"110100000",
  7279=>"011011011",
  7280=>"000111101",
  7281=>"001101111",
  7282=>"101001011",
  7283=>"111100010",
  7284=>"110101110",
  7285=>"010011101",
  7286=>"101001111",
  7287=>"111111001",
  7288=>"001001101",
  7289=>"100101111",
  7290=>"000110111",
  7291=>"000001011",
  7292=>"101001110",
  7293=>"001011110",
  7294=>"100110000",
  7295=>"100010110",
  7296=>"100110101",
  7297=>"010111001",
  7298=>"001101100",
  7299=>"100001001",
  7300=>"111101000",
  7301=>"001101100",
  7302=>"000001010",
  7303=>"101011111",
  7304=>"011010110",
  7305=>"100110001",
  7306=>"011000001",
  7307=>"101000000",
  7308=>"000111000",
  7309=>"010000010",
  7310=>"011000110",
  7311=>"010010101",
  7312=>"010100100",
  7313=>"011111001",
  7314=>"001101111",
  7315=>"110100010",
  7316=>"010100111",
  7317=>"110000011",
  7318=>"101000111",
  7319=>"110100001",
  7320=>"011011011",
  7321=>"000111001",
  7322=>"001101111",
  7323=>"101011000",
  7324=>"001101111",
  7325=>"001010110",
  7326=>"100000000",
  7327=>"010111110",
  7328=>"000100110",
  7329=>"111000010",
  7330=>"101110001",
  7331=>"000000001",
  7332=>"100111100",
  7333=>"001110111",
  7334=>"101001110",
  7335=>"001111011",
  7336=>"001001001",
  7337=>"000001010",
  7338=>"010011111",
  7339=>"110001001",
  7340=>"101101011",
  7341=>"010111101",
  7342=>"100010000",
  7343=>"001010010",
  7344=>"111011000",
  7345=>"000111110",
  7346=>"000010110",
  7347=>"010001001",
  7348=>"110001110",
  7349=>"010111010",
  7350=>"010110101",
  7351=>"001001111",
  7352=>"110000111",
  7353=>"111111010",
  7354=>"010101110",
  7355=>"111001111",
  7356=>"100101010",
  7357=>"111111011",
  7358=>"111101110",
  7359=>"001001010",
  7360=>"001010011",
  7361=>"111110011",
  7362=>"100010001",
  7363=>"000110000",
  7364=>"011000111",
  7365=>"000100010",
  7366=>"000111011",
  7367=>"000010011",
  7368=>"111101001",
  7369=>"001010001",
  7370=>"110011101",
  7371=>"101000111",
  7372=>"111011110",
  7373=>"011011011",
  7374=>"001100000",
  7375=>"011000000",
  7376=>"000010101",
  7377=>"101001000",
  7378=>"110010001",
  7379=>"111010000",
  7380=>"000010000",
  7381=>"101001011",
  7382=>"011111110",
  7383=>"001111111",
  7384=>"101100001",
  7385=>"110000011",
  7386=>"111111010",
  7387=>"010100010",
  7388=>"001100010",
  7389=>"010011011",
  7390=>"101101110",
  7391=>"001100000",
  7392=>"001000101",
  7393=>"011000000",
  7394=>"000001010",
  7395=>"001010111",
  7396=>"001010001",
  7397=>"001010101",
  7398=>"000001000",
  7399=>"001110100",
  7400=>"100111111",
  7401=>"011011101",
  7402=>"000111110",
  7403=>"000101010",
  7404=>"100001110",
  7405=>"001011111",
  7406=>"000110111",
  7407=>"110110011",
  7408=>"111000110",
  7409=>"111101111",
  7410=>"101001000",
  7411=>"100011000",
  7412=>"001001001",
  7413=>"010110011",
  7414=>"001011001",
  7415=>"010110000",
  7416=>"001110000",
  7417=>"101000001",
  7418=>"010101011",
  7419=>"100001000",
  7420=>"111101110",
  7421=>"110110110",
  7422=>"000110101",
  7423=>"101011100",
  7424=>"100111011",
  7425=>"001010111",
  7426=>"010100111",
  7427=>"000101101",
  7428=>"000010000",
  7429=>"001001000",
  7430=>"110001110",
  7431=>"010100000",
  7432=>"000000001",
  7433=>"110111000",
  7434=>"010001011",
  7435=>"001011000",
  7436=>"101101110",
  7437=>"100010001",
  7438=>"001110111",
  7439=>"001000010",
  7440=>"110101000",
  7441=>"010111010",
  7442=>"101100010",
  7443=>"001110111",
  7444=>"011000001",
  7445=>"010000011",
  7446=>"000001111",
  7447=>"100010011",
  7448=>"100101000",
  7449=>"110100011",
  7450=>"111010111",
  7451=>"100011111",
  7452=>"110011000",
  7453=>"001000100",
  7454=>"110011101",
  7455=>"110001110",
  7456=>"010101101",
  7457=>"110110011",
  7458=>"100000011",
  7459=>"010101000",
  7460=>"111101110",
  7461=>"101110011",
  7462=>"010100111",
  7463=>"111011101",
  7464=>"110111111",
  7465=>"011100011",
  7466=>"110010111",
  7467=>"001101011",
  7468=>"111010010",
  7469=>"000001000",
  7470=>"010010000",
  7471=>"100101011",
  7472=>"110001010",
  7473=>"000101100",
  7474=>"111010010",
  7475=>"001011111",
  7476=>"100001001",
  7477=>"110010100",
  7478=>"101011011",
  7479=>"011001100",
  7480=>"110011111",
  7481=>"100001011",
  7482=>"100001010",
  7483=>"101010111",
  7484=>"010111010",
  7485=>"011111000",
  7486=>"001000100",
  7487=>"000111110",
  7488=>"100100101",
  7489=>"001100010",
  7490=>"111111111",
  7491=>"110000011",
  7492=>"001000010",
  7493=>"000010001",
  7494=>"100001101",
  7495=>"110001000",
  7496=>"001101111",
  7497=>"111110000",
  7498=>"111100010",
  7499=>"001001010",
  7500=>"111011000",
  7501=>"000000001",
  7502=>"001101011",
  7503=>"011011010",
  7504=>"101010101",
  7505=>"011100010",
  7506=>"001001111",
  7507=>"000000010",
  7508=>"110011111",
  7509=>"000000011",
  7510=>"111011000",
  7511=>"101000000",
  7512=>"101110101",
  7513=>"010111110",
  7514=>"011011010",
  7515=>"101001010",
  7516=>"011110010",
  7517=>"111001010",
  7518=>"010011111",
  7519=>"010111111",
  7520=>"111110110",
  7521=>"101000110",
  7522=>"001101011",
  7523=>"000100001",
  7524=>"010010110",
  7525=>"001001100",
  7526=>"001010100",
  7527=>"111010001",
  7528=>"010010011",
  7529=>"110011100",
  7530=>"010000000",
  7531=>"000011101",
  7532=>"101110001",
  7533=>"101100011",
  7534=>"011000110",
  7535=>"100101011",
  7536=>"000110111",
  7537=>"001111000",
  7538=>"110010010",
  7539=>"110010101",
  7540=>"000111110",
  7541=>"010100101",
  7542=>"110000001",
  7543=>"100111011",
  7544=>"101110000",
  7545=>"011110000",
  7546=>"011000110",
  7547=>"000111110",
  7548=>"101100000",
  7549=>"000111010",
  7550=>"100000000",
  7551=>"111010101",
  7552=>"100111001",
  7553=>"001011111",
  7554=>"100110111",
  7555=>"101000101",
  7556=>"000000110",
  7557=>"001101001",
  7558=>"101010001",
  7559=>"101001100",
  7560=>"000000001",
  7561=>"001000110",
  7562=>"010100001",
  7563=>"101101010",
  7564=>"000000000",
  7565=>"000001011",
  7566=>"101000000",
  7567=>"110000101",
  7568=>"100011111",
  7569=>"000100011",
  7570=>"010010100",
  7571=>"110011110",
  7572=>"101100001",
  7573=>"000000111",
  7574=>"001110101",
  7575=>"111101110",
  7576=>"101010010",
  7577=>"010000011",
  7578=>"111101011",
  7579=>"101101001",
  7580=>"011100110",
  7581=>"110101110",
  7582=>"010000001",
  7583=>"100010010",
  7584=>"010011010",
  7585=>"001110011",
  7586=>"110111011",
  7587=>"000111010",
  7588=>"100100110",
  7589=>"100100100",
  7590=>"001000101",
  7591=>"100001111",
  7592=>"100001110",
  7593=>"101101000",
  7594=>"001110001",
  7595=>"110110010",
  7596=>"101010101",
  7597=>"111111010",
  7598=>"100000100",
  7599=>"000000010",
  7600=>"101111001",
  7601=>"101001110",
  7602=>"101000101",
  7603=>"000101010",
  7604=>"011111100",
  7605=>"011110101",
  7606=>"101110011",
  7607=>"010000110",
  7608=>"100110011",
  7609=>"110000101",
  7610=>"011111111",
  7611=>"110101010",
  7612=>"001010011",
  7613=>"001000111",
  7614=>"110111011",
  7615=>"110110101",
  7616=>"000001010",
  7617=>"111111110",
  7618=>"111010110",
  7619=>"100100011",
  7620=>"000010101",
  7621=>"001110010",
  7622=>"000101000",
  7623=>"001110000",
  7624=>"001110101",
  7625=>"000011111",
  7626=>"010000000",
  7627=>"001100100",
  7628=>"100001100",
  7629=>"110001111",
  7630=>"011100000",
  7631=>"110110100",
  7632=>"011110100",
  7633=>"110000010",
  7634=>"000110001",
  7635=>"001001100",
  7636=>"100011000",
  7637=>"001111011",
  7638=>"110010101",
  7639=>"010110100",
  7640=>"100111110",
  7641=>"110101101",
  7642=>"101111100",
  7643=>"111110000",
  7644=>"111011001",
  7645=>"010111100",
  7646=>"101100100",
  7647=>"100100000",
  7648=>"010000001",
  7649=>"100010110",
  7650=>"110011100",
  7651=>"111010111",
  7652=>"001010011",
  7653=>"011111110",
  7654=>"000100001",
  7655=>"000011010",
  7656=>"000101011",
  7657=>"010011100",
  7658=>"010100100",
  7659=>"000110110",
  7660=>"100001111",
  7661=>"001000101",
  7662=>"110011000",
  7663=>"010100110",
  7664=>"101101110",
  7665=>"011000000",
  7666=>"011010011",
  7667=>"110000100",
  7668=>"111000100",
  7669=>"001011101",
  7670=>"010110000",
  7671=>"000110100",
  7672=>"011101101",
  7673=>"001101001",
  7674=>"001111011",
  7675=>"111110101",
  7676=>"001100100",
  7677=>"001110001",
  7678=>"010101001",
  7679=>"111001100",
  7680=>"011100011",
  7681=>"000010100",
  7682=>"010100110",
  7683=>"100010100",
  7684=>"111111110",
  7685=>"001110011",
  7686=>"101111001",
  7687=>"011010110",
  7688=>"011000011",
  7689=>"010000110",
  7690=>"111000100",
  7691=>"001000010",
  7692=>"010000100",
  7693=>"111110010",
  7694=>"100011100",
  7695=>"010001110",
  7696=>"011101100",
  7697=>"010110000",
  7698=>"100110100",
  7699=>"100001111",
  7700=>"111100010",
  7701=>"001010110",
  7702=>"101001011",
  7703=>"001011011",
  7704=>"110100010",
  7705=>"011110011",
  7706=>"000011111",
  7707=>"010001010",
  7708=>"101011001",
  7709=>"100001100",
  7710=>"100010010",
  7711=>"100100101",
  7712=>"011100010",
  7713=>"101010101",
  7714=>"000100001",
  7715=>"111000101",
  7716=>"110101011",
  7717=>"011101000",
  7718=>"100010011",
  7719=>"101000100",
  7720=>"011111111",
  7721=>"111110101",
  7722=>"011110111",
  7723=>"000111111",
  7724=>"000110111",
  7725=>"110111010",
  7726=>"001110100",
  7727=>"101001001",
  7728=>"110011110",
  7729=>"111100110",
  7730=>"001000100",
  7731=>"100011100",
  7732=>"000000001",
  7733=>"110010001",
  7734=>"001110111",
  7735=>"111000110",
  7736=>"111010110",
  7737=>"110001111",
  7738=>"011001110",
  7739=>"001100010",
  7740=>"111101111",
  7741=>"000111110",
  7742=>"110110001",
  7743=>"100111000",
  7744=>"101110011",
  7745=>"001000110",
  7746=>"000100001",
  7747=>"010000100",
  7748=>"001011111",
  7749=>"100010110",
  7750=>"010010101",
  7751=>"010101000",
  7752=>"110011110",
  7753=>"011001111",
  7754=>"001001011",
  7755=>"110101111",
  7756=>"001100100",
  7757=>"011100001",
  7758=>"011111110",
  7759=>"101111000",
  7760=>"011110010",
  7761=>"101000001",
  7762=>"000011100",
  7763=>"111100000",
  7764=>"110000000",
  7765=>"101000100",
  7766=>"010111000",
  7767=>"000011100",
  7768=>"011111011",
  7769=>"110000011",
  7770=>"000100110",
  7771=>"110010011",
  7772=>"011110100",
  7773=>"000100110",
  7774=>"010010101",
  7775=>"101000010",
  7776=>"111111101",
  7777=>"000101000",
  7778=>"011011101",
  7779=>"111111111",
  7780=>"010111100",
  7781=>"100010110",
  7782=>"110100001",
  7783=>"010111100",
  7784=>"010111101",
  7785=>"011000100",
  7786=>"001100001",
  7787=>"001111010",
  7788=>"011111100",
  7789=>"010011011",
  7790=>"010001101",
  7791=>"101010110",
  7792=>"000100111",
  7793=>"111111111",
  7794=>"100101100",
  7795=>"101111000",
  7796=>"001111110",
  7797=>"000000000",
  7798=>"110000100",
  7799=>"100101000",
  7800=>"001000111",
  7801=>"011010010",
  7802=>"010011100",
  7803=>"111111100",
  7804=>"011001100",
  7805=>"100101110",
  7806=>"111011110",
  7807=>"111100100",
  7808=>"011000111",
  7809=>"111010110",
  7810=>"010101001",
  7811=>"111001110",
  7812=>"100111111",
  7813=>"100011010",
  7814=>"110100100",
  7815=>"010010010",
  7816=>"001000101",
  7817=>"101100110",
  7818=>"001000110",
  7819=>"000101111",
  7820=>"100100011",
  7821=>"011110001",
  7822=>"101111111",
  7823=>"000000110",
  7824=>"000001001",
  7825=>"101100101",
  7826=>"011001011",
  7827=>"011101010",
  7828=>"000111110",
  7829=>"110100011",
  7830=>"111011001",
  7831=>"011011100",
  7832=>"101101000",
  7833=>"100100001",
  7834=>"001000111",
  7835=>"100011011",
  7836=>"100000110",
  7837=>"111111001",
  7838=>"001010111",
  7839=>"011011011",
  7840=>"100000110",
  7841=>"111101111",
  7842=>"110101011",
  7843=>"111111000",
  7844=>"001001101",
  7845=>"001101101",
  7846=>"100100001",
  7847=>"001001111",
  7848=>"111010001",
  7849=>"101100000",
  7850=>"011011011",
  7851=>"110111011",
  7852=>"011110010",
  7853=>"111000110",
  7854=>"011011010",
  7855=>"101101100",
  7856=>"101001111",
  7857=>"010110011",
  7858=>"001011111",
  7859=>"000100001",
  7860=>"001011111",
  7861=>"100100001",
  7862=>"010110110",
  7863=>"111111011",
  7864=>"101101110",
  7865=>"010001011",
  7866=>"001001111",
  7867=>"001000110",
  7868=>"100111011",
  7869=>"011110100",
  7870=>"100000101",
  7871=>"011101101",
  7872=>"111111000",
  7873=>"011101110",
  7874=>"010010110",
  7875=>"000110101",
  7876=>"001010001",
  7877=>"001000111",
  7878=>"010100101",
  7879=>"010010100",
  7880=>"001001110",
  7881=>"100111000",
  7882=>"000011011",
  7883=>"011010000",
  7884=>"001101111",
  7885=>"101111010",
  7886=>"000101111",
  7887=>"001000110",
  7888=>"100000010",
  7889=>"010111111",
  7890=>"001001010",
  7891=>"001000000",
  7892=>"100010100",
  7893=>"111100101",
  7894=>"110111110",
  7895=>"001111010",
  7896=>"000101110",
  7897=>"111110101",
  7898=>"101101011",
  7899=>"100111001",
  7900=>"110010111",
  7901=>"110100010",
  7902=>"000100001",
  7903=>"100111001",
  7904=>"010011100",
  7905=>"110000010",
  7906=>"101101110",
  7907=>"110001110",
  7908=>"101101101",
  7909=>"001001110",
  7910=>"011110001",
  7911=>"111000000",
  7912=>"010100110",
  7913=>"110110011",
  7914=>"101111001",
  7915=>"001101001",
  7916=>"001000111",
  7917=>"111101011",
  7918=>"101110101",
  7919=>"010100011",
  7920=>"011010101",
  7921=>"011101100",
  7922=>"111101111",
  7923=>"100010011",
  7924=>"000111010",
  7925=>"001100110",
  7926=>"110111100",
  7927=>"010011111",
  7928=>"110100111",
  7929=>"110001000",
  7930=>"100011001",
  7931=>"010100100",
  7932=>"010101111",
  7933=>"100101000",
  7934=>"001100000",
  7935=>"010011010",
  7936=>"000001001",
  7937=>"000111101",
  7938=>"111010000",
  7939=>"010101001",
  7940=>"110110000",
  7941=>"000000101",
  7942=>"110000100",
  7943=>"001001000",
  7944=>"101110010",
  7945=>"011010011",
  7946=>"010001000",
  7947=>"110000000",
  7948=>"000001110",
  7949=>"011011110",
  7950=>"110101110",
  7951=>"010110101",
  7952=>"010000000",
  7953=>"101010001",
  7954=>"000011111",
  7955=>"001111011",
  7956=>"110010110",
  7957=>"001100010",
  7958=>"001100101",
  7959=>"011001000",
  7960=>"111101101",
  7961=>"000011000",
  7962=>"010000000",
  7963=>"111000001",
  7964=>"111010000",
  7965=>"100110001",
  7966=>"100100110",
  7967=>"011001011",
  7968=>"111110110",
  7969=>"100110110",
  7970=>"000101000",
  7971=>"111101101",
  7972=>"010010000",
  7973=>"010100100",
  7974=>"111000011",
  7975=>"110011110",
  7976=>"000010010",
  7977=>"011100000",
  7978=>"110111111",
  7979=>"001011101",
  7980=>"010011001",
  7981=>"010000001",
  7982=>"011000111",
  7983=>"100011011",
  7984=>"000110011",
  7985=>"100011000",
  7986=>"101111100",
  7987=>"001010001",
  7988=>"011010000",
  7989=>"011011100",
  7990=>"001000011",
  7991=>"000010110",
  7992=>"011100000",
  7993=>"111001100",
  7994=>"001111001",
  7995=>"000100110",
  7996=>"101011101",
  7997=>"000101000",
  7998=>"000111111",
  7999=>"011001101",
  8000=>"001111100",
  8001=>"000111111",
  8002=>"011110100",
  8003=>"100001000",
  8004=>"000011010",
  8005=>"110100110",
  8006=>"110101110",
  8007=>"010010101",
  8008=>"000100110",
  8009=>"000000000",
  8010=>"010011101",
  8011=>"111100010",
  8012=>"110111110",
  8013=>"100000010",
  8014=>"001000100",
  8015=>"010001010",
  8016=>"111000001",
  8017=>"000011011",
  8018=>"011110001",
  8019=>"001001000",
  8020=>"111100111",
  8021=>"001001001",
  8022=>"100011110",
  8023=>"100111000",
  8024=>"001010000",
  8025=>"110001110",
  8026=>"011000110",
  8027=>"100001000",
  8028=>"111110010",
  8029=>"101100111",
  8030=>"000010101",
  8031=>"000110011",
  8032=>"011011000",
  8033=>"111011010",
  8034=>"001110000",
  8035=>"111111111",
  8036=>"010011000",
  8037=>"110010110",
  8038=>"100001011",
  8039=>"100111111",
  8040=>"000011100",
  8041=>"000010110",
  8042=>"110010100",
  8043=>"011001011",
  8044=>"001100110",
  8045=>"000100110",
  8046=>"011010001",
  8047=>"010011101",
  8048=>"000011110",
  8049=>"011001011",
  8050=>"011000110",
  8051=>"111101001",
  8052=>"010010000",
  8053=>"111010001",
  8054=>"110111011",
  8055=>"001101011",
  8056=>"000001111",
  8057=>"001110001",
  8058=>"111001000",
  8059=>"100010011",
  8060=>"010101011",
  8061=>"010010010",
  8062=>"100011000",
  8063=>"110011001",
  8064=>"101111101",
  8065=>"100010100",
  8066=>"000000110",
  8067=>"000000010",
  8068=>"100000000",
  8069=>"100100100",
  8070=>"010000111",
  8071=>"011010111",
  8072=>"100011111",
  8073=>"111011101",
  8074=>"110101011",
  8075=>"001100100",
  8076=>"011010000",
  8077=>"010000111",
  8078=>"101111110",
  8079=>"111101001",
  8080=>"101101111",
  8081=>"000110111",
  8082=>"100010100",
  8083=>"011101110",
  8084=>"011110010",
  8085=>"011011111",
  8086=>"010101010",
  8087=>"101101101",
  8088=>"100100111",
  8089=>"111001000",
  8090=>"010000000",
  8091=>"000111110",
  8092=>"111101101",
  8093=>"010100001",
  8094=>"000000010",
  8095=>"100100111",
  8096=>"000001101",
  8097=>"111111111",
  8098=>"101000001",
  8099=>"101010101",
  8100=>"000011110",
  8101=>"001001000",
  8102=>"000101111",
  8103=>"010000000",
  8104=>"001110001",
  8105=>"001000010",
  8106=>"100100101",
  8107=>"110100000",
  8108=>"110111110",
  8109=>"000101110",
  8110=>"010100110",
  8111=>"000010101",
  8112=>"110100101",
  8113=>"010110010",
  8114=>"001011101",
  8115=>"100111010",
  8116=>"010111011",
  8117=>"010011101",
  8118=>"101011000",
  8119=>"011010010",
  8120=>"110011101",
  8121=>"010100010",
  8122=>"001110100",
  8123=>"011111111",
  8124=>"001001010",
  8125=>"110101010",
  8126=>"111101000",
  8127=>"000011101",
  8128=>"000000100",
  8129=>"000110100",
  8130=>"011001001",
  8131=>"001111000",
  8132=>"010100010",
  8133=>"011011101",
  8134=>"110111100",
  8135=>"010000010",
  8136=>"100101000",
  8137=>"101100111",
  8138=>"000001110",
  8139=>"111010110",
  8140=>"001110110",
  8141=>"110110100",
  8142=>"111101100",
  8143=>"111011111",
  8144=>"100010010",
  8145=>"100101100",
  8146=>"011110010",
  8147=>"001001101",
  8148=>"110110010",
  8149=>"100100001",
  8150=>"010111001",
  8151=>"010010011",
  8152=>"110111010",
  8153=>"010000010",
  8154=>"100000101",
  8155=>"101110000",
  8156=>"111001110",
  8157=>"111000000",
  8158=>"111011000",
  8159=>"100101001",
  8160=>"100000000",
  8161=>"001101010",
  8162=>"011101111",
  8163=>"001001101",
  8164=>"000111000",
  8165=>"110011000",
  8166=>"000110011",
  8167=>"000001000",
  8168=>"100001111",
  8169=>"000100111",
  8170=>"111011000",
  8171=>"100001011",
  8172=>"000111011",
  8173=>"001100010",
  8174=>"010010110",
  8175=>"100001100",
  8176=>"000001001",
  8177=>"000011110",
  8178=>"101101110",
  8179=>"001000000",
  8180=>"011110100",
  8181=>"010111101",
  8182=>"010111100",
  8183=>"111111010",
  8184=>"001010110",
  8185=>"000011111",
  8186=>"001010001",
  8187=>"001100011",
  8188=>"100000111",
  8189=>"101011011",
  8190=>"111000110",
  8191=>"000100001",
  8192=>"011001110",
  8193=>"111000011",
  8194=>"010110110",
  8195=>"010100011",
  8196=>"010100000",
  8197=>"100011110",
  8198=>"001001101",
  8199=>"110001111",
  8200=>"000111000",
  8201=>"100110001",
  8202=>"011111001",
  8203=>"111111110",
  8204=>"011000101",
  8205=>"011101111",
  8206=>"000110001",
  8207=>"101101010",
  8208=>"010110110",
  8209=>"100010000",
  8210=>"111010101",
  8211=>"111111010",
  8212=>"111110101",
  8213=>"110100110",
  8214=>"101010010",
  8215=>"111101000",
  8216=>"100111000",
  8217=>"111110011",
  8218=>"000000001",
  8219=>"010110100",
  8220=>"101011111",
  8221=>"111101100",
  8222=>"011100001",
  8223=>"010111111",
  8224=>"000101100",
  8225=>"011110010",
  8226=>"110101100",
  8227=>"101000110",
  8228=>"010001110",
  8229=>"100010000",
  8230=>"000110100",
  8231=>"110001111",
  8232=>"001011000",
  8233=>"010111010",
  8234=>"011001011",
  8235=>"111111001",
  8236=>"111010110",
  8237=>"010011000",
  8238=>"001001111",
  8239=>"100101101",
  8240=>"111010101",
  8241=>"011001110",
  8242=>"011010010",
  8243=>"000100010",
  8244=>"101000011",
  8245=>"100000101",
  8246=>"100001000",
  8247=>"101000111",
  8248=>"101000101",
  8249=>"001101000",
  8250=>"010010010",
  8251=>"111010101",
  8252=>"001111001",
  8253=>"011111000",
  8254=>"011100000",
  8255=>"101101001",
  8256=>"010111111",
  8257=>"010011011",
  8258=>"100100011",
  8259=>"000101011",
  8260=>"010011001",
  8261=>"001101010",
  8262=>"111011010",
  8263=>"110010010",
  8264=>"000001101",
  8265=>"101100011",
  8266=>"010111101",
  8267=>"011101100",
  8268=>"100010001",
  8269=>"001000000",
  8270=>"010101011",
  8271=>"010100111",
  8272=>"110000101",
  8273=>"000001001",
  8274=>"110101110",
  8275=>"101111100",
  8276=>"001010010",
  8277=>"010101000",
  8278=>"001111000",
  8279=>"101000011",
  8280=>"011100111",
  8281=>"111100011",
  8282=>"000110000",
  8283=>"001011001",
  8284=>"001110111",
  8285=>"100001111",
  8286=>"001011000",
  8287=>"100110100",
  8288=>"010011101",
  8289=>"011010111",
  8290=>"000100111",
  8291=>"011101110",
  8292=>"000001101",
  8293=>"101111111",
  8294=>"000110000",
  8295=>"001001111",
  8296=>"001001101",
  8297=>"001000111",
  8298=>"100000111",
  8299=>"000111110",
  8300=>"000110110",
  8301=>"101100000",
  8302=>"001001010",
  8303=>"001010001",
  8304=>"101000000",
  8305=>"001010001",
  8306=>"010100101",
  8307=>"001101001",
  8308=>"001010100",
  8309=>"010100000",
  8310=>"001000100",
  8311=>"000011010",
  8312=>"011101111",
  8313=>"101010000",
  8314=>"000010110",
  8315=>"001101111",
  8316=>"000001110",
  8317=>"001001111",
  8318=>"000010010",
  8319=>"111011010",
  8320=>"111111000",
  8321=>"001100000",
  8322=>"010001011",
  8323=>"101100110",
  8324=>"111101111",
  8325=>"000001110",
  8326=>"111011111",
  8327=>"101111001",
  8328=>"101101100",
  8329=>"111001001",
  8330=>"110010011",
  8331=>"110110110",
  8332=>"011000101",
  8333=>"010101000",
  8334=>"111011101",
  8335=>"000011000",
  8336=>"010110111",
  8337=>"100001010",
  8338=>"111000110",
  8339=>"010001101",
  8340=>"010111100",
  8341=>"100100000",
  8342=>"100110011",
  8343=>"111111011",
  8344=>"111001010",
  8345=>"110101010",
  8346=>"010100100",
  8347=>"111100010",
  8348=>"010001000",
  8349=>"001111000",
  8350=>"100111000",
  8351=>"110000010",
  8352=>"011111001",
  8353=>"011001011",
  8354=>"000000001",
  8355=>"010100010",
  8356=>"101100011",
  8357=>"101100101",
  8358=>"001011001",
  8359=>"011101010",
  8360=>"110110000",
  8361=>"001110110",
  8362=>"111010111",
  8363=>"100001011",
  8364=>"000111110",
  8365=>"100111111",
  8366=>"011110010",
  8367=>"100111110",
  8368=>"101111111",
  8369=>"001000000",
  8370=>"000100000",
  8371=>"001111001",
  8372=>"001011100",
  8373=>"000011000",
  8374=>"100111110",
  8375=>"110101000",
  8376=>"100101110",
  8377=>"011010111",
  8378=>"000110001",
  8379=>"110110110",
  8380=>"110000100",
  8381=>"111111011",
  8382=>"110001000",
  8383=>"111110011",
  8384=>"000001111",
  8385=>"100011100",
  8386=>"110000011",
  8387=>"100001110",
  8388=>"001110001",
  8389=>"111011111",
  8390=>"000001010",
  8391=>"001010011",
  8392=>"011101110",
  8393=>"011110000",
  8394=>"001010011",
  8395=>"010111111",
  8396=>"011111010",
  8397=>"001000011",
  8398=>"010010011",
  8399=>"000011001",
  8400=>"011110000",
  8401=>"000111011",
  8402=>"011000110",
  8403=>"000100011",
  8404=>"101010011",
  8405=>"110010001",
  8406=>"110110011",
  8407=>"100011010",
  8408=>"000100000",
  8409=>"110001101",
  8410=>"111101001",
  8411=>"100001000",
  8412=>"010001010",
  8413=>"111010111",
  8414=>"101000101",
  8415=>"101000001",
  8416=>"001000001",
  8417=>"000110000",
  8418=>"101111001",
  8419=>"100000100",
  8420=>"001001100",
  8421=>"111010000",
  8422=>"111110111",
  8423=>"111010001",
  8424=>"011111000",
  8425=>"101100010",
  8426=>"111001001",
  8427=>"101001001",
  8428=>"111000001",
  8429=>"111101111",
  8430=>"101011000",
  8431=>"111110111",
  8432=>"101110000",
  8433=>"011000001",
  8434=>"110100111",
  8435=>"001101010",
  8436=>"111011101",
  8437=>"110101110",
  8438=>"001000100",
  8439=>"110111111",
  8440=>"111111101",
  8441=>"110111010",
  8442=>"110010010",
  8443=>"111001010",
  8444=>"101101111",
  8445=>"100001111",
  8446=>"011000001",
  8447=>"110101001",
  8448=>"010001011",
  8449=>"110110001",
  8450=>"100011010",
  8451=>"011111011",
  8452=>"001000110",
  8453=>"010111010",
  8454=>"010111011",
  8455=>"111101001",
  8456=>"010000100",
  8457=>"010111001",
  8458=>"001111011",
  8459=>"001010110",
  8460=>"000011110",
  8461=>"111111111",
  8462=>"100101101",
  8463=>"010101111",
  8464=>"100110000",
  8465=>"001001101",
  8466=>"100001100",
  8467=>"001011011",
  8468=>"000011000",
  8469=>"011010010",
  8470=>"011001101",
  8471=>"100111100",
  8472=>"110110011",
  8473=>"110000000",
  8474=>"001100111",
  8475=>"000001100",
  8476=>"110000110",
  8477=>"011010000",
  8478=>"001010001",
  8479=>"100000001",
  8480=>"010110000",
  8481=>"111110111",
  8482=>"111101100",
  8483=>"010000100",
  8484=>"001000010",
  8485=>"011100110",
  8486=>"011110001",
  8487=>"101000110",
  8488=>"011000110",
  8489=>"010001001",
  8490=>"000000001",
  8491=>"100100000",
  8492=>"000101010",
  8493=>"000001010",
  8494=>"010111011",
  8495=>"000111011",
  8496=>"010010010",
  8497=>"111011000",
  8498=>"000011010",
  8499=>"111110010",
  8500=>"101001100",
  8501=>"110111011",
  8502=>"101100010",
  8503=>"111110010",
  8504=>"000011101",
  8505=>"111011101",
  8506=>"101111100",
  8507=>"111010011",
  8508=>"000100101",
  8509=>"011011100",
  8510=>"001000001",
  8511=>"011100101",
  8512=>"101011000",
  8513=>"010110101",
  8514=>"100100100",
  8515=>"100101011",
  8516=>"101000000",
  8517=>"110111111",
  8518=>"000000101",
  8519=>"111010010",
  8520=>"101001101",
  8521=>"010011000",
  8522=>"000111100",
  8523=>"010101111",
  8524=>"111000110",
  8525=>"101001001",
  8526=>"110001111",
  8527=>"111110010",
  8528=>"101111110",
  8529=>"010110100",
  8530=>"111010100",
  8531=>"100001011",
  8532=>"101010010",
  8533=>"000000011",
  8534=>"011000000",
  8535=>"100001000",
  8536=>"100111100",
  8537=>"101101110",
  8538=>"101011010",
  8539=>"101110011",
  8540=>"111110101",
  8541=>"010110010",
  8542=>"101010110",
  8543=>"101010001",
  8544=>"010101111",
  8545=>"010010010",
  8546=>"110000110",
  8547=>"101111100",
  8548=>"000000111",
  8549=>"011010111",
  8550=>"000001000",
  8551=>"010001101",
  8552=>"110111100",
  8553=>"010111110",
  8554=>"000010100",
  8555=>"110001001",
  8556=>"001100111",
  8557=>"101100011",
  8558=>"011011110",
  8559=>"001111101",
  8560=>"111011000",
  8561=>"001110011",
  8562=>"111001101",
  8563=>"011001011",
  8564=>"001010011",
  8565=>"010110101",
  8566=>"101010101",
  8567=>"100001001",
  8568=>"110000100",
  8569=>"111011100",
  8570=>"010111001",
  8571=>"000110010",
  8572=>"111101101",
  8573=>"001001101",
  8574=>"001111001",
  8575=>"000100000",
  8576=>"011110111",
  8577=>"100000001",
  8578=>"000111010",
  8579=>"010110010",
  8580=>"100001011",
  8581=>"110110000",
  8582=>"011000100",
  8583=>"011000110",
  8584=>"001001100",
  8585=>"101001111",
  8586=>"011000001",
  8587=>"011011000",
  8588=>"010111011",
  8589=>"010010101",
  8590=>"001011000",
  8591=>"110111110",
  8592=>"011000000",
  8593=>"000111010",
  8594=>"010011111",
  8595=>"010110111",
  8596=>"101111111",
  8597=>"010000011",
  8598=>"000010100",
  8599=>"110000000",
  8600=>"110100110",
  8601=>"111000001",
  8602=>"011011010",
  8603=>"000011011",
  8604=>"001111101",
  8605=>"101000011",
  8606=>"111001011",
  8607=>"110000011",
  8608=>"110000001",
  8609=>"110100011",
  8610=>"000110100",
  8611=>"000100010",
  8612=>"101001110",
  8613=>"011111011",
  8614=>"011110110",
  8615=>"110000010",
  8616=>"110011001",
  8617=>"001100010",
  8618=>"101000011",
  8619=>"000101100",
  8620=>"101100101",
  8621=>"101100111",
  8622=>"011101101",
  8623=>"000100101",
  8624=>"111000000",
  8625=>"000001100",
  8626=>"110110010",
  8627=>"000010000",
  8628=>"010000101",
  8629=>"101111110",
  8630=>"001111001",
  8631=>"101011000",
  8632=>"110110110",
  8633=>"011100101",
  8634=>"010101100",
  8635=>"110110000",
  8636=>"100001010",
  8637=>"010001010",
  8638=>"011001100",
  8639=>"101001000",
  8640=>"010011011",
  8641=>"101101111",
  8642=>"001100110",
  8643=>"111100101",
  8644=>"011001000",
  8645=>"100110100",
  8646=>"000011010",
  8647=>"000010100",
  8648=>"111010110",
  8649=>"111011001",
  8650=>"000011111",
  8651=>"110001010",
  8652=>"011011111",
  8653=>"111101000",
  8654=>"010001010",
  8655=>"010101101",
  8656=>"001101101",
  8657=>"000000011",
  8658=>"001100101",
  8659=>"001000101",
  8660=>"101001110",
  8661=>"000110101",
  8662=>"000110111",
  8663=>"101000000",
  8664=>"000100101",
  8665=>"110000011",
  8666=>"101001000",
  8667=>"010010001",
  8668=>"100010100",
  8669=>"010101101",
  8670=>"101110110",
  8671=>"111100110",
  8672=>"100000011",
  8673=>"001000000",
  8674=>"000011000",
  8675=>"111101010",
  8676=>"010011010",
  8677=>"110011000",
  8678=>"000011010",
  8679=>"111101011",
  8680=>"010001111",
  8681=>"111101011",
  8682=>"011010010",
  8683=>"111001000",
  8684=>"010100000",
  8685=>"001011110",
  8686=>"101011111",
  8687=>"001110111",
  8688=>"111111010",
  8689=>"100000001",
  8690=>"111111111",
  8691=>"010001110",
  8692=>"000100100",
  8693=>"111010001",
  8694=>"011011001",
  8695=>"100111101",
  8696=>"011111101",
  8697=>"011100100",
  8698=>"000110010",
  8699=>"110100011",
  8700=>"010110010",
  8701=>"000000100",
  8702=>"000001100",
  8703=>"000101010",
  8704=>"010010011",
  8705=>"110101100",
  8706=>"100101011",
  8707=>"110010001",
  8708=>"001010111",
  8709=>"100100000",
  8710=>"100010000",
  8711=>"100010000",
  8712=>"100011000",
  8713=>"010000100",
  8714=>"101101001",
  8715=>"010010100",
  8716=>"110010001",
  8717=>"100011011",
  8718=>"010100010",
  8719=>"110110011",
  8720=>"011111001",
  8721=>"111011011",
  8722=>"111100001",
  8723=>"000110111",
  8724=>"100100010",
  8725=>"001001110",
  8726=>"011110011",
  8727=>"001110001",
  8728=>"110110110",
  8729=>"110000101",
  8730=>"111001001",
  8731=>"000011011",
  8732=>"111000001",
  8733=>"101000100",
  8734=>"110101100",
  8735=>"110001100",
  8736=>"010111111",
  8737=>"011100100",
  8738=>"010000100",
  8739=>"101001110",
  8740=>"101100011",
  8741=>"011001110",
  8742=>"010011001",
  8743=>"101001110",
  8744=>"000101111",
  8745=>"011110000",
  8746=>"100001111",
  8747=>"101101100",
  8748=>"011000000",
  8749=>"000001100",
  8750=>"111001010",
  8751=>"110000110",
  8752=>"001100011",
  8753=>"010001000",
  8754=>"000111010",
  8755=>"011101000",
  8756=>"110111111",
  8757=>"101111000",
  8758=>"101101110",
  8759=>"100111101",
  8760=>"111101000",
  8761=>"000000111",
  8762=>"001000110",
  8763=>"010101010",
  8764=>"110000011",
  8765=>"000011001",
  8766=>"101110011",
  8767=>"000000001",
  8768=>"110001111",
  8769=>"101100010",
  8770=>"011010001",
  8771=>"101010111",
  8772=>"110001011",
  8773=>"010000100",
  8774=>"110001100",
  8775=>"010101111",
  8776=>"000000101",
  8777=>"111010111",
  8778=>"010111100",
  8779=>"000010111",
  8780=>"101100011",
  8781=>"001001001",
  8782=>"011000010",
  8783=>"100100101",
  8784=>"110101100",
  8785=>"010110101",
  8786=>"110000101",
  8787=>"010011110",
  8788=>"000111011",
  8789=>"010100011",
  8790=>"001111001",
  8791=>"111000000",
  8792=>"001000001",
  8793=>"111010010",
  8794=>"110111110",
  8795=>"101101011",
  8796=>"100101111",
  8797=>"101100000",
  8798=>"010000110",
  8799=>"001000001",
  8800=>"011111011",
  8801=>"010010000",
  8802=>"100111111",
  8803=>"000101010",
  8804=>"110100000",
  8805=>"000000100",
  8806=>"111001011",
  8807=>"011111010",
  8808=>"010010101",
  8809=>"000010101",
  8810=>"110110000",
  8811=>"011000000",
  8812=>"011011001",
  8813=>"101110111",
  8814=>"110110100",
  8815=>"001100110",
  8816=>"000110101",
  8817=>"100001101",
  8818=>"111100111",
  8819=>"000011000",
  8820=>"000110001",
  8821=>"000100110",
  8822=>"111111010",
  8823=>"011110111",
  8824=>"011110110",
  8825=>"000000101",
  8826=>"000010100",
  8827=>"111111101",
  8828=>"010011100",
  8829=>"010111000",
  8830=>"011010011",
  8831=>"001101011",
  8832=>"010011111",
  8833=>"111001011",
  8834=>"000001000",
  8835=>"101001111",
  8836=>"100010000",
  8837=>"000110010",
  8838=>"011011000",
  8839=>"111111111",
  8840=>"010010101",
  8841=>"011111001",
  8842=>"001011101",
  8843=>"100101111",
  8844=>"101111010",
  8845=>"101001010",
  8846=>"000010011",
  8847=>"010110111",
  8848=>"010111000",
  8849=>"100011001",
  8850=>"101001001",
  8851=>"011110010",
  8852=>"010011100",
  8853=>"110111010",
  8854=>"111010100",
  8855=>"111110101",
  8856=>"100110011",
  8857=>"101100111",
  8858=>"010110000",
  8859=>"100010110",
  8860=>"011010110",
  8861=>"111010001",
  8862=>"110100101",
  8863=>"010101010",
  8864=>"011110000",
  8865=>"110100110",
  8866=>"010001011",
  8867=>"101100100",
  8868=>"110001011",
  8869=>"011000011",
  8870=>"101111110",
  8871=>"000111110",
  8872=>"100111000",
  8873=>"101001011",
  8874=>"111100000",
  8875=>"011001000",
  8876=>"001000010",
  8877=>"010010100",
  8878=>"110110111",
  8879=>"001110101",
  8880=>"000000111",
  8881=>"011011000",
  8882=>"110100000",
  8883=>"000100010",
  8884=>"000000101",
  8885=>"110010001",
  8886=>"101111110",
  8887=>"011001111",
  8888=>"110100001",
  8889=>"010101000",
  8890=>"000010111",
  8891=>"010011111",
  8892=>"010011010",
  8893=>"110111000",
  8894=>"010000001",
  8895=>"001000000",
  8896=>"000111111",
  8897=>"111111001",
  8898=>"010000100",
  8899=>"100101110",
  8900=>"110101101",
  8901=>"000010010",
  8902=>"000101000",
  8903=>"101011000",
  8904=>"010011001",
  8905=>"000111100",
  8906=>"101111111",
  8907=>"000101001",
  8908=>"101110011",
  8909=>"101000000",
  8910=>"010010000",
  8911=>"100000000",
  8912=>"101000010",
  8913=>"000000001",
  8914=>"000100100",
  8915=>"110101110",
  8916=>"000000110",
  8917=>"001110111",
  8918=>"101111010",
  8919=>"000000001",
  8920=>"000101010",
  8921=>"101000100",
  8922=>"101110110",
  8923=>"001010010",
  8924=>"100010111",
  8925=>"011000001",
  8926=>"001100111",
  8927=>"011000110",
  8928=>"110011011",
  8929=>"011101011",
  8930=>"001001110",
  8931=>"011000000",
  8932=>"100100110",
  8933=>"000011011",
  8934=>"101110100",
  8935=>"010000100",
  8936=>"110100100",
  8937=>"001001110",
  8938=>"110111100",
  8939=>"110001011",
  8940=>"110110100",
  8941=>"000000110",
  8942=>"100000101",
  8943=>"111010000",
  8944=>"110000101",
  8945=>"101011100",
  8946=>"111011111",
  8947=>"100100011",
  8948=>"001101000",
  8949=>"010101011",
  8950=>"101111010",
  8951=>"010100111",
  8952=>"001100001",
  8953=>"010101100",
  8954=>"101001001",
  8955=>"010001100",
  8956=>"001100000",
  8957=>"000111010",
  8958=>"011100000",
  8959=>"000011000",
  8960=>"001011100",
  8961=>"110100011",
  8962=>"100001110",
  8963=>"111010100",
  8964=>"101011011",
  8965=>"000001011",
  8966=>"111000100",
  8967=>"011011111",
  8968=>"101011110",
  8969=>"101000001",
  8970=>"001101000",
  8971=>"000011000",
  8972=>"001111101",
  8973=>"001111100",
  8974=>"011110110",
  8975=>"111101000",
  8976=>"110001010",
  8977=>"001000000",
  8978=>"100110010",
  8979=>"110110110",
  8980=>"001100001",
  8981=>"100010010",
  8982=>"111111011",
  8983=>"001011001",
  8984=>"110001101",
  8985=>"101011100",
  8986=>"100001100",
  8987=>"111011100",
  8988=>"101001001",
  8989=>"110101111",
  8990=>"010100101",
  8991=>"001001010",
  8992=>"001110111",
  8993=>"010010111",
  8994=>"100100111",
  8995=>"010110000",
  8996=>"101111111",
  8997=>"100000001",
  8998=>"010111001",
  8999=>"111000101",
  9000=>"111111101",
  9001=>"000100011",
  9002=>"010100111",
  9003=>"001101000",
  9004=>"101101111",
  9005=>"110000101",
  9006=>"000100111",
  9007=>"010110111",
  9008=>"100100011",
  9009=>"111010101",
  9010=>"111111100",
  9011=>"011010100",
  9012=>"100111000",
  9013=>"100010101",
  9014=>"001001010",
  9015=>"010110100",
  9016=>"011111111",
  9017=>"000110001",
  9018=>"101000101",
  9019=>"110111000",
  9020=>"000101001",
  9021=>"101010111",
  9022=>"000001010",
  9023=>"100000001",
  9024=>"101001100",
  9025=>"100010111",
  9026=>"011011011",
  9027=>"011100110",
  9028=>"001100010",
  9029=>"001001100",
  9030=>"011011110",
  9031=>"011100100",
  9032=>"101010111",
  9033=>"111110110",
  9034=>"110101111",
  9035=>"100000001",
  9036=>"001110100",
  9037=>"000011100",
  9038=>"010011000",
  9039=>"101111011",
  9040=>"110010011",
  9041=>"111011001",
  9042=>"011010100",
  9043=>"110011010",
  9044=>"110011001",
  9045=>"011111110",
  9046=>"110001000",
  9047=>"011001001",
  9048=>"001010000",
  9049=>"110111100",
  9050=>"111011100",
  9051=>"101000101",
  9052=>"000010010",
  9053=>"010111101",
  9054=>"001010101",
  9055=>"011001111",
  9056=>"111100110",
  9057=>"100000011",
  9058=>"001111101",
  9059=>"110110011",
  9060=>"010001110",
  9061=>"111010010",
  9062=>"000010101",
  9063=>"111011011",
  9064=>"101010010",
  9065=>"011000000",
  9066=>"111001001",
  9067=>"000010100",
  9068=>"101111111",
  9069=>"000001000",
  9070=>"011111011",
  9071=>"101001000",
  9072=>"101011001",
  9073=>"100101100",
  9074=>"000101111",
  9075=>"111100011",
  9076=>"001100100",
  9077=>"001100111",
  9078=>"000111111",
  9079=>"111101010",
  9080=>"111100011",
  9081=>"111011010",
  9082=>"101101001",
  9083=>"101001110",
  9084=>"000110010",
  9085=>"010111000",
  9086=>"000101111",
  9087=>"101100101",
  9088=>"011111100",
  9089=>"111110011",
  9090=>"010000011",
  9091=>"000001001",
  9092=>"101010110",
  9093=>"001000000",
  9094=>"100010111",
  9095=>"011001101",
  9096=>"010010011",
  9097=>"110010000",
  9098=>"100001001",
  9099=>"111101100",
  9100=>"011101111",
  9101=>"001111101",
  9102=>"000100010",
  9103=>"111111111",
  9104=>"000101011",
  9105=>"100011001",
  9106=>"011010111",
  9107=>"111000111",
  9108=>"011000011",
  9109=>"110101111",
  9110=>"100001000",
  9111=>"000011110",
  9112=>"101011001",
  9113=>"011011111",
  9114=>"010001001",
  9115=>"001011000",
  9116=>"011111111",
  9117=>"111011111",
  9118=>"011001100",
  9119=>"111101100",
  9120=>"110001000",
  9121=>"111100000",
  9122=>"101111101",
  9123=>"110010101",
  9124=>"010111010",
  9125=>"100011111",
  9126=>"000010101",
  9127=>"110111101",
  9128=>"000101000",
  9129=>"101111110",
  9130=>"010100001",
  9131=>"110101011",
  9132=>"110111010",
  9133=>"110011110",
  9134=>"010000001",
  9135=>"101111011",
  9136=>"100111010",
  9137=>"101010000",
  9138=>"010111101",
  9139=>"000110010",
  9140=>"110010111",
  9141=>"111100101",
  9142=>"010010010",
  9143=>"100101111",
  9144=>"010110100",
  9145=>"111111111",
  9146=>"001011110",
  9147=>"010101001",
  9148=>"111110101",
  9149=>"110000100",
  9150=>"010000111",
  9151=>"111010000",
  9152=>"011101111",
  9153=>"010111110",
  9154=>"001111001",
  9155=>"001100111",
  9156=>"000101000",
  9157=>"000000110",
  9158=>"110000000",
  9159=>"110011110",
  9160=>"010100000",
  9161=>"000010100",
  9162=>"111000010",
  9163=>"010000000",
  9164=>"100011111",
  9165=>"001100000",
  9166=>"111010100",
  9167=>"010010110",
  9168=>"111010100",
  9169=>"011000010",
  9170=>"111110011",
  9171=>"111000101",
  9172=>"000111100",
  9173=>"001010111",
  9174=>"101101101",
  9175=>"000100110",
  9176=>"100111101",
  9177=>"010011001",
  9178=>"110110110",
  9179=>"111110111",
  9180=>"001111010",
  9181=>"010010101",
  9182=>"110100011",
  9183=>"000010000",
  9184=>"110010011",
  9185=>"101011011",
  9186=>"000011001",
  9187=>"101101100",
  9188=>"110110010",
  9189=>"111110011",
  9190=>"100010000",
  9191=>"101000110",
  9192=>"000011111",
  9193=>"110000010",
  9194=>"111011100",
  9195=>"011011101",
  9196=>"010100101",
  9197=>"111111011",
  9198=>"000010111",
  9199=>"100101111",
  9200=>"010000111",
  9201=>"101000001",
  9202=>"101111100",
  9203=>"100111110",
  9204=>"001011110",
  9205=>"100000011",
  9206=>"101011100",
  9207=>"101010010",
  9208=>"000001111",
  9209=>"110011110",
  9210=>"101011100",
  9211=>"101100110",
  9212=>"001100001",
  9213=>"101101000",
  9214=>"111111111",
  9215=>"000110110",
  9216=>"111101010",
  9217=>"010100001",
  9218=>"010001111",
  9219=>"000110000",
  9220=>"011111101",
  9221=>"000011101",
  9222=>"001001111",
  9223=>"100011011",
  9224=>"111111111",
  9225=>"000011111",
  9226=>"101100110",
  9227=>"101010011",
  9228=>"110101110",
  9229=>"010101000",
  9230=>"111110001",
  9231=>"111001111",
  9232=>"001110101",
  9233=>"110100100",
  9234=>"100111110",
  9235=>"000001100",
  9236=>"111011111",
  9237=>"011000100",
  9238=>"001010111",
  9239=>"110100000",
  9240=>"101111110",
  9241=>"011000001",
  9242=>"110101111",
  9243=>"100110111",
  9244=>"011010000",
  9245=>"011100001",
  9246=>"111111100",
  9247=>"101000110",
  9248=>"011000000",
  9249=>"100001011",
  9250=>"100100111",
  9251=>"010110111",
  9252=>"001011000",
  9253=>"001110111",
  9254=>"010101000",
  9255=>"110010110",
  9256=>"100111100",
  9257=>"000110100",
  9258=>"111000100",
  9259=>"101010011",
  9260=>"110010101",
  9261=>"100011101",
  9262=>"111110110",
  9263=>"011110101",
  9264=>"000110101",
  9265=>"110011001",
  9266=>"000000000",
  9267=>"010011011",
  9268=>"011000110",
  9269=>"111111010",
  9270=>"100100010",
  9271=>"000100010",
  9272=>"001001100",
  9273=>"110000101",
  9274=>"111011010",
  9275=>"100100100",
  9276=>"001100001",
  9277=>"011011100",
  9278=>"110100100",
  9279=>"110001001",
  9280=>"100101111",
  9281=>"001100010",
  9282=>"101001101",
  9283=>"011000001",
  9284=>"010001011",
  9285=>"100001111",
  9286=>"000010000",
  9287=>"010101001",
  9288=>"000011100",
  9289=>"010001000",
  9290=>"101010010",
  9291=>"111001001",
  9292=>"011101101",
  9293=>"010111111",
  9294=>"100010000",
  9295=>"111011001",
  9296=>"011001001",
  9297=>"010000100",
  9298=>"010000011",
  9299=>"110011010",
  9300=>"100101110",
  9301=>"011011000",
  9302=>"001111011",
  9303=>"110011001",
  9304=>"000000011",
  9305=>"110110010",
  9306=>"011110110",
  9307=>"010000101",
  9308=>"110111101",
  9309=>"001010100",
  9310=>"101111011",
  9311=>"100011110",
  9312=>"100001101",
  9313=>"010111010",
  9314=>"110110000",
  9315=>"111100011",
  9316=>"000011001",
  9317=>"001000001",
  9318=>"001111110",
  9319=>"111000101",
  9320=>"110011110",
  9321=>"100110110",
  9322=>"101111000",
  9323=>"000011101",
  9324=>"010010110",
  9325=>"101100100",
  9326=>"111101010",
  9327=>"001000000",
  9328=>"110100100",
  9329=>"000000100",
  9330=>"011110010",
  9331=>"000000101",
  9332=>"001000100",
  9333=>"111001101",
  9334=>"010011101",
  9335=>"111101010",
  9336=>"001101001",
  9337=>"101000111",
  9338=>"101011111",
  9339=>"100011011",
  9340=>"000100111",
  9341=>"100100100",
  9342=>"101110111",
  9343=>"111110110",
  9344=>"000001101",
  9345=>"010100110",
  9346=>"010011101",
  9347=>"010000001",
  9348=>"111101100",
  9349=>"001001010",
  9350=>"010010111",
  9351=>"101101110",
  9352=>"010110011",
  9353=>"100001110",
  9354=>"100000001",
  9355=>"010001110",
  9356=>"110011101",
  9357=>"101100000",
  9358=>"111010011",
  9359=>"000101111",
  9360=>"011000001",
  9361=>"110101111",
  9362=>"011100110",
  9363=>"110100111",
  9364=>"100011010",
  9365=>"000000101",
  9366=>"110010000",
  9367=>"111011000",
  9368=>"000000101",
  9369=>"101011100",
  9370=>"111000110",
  9371=>"100001001",
  9372=>"010111000",
  9373=>"010010001",
  9374=>"100010010",
  9375=>"001111000",
  9376=>"010000101",
  9377=>"110110110",
  9378=>"000010011",
  9379=>"110101011",
  9380=>"101100111",
  9381=>"010011101",
  9382=>"101100101",
  9383=>"110100111",
  9384=>"011110100",
  9385=>"110001001",
  9386=>"010101111",
  9387=>"010010101",
  9388=>"001011100",
  9389=>"110010110",
  9390=>"001100010",
  9391=>"001001011",
  9392=>"100011001",
  9393=>"010111110",
  9394=>"011100011",
  9395=>"000001011",
  9396=>"110001101",
  9397=>"010100111",
  9398=>"010100001",
  9399=>"000000001",
  9400=>"011000101",
  9401=>"100100010",
  9402=>"000101001",
  9403=>"110010011",
  9404=>"101000000",
  9405=>"000000101",
  9406=>"010001001",
  9407=>"001100101",
  9408=>"111011100",
  9409=>"110100100",
  9410=>"111010101",
  9411=>"001101011",
  9412=>"001100111",
  9413=>"001010011",
  9414=>"110011110",
  9415=>"111010100",
  9416=>"001100111",
  9417=>"101011101",
  9418=>"001000010",
  9419=>"011011000",
  9420=>"011010011",
  9421=>"110011100",
  9422=>"111110000",
  9423=>"000011000",
  9424=>"001000000",
  9425=>"000011101",
  9426=>"011000101",
  9427=>"011010000",
  9428=>"000100010",
  9429=>"001111001",
  9430=>"110000010",
  9431=>"010101110",
  9432=>"100101110",
  9433=>"101110101",
  9434=>"000011000",
  9435=>"011010010",
  9436=>"010101001",
  9437=>"101100100",
  9438=>"000111101",
  9439=>"001111000",
  9440=>"100000000",
  9441=>"011100001",
  9442=>"011000100",
  9443=>"101100001",
  9444=>"000110011",
  9445=>"011010000",
  9446=>"101000000",
  9447=>"101110000",
  9448=>"010100000",
  9449=>"110010011",
  9450=>"000101000",
  9451=>"101101100",
  9452=>"110111010",
  9453=>"001000100",
  9454=>"011101110",
  9455=>"000100011",
  9456=>"001011010",
  9457=>"010001011",
  9458=>"001010110",
  9459=>"010110101",
  9460=>"111100000",
  9461=>"110101111",
  9462=>"101010000",
  9463=>"001111010",
  9464=>"111010110",
  9465=>"010011100",
  9466=>"011100110",
  9467=>"110100010",
  9468=>"111010000",
  9469=>"001000001",
  9470=>"110111110",
  9471=>"110100100",
  9472=>"011011000",
  9473=>"001111011",
  9474=>"110011010",
  9475=>"110010101",
  9476=>"001110010",
  9477=>"011101000",
  9478=>"110011110",
  9479=>"011001101",
  9480=>"000001000",
  9481=>"101011001",
  9482=>"110100000",
  9483=>"001101101",
  9484=>"101101001",
  9485=>"111010010",
  9486=>"001111000",
  9487=>"101110000",
  9488=>"011011011",
  9489=>"101000101",
  9490=>"101011111",
  9491=>"110000111",
  9492=>"111101011",
  9493=>"001001101",
  9494=>"010110111",
  9495=>"100110100",
  9496=>"110010101",
  9497=>"110100001",
  9498=>"110011110",
  9499=>"101000000",
  9500=>"101010111",
  9501=>"101111001",
  9502=>"101101000",
  9503=>"110000110",
  9504=>"101000111",
  9505=>"110011101",
  9506=>"111110111",
  9507=>"000011011",
  9508=>"011011110",
  9509=>"011100001",
  9510=>"100001010",
  9511=>"101110000",
  9512=>"111010100",
  9513=>"010100010",
  9514=>"111010100",
  9515=>"111100011",
  9516=>"100100011",
  9517=>"101110101",
  9518=>"000110101",
  9519=>"100000101",
  9520=>"010001110",
  9521=>"011110001",
  9522=>"111000100",
  9523=>"001100000",
  9524=>"100010001",
  9525=>"001101111",
  9526=>"101000010",
  9527=>"001111000",
  9528=>"100001100",
  9529=>"101000000",
  9530=>"110101111",
  9531=>"001110111",
  9532=>"000000011",
  9533=>"000101001",
  9534=>"111001000",
  9535=>"010001001",
  9536=>"000110111",
  9537=>"110010011",
  9538=>"010000000",
  9539=>"010111000",
  9540=>"000000011",
  9541=>"110011001",
  9542=>"011111010",
  9543=>"101110100",
  9544=>"101000100",
  9545=>"011010100",
  9546=>"011110100",
  9547=>"101110100",
  9548=>"001110011",
  9549=>"111000011",
  9550=>"100110111",
  9551=>"110110100",
  9552=>"101100010",
  9553=>"010000000",
  9554=>"110101100",
  9555=>"000010000",
  9556=>"010100100",
  9557=>"011111100",
  9558=>"001101011",
  9559=>"010101011",
  9560=>"010110111",
  9561=>"110100111",
  9562=>"001000001",
  9563=>"000110000",
  9564=>"111000000",
  9565=>"010000111",
  9566=>"011111010",
  9567=>"011011111",
  9568=>"010101110",
  9569=>"000000011",
  9570=>"111000101",
  9571=>"100101110",
  9572=>"011111000",
  9573=>"111101011",
  9574=>"000000111",
  9575=>"000100000",
  9576=>"010001010",
  9577=>"110111111",
  9578=>"101000111",
  9579=>"000011001",
  9580=>"011000000",
  9581=>"111011111",
  9582=>"000011010",
  9583=>"101100010",
  9584=>"111111110",
  9585=>"011110010",
  9586=>"101000111",
  9587=>"001100001",
  9588=>"001011000",
  9589=>"000100100",
  9590=>"100101011",
  9591=>"000000111",
  9592=>"010101101",
  9593=>"010010100",
  9594=>"100111111",
  9595=>"011000011",
  9596=>"010010001",
  9597=>"100010000",
  9598=>"001001101",
  9599=>"011010010",
  9600=>"000100000",
  9601=>"111111111",
  9602=>"101110010",
  9603=>"010110110",
  9604=>"001111010",
  9605=>"010101110",
  9606=>"010001011",
  9607=>"111001011",
  9608=>"100011001",
  9609=>"000100110",
  9610=>"100111000",
  9611=>"000110010",
  9612=>"100101011",
  9613=>"000101111",
  9614=>"101111101",
  9615=>"011111100",
  9616=>"010010111",
  9617=>"010111000",
  9618=>"111011100",
  9619=>"000110110",
  9620=>"011111010",
  9621=>"000001000",
  9622=>"101010111",
  9623=>"110111111",
  9624=>"111110111",
  9625=>"010100110",
  9626=>"110011110",
  9627=>"010000010",
  9628=>"011100101",
  9629=>"100011001",
  9630=>"011000000",
  9631=>"101101001",
  9632=>"100110001",
  9633=>"100100011",
  9634=>"001111010",
  9635=>"000010000",
  9636=>"110011100",
  9637=>"101110100",
  9638=>"011100111",
  9639=>"011000111",
  9640=>"000101101",
  9641=>"111111100",
  9642=>"101101000",
  9643=>"011100000",
  9644=>"010111111",
  9645=>"100100001",
  9646=>"000000010",
  9647=>"101101001",
  9648=>"010111000",
  9649=>"010010001",
  9650=>"000111000",
  9651=>"110010111",
  9652=>"001110110",
  9653=>"001101010",
  9654=>"001010100",
  9655=>"011001111",
  9656=>"111111101",
  9657=>"011010000",
  9658=>"010100000",
  9659=>"001110011",
  9660=>"101110100",
  9661=>"001010111",
  9662=>"100100100",
  9663=>"011110101",
  9664=>"001000111",
  9665=>"000111110",
  9666=>"011010010",
  9667=>"000001010",
  9668=>"011100001",
  9669=>"111100000",
  9670=>"111110000",
  9671=>"000000010",
  9672=>"110110010",
  9673=>"101100110",
  9674=>"100010011",
  9675=>"100110100",
  9676=>"011111011",
  9677=>"001100101",
  9678=>"000101010",
  9679=>"110100100",
  9680=>"000011101",
  9681=>"000001101",
  9682=>"101001001",
  9683=>"110000000",
  9684=>"111011011",
  9685=>"000001000",
  9686=>"100100001",
  9687=>"111000111",
  9688=>"001010110",
  9689=>"011001100",
  9690=>"010000001",
  9691=>"010001100",
  9692=>"011101010",
  9693=>"001011100",
  9694=>"011111011",
  9695=>"110011101",
  9696=>"110111101",
  9697=>"000001100",
  9698=>"010111111",
  9699=>"110010110",
  9700=>"100110101",
  9701=>"111110101",
  9702=>"100101001",
  9703=>"001010101",
  9704=>"101110010",
  9705=>"111011100",
  9706=>"111111000",
  9707=>"001100110",
  9708=>"011000000",
  9709=>"011110001",
  9710=>"110010011",
  9711=>"001011000",
  9712=>"011111111",
  9713=>"111100000",
  9714=>"110011001",
  9715=>"101000010",
  9716=>"111000100",
  9717=>"011111110",
  9718=>"010110101",
  9719=>"001110000",
  9720=>"011101110",
  9721=>"111001011",
  9722=>"111110101",
  9723=>"111011110",
  9724=>"110110110",
  9725=>"010011000",
  9726=>"011011011",
  9727=>"110000101",
  9728=>"000100101",
  9729=>"000100111",
  9730=>"001111110",
  9731=>"000001010",
  9732=>"111011110",
  9733=>"111110111",
  9734=>"001000110",
  9735=>"100111111",
  9736=>"111100101",
  9737=>"010011010",
  9738=>"011101010",
  9739=>"110111010",
  9740=>"010011010",
  9741=>"010000001",
  9742=>"000100000",
  9743=>"011000111",
  9744=>"111010101",
  9745=>"111001011",
  9746=>"000100111",
  9747=>"100111001",
  9748=>"110011001",
  9749=>"001001001",
  9750=>"110111111",
  9751=>"011101001",
  9752=>"110111101",
  9753=>"001010100",
  9754=>"000001000",
  9755=>"000101111",
  9756=>"001010001",
  9757=>"111100001",
  9758=>"010010001",
  9759=>"111010101",
  9760=>"101101101",
  9761=>"100001100",
  9762=>"000111010",
  9763=>"000000011",
  9764=>"111100110",
  9765=>"101101001",
  9766=>"000010011",
  9767=>"011111000",
  9768=>"001100100",
  9769=>"111011001",
  9770=>"110010100",
  9771=>"111100000",
  9772=>"110000000",
  9773=>"000101110",
  9774=>"001011010",
  9775=>"000110000",
  9776=>"100101001",
  9777=>"110001100",
  9778=>"101101001",
  9779=>"010111110",
  9780=>"110100100",
  9781=>"001000111",
  9782=>"110100111",
  9783=>"110101001",
  9784=>"000011011",
  9785=>"010010100",
  9786=>"100010111",
  9787=>"010010101",
  9788=>"011010101",
  9789=>"010100010",
  9790=>"100001011",
  9791=>"100111001",
  9792=>"010001110",
  9793=>"101010110",
  9794=>"101100110",
  9795=>"110100110",
  9796=>"100100110",
  9797=>"101111101",
  9798=>"001001111",
  9799=>"100011001",
  9800=>"010110000",
  9801=>"001001100",
  9802=>"011100001",
  9803=>"111101110",
  9804=>"000001001",
  9805=>"111010110",
  9806=>"101100111",
  9807=>"001010100",
  9808=>"001100000",
  9809=>"010010011",
  9810=>"000010101",
  9811=>"111011101",
  9812=>"000100011",
  9813=>"101100000",
  9814=>"100000000",
  9815=>"001011001",
  9816=>"011011001",
  9817=>"010010000",
  9818=>"111111111",
  9819=>"000001111",
  9820=>"011000000",
  9821=>"010110001",
  9822=>"011111110",
  9823=>"110011111",
  9824=>"110000111",
  9825=>"100001011",
  9826=>"011100100",
  9827=>"111111110",
  9828=>"011110010",
  9829=>"000111101",
  9830=>"100111111",
  9831=>"111110010",
  9832=>"110010010",
  9833=>"100100100",
  9834=>"111110000",
  9835=>"010100000",
  9836=>"111111001",
  9837=>"001111100",
  9838=>"000010110",
  9839=>"010001100",
  9840=>"101111110",
  9841=>"000001100",
  9842=>"100101100",
  9843=>"000000110",
  9844=>"011111110",
  9845=>"111011101",
  9846=>"110111101",
  9847=>"000001111",
  9848=>"111000111",
  9849=>"001010000",
  9850=>"101001101",
  9851=>"001010011",
  9852=>"010010100",
  9853=>"101001000",
  9854=>"000100010",
  9855=>"010101101",
  9856=>"010110110",
  9857=>"001000100",
  9858=>"111001011",
  9859=>"101001001",
  9860=>"011000001",
  9861=>"101101101",
  9862=>"000100111",
  9863=>"111010000",
  9864=>"011101101",
  9865=>"110000001",
  9866=>"100011011",
  9867=>"000111010",
  9868=>"011000001",
  9869=>"111011101",
  9870=>"000011011",
  9871=>"010111010",
  9872=>"000000011",
  9873=>"100110110",
  9874=>"100000010",
  9875=>"011010111",
  9876=>"111010100",
  9877=>"001001000",
  9878=>"101001000",
  9879=>"010101110",
  9880=>"100011111",
  9881=>"101101100",
  9882=>"000110100",
  9883=>"100011000",
  9884=>"101010000",
  9885=>"110101011",
  9886=>"011100101",
  9887=>"110100111",
  9888=>"110111010",
  9889=>"000111101",
  9890=>"000011110",
  9891=>"000001001",
  9892=>"000000011",
  9893=>"000101010",
  9894=>"101111001",
  9895=>"000011000",
  9896=>"110010111",
  9897=>"111000011",
  9898=>"100001111",
  9899=>"100001010",
  9900=>"111001001",
  9901=>"000000001",
  9902=>"001001011",
  9903=>"110001001",
  9904=>"100010101",
  9905=>"010110010",
  9906=>"001100101",
  9907=>"010001111",
  9908=>"000001000",
  9909=>"000101101",
  9910=>"000111100",
  9911=>"110110111",
  9912=>"010100001",
  9913=>"010110011",
  9914=>"110001001",
  9915=>"111011111",
  9916=>"010011010",
  9917=>"010011011",
  9918=>"010101010",
  9919=>"111101111",
  9920=>"110000011",
  9921=>"111110101",
  9922=>"110110111",
  9923=>"001101000",
  9924=>"101010110",
  9925=>"110010110",
  9926=>"001100100",
  9927=>"000110010",
  9928=>"101101010",
  9929=>"110000111",
  9930=>"100001110",
  9931=>"000011011",
  9932=>"101101001",
  9933=>"000001101",
  9934=>"011010100",
  9935=>"100101011",
  9936=>"100010101",
  9937=>"101001111",
  9938=>"001100110",
  9939=>"100110100",
  9940=>"010000011",
  9941=>"011111110",
  9942=>"110000110",
  9943=>"100100000",
  9944=>"110100000",
  9945=>"110011110",
  9946=>"101000101",
  9947=>"101000001",
  9948=>"101101110",
  9949=>"101100000",
  9950=>"100111000",
  9951=>"100000010",
  9952=>"000011011",
  9953=>"000010000",
  9954=>"010011000",
  9955=>"111110110",
  9956=>"011001001",
  9957=>"110010111",
  9958=>"001100100",
  9959=>"000011110",
  9960=>"100001001",
  9961=>"011111100",
  9962=>"011011101",
  9963=>"001110110",
  9964=>"101000101",
  9965=>"001001111",
  9966=>"101111101",
  9967=>"101111000",
  9968=>"111001001",
  9969=>"001101111",
  9970=>"101011011",
  9971=>"101110000",
  9972=>"111010000",
  9973=>"101010011",
  9974=>"101111001",
  9975=>"100001010",
  9976=>"011001011",
  9977=>"111111000",
  9978=>"010001110",
  9979=>"011101010",
  9980=>"000110010",
  9981=>"110101110",
  9982=>"011000010",
  9983=>"100100010",
  9984=>"101111011",
  9985=>"000010001",
  9986=>"110000011",
  9987=>"000110000",
  9988=>"000010101",
  9989=>"001100000",
  9990=>"110100001",
  9991=>"010111101",
  9992=>"111001001",
  9993=>"110111000",
  9994=>"001010110",
  9995=>"100000111",
  9996=>"001000011",
  9997=>"010010100",
  9998=>"010001101",
  9999=>"001011010",
  10000=>"011000000",
  10001=>"100100000",
  10002=>"011010100",
  10003=>"100110100",
  10004=>"011010111",
  10005=>"111001100",
  10006=>"001110111",
  10007=>"100000111",
  10008=>"111100111",
  10009=>"100010101",
  10010=>"101111010",
  10011=>"010001100",
  10012=>"111001010",
  10013=>"001001111",
  10014=>"110000101",
  10015=>"101111011",
  10016=>"010001101",
  10017=>"110000110",
  10018=>"100110101",
  10019=>"010110000",
  10020=>"111000110",
  10021=>"100001000",
  10022=>"110101100",
  10023=>"000000011",
  10024=>"000110010",
  10025=>"111011001",
  10026=>"001111110",
  10027=>"011001100",
  10028=>"101001110",
  10029=>"000001101",
  10030=>"111101110",
  10031=>"110101110",
  10032=>"011110111",
  10033=>"010000001",
  10034=>"100101010",
  10035=>"101100101",
  10036=>"101010100",
  10037=>"000001001",
  10038=>"011000111",
  10039=>"101100100",
  10040=>"001010100",
  10041=>"001100011",
  10042=>"000101001",
  10043=>"110010110",
  10044=>"101001110",
  10045=>"010101010",
  10046=>"100001100",
  10047=>"001000111",
  10048=>"000010010",
  10049=>"011010000",
  10050=>"011111110",
  10051=>"111001111",
  10052=>"111111110",
  10053=>"100010101",
  10054=>"111100010",
  10055=>"001111000",
  10056=>"000101000",
  10057=>"011101000",
  10058=>"110010000",
  10059=>"111011000",
  10060=>"010110000",
  10061=>"101010011",
  10062=>"111111011",
  10063=>"011010110",
  10064=>"111011101",
  10065=>"011011010",
  10066=>"010101000",
  10067=>"001011111",
  10068=>"011000101",
  10069=>"001010011",
  10070=>"100010110",
  10071=>"011001101",
  10072=>"000000010",
  10073=>"101010000",
  10074=>"111111110",
  10075=>"111111110",
  10076=>"001000010",
  10077=>"000010011",
  10078=>"001001010",
  10079=>"110011001",
  10080=>"000011101",
  10081=>"110110100",
  10082=>"100101001",
  10083=>"111110101",
  10084=>"110111001",
  10085=>"001001001",
  10086=>"100000110",
  10087=>"110110111",
  10088=>"010010000",
  10089=>"011001001",
  10090=>"111001110",
  10091=>"100001101",
  10092=>"011101011",
  10093=>"010111000",
  10094=>"111001010",
  10095=>"000110110",
  10096=>"011101000",
  10097=>"010001010",
  10098=>"010100011",
  10099=>"000110000",
  10100=>"111011110",
  10101=>"000101101",
  10102=>"001111000",
  10103=>"111010011",
  10104=>"000100010",
  10105=>"010111110",
  10106=>"001100101",
  10107=>"111111101",
  10108=>"000010110",
  10109=>"000100000",
  10110=>"110100101",
  10111=>"111010100",
  10112=>"101011000",
  10113=>"000100011",
  10114=>"101101111",
  10115=>"010010111",
  10116=>"011100110",
  10117=>"100100011",
  10118=>"000110101",
  10119=>"000110001",
  10120=>"000100111",
  10121=>"001100000",
  10122=>"000100110",
  10123=>"000011101",
  10124=>"010010001",
  10125=>"011101111",
  10126=>"111101100",
  10127=>"011110011",
  10128=>"110001101",
  10129=>"111100010",
  10130=>"000110000",
  10131=>"011101111",
  10132=>"110001011",
  10133=>"001110100",
  10134=>"101000101",
  10135=>"001110000",
  10136=>"110100111",
  10137=>"000000111",
  10138=>"001001101",
  10139=>"100101001",
  10140=>"011010010",
  10141=>"010010101",
  10142=>"111101100",
  10143=>"100110111",
  10144=>"101001111",
  10145=>"000000001",
  10146=>"101010011",
  10147=>"101111100",
  10148=>"001000000",
  10149=>"111001011",
  10150=>"000011101",
  10151=>"011110000",
  10152=>"111001110",
  10153=>"100000101",
  10154=>"000111100",
  10155=>"001110111",
  10156=>"011100110",
  10157=>"111100101",
  10158=>"111000000",
  10159=>"010100101",
  10160=>"110011011",
  10161=>"011000011",
  10162=>"011101101",
  10163=>"111001010",
  10164=>"110011110",
  10165=>"011111111",
  10166=>"101100011",
  10167=>"000110110",
  10168=>"111100100",
  10169=>"111010101",
  10170=>"010010111",
  10171=>"101010010",
  10172=>"100001110",
  10173=>"001110110",
  10174=>"001000111",
  10175=>"011011110",
  10176=>"111001110",
  10177=>"010000100",
  10178=>"000100111",
  10179=>"011001001",
  10180=>"111111101",
  10181=>"000101001",
  10182=>"011000110",
  10183=>"100110110",
  10184=>"000010111",
  10185=>"011000101",
  10186=>"000011110",
  10187=>"001111110",
  10188=>"000101010",
  10189=>"110000110",
  10190=>"001110101",
  10191=>"100000011",
  10192=>"000001000",
  10193=>"111011000",
  10194=>"011111111",
  10195=>"011110000",
  10196=>"111111111",
  10197=>"000101100",
  10198=>"000000000",
  10199=>"000011011",
  10200=>"001111110",
  10201=>"100000011",
  10202=>"001010101",
  10203=>"001000101",
  10204=>"100010011",
  10205=>"010100110",
  10206=>"100111000",
  10207=>"000000100",
  10208=>"011101000",
  10209=>"101110010",
  10210=>"110001111",
  10211=>"001000000",
  10212=>"010001011",
  10213=>"000010101",
  10214=>"110010000",
  10215=>"111110011",
  10216=>"011111001",
  10217=>"000010000",
  10218=>"000100010",
  10219=>"101000101",
  10220=>"000110010",
  10221=>"001010110",
  10222=>"001011110",
  10223=>"010010000",
  10224=>"111010101",
  10225=>"010110100",
  10226=>"101101110",
  10227=>"011010011",
  10228=>"010001101",
  10229=>"110010011",
  10230=>"000110001",
  10231=>"001010001",
  10232=>"011111110",
  10233=>"011000110",
  10234=>"000001011",
  10235=>"001101110",
  10236=>"010001000",
  10237=>"001010101",
  10238=>"001011101",
  10239=>"010110101",
  10240=>"101010100",
  10241=>"100001110",
  10242=>"000110010",
  10243=>"100011101",
  10244=>"010001110",
  10245=>"101110010",
  10246=>"011110010",
  10247=>"000110001",
  10248=>"100011100",
  10249=>"001011010",
  10250=>"001000100",
  10251=>"001101101",
  10252=>"101000000",
  10253=>"111001110",
  10254=>"111111001",
  10255=>"010100000",
  10256=>"111101101",
  10257=>"011011110",
  10258=>"100110111",
  10259=>"101000011",
  10260=>"000101011",
  10261=>"000000111",
  10262=>"011011111",
  10263=>"101101000",
  10264=>"011010100",
  10265=>"101110011",
  10266=>"101001000",
  10267=>"111110110",
  10268=>"010001001",
  10269=>"010101000",
  10270=>"010101001",
  10271=>"101100011",
  10272=>"110011111",
  10273=>"100110111",
  10274=>"110010000",
  10275=>"000001011",
  10276=>"011101010",
  10277=>"110010101",
  10278=>"101000001",
  10279=>"010010110",
  10280=>"100011011",
  10281=>"101101101",
  10282=>"011110010",
  10283=>"011101001",
  10284=>"001110110",
  10285=>"000111100",
  10286=>"000000010",
  10287=>"001100101",
  10288=>"111110101",
  10289=>"110101110",
  10290=>"011111010",
  10291=>"000010101",
  10292=>"101101101",
  10293=>"010011001",
  10294=>"100010111",
  10295=>"110010001",
  10296=>"001100000",
  10297=>"101000010",
  10298=>"000001010",
  10299=>"010000110",
  10300=>"111110111",
  10301=>"001011011",
  10302=>"100100011",
  10303=>"111101100",
  10304=>"011100000",
  10305=>"001001100",
  10306=>"001100001",
  10307=>"101101101",
  10308=>"111010110",
  10309=>"010010011",
  10310=>"010000011",
  10311=>"000101101",
  10312=>"001111110",
  10313=>"100011001",
  10314=>"100111011",
  10315=>"101101110",
  10316=>"110000000",
  10317=>"101000011",
  10318=>"010010001",
  10319=>"101100000",
  10320=>"110001101",
  10321=>"011101101",
  10322=>"011000110",
  10323=>"011111110",
  10324=>"111111011",
  10325=>"111000000",
  10326=>"100000111",
  10327=>"001101001",
  10328=>"111010100",
  10329=>"001101100",
  10330=>"011000110",
  10331=>"001000111",
  10332=>"011100010",
  10333=>"101001010",
  10334=>"010100011",
  10335=>"111010000",
  10336=>"000011001",
  10337=>"101100001",
  10338=>"000100000",
  10339=>"110001010",
  10340=>"011001001",
  10341=>"101100000",
  10342=>"111111010",
  10343=>"100011010",
  10344=>"011110101",
  10345=>"110010011",
  10346=>"111010011",
  10347=>"111000010",
  10348=>"001001100",
  10349=>"111010110",
  10350=>"010010100",
  10351=>"100110001",
  10352=>"110100000",
  10353=>"001111011",
  10354=>"001010110",
  10355=>"010111000",
  10356=>"011110000",
  10357=>"001110100",
  10358=>"111011000",
  10359=>"111111011",
  10360=>"000100100",
  10361=>"110011011",
  10362=>"011010111",
  10363=>"110001011",
  10364=>"111101010",
  10365=>"110001001",
  10366=>"000000110",
  10367=>"010011010",
  10368=>"111001011",
  10369=>"010101101",
  10370=>"100010010",
  10371=>"101000110",
  10372=>"101101000",
  10373=>"101111100",
  10374=>"001000100",
  10375=>"001010010",
  10376=>"001001111",
  10377=>"001001001",
  10378=>"001001001",
  10379=>"111000100",
  10380=>"001010111",
  10381=>"110100110",
  10382=>"001011011",
  10383=>"011000100",
  10384=>"100010101",
  10385=>"011100001",
  10386=>"101001001",
  10387=>"101000010",
  10388=>"100110000",
  10389=>"000000011",
  10390=>"001001001",
  10391=>"000011111",
  10392=>"101011111",
  10393=>"101111110",
  10394=>"011100010",
  10395=>"010100101",
  10396=>"011001100",
  10397=>"000000101",
  10398=>"100001000",
  10399=>"110000001",
  10400=>"110101001",
  10401=>"000100000",
  10402=>"010010100",
  10403=>"111101101",
  10404=>"001101100",
  10405=>"010111111",
  10406=>"010101110",
  10407=>"000111100",
  10408=>"100000010",
  10409=>"011001010",
  10410=>"001010111",
  10411=>"000000001",
  10412=>"111100000",
  10413=>"010011110",
  10414=>"111111100",
  10415=>"001010111",
  10416=>"011010110",
  10417=>"011011101",
  10418=>"100101000",
  10419=>"100000001",
  10420=>"111111000",
  10421=>"000010001",
  10422=>"011101010",
  10423=>"010000100",
  10424=>"010010100",
  10425=>"001000100",
  10426=>"001100001",
  10427=>"001010110",
  10428=>"001010011",
  10429=>"110101010",
  10430=>"001100110",
  10431=>"001100011",
  10432=>"101111011",
  10433=>"101101100",
  10434=>"111100111",
  10435=>"110100110",
  10436=>"001010111",
  10437=>"001101001",
  10438=>"111000000",
  10439=>"100011011",
  10440=>"000110110",
  10441=>"000010011",
  10442=>"100000000",
  10443=>"101000000",
  10444=>"111001010",
  10445=>"100111110",
  10446=>"001001010",
  10447=>"010111001",
  10448=>"001011001",
  10449=>"000111000",
  10450=>"001111100",
  10451=>"111001011",
  10452=>"110011110",
  10453=>"100101011",
  10454=>"111101100",
  10455=>"111011000",
  10456=>"010000100",
  10457=>"100001000",
  10458=>"111010111",
  10459=>"101001010",
  10460=>"010101000",
  10461=>"000000001",
  10462=>"111000001",
  10463=>"100010011",
  10464=>"010011100",
  10465=>"001010011",
  10466=>"011110011",
  10467=>"010000110",
  10468=>"110101010",
  10469=>"011001100",
  10470=>"111101011",
  10471=>"001110001",
  10472=>"010000010",
  10473=>"100000110",
  10474=>"010000100",
  10475=>"001011110",
  10476=>"101001001",
  10477=>"110100101",
  10478=>"001100101",
  10479=>"001000100",
  10480=>"111101101",
  10481=>"111000000",
  10482=>"101100110",
  10483=>"110111110",
  10484=>"110010010",
  10485=>"001100011",
  10486=>"111101100",
  10487=>"011110111",
  10488=>"111010010",
  10489=>"110101110",
  10490=>"000010111",
  10491=>"001000110",
  10492=>"011001101",
  10493=>"010001100",
  10494=>"000111111",
  10495=>"111001111",
  10496=>"000100010",
  10497=>"110000011",
  10498=>"110111010",
  10499=>"101111111",
  10500=>"110000010",
  10501=>"110011111",
  10502=>"010011100",
  10503=>"100000101",
  10504=>"111101010",
  10505=>"101000000",
  10506=>"100111001",
  10507=>"101100000",
  10508=>"000100011",
  10509=>"000010010",
  10510=>"100101000",
  10511=>"000011111",
  10512=>"111010000",
  10513=>"100110010",
  10514=>"010011101",
  10515=>"011010101",
  10516=>"010000000",
  10517=>"011111000",
  10518=>"010000110",
  10519=>"000001010",
  10520=>"101100001",
  10521=>"001111011",
  10522=>"110111101",
  10523=>"101011110",
  10524=>"101100101",
  10525=>"100010000",
  10526=>"110100110",
  10527=>"000101010",
  10528=>"000001101",
  10529=>"100001000",
  10530=>"101010110",
  10531=>"010001101",
  10532=>"000101001",
  10533=>"000011010",
  10534=>"001001000",
  10535=>"101000100",
  10536=>"000010011",
  10537=>"110001011",
  10538=>"000111111",
  10539=>"110110010",
  10540=>"000110100",
  10541=>"101001000",
  10542=>"100001001",
  10543=>"011101111",
  10544=>"010100000",
  10545=>"010110001",
  10546=>"011101111",
  10547=>"011111111",
  10548=>"110010011",
  10549=>"001100101",
  10550=>"100010100",
  10551=>"000110000",
  10552=>"001000110",
  10553=>"011101001",
  10554=>"011001000",
  10555=>"011001000",
  10556=>"010111111",
  10557=>"011001010",
  10558=>"010101110",
  10559=>"010100101",
  10560=>"111011001",
  10561=>"011011100",
  10562=>"011001110",
  10563=>"010001011",
  10564=>"110101111",
  10565=>"100100000",
  10566=>"110000010",
  10567=>"010110000",
  10568=>"101011100",
  10569=>"101000001",
  10570=>"010100000",
  10571=>"000000000",
  10572=>"011000101",
  10573=>"010000000",
  10574=>"000011101",
  10575=>"010011111",
  10576=>"010111000",
  10577=>"100111110",
  10578=>"000101000",
  10579=>"100000101",
  10580=>"000110110",
  10581=>"000111111",
  10582=>"110011100",
  10583=>"111110000",
  10584=>"110101010",
  10585=>"001011110",
  10586=>"001101001",
  10587=>"101101011",
  10588=>"100100001",
  10589=>"111010110",
  10590=>"001011011",
  10591=>"101111000",
  10592=>"010000010",
  10593=>"001011111",
  10594=>"011011110",
  10595=>"001110000",
  10596=>"001000111",
  10597=>"101111110",
  10598=>"111011011",
  10599=>"111100100",
  10600=>"000001100",
  10601=>"111110100",
  10602=>"001000101",
  10603=>"011111000",
  10604=>"110000101",
  10605=>"111100100",
  10606=>"001110000",
  10607=>"000000000",
  10608=>"101101001",
  10609=>"110111100",
  10610=>"011110001",
  10611=>"110000101",
  10612=>"111100100",
  10613=>"010111010",
  10614=>"111001110",
  10615=>"001110100",
  10616=>"100101001",
  10617=>"100001100",
  10618=>"101101101",
  10619=>"000000000",
  10620=>"101000010",
  10621=>"001011101",
  10622=>"100100111",
  10623=>"100001010",
  10624=>"001000111",
  10625=>"010010101",
  10626=>"000010001",
  10627=>"000111100",
  10628=>"111110101",
  10629=>"110000000",
  10630=>"011000101",
  10631=>"011001001",
  10632=>"001011110",
  10633=>"111101111",
  10634=>"100111000",
  10635=>"001100111",
  10636=>"000010110",
  10637=>"001000010",
  10638=>"101001000",
  10639=>"010110000",
  10640=>"000101101",
  10641=>"000001110",
  10642=>"010011111",
  10643=>"010100101",
  10644=>"110011011",
  10645=>"011001000",
  10646=>"000010010",
  10647=>"110000000",
  10648=>"111111111",
  10649=>"100000101",
  10650=>"110000010",
  10651=>"010111110",
  10652=>"010110101",
  10653=>"010110010",
  10654=>"000011101",
  10655=>"111000001",
  10656=>"100011000",
  10657=>"100100111",
  10658=>"110010000",
  10659=>"001110101",
  10660=>"100000011",
  10661=>"010000111",
  10662=>"100000000",
  10663=>"111010100",
  10664=>"001001000",
  10665=>"100100100",
  10666=>"011001010",
  10667=>"000011011",
  10668=>"101011011",
  10669=>"000111000",
  10670=>"101010111",
  10671=>"011011011",
  10672=>"000001000",
  10673=>"010000011",
  10674=>"000000101",
  10675=>"011011011",
  10676=>"100011101",
  10677=>"000010011",
  10678=>"001011000",
  10679=>"100101110",
  10680=>"100000000",
  10681=>"111000010",
  10682=>"010000000",
  10683=>"011001100",
  10684=>"010000011",
  10685=>"001100001",
  10686=>"110101111",
  10687=>"000111010",
  10688=>"010001110",
  10689=>"000000010",
  10690=>"011000011",
  10691=>"010000110",
  10692=>"000010100",
  10693=>"100101101",
  10694=>"100100011",
  10695=>"011011001",
  10696=>"111000011",
  10697=>"001011111",
  10698=>"011110010",
  10699=>"111111011",
  10700=>"000101111",
  10701=>"000101111",
  10702=>"010010011",
  10703=>"001011100",
  10704=>"011001000",
  10705=>"011101011",
  10706=>"010000111",
  10707=>"100000110",
  10708=>"100100100",
  10709=>"000000110",
  10710=>"111110111",
  10711=>"010000001",
  10712=>"101010001",
  10713=>"010011000",
  10714=>"111111010",
  10715=>"001101101",
  10716=>"111110101",
  10717=>"100011110",
  10718=>"000101001",
  10719=>"100000110",
  10720=>"110111101",
  10721=>"101111010",
  10722=>"110100111",
  10723=>"011000111",
  10724=>"010011101",
  10725=>"000001010",
  10726=>"110110001",
  10727=>"011001100",
  10728=>"001111100",
  10729=>"101010000",
  10730=>"100110001",
  10731=>"011011100",
  10732=>"100100110",
  10733=>"110001011",
  10734=>"101000010",
  10735=>"010101100",
  10736=>"001001101",
  10737=>"111010001",
  10738=>"111011000",
  10739=>"111101111",
  10740=>"010001010",
  10741=>"000010011",
  10742=>"011011001",
  10743=>"000011010",
  10744=>"111101001",
  10745=>"110010101",
  10746=>"010010111",
  10747=>"000110100",
  10748=>"001010111",
  10749=>"111010111",
  10750=>"100111001",
  10751=>"001010111",
  10752=>"101100100",
  10753=>"111110111",
  10754=>"111000011",
  10755=>"001000000",
  10756=>"001101011",
  10757=>"010101010",
  10758=>"101000010",
  10759=>"100100011",
  10760=>"000001100",
  10761=>"010000010",
  10762=>"100110101",
  10763=>"010110101",
  10764=>"011101001",
  10765=>"111111100",
  10766=>"100000100",
  10767=>"010010010",
  10768=>"111101011",
  10769=>"100000100",
  10770=>"111100000",
  10771=>"011101101",
  10772=>"101001000",
  10773=>"100010111",
  10774=>"000011100",
  10775=>"000011000",
  10776=>"101001001",
  10777=>"001111100",
  10778=>"001111001",
  10779=>"011000011",
  10780=>"111100101",
  10781=>"010111011",
  10782=>"111110111",
  10783=>"100001000",
  10784=>"110010011",
  10785=>"010010000",
  10786=>"011111110",
  10787=>"101110000",
  10788=>"000110000",
  10789=>"000000101",
  10790=>"101100001",
  10791=>"000001000",
  10792=>"111111100",
  10793=>"000111111",
  10794=>"111001100",
  10795=>"001111001",
  10796=>"110010011",
  10797=>"100101011",
  10798=>"011010111",
  10799=>"111011111",
  10800=>"100101010",
  10801=>"110111110",
  10802=>"100001001",
  10803=>"101111011",
  10804=>"111000010",
  10805=>"110001011",
  10806=>"010111110",
  10807=>"001000110",
  10808=>"010100111",
  10809=>"111100000",
  10810=>"111001001",
  10811=>"100110100",
  10812=>"001011101",
  10813=>"111000000",
  10814=>"101110001",
  10815=>"101101001",
  10816=>"001101011",
  10817=>"111000011",
  10818=>"001111110",
  10819=>"111001010",
  10820=>"100000011",
  10821=>"000100000",
  10822=>"001010000",
  10823=>"000010101",
  10824=>"000000101",
  10825=>"010010100",
  10826=>"010110000",
  10827=>"010101010",
  10828=>"010110000",
  10829=>"111000100",
  10830=>"010010110",
  10831=>"101101000",
  10832=>"000000111",
  10833=>"011010000",
  10834=>"100110101",
  10835=>"000111000",
  10836=>"101001111",
  10837=>"010011010",
  10838=>"101111101",
  10839=>"111101100",
  10840=>"001101000",
  10841=>"001001000",
  10842=>"001110110",
  10843=>"100111101",
  10844=>"001110011",
  10845=>"001110011",
  10846=>"101100011",
  10847=>"110011000",
  10848=>"011001011",
  10849=>"110101011",
  10850=>"001010000",
  10851=>"100010001",
  10852=>"011101011",
  10853=>"001001101",
  10854=>"010010100",
  10855=>"001101000",
  10856=>"010010110",
  10857=>"111101111",
  10858=>"000001011",
  10859=>"101000000",
  10860=>"010111101",
  10861=>"110110000",
  10862=>"000101100",
  10863=>"001010101",
  10864=>"001001001",
  10865=>"000100001",
  10866=>"100000110",
  10867=>"001101111",
  10868=>"011001001",
  10869=>"100100100",
  10870=>"000101001",
  10871=>"010100010",
  10872=>"011111100",
  10873=>"001101011",
  10874=>"101001100",
  10875=>"001111010",
  10876=>"001011100",
  10877=>"111010001",
  10878=>"101100111",
  10879=>"010001011",
  10880=>"100100100",
  10881=>"111011011",
  10882=>"001001011",
  10883=>"010011011",
  10884=>"110110010",
  10885=>"100100000",
  10886=>"010100100",
  10887=>"111101000",
  10888=>"000100000",
  10889=>"011111101",
  10890=>"011000011",
  10891=>"111000010",
  10892=>"010001010",
  10893=>"111100000",
  10894=>"010010010",
  10895=>"001001001",
  10896=>"011110101",
  10897=>"100011011",
  10898=>"111111111",
  10899=>"000010001",
  10900=>"100000011",
  10901=>"001010101",
  10902=>"011000101",
  10903=>"011001010",
  10904=>"101110011",
  10905=>"110100011",
  10906=>"011000100",
  10907=>"101100111",
  10908=>"101101011",
  10909=>"011101100",
  10910=>"000011011",
  10911=>"011011100",
  10912=>"100011001",
  10913=>"000010011",
  10914=>"010101000",
  10915=>"101110101",
  10916=>"000010111",
  10917=>"101101001",
  10918=>"100100110",
  10919=>"000011100",
  10920=>"100010110",
  10921=>"100011011",
  10922=>"101000011",
  10923=>"000000101",
  10924=>"100010000",
  10925=>"000000100",
  10926=>"100101001",
  10927=>"011110110",
  10928=>"100101100",
  10929=>"001101110",
  10930=>"001100100",
  10931=>"000010000",
  10932=>"101011101",
  10933=>"011111010",
  10934=>"111011010",
  10935=>"001101100",
  10936=>"111100001",
  10937=>"010100101",
  10938=>"011101011",
  10939=>"100100000",
  10940=>"111100101",
  10941=>"000011011",
  10942=>"101101000",
  10943=>"001101000",
  10944=>"000011000",
  10945=>"100100001",
  10946=>"000101111",
  10947=>"101110110",
  10948=>"010100101",
  10949=>"001001111",
  10950=>"111101000",
  10951=>"110101110",
  10952=>"001111101",
  10953=>"011000110",
  10954=>"000001011",
  10955=>"111101001",
  10956=>"001010111",
  10957=>"111110110",
  10958=>"010000110",
  10959=>"001101000",
  10960=>"100110101",
  10961=>"111100010",
  10962=>"000010111",
  10963=>"101011011",
  10964=>"100010010",
  10965=>"010100100",
  10966=>"000110100",
  10967=>"111000110",
  10968=>"001001001",
  10969=>"110100010",
  10970=>"000000111",
  10971=>"111101111",
  10972=>"101101101",
  10973=>"100001000",
  10974=>"111000100",
  10975=>"010001011",
  10976=>"010000001",
  10977=>"011000000",
  10978=>"101100111",
  10979=>"000001110",
  10980=>"101110000",
  10981=>"101000100",
  10982=>"010100001",
  10983=>"001011110",
  10984=>"111010111",
  10985=>"011100000",
  10986=>"111011111",
  10987=>"110000101",
  10988=>"001010101",
  10989=>"101111100",
  10990=>"100111000",
  10991=>"010000101",
  10992=>"111000001",
  10993=>"100011011",
  10994=>"011010101",
  10995=>"011000110",
  10996=>"001001011",
  10997=>"000100010",
  10998=>"100011110",
  10999=>"110011011",
  11000=>"111100001",
  11001=>"001000101",
  11002=>"011011001",
  11003=>"001000111",
  11004=>"001101111",
  11005=>"101111110",
  11006=>"001101110",
  11007=>"100100001",
  11008=>"010000110",
  11009=>"111001110",
  11010=>"101111010",
  11011=>"000111110",
  11012=>"001001000",
  11013=>"110000101",
  11014=>"101111010",
  11015=>"000111101",
  11016=>"100000001",
  11017=>"000001101",
  11018=>"100011100",
  11019=>"011001111",
  11020=>"110101110",
  11021=>"000101000",
  11022=>"100110001",
  11023=>"011011101",
  11024=>"010001100",
  11025=>"101111110",
  11026=>"101100001",
  11027=>"111001101",
  11028=>"100100100",
  11029=>"011110000",
  11030=>"001010100",
  11031=>"111110111",
  11032=>"101011110",
  11033=>"011001100",
  11034=>"000110100",
  11035=>"111101101",
  11036=>"010011110",
  11037=>"011101011",
  11038=>"101100001",
  11039=>"110011000",
  11040=>"000111111",
  11041=>"101000011",
  11042=>"111110110",
  11043=>"101001001",
  11044=>"111000010",
  11045=>"000110101",
  11046=>"111001101",
  11047=>"000001111",
  11048=>"010001000",
  11049=>"101010111",
  11050=>"011110011",
  11051=>"110010100",
  11052=>"000101110",
  11053=>"100010000",
  11054=>"000001101",
  11055=>"100011010",
  11056=>"100100110",
  11057=>"011100110",
  11058=>"010011111",
  11059=>"100110111",
  11060=>"011010000",
  11061=>"100011000",
  11062=>"100111000",
  11063=>"011001010",
  11064=>"111111111",
  11065=>"001100001",
  11066=>"101001000",
  11067=>"111101111",
  11068=>"110100100",
  11069=>"000100101",
  11070=>"000101000",
  11071=>"011101001",
  11072=>"001001110",
  11073=>"111000010",
  11074=>"101110011",
  11075=>"111010100",
  11076=>"100101010",
  11077=>"110101111",
  11078=>"000101111",
  11079=>"110011010",
  11080=>"010111111",
  11081=>"001100100",
  11082=>"010010011",
  11083=>"110000011",
  11084=>"100110001",
  11085=>"011000001",
  11086=>"101100001",
  11087=>"000001100",
  11088=>"111000100",
  11089=>"001000111",
  11090=>"011110101",
  11091=>"101000110",
  11092=>"000101001",
  11093=>"010010011",
  11094=>"001101100",
  11095=>"101001010",
  11096=>"000100011",
  11097=>"011100111",
  11098=>"001100000",
  11099=>"000000100",
  11100=>"010100000",
  11101=>"011100111",
  11102=>"101011010",
  11103=>"001000001",
  11104=>"011000000",
  11105=>"110010001",
  11106=>"111101100",
  11107=>"000010000",
  11108=>"111101111",
  11109=>"001110000",
  11110=>"101101111",
  11111=>"101000101",
  11112=>"000001001",
  11113=>"110000111",
  11114=>"101001000",
  11115=>"100011111",
  11116=>"101001111",
  11117=>"111101001",
  11118=>"000100011",
  11119=>"101001001",
  11120=>"010111001",
  11121=>"110101110",
  11122=>"011100110",
  11123=>"101001000",
  11124=>"101101010",
  11125=>"000011000",
  11126=>"100011110",
  11127=>"100101001",
  11128=>"100001010",
  11129=>"001100101",
  11130=>"011000100",
  11131=>"000101010",
  11132=>"000011001",
  11133=>"011001000",
  11134=>"000001100",
  11135=>"110110001",
  11136=>"111011011",
  11137=>"000001010",
  11138=>"011111110",
  11139=>"000010101",
  11140=>"011111010",
  11141=>"101011111",
  11142=>"000000100",
  11143=>"110111110",
  11144=>"100010000",
  11145=>"110010001",
  11146=>"100101111",
  11147=>"000101011",
  11148=>"101011110",
  11149=>"001001011",
  11150=>"011111001",
  11151=>"111111011",
  11152=>"001101101",
  11153=>"011010000",
  11154=>"001101001",
  11155=>"000110111",
  11156=>"001010011",
  11157=>"100101010",
  11158=>"000000100",
  11159=>"010000100",
  11160=>"000110100",
  11161=>"100100001",
  11162=>"111101011",
  11163=>"010110110",
  11164=>"111111100",
  11165=>"111100001",
  11166=>"101011100",
  11167=>"011010000",
  11168=>"011011001",
  11169=>"010001010",
  11170=>"111011100",
  11171=>"101000000",
  11172=>"101110110",
  11173=>"010111111",
  11174=>"000111000",
  11175=>"101010111",
  11176=>"111001010",
  11177=>"000000011",
  11178=>"111111011",
  11179=>"100001001",
  11180=>"111000001",
  11181=>"110111110",
  11182=>"011111111",
  11183=>"110110111",
  11184=>"011100010",
  11185=>"111110111",
  11186=>"001001100",
  11187=>"001100011",
  11188=>"100011111",
  11189=>"000000101",
  11190=>"111010110",
  11191=>"110100100",
  11192=>"111100001",
  11193=>"001110100",
  11194=>"110011010",
  11195=>"101110001",
  11196=>"111010011",
  11197=>"110000010",
  11198=>"111101001",
  11199=>"100001011",
  11200=>"010001100",
  11201=>"111101000",
  11202=>"000100011",
  11203=>"100111110",
  11204=>"110100101",
  11205=>"101110011",
  11206=>"010111100",
  11207=>"100111010",
  11208=>"100000010",
  11209=>"110001111",
  11210=>"000110110",
  11211=>"001010100",
  11212=>"010110111",
  11213=>"101100100",
  11214=>"010000111",
  11215=>"000101000",
  11216=>"011101101",
  11217=>"000110111",
  11218=>"010000011",
  11219=>"011001110",
  11220=>"100011101",
  11221=>"011110110",
  11222=>"010010000",
  11223=>"100110101",
  11224=>"100001110",
  11225=>"111011111",
  11226=>"100001000",
  11227=>"111101011",
  11228=>"101000001",
  11229=>"011011101",
  11230=>"010100000",
  11231=>"101010000",
  11232=>"101111000",
  11233=>"010010000",
  11234=>"011111111",
  11235=>"111100101",
  11236=>"001001111",
  11237=>"010100010",
  11238=>"100000101",
  11239=>"111110100",
  11240=>"001001011",
  11241=>"010110011",
  11242=>"101001101",
  11243=>"010011010",
  11244=>"101111000",
  11245=>"011101000",
  11246=>"000000011",
  11247=>"000011000",
  11248=>"001010100",
  11249=>"010111100",
  11250=>"000110001",
  11251=>"100000101",
  11252=>"000110101",
  11253=>"010010010",
  11254=>"110111101",
  11255=>"100100101",
  11256=>"100111101",
  11257=>"011111111",
  11258=>"000010001",
  11259=>"110101110",
  11260=>"011011000",
  11261=>"100000100",
  11262=>"011000001",
  11263=>"000110100",
  11264=>"000000000",
  11265=>"100011111",
  11266=>"011111011",
  11267=>"001110011",
  11268=>"101100100",
  11269=>"110010001",
  11270=>"001111100",
  11271=>"110011010",
  11272=>"101110000",
  11273=>"001001110",
  11274=>"101100101",
  11275=>"101111111",
  11276=>"111100100",
  11277=>"110101110",
  11278=>"010101111",
  11279=>"110100001",
  11280=>"011001001",
  11281=>"011000011",
  11282=>"000000010",
  11283=>"010000110",
  11284=>"111011111",
  11285=>"000000000",
  11286=>"110110000",
  11287=>"111100001",
  11288=>"100011110",
  11289=>"111101011",
  11290=>"001101011",
  11291=>"000011111",
  11292=>"000011011",
  11293=>"011111100",
  11294=>"110100100",
  11295=>"111111001",
  11296=>"100001001",
  11297=>"001011101",
  11298=>"001011110",
  11299=>"100010100",
  11300=>"111111101",
  11301=>"011110100",
  11302=>"000000011",
  11303=>"000000110",
  11304=>"000100110",
  11305=>"000100111",
  11306=>"111100001",
  11307=>"010000110",
  11308=>"100111000",
  11309=>"101110101",
  11310=>"001101000",
  11311=>"001111010",
  11312=>"111101011",
  11313=>"010010010",
  11314=>"011001101",
  11315=>"000101111",
  11316=>"000100111",
  11317=>"011010011",
  11318=>"010100111",
  11319=>"001011111",
  11320=>"101110010",
  11321=>"100101111",
  11322=>"001111000",
  11323=>"010011000",
  11324=>"110010000",
  11325=>"100111000",
  11326=>"000100110",
  11327=>"000110110",
  11328=>"101001010",
  11329=>"000110000",
  11330=>"000010000",
  11331=>"100000000",
  11332=>"110100011",
  11333=>"111111001",
  11334=>"000111101",
  11335=>"000001100",
  11336=>"111101000",
  11337=>"000111000",
  11338=>"110011001",
  11339=>"000001010",
  11340=>"000101011",
  11341=>"000111110",
  11342=>"111001011",
  11343=>"011001101",
  11344=>"001001000",
  11345=>"110100101",
  11346=>"001110110",
  11347=>"010001000",
  11348=>"111000110",
  11349=>"101000001",
  11350=>"010101000",
  11351=>"001001001",
  11352=>"000110001",
  11353=>"001111011",
  11354=>"010001111",
  11355=>"010100000",
  11356=>"000010011",
  11357=>"101011011",
  11358=>"100000001",
  11359=>"001000100",
  11360=>"100110111",
  11361=>"100010000",
  11362=>"011110100",
  11363=>"110011001",
  11364=>"010000000",
  11365=>"010010111",
  11366=>"001001100",
  11367=>"000111010",
  11368=>"100000111",
  11369=>"111111110",
  11370=>"000011101",
  11371=>"000101100",
  11372=>"101111010",
  11373=>"000011101",
  11374=>"010000001",
  11375=>"000101101",
  11376=>"000111100",
  11377=>"011000011",
  11378=>"111111011",
  11379=>"001000011",
  11380=>"011101000",
  11381=>"101100111",
  11382=>"011111110",
  11383=>"100001010",
  11384=>"010010001",
  11385=>"111000101",
  11386=>"010000111",
  11387=>"001000110",
  11388=>"000000010",
  11389=>"001010000",
  11390=>"000100010",
  11391=>"011001001",
  11392=>"000001100",
  11393=>"110010111",
  11394=>"001100000",
  11395=>"101111001",
  11396=>"110010101",
  11397=>"011001101",
  11398=>"000001100",
  11399=>"001100010",
  11400=>"100110010",
  11401=>"100101100",
  11402=>"110110010",
  11403=>"111100011",
  11404=>"010101000",
  11405=>"000010010",
  11406=>"101011111",
  11407=>"011011110",
  11408=>"010101001",
  11409=>"111101001",
  11410=>"100100001",
  11411=>"001001101",
  11412=>"101110100",
  11413=>"001000111",
  11414=>"100101001",
  11415=>"010101111",
  11416=>"101010110",
  11417=>"001011001",
  11418=>"110011100",
  11419=>"100101110",
  11420=>"101100111",
  11421=>"110000111",
  11422=>"000011111",
  11423=>"011011101",
  11424=>"110100010",
  11425=>"000011111",
  11426=>"001010011",
  11427=>"011011110",
  11428=>"011100010",
  11429=>"101110011",
  11430=>"110000010",
  11431=>"101000001",
  11432=>"000000011",
  11433=>"011101000",
  11434=>"111100010",
  11435=>"111100000",
  11436=>"010011000",
  11437=>"111100110",
  11438=>"101101101",
  11439=>"010101100",
  11440=>"100000110",
  11441=>"010000011",
  11442=>"000110010",
  11443=>"101100100",
  11444=>"100010100",
  11445=>"000001001",
  11446=>"100011010",
  11447=>"100000101",
  11448=>"001110000",
  11449=>"011111111",
  11450=>"000001100",
  11451=>"101100111",
  11452=>"111100011",
  11453=>"010110111",
  11454=>"010110011",
  11455=>"000001110",
  11456=>"010011111",
  11457=>"110101111",
  11458=>"001001110",
  11459=>"001011101",
  11460=>"100010010",
  11461=>"000010111",
  11462=>"100001111",
  11463=>"101111000",
  11464=>"010110100",
  11465=>"101111110",
  11466=>"110001101",
  11467=>"001111100",
  11468=>"011001001",
  11469=>"011001101",
  11470=>"010000001",
  11471=>"101011111",
  11472=>"100000000",
  11473=>"101001011",
  11474=>"100111100",
  11475=>"100010000",
  11476=>"101001010",
  11477=>"100011111",
  11478=>"001101000",
  11479=>"101011011",
  11480=>"111011110",
  11481=>"010111011",
  11482=>"011111011",
  11483=>"111010110",
  11484=>"110010010",
  11485=>"101000001",
  11486=>"001010110",
  11487=>"001000000",
  11488=>"101000101",
  11489=>"000010110",
  11490=>"010011001",
  11491=>"000101111",
  11492=>"101110110",
  11493=>"001110000",
  11494=>"111110111",
  11495=>"101100000",
  11496=>"000111110",
  11497=>"000000000",
  11498=>"010100100",
  11499=>"101100100",
  11500=>"001001100",
  11501=>"000010110",
  11502=>"001100110",
  11503=>"101001011",
  11504=>"100011001",
  11505=>"100111100",
  11506=>"111000011",
  11507=>"110111010",
  11508=>"001110011",
  11509=>"101100101",
  11510=>"100000100",
  11511=>"001000000",
  11512=>"000010010",
  11513=>"001000110",
  11514=>"001011001",
  11515=>"011011101",
  11516=>"101010001",
  11517=>"100001010",
  11518=>"011111100",
  11519=>"100101111",
  11520=>"001111010",
  11521=>"000101101",
  11522=>"001110010",
  11523=>"100000101",
  11524=>"000111000",
  11525=>"100010000",
  11526=>"011110111",
  11527=>"001001110",
  11528=>"011111101",
  11529=>"000011001",
  11530=>"100111111",
  11531=>"001011100",
  11532=>"000001010",
  11533=>"000110011",
  11534=>"100001000",
  11535=>"010101000",
  11536=>"111100110",
  11537=>"111000011",
  11538=>"110110001",
  11539=>"000000011",
  11540=>"001000000",
  11541=>"110110001",
  11542=>"000111111",
  11543=>"101010000",
  11544=>"001101110",
  11545=>"010001010",
  11546=>"010101110",
  11547=>"111100011",
  11548=>"011110110",
  11549=>"110111010",
  11550=>"111001101",
  11551=>"011111000",
  11552=>"001001010",
  11553=>"010001110",
  11554=>"000001110",
  11555=>"011100010",
  11556=>"001111000",
  11557=>"111011011",
  11558=>"000000011",
  11559=>"001100101",
  11560=>"001000101",
  11561=>"110101001",
  11562=>"111101010",
  11563=>"000100110",
  11564=>"111000111",
  11565=>"101010011",
  11566=>"000011111",
  11567=>"001100011",
  11568=>"111001101",
  11569=>"010110101",
  11570=>"011000111",
  11571=>"000110010",
  11572=>"011100010",
  11573=>"010011101",
  11574=>"001100001",
  11575=>"111111111",
  11576=>"111100110",
  11577=>"000000001",
  11578=>"001111110",
  11579=>"000101011",
  11580=>"011001110",
  11581=>"110111111",
  11582=>"101000001",
  11583=>"000010101",
  11584=>"110111000",
  11585=>"010110111",
  11586=>"000101001",
  11587=>"111101010",
  11588=>"100000000",
  11589=>"110110110",
  11590=>"111000000",
  11591=>"000101101",
  11592=>"011011000",
  11593=>"000111100",
  11594=>"100011011",
  11595=>"100000011",
  11596=>"010000010",
  11597=>"001101100",
  11598=>"110001111",
  11599=>"000010010",
  11600=>"101011010",
  11601=>"101010101",
  11602=>"000001000",
  11603=>"100000101",
  11604=>"000101000",
  11605=>"101011111",
  11606=>"010101101",
  11607=>"100011110",
  11608=>"001010100",
  11609=>"110101100",
  11610=>"010010000",
  11611=>"000111011",
  11612=>"011111000",
  11613=>"100110011",
  11614=>"100001110",
  11615=>"010010100",
  11616=>"110101100",
  11617=>"000000000",
  11618=>"100001000",
  11619=>"001000110",
  11620=>"110011011",
  11621=>"110000011",
  11622=>"110011111",
  11623=>"011110110",
  11624=>"100111111",
  11625=>"110000101",
  11626=>"000000110",
  11627=>"011110000",
  11628=>"110111011",
  11629=>"111110110",
  11630=>"010000001",
  11631=>"001000001",
  11632=>"000001010",
  11633=>"000111110",
  11634=>"111101010",
  11635=>"111010110",
  11636=>"111010001",
  11637=>"000000110",
  11638=>"111011111",
  11639=>"100101001",
  11640=>"110011101",
  11641=>"101100101",
  11642=>"111110101",
  11643=>"010000000",
  11644=>"001000010",
  11645=>"111100111",
  11646=>"110101110",
  11647=>"111100110",
  11648=>"100111000",
  11649=>"110010100",
  11650=>"011010011",
  11651=>"001111110",
  11652=>"101111101",
  11653=>"001101101",
  11654=>"100110000",
  11655=>"100010110",
  11656=>"101110111",
  11657=>"001010101",
  11658=>"000000000",
  11659=>"100010000",
  11660=>"011010001",
  11661=>"000011111",
  11662=>"001000000",
  11663=>"011111000",
  11664=>"111111110",
  11665=>"101000010",
  11666=>"111011101",
  11667=>"011100111",
  11668=>"001011000",
  11669=>"100001001",
  11670=>"100011101",
  11671=>"001101001",
  11672=>"011111010",
  11673=>"000111110",
  11674=>"010010011",
  11675=>"100110001",
  11676=>"011111001",
  11677=>"001010000",
  11678=>"101000111",
  11679=>"100011101",
  11680=>"110110111",
  11681=>"101100100",
  11682=>"111111010",
  11683=>"010100101",
  11684=>"111110100",
  11685=>"101000011",
  11686=>"100001010",
  11687=>"000100001",
  11688=>"010111111",
  11689=>"001111001",
  11690=>"011110111",
  11691=>"001101111",
  11692=>"010011010",
  11693=>"101111000",
  11694=>"111101011",
  11695=>"011100101",
  11696=>"111100111",
  11697=>"000101101",
  11698=>"001000110",
  11699=>"101101000",
  11700=>"000000101",
  11701=>"101000110",
  11702=>"100011111",
  11703=>"101010001",
  11704=>"101111101",
  11705=>"001010110",
  11706=>"001001010",
  11707=>"000000111",
  11708=>"000000011",
  11709=>"111100110",
  11710=>"100011000",
  11711=>"111101110",
  11712=>"100101110",
  11713=>"000010010",
  11714=>"011010101",
  11715=>"110001001",
  11716=>"110100001",
  11717=>"111110110",
  11718=>"010111111",
  11719=>"000001000",
  11720=>"100110101",
  11721=>"111111000",
  11722=>"001101011",
  11723=>"000000001",
  11724=>"100100001",
  11725=>"100100101",
  11726=>"001000101",
  11727=>"100110001",
  11728=>"100011000",
  11729=>"010000100",
  11730=>"001001011",
  11731=>"101010101",
  11732=>"111110100",
  11733=>"001101000",
  11734=>"010111100",
  11735=>"110101001",
  11736=>"010010001",
  11737=>"010000001",
  11738=>"100010111",
  11739=>"111011111",
  11740=>"010110001",
  11741=>"111011011",
  11742=>"001010100",
  11743=>"111101100",
  11744=>"001000001",
  11745=>"011001001",
  11746=>"100011101",
  11747=>"001100010",
  11748=>"001011111",
  11749=>"100100100",
  11750=>"010010001",
  11751=>"001110100",
  11752=>"001010000",
  11753=>"100011111",
  11754=>"101000000",
  11755=>"111101100",
  11756=>"111111111",
  11757=>"010001000",
  11758=>"000001001",
  11759=>"110000110",
  11760=>"001001101",
  11761=>"000011000",
  11762=>"010010110",
  11763=>"110100110",
  11764=>"011010001",
  11765=>"111111000",
  11766=>"010111000",
  11767=>"000111011",
  11768=>"011000100",
  11769=>"111100000",
  11770=>"111011010",
  11771=>"011111100",
  11772=>"001000001",
  11773=>"101100010",
  11774=>"100000100",
  11775=>"000000001",
  11776=>"100111000",
  11777=>"111010110",
  11778=>"111000010",
  11779=>"110110001",
  11780=>"111011010",
  11781=>"010111111",
  11782=>"111011001",
  11783=>"001001110",
  11784=>"010111110",
  11785=>"101101001",
  11786=>"101010110",
  11787=>"011000000",
  11788=>"011101101",
  11789=>"001100100",
  11790=>"110001100",
  11791=>"010000101",
  11792=>"000111101",
  11793=>"011011011",
  11794=>"010100100",
  11795=>"011011010",
  11796=>"011010110",
  11797=>"110110101",
  11798=>"001011011",
  11799=>"010000000",
  11800=>"110101000",
  11801=>"100001011",
  11802=>"010100001",
  11803=>"110001000",
  11804=>"001001000",
  11805=>"001001101",
  11806=>"101111001",
  11807=>"010010101",
  11808=>"110101001",
  11809=>"111011101",
  11810=>"000110110",
  11811=>"001110100",
  11812=>"111001011",
  11813=>"100111110",
  11814=>"111110001",
  11815=>"000100010",
  11816=>"110010011",
  11817=>"111000011",
  11818=>"100000101",
  11819=>"101001011",
  11820=>"010010010",
  11821=>"000000011",
  11822=>"110110111",
  11823=>"000010101",
  11824=>"101001010",
  11825=>"100101111",
  11826=>"111111000",
  11827=>"000010010",
  11828=>"000101111",
  11829=>"000011101",
  11830=>"001010001",
  11831=>"100011001",
  11832=>"011001010",
  11833=>"001000011",
  11834=>"100100101",
  11835=>"101011111",
  11836=>"100010111",
  11837=>"100110101",
  11838=>"011010000",
  11839=>"011000100",
  11840=>"010110011",
  11841=>"111001001",
  11842=>"101101110",
  11843=>"000010110",
  11844=>"111101011",
  11845=>"111000100",
  11846=>"000000010",
  11847=>"000011001",
  11848=>"100000111",
  11849=>"011010011",
  11850=>"111101100",
  11851=>"111111101",
  11852=>"010101000",
  11853=>"100000100",
  11854=>"110010100",
  11855=>"001100011",
  11856=>"100000110",
  11857=>"111101110",
  11858=>"110110100",
  11859=>"110111110",
  11860=>"110100101",
  11861=>"000001111",
  11862=>"010011011",
  11863=>"100010010",
  11864=>"101000110",
  11865=>"101111110",
  11866=>"100000100",
  11867=>"110011111",
  11868=>"100101110",
  11869=>"101000000",
  11870=>"111001000",
  11871=>"011111101",
  11872=>"001000011",
  11873=>"010110111",
  11874=>"100100000",
  11875=>"000101001",
  11876=>"110100100",
  11877=>"100111110",
  11878=>"111011100",
  11879=>"010010001",
  11880=>"000000010",
  11881=>"000001111",
  11882=>"100000001",
  11883=>"001100001",
  11884=>"101010011",
  11885=>"110100111",
  11886=>"110100010",
  11887=>"000110101",
  11888=>"101010100",
  11889=>"000000000",
  11890=>"110010000",
  11891=>"000101110",
  11892=>"110000001",
  11893=>"001101110",
  11894=>"001101101",
  11895=>"100010000",
  11896=>"111001010",
  11897=>"111100111",
  11898=>"111000101",
  11899=>"100111000",
  11900=>"000011011",
  11901=>"001110110",
  11902=>"100101100",
  11903=>"101110110",
  11904=>"101000001",
  11905=>"010110100",
  11906=>"100101110",
  11907=>"110110100",
  11908=>"000110001",
  11909=>"100111001",
  11910=>"110010001",
  11911=>"001000001",
  11912=>"011101001",
  11913=>"100010111",
  11914=>"000111101",
  11915=>"011111110",
  11916=>"110110100",
  11917=>"110110110",
  11918=>"011100101",
  11919=>"100111100",
  11920=>"010110101",
  11921=>"010101010",
  11922=>"011001110",
  11923=>"011100100",
  11924=>"100101001",
  11925=>"011100010",
  11926=>"110000011",
  11927=>"111110110",
  11928=>"011100111",
  11929=>"010010000",
  11930=>"110000000",
  11931=>"111001111",
  11932=>"111011011",
  11933=>"100100000",
  11934=>"000000010",
  11935=>"110101001",
  11936=>"011101100",
  11937=>"111110101",
  11938=>"001011010",
  11939=>"011100011",
  11940=>"000010101",
  11941=>"001001011",
  11942=>"100011111",
  11943=>"000101110",
  11944=>"110001001",
  11945=>"011100101",
  11946=>"101001101",
  11947=>"010110100",
  11948=>"000011110",
  11949=>"110110000",
  11950=>"011110010",
  11951=>"010010111",
  11952=>"110101011",
  11953=>"100111011",
  11954=>"110011010",
  11955=>"011010100",
  11956=>"000001000",
  11957=>"111111011",
  11958=>"111001010",
  11959=>"001010000",
  11960=>"000011000",
  11961=>"111100001",
  11962=>"000001010",
  11963=>"010011000",
  11964=>"000111100",
  11965=>"110011100",
  11966=>"101101100",
  11967=>"001111001",
  11968=>"110101111",
  11969=>"011110010",
  11970=>"000010000",
  11971=>"010010011",
  11972=>"010100111",
  11973=>"100001001",
  11974=>"100000101",
  11975=>"110110001",
  11976=>"011011000",
  11977=>"010100000",
  11978=>"000100000",
  11979=>"100000100",
  11980=>"010101110",
  11981=>"000100101",
  11982=>"011000101",
  11983=>"010011110",
  11984=>"000110111",
  11985=>"000001010",
  11986=>"010110100",
  11987=>"111100110",
  11988=>"011101110",
  11989=>"110011011",
  11990=>"011100000",
  11991=>"000100101",
  11992=>"110110001",
  11993=>"101010001",
  11994=>"000010001",
  11995=>"101001101",
  11996=>"101111000",
  11997=>"101001101",
  11998=>"000001011",
  11999=>"110000000",
  12000=>"111111110",
  12001=>"100011101",
  12002=>"101101100",
  12003=>"110110011",
  12004=>"011011010",
  12005=>"111101111",
  12006=>"000001111",
  12007=>"001100111",
  12008=>"111011111",
  12009=>"110000110",
  12010=>"111110100",
  12011=>"000011110",
  12012=>"000011001",
  12013=>"000000001",
  12014=>"010110110",
  12015=>"000100100",
  12016=>"001001111",
  12017=>"010010010",
  12018=>"101110011",
  12019=>"001100011",
  12020=>"100010001",
  12021=>"011001110",
  12022=>"010000001",
  12023=>"110001110",
  12024=>"000001100",
  12025=>"010111100",
  12026=>"000001000",
  12027=>"110000011",
  12028=>"011101101",
  12029=>"111100100",
  12030=>"011110110",
  12031=>"001010100",
  12032=>"111101101",
  12033=>"000000110",
  12034=>"111000111",
  12035=>"000010101",
  12036=>"001000000",
  12037=>"110000000",
  12038=>"000111010",
  12039=>"000011111",
  12040=>"000001000",
  12041=>"111110000",
  12042=>"110010011",
  12043=>"001000000",
  12044=>"010101000",
  12045=>"101001100",
  12046=>"111100110",
  12047=>"111100110",
  12048=>"100001111",
  12049=>"101100111",
  12050=>"000010110",
  12051=>"110100001",
  12052=>"000001111",
  12053=>"010001101",
  12054=>"100001000",
  12055=>"011011000",
  12056=>"110001100",
  12057=>"110011011",
  12058=>"000000100",
  12059=>"110110101",
  12060=>"101110111",
  12061=>"111000000",
  12062=>"101011111",
  12063=>"010000001",
  12064=>"000010000",
  12065=>"111111111",
  12066=>"111100111",
  12067=>"011010111",
  12068=>"000011010",
  12069=>"101111110",
  12070=>"110010000",
  12071=>"011001001",
  12072=>"000000110",
  12073=>"000000000",
  12074=>"100011000",
  12075=>"011111101",
  12076=>"001011100",
  12077=>"000010010",
  12078=>"001100010",
  12079=>"110111011",
  12080=>"000000110",
  12081=>"000100010",
  12082=>"101001110",
  12083=>"100101110",
  12084=>"000010000",
  12085=>"010111101",
  12086=>"001011111",
  12087=>"010110001",
  12088=>"100011100",
  12089=>"111011001",
  12090=>"110101111",
  12091=>"001010001",
  12092=>"000010000",
  12093=>"000000010",
  12094=>"111011001",
  12095=>"110110111",
  12096=>"111111011",
  12097=>"000010110",
  12098=>"110000101",
  12099=>"111101000",
  12100=>"101100101",
  12101=>"010000010",
  12102=>"111111100",
  12103=>"011010001",
  12104=>"101000101",
  12105=>"010100011",
  12106=>"001101010",
  12107=>"100011000",
  12108=>"001000010",
  12109=>"101001011",
  12110=>"101110100",
  12111=>"000110010",
  12112=>"100010100",
  12113=>"000000111",
  12114=>"000010101",
  12115=>"111001101",
  12116=>"110010000",
  12117=>"110011001",
  12118=>"110111111",
  12119=>"000000011",
  12120=>"101000100",
  12121=>"100110101",
  12122=>"111000111",
  12123=>"111010001",
  12124=>"111001110",
  12125=>"111110101",
  12126=>"010100100",
  12127=>"101000000",
  12128=>"100101101",
  12129=>"000000000",
  12130=>"001000010",
  12131=>"111100000",
  12132=>"111000101",
  12133=>"001110001",
  12134=>"000101100",
  12135=>"100101010",
  12136=>"001101101",
  12137=>"001111011",
  12138=>"101100000",
  12139=>"011010110",
  12140=>"011100111",
  12141=>"011111111",
  12142=>"110011011",
  12143=>"011110000",
  12144=>"100000101",
  12145=>"001110110",
  12146=>"100111111",
  12147=>"111001011",
  12148=>"101001100",
  12149=>"010110110",
  12150=>"111010111",
  12151=>"000000000",
  12152=>"101011100",
  12153=>"100000011",
  12154=>"111011110",
  12155=>"000011000",
  12156=>"101100110",
  12157=>"010100110",
  12158=>"101101111",
  12159=>"111011001",
  12160=>"000101100",
  12161=>"011100011",
  12162=>"010101101",
  12163=>"001011111",
  12164=>"100101110",
  12165=>"100011100",
  12166=>"011001111",
  12167=>"110100101",
  12168=>"111001001",
  12169=>"000110011",
  12170=>"010110110",
  12171=>"000110011",
  12172=>"101011000",
  12173=>"001110011",
  12174=>"111111011",
  12175=>"000110001",
  12176=>"110111110",
  12177=>"101010101",
  12178=>"100001111",
  12179=>"111000010",
  12180=>"110101110",
  12181=>"001010110",
  12182=>"001000001",
  12183=>"101000101",
  12184=>"010100110",
  12185=>"111001111",
  12186=>"011010111",
  12187=>"011111110",
  12188=>"000001000",
  12189=>"100000011",
  12190=>"000101101",
  12191=>"111000001",
  12192=>"000001010",
  12193=>"111000101",
  12194=>"101011001",
  12195=>"111111011",
  12196=>"100010101",
  12197=>"101110100",
  12198=>"010000011",
  12199=>"000000000",
  12200=>"111001110",
  12201=>"000010010",
  12202=>"111000111",
  12203=>"010111011",
  12204=>"101001101",
  12205=>"110000101",
  12206=>"000011000",
  12207=>"101000011",
  12208=>"010101001",
  12209=>"000011110",
  12210=>"000100111",
  12211=>"101000101",
  12212=>"001110001",
  12213=>"111101001",
  12214=>"010110011",
  12215=>"111111001",
  12216=>"000100110",
  12217=>"000110001",
  12218=>"111000111",
  12219=>"100001101",
  12220=>"011100111",
  12221=>"001100100",
  12222=>"100000111",
  12223=>"011001001",
  12224=>"000001001",
  12225=>"010110000",
  12226=>"110001011",
  12227=>"111111000",
  12228=>"000011110",
  12229=>"110000001",
  12230=>"000101100",
  12231=>"000110011",
  12232=>"100100000",
  12233=>"100001011",
  12234=>"101010100",
  12235=>"111100000",
  12236=>"111011001",
  12237=>"100111110",
  12238=>"111101111",
  12239=>"011000110",
  12240=>"010100100",
  12241=>"110011011",
  12242=>"001000000",
  12243=>"000000001",
  12244=>"110101111",
  12245=>"111001010",
  12246=>"101111000",
  12247=>"111100111",
  12248=>"010010100",
  12249=>"111000101",
  12250=>"110001111",
  12251=>"011000100",
  12252=>"100101000",
  12253=>"000001010",
  12254=>"100111010",
  12255=>"111100000",
  12256=>"001110011",
  12257=>"001011010",
  12258=>"011010011",
  12259=>"010101111",
  12260=>"111010100",
  12261=>"001100101",
  12262=>"010100010",
  12263=>"110111011",
  12264=>"100010101",
  12265=>"011001111",
  12266=>"100101100",
  12267=>"110110110",
  12268=>"010000110",
  12269=>"100110011",
  12270=>"110100001",
  12271=>"001001010",
  12272=>"100101011",
  12273=>"111101011",
  12274=>"000100001",
  12275=>"010010110",
  12276=>"110110110",
  12277=>"000001000",
  12278=>"011011001",
  12279=>"100111011",
  12280=>"000110001",
  12281=>"101010010",
  12282=>"101011001",
  12283=>"000001011",
  12284=>"101100110",
  12285=>"101000001",
  12286=>"000110010",
  12287=>"010110000",
  12288=>"111111111",
  12289=>"100000001",
  12290=>"011000000",
  12291=>"010101001",
  12292=>"010011001",
  12293=>"100000111",
  12294=>"001001100",
  12295=>"110011111",
  12296=>"001111100",
  12297=>"000010011",
  12298=>"100101000",
  12299=>"010110001",
  12300=>"110110110",
  12301=>"000011011",
  12302=>"001000011",
  12303=>"100111100",
  12304=>"100010010",
  12305=>"000110010",
  12306=>"101100111",
  12307=>"001110111",
  12308=>"001001010",
  12309=>"000110111",
  12310=>"101010001",
  12311=>"001001100",
  12312=>"111100110",
  12313=>"000010101",
  12314=>"110010010",
  12315=>"111100110",
  12316=>"010010101",
  12317=>"001110101",
  12318=>"001100000",
  12319=>"110001000",
  12320=>"000010001",
  12321=>"000000111",
  12322=>"101111101",
  12323=>"100011011",
  12324=>"011001000",
  12325=>"101001001",
  12326=>"001010011",
  12327=>"100100100",
  12328=>"111100011",
  12329=>"100000010",
  12330=>"010110000",
  12331=>"101010011",
  12332=>"101010101",
  12333=>"000010011",
  12334=>"001101100",
  12335=>"101100101",
  12336=>"100001110",
  12337=>"110100000",
  12338=>"111010100",
  12339=>"111110111",
  12340=>"000100110",
  12341=>"010010011",
  12342=>"111101000",
  12343=>"100001001",
  12344=>"000000010",
  12345=>"011100111",
  12346=>"101010010",
  12347=>"110100110",
  12348=>"111110010",
  12349=>"011100111",
  12350=>"011001011",
  12351=>"010000010",
  12352=>"000101000",
  12353=>"111010011",
  12354=>"001111000",
  12355=>"110100011",
  12356=>"101010100",
  12357=>"001000000",
  12358=>"011111111",
  12359=>"010100011",
  12360=>"111110101",
  12361=>"011000010",
  12362=>"111000011",
  12363=>"000000011",
  12364=>"110111101",
  12365=>"011101011",
  12366=>"011101000",
  12367=>"100011001",
  12368=>"000011011",
  12369=>"100000001",
  12370=>"001100110",
  12371=>"101010001",
  12372=>"101101000",
  12373=>"100011001",
  12374=>"101111111",
  12375=>"101010111",
  12376=>"111100110",
  12377=>"101111011",
  12378=>"100010010",
  12379=>"011001010",
  12380=>"010000110",
  12381=>"010110110",
  12382=>"000001110",
  12383=>"111111001",
  12384=>"111100101",
  12385=>"000000001",
  12386=>"000000000",
  12387=>"100110111",
  12388=>"001100010",
  12389=>"111000001",
  12390=>"000101110",
  12391=>"011110101",
  12392=>"000100110",
  12393=>"110001111",
  12394=>"010000101",
  12395=>"001100111",
  12396=>"000000110",
  12397=>"110001100",
  12398=>"100000010",
  12399=>"110011000",
  12400=>"010101100",
  12401=>"100111010",
  12402=>"000111011",
  12403=>"100011010",
  12404=>"100101000",
  12405=>"000111111",
  12406=>"110010010",
  12407=>"111100000",
  12408=>"110011101",
  12409=>"010001111",
  12410=>"001101001",
  12411=>"000001100",
  12412=>"111010101",
  12413=>"010000111",
  12414=>"011011001",
  12415=>"100001101",
  12416=>"001001101",
  12417=>"101110010",
  12418=>"011001000",
  12419=>"011111000",
  12420=>"010011101",
  12421=>"010011110",
  12422=>"101101010",
  12423=>"101100010",
  12424=>"011111010",
  12425=>"011011110",
  12426=>"111011110",
  12427=>"001100101",
  12428=>"101111110",
  12429=>"111111010",
  12430=>"010101011",
  12431=>"100011110",
  12432=>"011011001",
  12433=>"111001011",
  12434=>"100110110",
  12435=>"111000111",
  12436=>"110101100",
  12437=>"001101010",
  12438=>"110100000",
  12439=>"111000100",
  12440=>"001000000",
  12441=>"000111100",
  12442=>"110000111",
  12443=>"111001010",
  12444=>"000000100",
  12445=>"101100101",
  12446=>"100010000",
  12447=>"001010101",
  12448=>"100010001",
  12449=>"101001011",
  12450=>"000111100",
  12451=>"000010010",
  12452=>"110001010",
  12453=>"010100010",
  12454=>"110100100",
  12455=>"011001000",
  12456=>"010110110",
  12457=>"011001110",
  12458=>"011010011",
  12459=>"110011011",
  12460=>"000110011",
  12461=>"011110010",
  12462=>"110110010",
  12463=>"001100011",
  12464=>"001100010",
  12465=>"101101010",
  12466=>"010010011",
  12467=>"010000000",
  12468=>"001000000",
  12469=>"101100100",
  12470=>"000010110",
  12471=>"111001110",
  12472=>"100111111",
  12473=>"001010001",
  12474=>"001110001",
  12475=>"011011001",
  12476=>"000101111",
  12477=>"111100101",
  12478=>"000000101",
  12479=>"100000001",
  12480=>"010010000",
  12481=>"001100000",
  12482=>"100010010",
  12483=>"101101110",
  12484=>"010110010",
  12485=>"001101010",
  12486=>"100000111",
  12487=>"110011001",
  12488=>"011111111",
  12489=>"001101101",
  12490=>"001100001",
  12491=>"010101110",
  12492=>"100011101",
  12493=>"000000100",
  12494=>"101100100",
  12495=>"010111110",
  12496=>"111001101",
  12497=>"100010101",
  12498=>"101001101",
  12499=>"011100010",
  12500=>"100101100",
  12501=>"011111100",
  12502=>"110010101",
  12503=>"100011001",
  12504=>"001001011",
  12505=>"001000100",
  12506=>"000100000",
  12507=>"110011101",
  12508=>"010011010",
  12509=>"111111110",
  12510=>"000110000",
  12511=>"111100100",
  12512=>"101010001",
  12513=>"000111011",
  12514=>"011110001",
  12515=>"001000000",
  12516=>"011011001",
  12517=>"100110011",
  12518=>"111110000",
  12519=>"111111011",
  12520=>"000100010",
  12521=>"001111101",
  12522=>"001010000",
  12523=>"100110111",
  12524=>"010110110",
  12525=>"010110101",
  12526=>"010001101",
  12527=>"110101001",
  12528=>"110010011",
  12529=>"000000011",
  12530=>"000100100",
  12531=>"100000101",
  12532=>"101010111",
  12533=>"010001011",
  12534=>"000100000",
  12535=>"000010101",
  12536=>"111001100",
  12537=>"010011111",
  12538=>"111010111",
  12539=>"100000100",
  12540=>"001110101",
  12541=>"100001100",
  12542=>"110101011",
  12543=>"011011011",
  12544=>"011011101",
  12545=>"111011010",
  12546=>"111100010",
  12547=>"010101011",
  12548=>"111101101",
  12549=>"000000000",
  12550=>"000010001",
  12551=>"100001100",
  12552=>"110001010",
  12553=>"100010000",
  12554=>"101000101",
  12555=>"111011100",
  12556=>"000000010",
  12557=>"101001101",
  12558=>"110000000",
  12559=>"001000000",
  12560=>"010010111",
  12561=>"100001010",
  12562=>"000000101",
  12563=>"111011000",
  12564=>"100010101",
  12565=>"001100101",
  12566=>"101100100",
  12567=>"010110101",
  12568=>"011000010",
  12569=>"010110100",
  12570=>"011001100",
  12571=>"011000001",
  12572=>"111111010",
  12573=>"011110000",
  12574=>"101001111",
  12575=>"010101000",
  12576=>"000000100",
  12577=>"001111010",
  12578=>"111110111",
  12579=>"011110101",
  12580=>"011101011",
  12581=>"001001010",
  12582=>"110101111",
  12583=>"101011001",
  12584=>"010101110",
  12585=>"101011001",
  12586=>"100011001",
  12587=>"010010110",
  12588=>"110000010",
  12589=>"101011101",
  12590=>"110011011",
  12591=>"111110100",
  12592=>"100110011",
  12593=>"000111100",
  12594=>"111110110",
  12595=>"100000001",
  12596=>"011010011",
  12597=>"101000000",
  12598=>"011111100",
  12599=>"100111000",
  12600=>"001000001",
  12601=>"010000011",
  12602=>"111010011",
  12603=>"011110010",
  12604=>"111101111",
  12605=>"111111010",
  12606=>"001001110",
  12607=>"001111111",
  12608=>"100110001",
  12609=>"101011111",
  12610=>"111111111",
  12611=>"010110010",
  12612=>"000000100",
  12613=>"011001011",
  12614=>"000001101",
  12615=>"100001011",
  12616=>"000010111",
  12617=>"111011010",
  12618=>"000101011",
  12619=>"010100011",
  12620=>"111011111",
  12621=>"111101110",
  12622=>"001100100",
  12623=>"000011100",
  12624=>"110010110",
  12625=>"100001101",
  12626=>"110010010",
  12627=>"110000001",
  12628=>"100110111",
  12629=>"011010010",
  12630=>"000000110",
  12631=>"100110100",
  12632=>"000101000",
  12633=>"100011100",
  12634=>"111011001",
  12635=>"111010010",
  12636=>"001000001",
  12637=>"100011101",
  12638=>"110001000",
  12639=>"010010000",
  12640=>"101001001",
  12641=>"110011111",
  12642=>"000110000",
  12643=>"010100110",
  12644=>"101111101",
  12645=>"110001100",
  12646=>"000110011",
  12647=>"001100111",
  12648=>"000111000",
  12649=>"010101100",
  12650=>"000100001",
  12651=>"110010011",
  12652=>"011001000",
  12653=>"100011001",
  12654=>"001010000",
  12655=>"101001011",
  12656=>"110110101",
  12657=>"001000001",
  12658=>"011100111",
  12659=>"010010000",
  12660=>"000100010",
  12661=>"111100100",
  12662=>"010100011",
  12663=>"011010011",
  12664=>"100001110",
  12665=>"001110101",
  12666=>"101011011",
  12667=>"100101101",
  12668=>"100011100",
  12669=>"001111110",
  12670=>"101011101",
  12671=>"000100000",
  12672=>"001011111",
  12673=>"100001100",
  12674=>"101001101",
  12675=>"100001111",
  12676=>"111100011",
  12677=>"110100010",
  12678=>"100111001",
  12679=>"100010001",
  12680=>"110000000",
  12681=>"100100000",
  12682=>"000000111",
  12683=>"100011000",
  12684=>"110111100",
  12685=>"010011001",
  12686=>"111111111",
  12687=>"010001100",
  12688=>"010010000",
  12689=>"010000100",
  12690=>"110000000",
  12691=>"000000110",
  12692=>"000011111",
  12693=>"100100000",
  12694=>"111111110",
  12695=>"111010111",
  12696=>"010001001",
  12697=>"100100100",
  12698=>"001001000",
  12699=>"010001000",
  12700=>"111001110",
  12701=>"100100001",
  12702=>"010100000",
  12703=>"011000100",
  12704=>"101100100",
  12705=>"001001011",
  12706=>"000100111",
  12707=>"100000001",
  12708=>"011100010",
  12709=>"011011011",
  12710=>"100001000",
  12711=>"110110011",
  12712=>"010010011",
  12713=>"000110000",
  12714=>"100000010",
  12715=>"010100001",
  12716=>"011110001",
  12717=>"010110011",
  12718=>"011001101",
  12719=>"111111110",
  12720=>"111110111",
  12721=>"010100010",
  12722=>"001100001",
  12723=>"101100000",
  12724=>"001000101",
  12725=>"011110010",
  12726=>"101110100",
  12727=>"101111101",
  12728=>"010001110",
  12729=>"001010101",
  12730=>"111010111",
  12731=>"001011011",
  12732=>"101001010",
  12733=>"101001000",
  12734=>"000001010",
  12735=>"111111000",
  12736=>"110000111",
  12737=>"010010100",
  12738=>"000010111",
  12739=>"110011010",
  12740=>"111111000",
  12741=>"010110100",
  12742=>"110111011",
  12743=>"000010000",
  12744=>"111100000",
  12745=>"100000000",
  12746=>"000110010",
  12747=>"010100101",
  12748=>"011000100",
  12749=>"011010001",
  12750=>"111110011",
  12751=>"110011000",
  12752=>"111001101",
  12753=>"110101011",
  12754=>"001110110",
  12755=>"110000000",
  12756=>"101000111",
  12757=>"011011001",
  12758=>"100101000",
  12759=>"001100010",
  12760=>"001111010",
  12761=>"000111111",
  12762=>"111000110",
  12763=>"010000100",
  12764=>"110110010",
  12765=>"101100000",
  12766=>"100101100",
  12767=>"111010010",
  12768=>"111111010",
  12769=>"000101111",
  12770=>"110010110",
  12771=>"001011001",
  12772=>"011001001",
  12773=>"001100101",
  12774=>"001011001",
  12775=>"100100011",
  12776=>"000000110",
  12777=>"011110011",
  12778=>"011010111",
  12779=>"101101111",
  12780=>"011010000",
  12781=>"011011101",
  12782=>"011110101",
  12783=>"110111101",
  12784=>"111111111",
  12785=>"111100100",
  12786=>"100000000",
  12787=>"011110100",
  12788=>"011001101",
  12789=>"011000011",
  12790=>"100011100",
  12791=>"000001000",
  12792=>"100110110",
  12793=>"001000011",
  12794=>"000000111",
  12795=>"010111010",
  12796=>"100111010",
  12797=>"101000011",
  12798=>"110000111",
  12799=>"011010101",
  12800=>"111010110",
  12801=>"000111101",
  12802=>"011100010",
  12803=>"110110010",
  12804=>"011110100",
  12805=>"100000000",
  12806=>"110101011",
  12807=>"100101100",
  12808=>"001010101",
  12809=>"010101110",
  12810=>"111010101",
  12811=>"010110100",
  12812=>"101100110",
  12813=>"110100111",
  12814=>"111101111",
  12815=>"110010100",
  12816=>"010111101",
  12817=>"010010000",
  12818=>"010111000",
  12819=>"001100110",
  12820=>"010000111",
  12821=>"111111011",
  12822=>"111001010",
  12823=>"010001001",
  12824=>"010100101",
  12825=>"001000101",
  12826=>"111110111",
  12827=>"000001000",
  12828=>"101111110",
  12829=>"100011111",
  12830=>"000100111",
  12831=>"111000111",
  12832=>"110100100",
  12833=>"101011001",
  12834=>"100111001",
  12835=>"001110011",
  12836=>"111100011",
  12837=>"001010101",
  12838=>"101111011",
  12839=>"010110100",
  12840=>"110010000",
  12841=>"110001001",
  12842=>"000100000",
  12843=>"001100110",
  12844=>"000011000",
  12845=>"000011110",
  12846=>"011000100",
  12847=>"101001101",
  12848=>"010101000",
  12849=>"011011110",
  12850=>"111001110",
  12851=>"101111111",
  12852=>"001001000",
  12853=>"000001100",
  12854=>"101101000",
  12855=>"110000010",
  12856=>"100001111",
  12857=>"000011100",
  12858=>"110001010",
  12859=>"111110010",
  12860=>"001000110",
  12861=>"011000011",
  12862=>"001010000",
  12863=>"111010110",
  12864=>"001010111",
  12865=>"000011100",
  12866=>"011111011",
  12867=>"001110111",
  12868=>"111011101",
  12869=>"011001010",
  12870=>"001110111",
  12871=>"010001101",
  12872=>"101001110",
  12873=>"101100110",
  12874=>"110011110",
  12875=>"111101101",
  12876=>"101011100",
  12877=>"010000010",
  12878=>"000001111",
  12879=>"001001001",
  12880=>"011011000",
  12881=>"110011000",
  12882=>"001111110",
  12883=>"000001001",
  12884=>"110011001",
  12885=>"110110101",
  12886=>"101101111",
  12887=>"110010110",
  12888=>"100101111",
  12889=>"110100001",
  12890=>"111111000",
  12891=>"010101111",
  12892=>"101010001",
  12893=>"111010000",
  12894=>"110110010",
  12895=>"100100010",
  12896=>"001010111",
  12897=>"110101101",
  12898=>"100001010",
  12899=>"111100100",
  12900=>"001110001",
  12901=>"101100000",
  12902=>"111011010",
  12903=>"001001101",
  12904=>"000101111",
  12905=>"100011000",
  12906=>"001000110",
  12907=>"110111101",
  12908=>"011011011",
  12909=>"000000000",
  12910=>"101100011",
  12911=>"110010011",
  12912=>"101001011",
  12913=>"000110101",
  12914=>"000001001",
  12915=>"101101010",
  12916=>"011000001",
  12917=>"110011011",
  12918=>"000110001",
  12919=>"010010011",
  12920=>"001011011",
  12921=>"000101001",
  12922=>"000011111",
  12923=>"101001001",
  12924=>"111011010",
  12925=>"110100111",
  12926=>"111001101",
  12927=>"100001111",
  12928=>"010111000",
  12929=>"000011110",
  12930=>"110101101",
  12931=>"011000001",
  12932=>"000110111",
  12933=>"101110000",
  12934=>"111101110",
  12935=>"110101110",
  12936=>"010011111",
  12937=>"011111001",
  12938=>"100110010",
  12939=>"000110111",
  12940=>"100010100",
  12941=>"101001101",
  12942=>"000100100",
  12943=>"111100010",
  12944=>"111001110",
  12945=>"101001000",
  12946=>"100100101",
  12947=>"001000011",
  12948=>"000000101",
  12949=>"110011101",
  12950=>"001010101",
  12951=>"001000000",
  12952=>"100100011",
  12953=>"000000001",
  12954=>"100100100",
  12955=>"111010101",
  12956=>"100010000",
  12957=>"101101100",
  12958=>"110010010",
  12959=>"001101111",
  12960=>"011111000",
  12961=>"010000110",
  12962=>"110001111",
  12963=>"110100011",
  12964=>"001100011",
  12965=>"100100110",
  12966=>"100110100",
  12967=>"000010101",
  12968=>"011000101",
  12969=>"101010001",
  12970=>"000000001",
  12971=>"100110000",
  12972=>"101011010",
  12973=>"000000110",
  12974=>"101100110",
  12975=>"000000110",
  12976=>"010100111",
  12977=>"100010100",
  12978=>"000001010",
  12979=>"110100111",
  12980=>"001110101",
  12981=>"000001101",
  12982=>"011111001",
  12983=>"000100100",
  12984=>"111111100",
  12985=>"010110010",
  12986=>"110001110",
  12987=>"010100001",
  12988=>"000010101",
  12989=>"010010100",
  12990=>"111100000",
  12991=>"011011001",
  12992=>"101000101",
  12993=>"101111110",
  12994=>"010001111",
  12995=>"110000011",
  12996=>"111000001",
  12997=>"010010000",
  12998=>"001011010",
  12999=>"101010010",
  13000=>"101000100",
  13001=>"111001010",
  13002=>"010000111",
  13003=>"001111101",
  13004=>"011011110",
  13005=>"011111100",
  13006=>"001100110",
  13007=>"010100111",
  13008=>"110110010",
  13009=>"111110111",
  13010=>"001101111",
  13011=>"101000110",
  13012=>"111010111",
  13013=>"011111101",
  13014=>"011010110",
  13015=>"111001011",
  13016=>"100111000",
  13017=>"001110110",
  13018=>"110011010",
  13019=>"000101010",
  13020=>"111110001",
  13021=>"110110011",
  13022=>"000001011",
  13023=>"001110110",
  13024=>"111100000",
  13025=>"000000010",
  13026=>"000110100",
  13027=>"001110111",
  13028=>"000011000",
  13029=>"110111010",
  13030=>"110111111",
  13031=>"111111111",
  13032=>"000111111",
  13033=>"101110000",
  13034=>"111100001",
  13035=>"011111101",
  13036=>"100111010",
  13037=>"010011010",
  13038=>"111110010",
  13039=>"000110000",
  13040=>"111111001",
  13041=>"000101011",
  13042=>"110101110",
  13043=>"101100100",
  13044=>"100001011",
  13045=>"000010100",
  13046=>"101001001",
  13047=>"011100111",
  13048=>"010001110",
  13049=>"011101010",
  13050=>"110100010",
  13051=>"110000101",
  13052=>"000001100",
  13053=>"101101011",
  13054=>"001000001",
  13055=>"110000101",
  13056=>"000011001",
  13057=>"101110100",
  13058=>"101010000",
  13059=>"001110001",
  13060=>"010111101",
  13061=>"100000110",
  13062=>"010100100",
  13063=>"111011110",
  13064=>"000000100",
  13065=>"000011010",
  13066=>"100011000",
  13067=>"111001100",
  13068=>"111011001",
  13069=>"000000010",
  13070=>"000011110",
  13071=>"110100010",
  13072=>"010100001",
  13073=>"000011010",
  13074=>"110100100",
  13075=>"111111011",
  13076=>"110001110",
  13077=>"000111000",
  13078=>"000101101",
  13079=>"000010010",
  13080=>"000000001",
  13081=>"000011111",
  13082=>"001100000",
  13083=>"111101001",
  13084=>"011010100",
  13085=>"011010011",
  13086=>"000111001",
  13087=>"100111011",
  13088=>"011010011",
  13089=>"111001010",
  13090=>"001100001",
  13091=>"111111000",
  13092=>"010000100",
  13093=>"110110111",
  13094=>"111110100",
  13095=>"000010110",
  13096=>"111000100",
  13097=>"011111100",
  13098=>"001101011",
  13099=>"000000101",
  13100=>"011011010",
  13101=>"111101010",
  13102=>"011101000",
  13103=>"101111110",
  13104=>"010101101",
  13105=>"011011111",
  13106=>"101100101",
  13107=>"100000101",
  13108=>"001110000",
  13109=>"100100111",
  13110=>"100100111",
  13111=>"001110000",
  13112=>"110011001",
  13113=>"110011001",
  13114=>"000111100",
  13115=>"111101010",
  13116=>"110011110",
  13117=>"000100010",
  13118=>"100000111",
  13119=>"010110010",
  13120=>"101000100",
  13121=>"111100000",
  13122=>"111101010",
  13123=>"100110101",
  13124=>"111100100",
  13125=>"111110111",
  13126=>"111011001",
  13127=>"000100100",
  13128=>"111010100",
  13129=>"001111010",
  13130=>"101001000",
  13131=>"110010111",
  13132=>"010010001",
  13133=>"111011000",
  13134=>"000010010",
  13135=>"110011101",
  13136=>"101100000",
  13137=>"010000000",
  13138=>"110111000",
  13139=>"001000101",
  13140=>"011000011",
  13141=>"011101100",
  13142=>"010111100",
  13143=>"111110010",
  13144=>"001111101",
  13145=>"000111100",
  13146=>"101000110",
  13147=>"000000010",
  13148=>"000111000",
  13149=>"101001101",
  13150=>"011010100",
  13151=>"111101000",
  13152=>"011101110",
  13153=>"000001100",
  13154=>"110011110",
  13155=>"001100010",
  13156=>"001000010",
  13157=>"111001110",
  13158=>"100010001",
  13159=>"001011000",
  13160=>"001001011",
  13161=>"111101100",
  13162=>"011100101",
  13163=>"000101011",
  13164=>"110111001",
  13165=>"010101011",
  13166=>"001010000",
  13167=>"111001100",
  13168=>"001011101",
  13169=>"000001010",
  13170=>"010011000",
  13171=>"010110010",
  13172=>"100111001",
  13173=>"101010110",
  13174=>"000000011",
  13175=>"101110010",
  13176=>"110111011",
  13177=>"110010101",
  13178=>"100000000",
  13179=>"111100011",
  13180=>"101110101",
  13181=>"111100110",
  13182=>"101010110",
  13183=>"010010000",
  13184=>"000011000",
  13185=>"000010000",
  13186=>"000111111",
  13187=>"000110110",
  13188=>"110000010",
  13189=>"101101110",
  13190=>"101000010",
  13191=>"110111010",
  13192=>"110000101",
  13193=>"101111000",
  13194=>"101111101",
  13195=>"100000101",
  13196=>"001111001",
  13197=>"010000001",
  13198=>"000100100",
  13199=>"001101101",
  13200=>"001011111",
  13201=>"110111001",
  13202=>"000100001",
  13203=>"011100100",
  13204=>"010011110",
  13205=>"111000010",
  13206=>"101100001",
  13207=>"100010001",
  13208=>"110000101",
  13209=>"100000001",
  13210=>"000000001",
  13211=>"001111001",
  13212=>"100001100",
  13213=>"010111101",
  13214=>"001100101",
  13215=>"110000000",
  13216=>"011010010",
  13217=>"110100001",
  13218=>"011000010",
  13219=>"000101011",
  13220=>"111100100",
  13221=>"001111010",
  13222=>"000010001",
  13223=>"111100011",
  13224=>"010110010",
  13225=>"100000000",
  13226=>"111001101",
  13227=>"011010000",
  13228=>"101010010",
  13229=>"111000111",
  13230=>"111010001",
  13231=>"111101100",
  13232=>"111010000",
  13233=>"011101110",
  13234=>"110011010",
  13235=>"111111110",
  13236=>"011101111",
  13237=>"100010110",
  13238=>"100011110",
  13239=>"110110100",
  13240=>"110010111",
  13241=>"011001101",
  13242=>"001010100",
  13243=>"110110101",
  13244=>"011101100",
  13245=>"000010000",
  13246=>"110100000",
  13247=>"011111001",
  13248=>"000011101",
  13249=>"000011100",
  13250=>"111100101",
  13251=>"000001110",
  13252=>"100101110",
  13253=>"101010010",
  13254=>"100011110",
  13255=>"101000101",
  13256=>"000010000",
  13257=>"010100010",
  13258=>"010000001",
  13259=>"001101111",
  13260=>"000101101",
  13261=>"010111101",
  13262=>"101110000",
  13263=>"000011000",
  13264=>"110111001",
  13265=>"011011001",
  13266=>"011110111",
  13267=>"010011001",
  13268=>"010101101",
  13269=>"101100110",
  13270=>"101101000",
  13271=>"011101111",
  13272=>"111010010",
  13273=>"100000001",
  13274=>"101000000",
  13275=>"101001011",
  13276=>"000101100",
  13277=>"111111010",
  13278=>"101100010",
  13279=>"010010001",
  13280=>"100011000",
  13281=>"001001011",
  13282=>"001100110",
  13283=>"001001101",
  13284=>"001100011",
  13285=>"001001110",
  13286=>"001011011",
  13287=>"110101100",
  13288=>"000110110",
  13289=>"111110010",
  13290=>"011110100",
  13291=>"010011111",
  13292=>"110000001",
  13293=>"011000010",
  13294=>"111011101",
  13295=>"111000100",
  13296=>"111110001",
  13297=>"111100011",
  13298=>"000011100",
  13299=>"011010000",
  13300=>"111001100",
  13301=>"111111001",
  13302=>"001101011",
  13303=>"110101010",
  13304=>"101110010",
  13305=>"000111101",
  13306=>"111111110",
  13307=>"111000110",
  13308=>"011001101",
  13309=>"001010011",
  13310=>"110010110",
  13311=>"011011100",
  13312=>"110000110",
  13313=>"001100010",
  13314=>"001001010",
  13315=>"000010010",
  13316=>"010111010",
  13317=>"111110100",
  13318=>"001101001",
  13319=>"001011100",
  13320=>"111001000",
  13321=>"110010001",
  13322=>"001000111",
  13323=>"010101000",
  13324=>"100011110",
  13325=>"001110111",
  13326=>"111110111",
  13327=>"100101001",
  13328=>"111010010",
  13329=>"100111001",
  13330=>"110000000",
  13331=>"101001011",
  13332=>"100110100",
  13333=>"100000001",
  13334=>"101010111",
  13335=>"111001000",
  13336=>"101110110",
  13337=>"100011010",
  13338=>"010000101",
  13339=>"010110100",
  13340=>"111110010",
  13341=>"111001111",
  13342=>"100110111",
  13343=>"011111000",
  13344=>"110111110",
  13345=>"000000000",
  13346=>"011100110",
  13347=>"001100111",
  13348=>"101010011",
  13349=>"111100011",
  13350=>"111110000",
  13351=>"101110110",
  13352=>"100011101",
  13353=>"001000010",
  13354=>"000000010",
  13355=>"000100111",
  13356=>"000010000",
  13357=>"100000000",
  13358=>"100101000",
  13359=>"011001011",
  13360=>"111011011",
  13361=>"100011110",
  13362=>"010001100",
  13363=>"101100001",
  13364=>"000011001",
  13365=>"010010100",
  13366=>"100101011",
  13367=>"111010110",
  13368=>"000001011",
  13369=>"010100000",
  13370=>"100101111",
  13371=>"100111010",
  13372=>"101100110",
  13373=>"000110011",
  13374=>"000001101",
  13375=>"001000010",
  13376=>"010000010",
  13377=>"001000110",
  13378=>"110000001",
  13379=>"001001001",
  13380=>"001111001",
  13381=>"101010100",
  13382=>"011011110",
  13383=>"100111101",
  13384=>"011001111",
  13385=>"100101000",
  13386=>"001011100",
  13387=>"101111110",
  13388=>"111001111",
  13389=>"000000111",
  13390=>"110110011",
  13391=>"101111101",
  13392=>"010110001",
  13393=>"001010001",
  13394=>"000001100",
  13395=>"010110111",
  13396=>"011101001",
  13397=>"000010011",
  13398=>"000111001",
  13399=>"000000110",
  13400=>"101110111",
  13401=>"011111110",
  13402=>"110010111",
  13403=>"010011000",
  13404=>"011000100",
  13405=>"101010100",
  13406=>"001101010",
  13407=>"110110111",
  13408=>"101011101",
  13409=>"011001010",
  13410=>"101010111",
  13411=>"001100100",
  13412=>"010000000",
  13413=>"110010110",
  13414=>"101100100",
  13415=>"110001000",
  13416=>"100000101",
  13417=>"001010011",
  13418=>"000000000",
  13419=>"000011100",
  13420=>"100110010",
  13421=>"100001010",
  13422=>"101101011",
  13423=>"101000001",
  13424=>"001011101",
  13425=>"010100011",
  13426=>"000111001",
  13427=>"011010010",
  13428=>"010101110",
  13429=>"101001011",
  13430=>"111100111",
  13431=>"011000011",
  13432=>"001001000",
  13433=>"101101100",
  13434=>"111110111",
  13435=>"011010110",
  13436=>"110111111",
  13437=>"000001011",
  13438=>"011010111",
  13439=>"110000010",
  13440=>"000110000",
  13441=>"100111111",
  13442=>"001000100",
  13443=>"011111111",
  13444=>"111010001",
  13445=>"010111001",
  13446=>"010111110",
  13447=>"010011010",
  13448=>"000000011",
  13449=>"000101000",
  13450=>"111001001",
  13451=>"100011111",
  13452=>"101100101",
  13453=>"011100101",
  13454=>"101010001",
  13455=>"011001000",
  13456=>"111011110",
  13457=>"010110100",
  13458=>"110110101",
  13459=>"110110100",
  13460=>"101100110",
  13461=>"100011101",
  13462=>"100001101",
  13463=>"101000110",
  13464=>"000100110",
  13465=>"101100100",
  13466=>"100001000",
  13467=>"001001110",
  13468=>"111011001",
  13469=>"000010100",
  13470=>"100010011",
  13471=>"011010111",
  13472=>"111101111",
  13473=>"101001011",
  13474=>"100100001",
  13475=>"010110111",
  13476=>"101000000",
  13477=>"011001101",
  13478=>"101001100",
  13479=>"000111101",
  13480=>"101000111",
  13481=>"011111100",
  13482=>"101000000",
  13483=>"110001000",
  13484=>"001101000",
  13485=>"001011010",
  13486=>"100111101",
  13487=>"100110101",
  13488=>"000110011",
  13489=>"101111001",
  13490=>"100111010",
  13491=>"100001100",
  13492=>"110110000",
  13493=>"011000101",
  13494=>"011101111",
  13495=>"100011000",
  13496=>"111010101",
  13497=>"111111001",
  13498=>"100010101",
  13499=>"000101001",
  13500=>"000111111",
  13501=>"001110100",
  13502=>"010001001",
  13503=>"010010000",
  13504=>"100000001",
  13505=>"100100000",
  13506=>"111100101",
  13507=>"000100111",
  13508=>"101100010",
  13509=>"001011101",
  13510=>"000111110",
  13511=>"101100100",
  13512=>"100010110",
  13513=>"111010111",
  13514=>"001001000",
  13515=>"110111010",
  13516=>"010001001",
  13517=>"011000000",
  13518=>"000000101",
  13519=>"001111101",
  13520=>"100100000",
  13521=>"011000110",
  13522=>"100100110",
  13523=>"010000010",
  13524=>"101100010",
  13525=>"110111011",
  13526=>"101110111",
  13527=>"000000001",
  13528=>"011100001",
  13529=>"100011111",
  13530=>"110011101",
  13531=>"001010111",
  13532=>"011000000",
  13533=>"001100111",
  13534=>"011010111",
  13535=>"011111010",
  13536=>"100110100",
  13537=>"100101010",
  13538=>"111010100",
  13539=>"111100100",
  13540=>"111101010",
  13541=>"101010000",
  13542=>"011110011",
  13543=>"001110010",
  13544=>"010111001",
  13545=>"001101010",
  13546=>"001100101",
  13547=>"101000111",
  13548=>"001011100",
  13549=>"110010110",
  13550=>"100100011",
  13551=>"101000010",
  13552=>"111010011",
  13553=>"011000100",
  13554=>"100010100",
  13555=>"100110101",
  13556=>"110101000",
  13557=>"010101110",
  13558=>"010001101",
  13559=>"101000110",
  13560=>"010100110",
  13561=>"110110001",
  13562=>"010110000",
  13563=>"011000011",
  13564=>"111101100",
  13565=>"011101100",
  13566=>"111101101",
  13567=>"011110110",
  13568=>"100111100",
  13569=>"010111001",
  13570=>"101000110",
  13571=>"110110011",
  13572=>"100110000",
  13573=>"111101101",
  13574=>"010100111",
  13575=>"010001100",
  13576=>"100011001",
  13577=>"001001110",
  13578=>"011100011",
  13579=>"111011111",
  13580=>"110101001",
  13581=>"011110011",
  13582=>"100000101",
  13583=>"101000101",
  13584=>"010001111",
  13585=>"001001001",
  13586=>"000000000",
  13587=>"100001001",
  13588=>"101001011",
  13589=>"010001001",
  13590=>"100111101",
  13591=>"110111010",
  13592=>"101000100",
  13593=>"001000111",
  13594=>"110100001",
  13595=>"101110001",
  13596=>"111010110",
  13597=>"101101000",
  13598=>"110011100",
  13599=>"100010100",
  13600=>"010010011",
  13601=>"100111100",
  13602=>"111001111",
  13603=>"101101111",
  13604=>"011001001",
  13605=>"111010111",
  13606=>"100001000",
  13607=>"001100101",
  13608=>"001101000",
  13609=>"100011101",
  13610=>"011011010",
  13611=>"000001001",
  13612=>"100000111",
  13613=>"000101111",
  13614=>"110111010",
  13615=>"011110100",
  13616=>"000011000",
  13617=>"001111000",
  13618=>"011011011",
  13619=>"011110001",
  13620=>"010000001",
  13621=>"100111101",
  13622=>"110011000",
  13623=>"110011100",
  13624=>"100010110",
  13625=>"110011101",
  13626=>"100110100",
  13627=>"110110100",
  13628=>"001010110",
  13629=>"100011111",
  13630=>"111110111",
  13631=>"011001011",
  13632=>"100001010",
  13633=>"000000010",
  13634=>"111010011",
  13635=>"110111010",
  13636=>"101001111",
  13637=>"111000110",
  13638=>"011101001",
  13639=>"000010100",
  13640=>"110011010",
  13641=>"111110011",
  13642=>"001100000",
  13643=>"000110100",
  13644=>"001111001",
  13645=>"001011110",
  13646=>"111111001",
  13647=>"001000001",
  13648=>"101010010",
  13649=>"101100001",
  13650=>"000010101",
  13651=>"001010100",
  13652=>"101100111",
  13653=>"110111110",
  13654=>"011100101",
  13655=>"001000000",
  13656=>"000001011",
  13657=>"111010111",
  13658=>"001111100",
  13659=>"000000001",
  13660=>"011110110",
  13661=>"010111111",
  13662=>"011101100",
  13663=>"011000000",
  13664=>"110011011",
  13665=>"011001101",
  13666=>"100000110",
  13667=>"111110010",
  13668=>"011000101",
  13669=>"000000001",
  13670=>"010110001",
  13671=>"100011110",
  13672=>"011111101",
  13673=>"001111110",
  13674=>"111010111",
  13675=>"000111001",
  13676=>"011110100",
  13677=>"111011101",
  13678=>"000101010",
  13679=>"010011010",
  13680=>"000000000",
  13681=>"010111111",
  13682=>"100000000",
  13683=>"001010101",
  13684=>"111011001",
  13685=>"000101011",
  13686=>"110111101",
  13687=>"011111011",
  13688=>"001100100",
  13689=>"001000000",
  13690=>"011100100",
  13691=>"011110100",
  13692=>"100011011",
  13693=>"111011100",
  13694=>"000001000",
  13695=>"111111000",
  13696=>"110111110",
  13697=>"010010001",
  13698=>"010010110",
  13699=>"110100100",
  13700=>"010001111",
  13701=>"001000110",
  13702=>"110101100",
  13703=>"010100111",
  13704=>"100011000",
  13705=>"110010001",
  13706=>"101001011",
  13707=>"010001111",
  13708=>"000010000",
  13709=>"011111110",
  13710=>"000111010",
  13711=>"111001111",
  13712=>"111000110",
  13713=>"001001111",
  13714=>"011001000",
  13715=>"101111101",
  13716=>"011000111",
  13717=>"100011100",
  13718=>"111111000",
  13719=>"010100000",
  13720=>"110001101",
  13721=>"000011110",
  13722=>"011111110",
  13723=>"110011011",
  13724=>"100010000",
  13725=>"011110101",
  13726=>"100100001",
  13727=>"011010001",
  13728=>"111001000",
  13729=>"000000011",
  13730=>"101011010",
  13731=>"000010100",
  13732=>"001001011",
  13733=>"111011111",
  13734=>"011101101",
  13735=>"001101000",
  13736=>"011001001",
  13737=>"000010000",
  13738=>"100101110",
  13739=>"001000001",
  13740=>"010100010",
  13741=>"111101100",
  13742=>"001110011",
  13743=>"010101000",
  13744=>"101110011",
  13745=>"101111110",
  13746=>"001101100",
  13747=>"100011110",
  13748=>"010110111",
  13749=>"001110100",
  13750=>"000101101",
  13751=>"111111110",
  13752=>"110111000",
  13753=>"111101011",
  13754=>"111101010",
  13755=>"110001010",
  13756=>"111010101",
  13757=>"001000011",
  13758=>"110011010",
  13759=>"111011010",
  13760=>"100100010",
  13761=>"110011111",
  13762=>"100100000",
  13763=>"011000101",
  13764=>"111001010",
  13765=>"000101011",
  13766=>"100110101",
  13767=>"111100000",
  13768=>"111010011",
  13769=>"100111011",
  13770=>"001101110",
  13771=>"001101101",
  13772=>"010100000",
  13773=>"101101000",
  13774=>"110000110",
  13775=>"001101010",
  13776=>"110111111",
  13777=>"100111100",
  13778=>"011101100",
  13779=>"000010010",
  13780=>"101111111",
  13781=>"111110001",
  13782=>"011111111",
  13783=>"101100110",
  13784=>"001100111",
  13785=>"011110010",
  13786=>"010000100",
  13787=>"110100101",
  13788=>"111111110",
  13789=>"011010010",
  13790=>"111111011",
  13791=>"101101111",
  13792=>"101011110",
  13793=>"000110011",
  13794=>"110111101",
  13795=>"011110110",
  13796=>"010101110",
  13797=>"110010101",
  13798=>"001011100",
  13799=>"110000110",
  13800=>"010111001",
  13801=>"010000001",
  13802=>"110000110",
  13803=>"001001010",
  13804=>"000001001",
  13805=>"100001011",
  13806=>"101101111",
  13807=>"001001100",
  13808=>"111100110",
  13809=>"001011100",
  13810=>"111101110",
  13811=>"111100111",
  13812=>"010110000",
  13813=>"000010010",
  13814=>"100111001",
  13815=>"111000100",
  13816=>"010101111",
  13817=>"111000001",
  13818=>"110011000",
  13819=>"001010101",
  13820=>"010111110",
  13821=>"101010101",
  13822=>"010111000",
  13823=>"100000111",
  13824=>"101001111",
  13825=>"010011011",
  13826=>"100110001",
  13827=>"000011100",
  13828=>"111110100",
  13829=>"111000011",
  13830=>"000101011",
  13831=>"111100110",
  13832=>"111111101",
  13833=>"001011111",
  13834=>"111010111",
  13835=>"001110000",
  13836=>"001011110",
  13837=>"101000110",
  13838=>"001110000",
  13839=>"101101101",
  13840=>"001111001",
  13841=>"100001101",
  13842=>"010000011",
  13843=>"111001011",
  13844=>"000100000",
  13845=>"111000010",
  13846=>"110110000",
  13847=>"000001001",
  13848=>"101001111",
  13849=>"100010000",
  13850=>"000111010",
  13851=>"111001101",
  13852=>"000010110",
  13853=>"100101000",
  13854=>"101111001",
  13855=>"010000000",
  13856=>"011110000",
  13857=>"111000110",
  13858=>"000001000",
  13859=>"110110111",
  13860=>"110011011",
  13861=>"011011010",
  13862=>"001000111",
  13863=>"100101011",
  13864=>"110101011",
  13865=>"011100010",
  13866=>"101001111",
  13867=>"101010001",
  13868=>"110001010",
  13869=>"000011001",
  13870=>"111001111",
  13871=>"001001010",
  13872=>"011011100",
  13873=>"010000110",
  13874=>"011111110",
  13875=>"100101001",
  13876=>"001110011",
  13877=>"110111001",
  13878=>"001111100",
  13879=>"010101110",
  13880=>"011110101",
  13881=>"010010100",
  13882=>"011000001",
  13883=>"110101111",
  13884=>"100111111",
  13885=>"010100010",
  13886=>"110010000",
  13887=>"001010010",
  13888=>"011011011",
  13889=>"111100001",
  13890=>"010100100",
  13891=>"011000011",
  13892=>"101010111",
  13893=>"010101000",
  13894=>"011111111",
  13895=>"110000010",
  13896=>"011111111",
  13897=>"111001100",
  13898=>"010011100",
  13899=>"000011111",
  13900=>"011100101",
  13901=>"001000011",
  13902=>"001110011",
  13903=>"011100111",
  13904=>"000010101",
  13905=>"010001100",
  13906=>"000110100",
  13907=>"000111100",
  13908=>"010110000",
  13909=>"000101110",
  13910=>"000011001",
  13911=>"101001011",
  13912=>"101100011",
  13913=>"010000101",
  13914=>"000100100",
  13915=>"000100001",
  13916=>"100110010",
  13917=>"001111011",
  13918=>"000011111",
  13919=>"110010101",
  13920=>"011111011",
  13921=>"010011000",
  13922=>"011111110",
  13923=>"001000101",
  13924=>"111001101",
  13925=>"001010010",
  13926=>"111110001",
  13927=>"010011011",
  13928=>"100011000",
  13929=>"111100000",
  13930=>"111010001",
  13931=>"111100110",
  13932=>"110111110",
  13933=>"000110110",
  13934=>"011111110",
  13935=>"111100000",
  13936=>"011001010",
  13937=>"100100010",
  13938=>"001110010",
  13939=>"100100100",
  13940=>"001100111",
  13941=>"000010100",
  13942=>"110000101",
  13943=>"111100100",
  13944=>"011010110",
  13945=>"110011110",
  13946=>"110000100",
  13947=>"110110100",
  13948=>"000001111",
  13949=>"100101001",
  13950=>"101111111",
  13951=>"011000101",
  13952=>"101001110",
  13953=>"100000000",
  13954=>"100000010",
  13955=>"001001101",
  13956=>"111100011",
  13957=>"111001110",
  13958=>"110101001",
  13959=>"000010010",
  13960=>"010111100",
  13961=>"110111100",
  13962=>"101001010",
  13963=>"110110111",
  13964=>"110101111",
  13965=>"110000110",
  13966=>"010101011",
  13967=>"111000010",
  13968=>"010110110",
  13969=>"101011001",
  13970=>"011110100",
  13971=>"101011110",
  13972=>"101010001",
  13973=>"101011010",
  13974=>"000001001",
  13975=>"110000000",
  13976=>"000001010",
  13977=>"101100000",
  13978=>"111100011",
  13979=>"110101010",
  13980=>"110000100",
  13981=>"011110001",
  13982=>"111101101",
  13983=>"000100100",
  13984=>"101100011",
  13985=>"101010001",
  13986=>"100111001",
  13987=>"010000000",
  13988=>"111111101",
  13989=>"011000111",
  13990=>"111001001",
  13991=>"100010011",
  13992=>"010101101",
  13993=>"101111011",
  13994=>"000001101",
  13995=>"101100100",
  13996=>"101011000",
  13997=>"010001111",
  13998=>"100010111",
  13999=>"001111001",
  14000=>"000000001",
  14001=>"110110110",
  14002=>"011100010",
  14003=>"011100110",
  14004=>"011011000",
  14005=>"100101111",
  14006=>"010010011",
  14007=>"111000101",
  14008=>"110100100",
  14009=>"101101001",
  14010=>"101110010",
  14011=>"011000010",
  14012=>"111101100",
  14013=>"110001100",
  14014=>"100001010",
  14015=>"001110100",
  14016=>"000111110",
  14017=>"010100011",
  14018=>"111111100",
  14019=>"011101110",
  14020=>"110001000",
  14021=>"001001100",
  14022=>"011000011",
  14023=>"101001000",
  14024=>"111011111",
  14025=>"110010100",
  14026=>"001110001",
  14027=>"011000110",
  14028=>"110001000",
  14029=>"110110110",
  14030=>"000101000",
  14031=>"110001000",
  14032=>"111110100",
  14033=>"000000100",
  14034=>"110000010",
  14035=>"011001100",
  14036=>"001001000",
  14037=>"010001111",
  14038=>"001100001",
  14039=>"010010000",
  14040=>"111000011",
  14041=>"111101101",
  14042=>"110010101",
  14043=>"100001100",
  14044=>"000001111",
  14045=>"010010001",
  14046=>"111011010",
  14047=>"101100111",
  14048=>"100110101",
  14049=>"100111011",
  14050=>"000101110",
  14051=>"011100111",
  14052=>"111110000",
  14053=>"000010001",
  14054=>"001000000",
  14055=>"011001010",
  14056=>"110111011",
  14057=>"000100011",
  14058=>"011101110",
  14059=>"010000100",
  14060=>"000010011",
  14061=>"100000110",
  14062=>"001101110",
  14063=>"000111011",
  14064=>"111011001",
  14065=>"111000011",
  14066=>"100100010",
  14067=>"001111000",
  14068=>"010101111",
  14069=>"110000101",
  14070=>"001111100",
  14071=>"110010110",
  14072=>"001101111",
  14073=>"100111110",
  14074=>"011100011",
  14075=>"000111100",
  14076=>"001001010",
  14077=>"010001100",
  14078=>"101101001",
  14079=>"111101000",
  14080=>"010010100",
  14081=>"010011010",
  14082=>"010100110",
  14083=>"110110000",
  14084=>"010001100",
  14085=>"000101100",
  14086=>"011000100",
  14087=>"101100010",
  14088=>"011100110",
  14089=>"110110101",
  14090=>"011010111",
  14091=>"010000010",
  14092=>"110101001",
  14093=>"110101111",
  14094=>"101011101",
  14095=>"100000010",
  14096=>"000010001",
  14097=>"000011100",
  14098=>"100011101",
  14099=>"101011110",
  14100=>"001101111",
  14101=>"000010000",
  14102=>"010011110",
  14103=>"100000001",
  14104=>"100101100",
  14105=>"111011010",
  14106=>"011110011",
  14107=>"101110010",
  14108=>"010110111",
  14109=>"011101001",
  14110=>"110101000",
  14111=>"100101000",
  14112=>"001000001",
  14113=>"110001110",
  14114=>"010100101",
  14115=>"100100110",
  14116=>"011110010",
  14117=>"010011010",
  14118=>"111111111",
  14119=>"101100001",
  14120=>"001101111",
  14121=>"110111100",
  14122=>"000000110",
  14123=>"101100101",
  14124=>"110001001",
  14125=>"100001001",
  14126=>"001111110",
  14127=>"100010011",
  14128=>"001110000",
  14129=>"101011111",
  14130=>"100111111",
  14131=>"011111111",
  14132=>"111000111",
  14133=>"111001110",
  14134=>"110010010",
  14135=>"101101100",
  14136=>"101111001",
  14137=>"100010110",
  14138=>"111100100",
  14139=>"010110000",
  14140=>"001101011",
  14141=>"110000101",
  14142=>"011001010",
  14143=>"111110110",
  14144=>"011110110",
  14145=>"011010011",
  14146=>"101100111",
  14147=>"101111111",
  14148=>"110011101",
  14149=>"001011111",
  14150=>"001000111",
  14151=>"001100101",
  14152=>"100110000",
  14153=>"111000001",
  14154=>"100011101",
  14155=>"110111111",
  14156=>"110100101",
  14157=>"001010110",
  14158=>"000000110",
  14159=>"011100000",
  14160=>"101000011",
  14161=>"001110101",
  14162=>"110000101",
  14163=>"001100110",
  14164=>"101010011",
  14165=>"000111000",
  14166=>"110001010",
  14167=>"000010001",
  14168=>"111011011",
  14169=>"001010111",
  14170=>"001101111",
  14171=>"100111011",
  14172=>"000100010",
  14173=>"101000101",
  14174=>"111011010",
  14175=>"100000101",
  14176=>"100110111",
  14177=>"011111000",
  14178=>"101010111",
  14179=>"110001001",
  14180=>"101000010",
  14181=>"110101110",
  14182=>"110010111",
  14183=>"000110011",
  14184=>"101010111",
  14185=>"000000111",
  14186=>"001111010",
  14187=>"000010010",
  14188=>"111110011",
  14189=>"100101000",
  14190=>"101011110",
  14191=>"000001111",
  14192=>"000010001",
  14193=>"011000111",
  14194=>"111010111",
  14195=>"110011101",
  14196=>"011010101",
  14197=>"001110101",
  14198=>"111000110",
  14199=>"001011111",
  14200=>"010010011",
  14201=>"001000011",
  14202=>"110111011",
  14203=>"111000100",
  14204=>"010101010",
  14205=>"000000011",
  14206=>"000101101",
  14207=>"110011111",
  14208=>"010100100",
  14209=>"100000100",
  14210=>"011010010",
  14211=>"000010100",
  14212=>"111011011",
  14213=>"111010000",
  14214=>"111110000",
  14215=>"110011010",
  14216=>"111110110",
  14217=>"000001001",
  14218=>"011001101",
  14219=>"110000111",
  14220=>"111101001",
  14221=>"101111001",
  14222=>"010101011",
  14223=>"101001001",
  14224=>"101101110",
  14225=>"001010011",
  14226=>"000100011",
  14227=>"111011000",
  14228=>"011100000",
  14229=>"100000110",
  14230=>"100010001",
  14231=>"001011001",
  14232=>"111001010",
  14233=>"000100010",
  14234=>"010110110",
  14235=>"101011111",
  14236=>"111000000",
  14237=>"100111111",
  14238=>"001111010",
  14239=>"000000000",
  14240=>"101010111",
  14241=>"101001101",
  14242=>"000101111",
  14243=>"100000110",
  14244=>"101010110",
  14245=>"111010100",
  14246=>"000011011",
  14247=>"100001010",
  14248=>"000101101",
  14249=>"110000011",
  14250=>"011000010",
  14251=>"011001011",
  14252=>"110000010",
  14253=>"000000101",
  14254=>"110010100",
  14255=>"001000001",
  14256=>"111001000",
  14257=>"111011110",
  14258=>"100111101",
  14259=>"010000101",
  14260=>"100101000",
  14261=>"111000111",
  14262=>"000001001",
  14263=>"101010000",
  14264=>"111011011",
  14265=>"001010111",
  14266=>"011101101",
  14267=>"011111000",
  14268=>"100111100",
  14269=>"101101101",
  14270=>"101001010",
  14271=>"110011101",
  14272=>"110110111",
  14273=>"011101000",
  14274=>"101000111",
  14275=>"001110100",
  14276=>"010011001",
  14277=>"110111101",
  14278=>"011111111",
  14279=>"011011101",
  14280=>"000001111",
  14281=>"011010110",
  14282=>"101010011",
  14283=>"100011011",
  14284=>"001000110",
  14285=>"000001100",
  14286=>"110100010",
  14287=>"100111010",
  14288=>"101100100",
  14289=>"101100100",
  14290=>"000110101",
  14291=>"111100110",
  14292=>"111111001",
  14293=>"101110101",
  14294=>"100011011",
  14295=>"011011010",
  14296=>"111101001",
  14297=>"001010101",
  14298=>"000010011",
  14299=>"001011001",
  14300=>"010100101",
  14301=>"100110110",
  14302=>"000000111",
  14303=>"100101101",
  14304=>"110110111",
  14305=>"011111111",
  14306=>"111101100",
  14307=>"100010011",
  14308=>"011101111",
  14309=>"000001110",
  14310=>"110110100",
  14311=>"100111011",
  14312=>"100101011",
  14313=>"001000110",
  14314=>"010111101",
  14315=>"000001110",
  14316=>"001100001",
  14317=>"100100000",
  14318=>"011100000",
  14319=>"000100110",
  14320=>"101111110",
  14321=>"110000010",
  14322=>"000110111",
  14323=>"101011101",
  14324=>"100010000",
  14325=>"100011101",
  14326=>"101001001",
  14327=>"100000100",
  14328=>"111100101",
  14329=>"110100111",
  14330=>"111110100",
  14331=>"010111111",
  14332=>"000010010",
  14333=>"111001010",
  14334=>"000000011",
  14335=>"110001000",
  14336=>"110111101",
  14337=>"001100011",
  14338=>"001001001",
  14339=>"100001011",
  14340=>"111101110",
  14341=>"110010011",
  14342=>"101110101",
  14343=>"000001111",
  14344=>"000100110",
  14345=>"010010110",
  14346=>"000110010",
  14347=>"110100111",
  14348=>"110100011",
  14349=>"001001101",
  14350=>"001000100",
  14351=>"010111110",
  14352=>"111111000",
  14353=>"110110000",
  14354=>"010100001",
  14355=>"000011100",
  14356=>"001101110",
  14357=>"001111111",
  14358=>"100001000",
  14359=>"100010000",
  14360=>"100001001",
  14361=>"010101101",
  14362=>"110110101",
  14363=>"000100111",
  14364=>"100011100",
  14365=>"011000010",
  14366=>"100001011",
  14367=>"111001010",
  14368=>"000010111",
  14369=>"010001010",
  14370=>"100110001",
  14371=>"010001110",
  14372=>"001101010",
  14373=>"010010110",
  14374=>"111110111",
  14375=>"000110001",
  14376=>"110010001",
  14377=>"011110000",
  14378=>"101000111",
  14379=>"111010100",
  14380=>"100111011",
  14381=>"101011000",
  14382=>"010100010",
  14383=>"110001011",
  14384=>"010110110",
  14385=>"110011010",
  14386=>"001000001",
  14387=>"010110001",
  14388=>"000010100",
  14389=>"111100100",
  14390=>"011011010",
  14391=>"011011000",
  14392=>"100000110",
  14393=>"011010110",
  14394=>"101000010",
  14395=>"001110100",
  14396=>"110001111",
  14397=>"000100011",
  14398=>"100001011",
  14399=>"000100110",
  14400=>"101000011",
  14401=>"000010000",
  14402=>"101010011",
  14403=>"000101100",
  14404=>"110000000",
  14405=>"100111101",
  14406=>"000101110",
  14407=>"111100111",
  14408=>"011100000",
  14409=>"000101001",
  14410=>"111110001",
  14411=>"001111101",
  14412=>"110110010",
  14413=>"110010001",
  14414=>"100000100",
  14415=>"101000000",
  14416=>"100011101",
  14417=>"000000001",
  14418=>"100110011",
  14419=>"101011011",
  14420=>"011010110",
  14421=>"101011110",
  14422=>"000000110",
  14423=>"010011101",
  14424=>"010111011",
  14425=>"100011111",
  14426=>"100001000",
  14427=>"101001100",
  14428=>"001100110",
  14429=>"111110010",
  14430=>"101011100",
  14431=>"100101111",
  14432=>"111111100",
  14433=>"100000100",
  14434=>"111100111",
  14435=>"001111110",
  14436=>"100101001",
  14437=>"000001110",
  14438=>"001101101",
  14439=>"000000111",
  14440=>"100010111",
  14441=>"101100101",
  14442=>"011011101",
  14443=>"000111000",
  14444=>"011010000",
  14445=>"000100101",
  14446=>"010000001",
  14447=>"000011010",
  14448=>"011100000",
  14449=>"111001101",
  14450=>"011011001",
  14451=>"100010010",
  14452=>"010100111",
  14453=>"010010010",
  14454=>"010111001",
  14455=>"100100011",
  14456=>"111100101",
  14457=>"000011100",
  14458=>"101011011",
  14459=>"111100011",
  14460=>"001010111",
  14461=>"110111000",
  14462=>"101101000",
  14463=>"001111100",
  14464=>"100111101",
  14465=>"001001000",
  14466=>"110111101",
  14467=>"100110011",
  14468=>"000001000",
  14469=>"110101001",
  14470=>"100010110",
  14471=>"001110011",
  14472=>"111110011",
  14473=>"110010111",
  14474=>"111001110",
  14475=>"101001001",
  14476=>"101110101",
  14477=>"101101101",
  14478=>"011111001",
  14479=>"111100110",
  14480=>"001001101",
  14481=>"111011100",
  14482=>"010111111",
  14483=>"111110011",
  14484=>"111101001",
  14485=>"101010101",
  14486=>"011000010",
  14487=>"010111000",
  14488=>"000100000",
  14489=>"010111000",
  14490=>"111111100",
  14491=>"101111001",
  14492=>"110111111",
  14493=>"101110111",
  14494=>"110000100",
  14495=>"111110100",
  14496=>"000100010",
  14497=>"011100101",
  14498=>"110111101",
  14499=>"011110110",
  14500=>"000011011",
  14501=>"000001110",
  14502=>"111010000",
  14503=>"010010101",
  14504=>"101101111",
  14505=>"101010100",
  14506=>"000000000",
  14507=>"111000000",
  14508=>"011010110",
  14509=>"000011110",
  14510=>"000010111",
  14511=>"111011011",
  14512=>"010001100",
  14513=>"001000010",
  14514=>"001000010",
  14515=>"000110100",
  14516=>"111100101",
  14517=>"010101101",
  14518=>"101101011",
  14519=>"011111001",
  14520=>"011110100",
  14521=>"101011110",
  14522=>"111001010",
  14523=>"110000110",
  14524=>"010100000",
  14525=>"001011001",
  14526=>"100010010",
  14527=>"010101101",
  14528=>"000010110",
  14529=>"110110001",
  14530=>"001011010",
  14531=>"000001001",
  14532=>"101100011",
  14533=>"010000010",
  14534=>"111101100",
  14535=>"001000000",
  14536=>"100001000",
  14537=>"001001001",
  14538=>"010011001",
  14539=>"101001000",
  14540=>"101010000",
  14541=>"101101001",
  14542=>"111100100",
  14543=>"001101101",
  14544=>"011001101",
  14545=>"100001010",
  14546=>"000110111",
  14547=>"100011000",
  14548=>"100111111",
  14549=>"101100111",
  14550=>"111010100",
  14551=>"010010100",
  14552=>"000010101",
  14553=>"111100101",
  14554=>"110001100",
  14555=>"001001000",
  14556=>"101100110",
  14557=>"011000100",
  14558=>"011010110",
  14559=>"101110000",
  14560=>"110111000",
  14561=>"110010011",
  14562=>"011101101",
  14563=>"111101111",
  14564=>"111001010",
  14565=>"011010111",
  14566=>"010010100",
  14567=>"011001110",
  14568=>"111011010",
  14569=>"101010110",
  14570=>"110110101",
  14571=>"000000000",
  14572=>"111100010",
  14573=>"001000100",
  14574=>"010100110",
  14575=>"111111010",
  14576=>"001010000",
  14577=>"111010111",
  14578=>"110010111",
  14579=>"111001110",
  14580=>"001110010",
  14581=>"000101101",
  14582=>"000111110",
  14583=>"011011000",
  14584=>"110001011",
  14585=>"111100101",
  14586=>"101110111",
  14587=>"000011011",
  14588=>"101001000",
  14589=>"001000110",
  14590=>"000010100",
  14591=>"010011000",
  14592=>"111110010",
  14593=>"000111101",
  14594=>"010000110",
  14595=>"110011001",
  14596=>"000101100",
  14597=>"001101111",
  14598=>"111110111",
  14599=>"111000010",
  14600=>"010101000",
  14601=>"010101010",
  14602=>"010100101",
  14603=>"010010000",
  14604=>"010011010",
  14605=>"000001000",
  14606=>"000100011",
  14607=>"000100000",
  14608=>"011011000",
  14609=>"010000001",
  14610=>"000001111",
  14611=>"111111100",
  14612=>"101110001",
  14613=>"101110011",
  14614=>"000001001",
  14615=>"111010111",
  14616=>"100000011",
  14617=>"111101011",
  14618=>"111111011",
  14619=>"110100110",
  14620=>"010011111",
  14621=>"011011001",
  14622=>"010001110",
  14623=>"011010000",
  14624=>"101110101",
  14625=>"001000111",
  14626=>"010110000",
  14627=>"010011011",
  14628=>"000110001",
  14629=>"111000100",
  14630=>"011111000",
  14631=>"001101011",
  14632=>"001111100",
  14633=>"101010110",
  14634=>"010011101",
  14635=>"111110010",
  14636=>"000101000",
  14637=>"101101101",
  14638=>"001000100",
  14639=>"101100001",
  14640=>"101000000",
  14641=>"111100110",
  14642=>"011001000",
  14643=>"000111110",
  14644=>"000010100",
  14645=>"001100111",
  14646=>"011011010",
  14647=>"001001001",
  14648=>"010111010",
  14649=>"101000010",
  14650=>"101000100",
  14651=>"110110111",
  14652=>"100111000",
  14653=>"111011010",
  14654=>"010101001",
  14655=>"010010100",
  14656=>"111110110",
  14657=>"110100010",
  14658=>"111001111",
  14659=>"100101001",
  14660=>"100011111",
  14661=>"111000101",
  14662=>"000011001",
  14663=>"000010000",
  14664=>"011011111",
  14665=>"111001101",
  14666=>"010010010",
  14667=>"000000011",
  14668=>"000010100",
  14669=>"101110110",
  14670=>"111101011",
  14671=>"110101001",
  14672=>"111110001",
  14673=>"110111100",
  14674=>"111100111",
  14675=>"001001000",
  14676=>"000010101",
  14677=>"110101110",
  14678=>"110110011",
  14679=>"010111011",
  14680=>"000011010",
  14681=>"000010000",
  14682=>"010000110",
  14683=>"111001001",
  14684=>"010100100",
  14685=>"111111111",
  14686=>"011011101",
  14687=>"110000110",
  14688=>"111011100",
  14689=>"100100011",
  14690=>"100111000",
  14691=>"001001010",
  14692=>"111000011",
  14693=>"001010011",
  14694=>"010011010",
  14695=>"110000000",
  14696=>"110100110",
  14697=>"111110111",
  14698=>"110110001",
  14699=>"010100100",
  14700=>"000000110",
  14701=>"011001000",
  14702=>"101000000",
  14703=>"001100010",
  14704=>"111111101",
  14705=>"000101010",
  14706=>"100111111",
  14707=>"110110100",
  14708=>"010101100",
  14709=>"111111111",
  14710=>"110000101",
  14711=>"110100010",
  14712=>"100110000",
  14713=>"000001001",
  14714=>"011011011",
  14715=>"011010100",
  14716=>"101001000",
  14717=>"011111000",
  14718=>"101101000",
  14719=>"101011100",
  14720=>"101111111",
  14721=>"110110111",
  14722=>"010000010",
  14723=>"010001000",
  14724=>"101011100",
  14725=>"000101100",
  14726=>"111110010",
  14727=>"100111111",
  14728=>"000110111",
  14729=>"111010111",
  14730=>"111011101",
  14731=>"011101110",
  14732=>"011111111",
  14733=>"110001010",
  14734=>"000100000",
  14735=>"110001101",
  14736=>"011100111",
  14737=>"110001010",
  14738=>"000000110",
  14739=>"101010111",
  14740=>"000100000",
  14741=>"110101010",
  14742=>"111100110",
  14743=>"001100000",
  14744=>"101101001",
  14745=>"100010110",
  14746=>"001010101",
  14747=>"011101001",
  14748=>"101100000",
  14749=>"001000001",
  14750=>"010000010",
  14751=>"101010100",
  14752=>"101000011",
  14753=>"100001111",
  14754=>"111111111",
  14755=>"110111111",
  14756=>"100101111",
  14757=>"001110110",
  14758=>"101000101",
  14759=>"011011000",
  14760=>"000110010",
  14761=>"111100111",
  14762=>"001011010",
  14763=>"100000001",
  14764=>"101110110",
  14765=>"101000111",
  14766=>"111010110",
  14767=>"111111001",
  14768=>"100111000",
  14769=>"111011011",
  14770=>"000001000",
  14771=>"011101000",
  14772=>"000010001",
  14773=>"100100011",
  14774=>"101001111",
  14775=>"010000100",
  14776=>"111101010",
  14777=>"000100100",
  14778=>"010001010",
  14779=>"100001011",
  14780=>"111011010",
  14781=>"110111100",
  14782=>"111111111",
  14783=>"000001101",
  14784=>"110101011",
  14785=>"010011111",
  14786=>"010110011",
  14787=>"110111010",
  14788=>"110011110",
  14789=>"101000000",
  14790=>"110111100",
  14791=>"001000000",
  14792=>"010001011",
  14793=>"000101110",
  14794=>"000111111",
  14795=>"000101110",
  14796=>"111100010",
  14797=>"110000100",
  14798=>"111000111",
  14799=>"100000010",
  14800=>"100111000",
  14801=>"000111100",
  14802=>"001000000",
  14803=>"010100100",
  14804=>"000101101",
  14805=>"100000101",
  14806=>"011001010",
  14807=>"111101100",
  14808=>"000001000",
  14809=>"001100101",
  14810=>"010110011",
  14811=>"000011110",
  14812=>"101101001",
  14813=>"110000110",
  14814=>"001101001",
  14815=>"100011101",
  14816=>"111101101",
  14817=>"001001001",
  14818=>"101111101",
  14819=>"101000111",
  14820=>"110010101",
  14821=>"101100010",
  14822=>"000011101",
  14823=>"000110010",
  14824=>"010001111",
  14825=>"001011111",
  14826=>"110010011",
  14827=>"110100001",
  14828=>"110111000",
  14829=>"011001000",
  14830=>"110011110",
  14831=>"011100010",
  14832=>"100111110",
  14833=>"001111100",
  14834=>"101000110",
  14835=>"010001001",
  14836=>"000101001",
  14837=>"010000011",
  14838=>"001111010",
  14839=>"000111001",
  14840=>"111111000",
  14841=>"001010110",
  14842=>"001000110",
  14843=>"000000111",
  14844=>"110011111",
  14845=>"001011010",
  14846=>"000110010",
  14847=>"011001000",
  14848=>"100001110",
  14849=>"101011000",
  14850=>"011010001",
  14851=>"000000001",
  14852=>"001001001",
  14853=>"111010101",
  14854=>"011110111",
  14855=>"011000000",
  14856=>"001110011",
  14857=>"010010001",
  14858=>"100000100",
  14859=>"110000101",
  14860=>"011101110",
  14861=>"011001000",
  14862=>"100110101",
  14863=>"001000101",
  14864=>"110101110",
  14865=>"011101100",
  14866=>"100000000",
  14867=>"010010011",
  14868=>"010001010",
  14869=>"000110000",
  14870=>"100000100",
  14871=>"111011011",
  14872=>"011001000",
  14873=>"000001111",
  14874=>"110001000",
  14875=>"011011100",
  14876=>"001010011",
  14877=>"100100110",
  14878=>"001000000",
  14879=>"100011111",
  14880=>"100111001",
  14881=>"001111011",
  14882=>"000101100",
  14883=>"101101111",
  14884=>"010000001",
  14885=>"100111110",
  14886=>"000101011",
  14887=>"100100111",
  14888=>"011100111",
  14889=>"010001110",
  14890=>"111010011",
  14891=>"110111000",
  14892=>"010001100",
  14893=>"101111111",
  14894=>"100001111",
  14895=>"111100100",
  14896=>"111100101",
  14897=>"111110000",
  14898=>"000000000",
  14899=>"010100000",
  14900=>"101010001",
  14901=>"011111001",
  14902=>"001010011",
  14903=>"100010110",
  14904=>"011100010",
  14905=>"110111101",
  14906=>"010100010",
  14907=>"011110010",
  14908=>"110110000",
  14909=>"010111010",
  14910=>"110101111",
  14911=>"100111111",
  14912=>"101101110",
  14913=>"100100100",
  14914=>"100000010",
  14915=>"001101100",
  14916=>"001110111",
  14917=>"011110110",
  14918=>"011010000",
  14919=>"001000011",
  14920=>"011001110",
  14921=>"011001011",
  14922=>"010000001",
  14923=>"111011101",
  14924=>"000000000",
  14925=>"111101101",
  14926=>"110111111",
  14927=>"011100110",
  14928=>"111110111",
  14929=>"001110010",
  14930=>"100111110",
  14931=>"011101101",
  14932=>"010101101",
  14933=>"001000011",
  14934=>"001100001",
  14935=>"010001010",
  14936=>"010111111",
  14937=>"100010101",
  14938=>"000110110",
  14939=>"000101001",
  14940=>"001011111",
  14941=>"001100100",
  14942=>"000011101",
  14943=>"000000100",
  14944=>"011011010",
  14945=>"110110001",
  14946=>"111111111",
  14947=>"001111011",
  14948=>"011011101",
  14949=>"111001000",
  14950=>"111011111",
  14951=>"110010101",
  14952=>"011000000",
  14953=>"010011111",
  14954=>"110001011",
  14955=>"100000000",
  14956=>"110011111",
  14957=>"001000001",
  14958=>"110010111",
  14959=>"110011010",
  14960=>"000100001",
  14961=>"111011011",
  14962=>"111011111",
  14963=>"001101101",
  14964=>"001101101",
  14965=>"000010101",
  14966=>"011011100",
  14967=>"000010011",
  14968=>"111100001",
  14969=>"010101001",
  14970=>"101101101",
  14971=>"001001110",
  14972=>"000100000",
  14973=>"111011001",
  14974=>"100001011",
  14975=>"001001001",
  14976=>"101101100",
  14977=>"011011110",
  14978=>"011110011",
  14979=>"000010000",
  14980=>"100001110",
  14981=>"001111111",
  14982=>"100010000",
  14983=>"101001101",
  14984=>"000001110",
  14985=>"000010000",
  14986=>"010001011",
  14987=>"001000101",
  14988=>"111011011",
  14989=>"100101011",
  14990=>"111111000",
  14991=>"101010111",
  14992=>"101010011",
  14993=>"010010000",
  14994=>"000101101",
  14995=>"111101100",
  14996=>"111010111",
  14997=>"101000110",
  14998=>"110000001",
  14999=>"011111000",
  15000=>"101101101",
  15001=>"111000011",
  15002=>"111101000",
  15003=>"001011011",
  15004=>"000001111",
  15005=>"000110110",
  15006=>"010111101",
  15007=>"001000101",
  15008=>"100101101",
  15009=>"110001001",
  15010=>"011000011",
  15011=>"101010101",
  15012=>"001101100",
  15013=>"111011001",
  15014=>"110000110",
  15015=>"011111001",
  15016=>"110101111",
  15017=>"111100001",
  15018=>"110111011",
  15019=>"110110101",
  15020=>"111011000",
  15021=>"000101110",
  15022=>"110011010",
  15023=>"111010011",
  15024=>"110100110",
  15025=>"010000101",
  15026=>"001100001",
  15027=>"101100101",
  15028=>"010110100",
  15029=>"001000101",
  15030=>"101110100",
  15031=>"010101011",
  15032=>"011111010",
  15033=>"111101111",
  15034=>"010010110",
  15035=>"011101110",
  15036=>"100100110",
  15037=>"000001001",
  15038=>"000100110",
  15039=>"010101101",
  15040=>"110000000",
  15041=>"010111001",
  15042=>"111000101",
  15043=>"001011001",
  15044=>"111000010",
  15045=>"101100110",
  15046=>"011111111",
  15047=>"001101101",
  15048=>"001010111",
  15049=>"000101001",
  15050=>"011111111",
  15051=>"000000010",
  15052=>"000100001",
  15053=>"011111101",
  15054=>"000000011",
  15055=>"100000001",
  15056=>"111111010",
  15057=>"000100000",
  15058=>"011111010",
  15059=>"001010010",
  15060=>"001000110",
  15061=>"000000001",
  15062=>"000010010",
  15063=>"011100110",
  15064=>"100011111",
  15065=>"000100011",
  15066=>"110010010",
  15067=>"011110110",
  15068=>"011011110",
  15069=>"001001101",
  15070=>"010111000",
  15071=>"101100110",
  15072=>"110100110",
  15073=>"110000111",
  15074=>"000010011",
  15075=>"011100100",
  15076=>"101011101",
  15077=>"110101111",
  15078=>"011000110",
  15079=>"001011011",
  15080=>"001001100",
  15081=>"101000100",
  15082=>"000011010",
  15083=>"100000001",
  15084=>"010001010",
  15085=>"111110101",
  15086=>"000010100",
  15087=>"100010001",
  15088=>"100011101",
  15089=>"101011101",
  15090=>"011111000",
  15091=>"001000001",
  15092=>"011010100",
  15093=>"100101110",
  15094=>"110110100",
  15095=>"011101111",
  15096=>"001011001",
  15097=>"110111001",
  15098=>"111100011",
  15099=>"110010110",
  15100=>"111000001",
  15101=>"001011111",
  15102=>"001000000",
  15103=>"000000101",
  15104=>"010101100",
  15105=>"100100011",
  15106=>"101011101",
  15107=>"110111110",
  15108=>"010110100",
  15109=>"010110110",
  15110=>"100000010",
  15111=>"000001000",
  15112=>"101100000",
  15113=>"000111101",
  15114=>"100100001",
  15115=>"110010111",
  15116=>"011100111",
  15117=>"101000010",
  15118=>"110111111",
  15119=>"000111111",
  15120=>"110101001",
  15121=>"100000010",
  15122=>"010110011",
  15123=>"001010100",
  15124=>"010100011",
  15125=>"101001100",
  15126=>"111111011",
  15127=>"001000001",
  15128=>"100100010",
  15129=>"000000001",
  15130=>"000001010",
  15131=>"110111011",
  15132=>"000000100",
  15133=>"110000111",
  15134=>"110110001",
  15135=>"101111110",
  15136=>"100100100",
  15137=>"010110000",
  15138=>"001010101",
  15139=>"001111111",
  15140=>"110011111",
  15141=>"001101001",
  15142=>"100010011",
  15143=>"110000110",
  15144=>"000011111",
  15145=>"101111110",
  15146=>"100101010",
  15147=>"100100010",
  15148=>"111111001",
  15149=>"110011100",
  15150=>"001101100",
  15151=>"000101010",
  15152=>"111110011",
  15153=>"000011101",
  15154=>"101010000",
  15155=>"101101010",
  15156=>"011010101",
  15157=>"110111111",
  15158=>"111011011",
  15159=>"110110110",
  15160=>"000100011",
  15161=>"111101110",
  15162=>"111100000",
  15163=>"010110011",
  15164=>"100011100",
  15165=>"001010101",
  15166=>"001110100",
  15167=>"110000111",
  15168=>"001110001",
  15169=>"101000000",
  15170=>"101111111",
  15171=>"000101111",
  15172=>"101000000",
  15173=>"010101000",
  15174=>"100100100",
  15175=>"101111101",
  15176=>"100010000",
  15177=>"111111001",
  15178=>"100111000",
  15179=>"110111101",
  15180=>"000101011",
  15181=>"101011110",
  15182=>"010000100",
  15183=>"000001010",
  15184=>"011001000",
  15185=>"000011100",
  15186=>"001111010",
  15187=>"111101110",
  15188=>"000100100",
  15189=>"100011110",
  15190=>"110110100",
  15191=>"001101001",
  15192=>"000000100",
  15193=>"001000111",
  15194=>"110110111",
  15195=>"010011101",
  15196=>"110111101",
  15197=>"110100111",
  15198=>"111011101",
  15199=>"010010011",
  15200=>"100001110",
  15201=>"110111110",
  15202=>"100010011",
  15203=>"011011001",
  15204=>"011110010",
  15205=>"000011100",
  15206=>"101101000",
  15207=>"011101111",
  15208=>"100000010",
  15209=>"100101111",
  15210=>"000100100",
  15211=>"010111111",
  15212=>"001011111",
  15213=>"111001110",
  15214=>"100010100",
  15215=>"010000110",
  15216=>"000001011",
  15217=>"000010100",
  15218=>"001001011",
  15219=>"001110110",
  15220=>"000000100",
  15221=>"001011010",
  15222=>"111100011",
  15223=>"010010101",
  15224=>"110111100",
  15225=>"001100101",
  15226=>"100011101",
  15227=>"010000001",
  15228=>"010001001",
  15229=>"101010101",
  15230=>"001001110",
  15231=>"100100011",
  15232=>"110101110",
  15233=>"111111110",
  15234=>"101000100",
  15235=>"100110000",
  15236=>"110010110",
  15237=>"011110111",
  15238=>"100001010",
  15239=>"101111111",
  15240=>"010011011",
  15241=>"000010101",
  15242=>"000011110",
  15243=>"101000000",
  15244=>"010100011",
  15245=>"011110000",
  15246=>"010100111",
  15247=>"100010100",
  15248=>"101101101",
  15249=>"001010101",
  15250=>"010110000",
  15251=>"011010001",
  15252=>"011110111",
  15253=>"100100001",
  15254=>"001010000",
  15255=>"001011011",
  15256=>"010010111",
  15257=>"000011100",
  15258=>"000011111",
  15259=>"101001011",
  15260=>"111110000",
  15261=>"000100010",
  15262=>"110010111",
  15263=>"001000000",
  15264=>"010101110",
  15265=>"011111110",
  15266=>"011011110",
  15267=>"001000101",
  15268=>"100110111",
  15269=>"001111010",
  15270=>"000000011",
  15271=>"110000100",
  15272=>"000011001",
  15273=>"110011000",
  15274=>"100100011",
  15275=>"110110010",
  15276=>"110100110",
  15277=>"100100000",
  15278=>"000010000",
  15279=>"011101110",
  15280=>"011000000",
  15281=>"110001010",
  15282=>"101100111",
  15283=>"011010001",
  15284=>"010101100",
  15285=>"010100101",
  15286=>"001000100",
  15287=>"000010000",
  15288=>"010011110",
  15289=>"111011000",
  15290=>"100111010",
  15291=>"011100100",
  15292=>"100111101",
  15293=>"101010000",
  15294=>"110000101",
  15295=>"101110111",
  15296=>"001001100",
  15297=>"100101110",
  15298=>"100011101",
  15299=>"110100000",
  15300=>"001000010",
  15301=>"000100100",
  15302=>"000111101",
  15303=>"010111000",
  15304=>"011100110",
  15305=>"011001011",
  15306=>"010010101",
  15307=>"100110100",
  15308=>"010101110",
  15309=>"111000110",
  15310=>"111101111",
  15311=>"101011011",
  15312=>"000011000",
  15313=>"011101001",
  15314=>"011110111",
  15315=>"010110000",
  15316=>"000110011",
  15317=>"110100001",
  15318=>"110001101",
  15319=>"001000101",
  15320=>"100100111",
  15321=>"101001000",
  15322=>"110011000",
  15323=>"000101000",
  15324=>"110111111",
  15325=>"101110000",
  15326=>"000011100",
  15327=>"110100101",
  15328=>"001110110",
  15329=>"100101111",
  15330=>"001110011",
  15331=>"001001011",
  15332=>"111101101",
  15333=>"000111101",
  15334=>"000111100",
  15335=>"100000001",
  15336=>"111111010",
  15337=>"000111011",
  15338=>"011000010",
  15339=>"111001001",
  15340=>"011110110",
  15341=>"101011111",
  15342=>"101110000",
  15343=>"110000010",
  15344=>"010001011",
  15345=>"100110000",
  15346=>"101101011",
  15347=>"111001101",
  15348=>"001101011",
  15349=>"000110101",
  15350=>"010101011",
  15351=>"000011000",
  15352=>"000110110",
  15353=>"000100000",
  15354=>"010000001",
  15355=>"010111110",
  15356=>"001010010",
  15357=>"011001000",
  15358=>"100010100",
  15359=>"011010000",
  15360=>"010100101",
  15361=>"010001001",
  15362=>"111001111",
  15363=>"001100000",
  15364=>"010111010",
  15365=>"100010100",
  15366=>"010000100",
  15367=>"101110000",
  15368=>"010000110",
  15369=>"110000001",
  15370=>"001110010",
  15371=>"111010001",
  15372=>"110111010",
  15373=>"100000000",
  15374=>"111101001",
  15375=>"110001001",
  15376=>"000001101",
  15377=>"010001010",
  15378=>"001111101",
  15379=>"110011001",
  15380=>"100111110",
  15381=>"001110011",
  15382=>"010111101",
  15383=>"101110101",
  15384=>"111111111",
  15385=>"100101110",
  15386=>"010110110",
  15387=>"110001111",
  15388=>"110011111",
  15389=>"011111001",
  15390=>"101101101",
  15391=>"100000101",
  15392=>"001100001",
  15393=>"100111101",
  15394=>"001110110",
  15395=>"011110000",
  15396=>"101011111",
  15397=>"001100111",
  15398=>"011100111",
  15399=>"100011101",
  15400=>"110000001",
  15401=>"000010100",
  15402=>"010010010",
  15403=>"110000000",
  15404=>"101001100",
  15405=>"001110110",
  15406=>"011010001",
  15407=>"111000111",
  15408=>"100011111",
  15409=>"010010011",
  15410=>"001110111",
  15411=>"110000011",
  15412=>"101000111",
  15413=>"110001001",
  15414=>"111000001",
  15415=>"010100011",
  15416=>"111001101",
  15417=>"100011010",
  15418=>"100001100",
  15419=>"010001100",
  15420=>"000001111",
  15421=>"111011000",
  15422=>"111010000",
  15423=>"010000010",
  15424=>"010000101",
  15425=>"001111001",
  15426=>"101111000",
  15427=>"000100000",
  15428=>"111001001",
  15429=>"110101100",
  15430=>"011000011",
  15431=>"100001101",
  15432=>"011100001",
  15433=>"001011001",
  15434=>"010010001",
  15435=>"010101100",
  15436=>"000001011",
  15437=>"111001101",
  15438=>"011011010",
  15439=>"110110001",
  15440=>"101011001",
  15441=>"110101101",
  15442=>"010001001",
  15443=>"101101011",
  15444=>"101101000",
  15445=>"110001101",
  15446=>"010010100",
  15447=>"101100000",
  15448=>"001101011",
  15449=>"100111110",
  15450=>"110001010",
  15451=>"000001010",
  15452=>"011010001",
  15453=>"001000101",
  15454=>"101110000",
  15455=>"011001001",
  15456=>"110011011",
  15457=>"010001100",
  15458=>"111011001",
  15459=>"000101000",
  15460=>"100110000",
  15461=>"011110100",
  15462=>"001000100",
  15463=>"011000100",
  15464=>"110000010",
  15465=>"110000101",
  15466=>"011100001",
  15467=>"100101001",
  15468=>"011000000",
  15469=>"101101011",
  15470=>"100111011",
  15471=>"110111100",
  15472=>"010101100",
  15473=>"001000100",
  15474=>"111001100",
  15475=>"011110111",
  15476=>"101010001",
  15477=>"110101110",
  15478=>"010110100",
  15479=>"101111101",
  15480=>"111111010",
  15481=>"011010110",
  15482=>"101110011",
  15483=>"000101001",
  15484=>"100111110",
  15485=>"010100000",
  15486=>"111110111",
  15487=>"110010011",
  15488=>"001110101",
  15489=>"101011010",
  15490=>"001010011",
  15491=>"000101111",
  15492=>"100100001",
  15493=>"101101001",
  15494=>"100101001",
  15495=>"110100110",
  15496=>"101111110",
  15497=>"000000011",
  15498=>"001110001",
  15499=>"001101111",
  15500=>"000011111",
  15501=>"000100101",
  15502=>"001110110",
  15503=>"000101011",
  15504=>"110111111",
  15505=>"001110111",
  15506=>"000000111",
  15507=>"011100011",
  15508=>"111000011",
  15509=>"010011000",
  15510=>"101000001",
  15511=>"011010010",
  15512=>"001010110",
  15513=>"100110100",
  15514=>"001011000",
  15515=>"100010011",
  15516=>"110101010",
  15517=>"111110100",
  15518=>"100111010",
  15519=>"110001101",
  15520=>"001100100",
  15521=>"111001001",
  15522=>"011010100",
  15523=>"010101001",
  15524=>"111011111",
  15525=>"100111010",
  15526=>"000000011",
  15527=>"001101001",
  15528=>"100111000",
  15529=>"101000010",
  15530=>"100001011",
  15531=>"100111110",
  15532=>"010011010",
  15533=>"001101110",
  15534=>"011000000",
  15535=>"001101111",
  15536=>"010011011",
  15537=>"000010010",
  15538=>"000011010",
  15539=>"111000110",
  15540=>"011010001",
  15541=>"001101100",
  15542=>"000101011",
  15543=>"111101101",
  15544=>"101101000",
  15545=>"110001000",
  15546=>"100101011",
  15547=>"111000111",
  15548=>"011011010",
  15549=>"000011111",
  15550=>"001100100",
  15551=>"100010000",
  15552=>"101100010",
  15553=>"101000100",
  15554=>"110011001",
  15555=>"101100101",
  15556=>"101011100",
  15557=>"001000100",
  15558=>"111010010",
  15559=>"100100111",
  15560=>"001100010",
  15561=>"100000110",
  15562=>"111011111",
  15563=>"011001100",
  15564=>"010011110",
  15565=>"111011111",
  15566=>"000010110",
  15567=>"111010011",
  15568=>"001000000",
  15569=>"100111100",
  15570=>"010001111",
  15571=>"000100100",
  15572=>"011010100",
  15573=>"010110111",
  15574=>"110011110",
  15575=>"001010000",
  15576=>"110100010",
  15577=>"011100010",
  15578=>"011010100",
  15579=>"000000001",
  15580=>"001010001",
  15581=>"001100100",
  15582=>"000000111",
  15583=>"110010100",
  15584=>"000011101",
  15585=>"010100000",
  15586=>"111011000",
  15587=>"100100010",
  15588=>"011110011",
  15589=>"110110101",
  15590=>"000000001",
  15591=>"111111011",
  15592=>"100010001",
  15593=>"110001111",
  15594=>"010000000",
  15595=>"100110001",
  15596=>"000000000",
  15597=>"100110001",
  15598=>"001100011",
  15599=>"100100010",
  15600=>"001111010",
  15601=>"011001011",
  15602=>"111001100",
  15603=>"100100000",
  15604=>"001001000",
  15605=>"110111111",
  15606=>"101011010",
  15607=>"000100110",
  15608=>"111111100",
  15609=>"000001100",
  15610=>"110000110",
  15611=>"100011100",
  15612=>"101000010",
  15613=>"011000100",
  15614=>"001100111",
  15615=>"000101100",
  15616=>"011100011",
  15617=>"100011001",
  15618=>"011000000",
  15619=>"101101001",
  15620=>"110001110",
  15621=>"111100001",
  15622=>"001000010",
  15623=>"100000011",
  15624=>"010001010",
  15625=>"000000011",
  15626=>"010111011",
  15627=>"011100100",
  15628=>"100110101",
  15629=>"000100010",
  15630=>"011001111",
  15631=>"000000000",
  15632=>"100111010",
  15633=>"100100100",
  15634=>"011100011",
  15635=>"100010101",
  15636=>"110111001",
  15637=>"011011110",
  15638=>"011011011",
  15639=>"010001100",
  15640=>"000100111",
  15641=>"011011000",
  15642=>"100011110",
  15643=>"011111010",
  15644=>"000011001",
  15645=>"101100001",
  15646=>"111000111",
  15647=>"111000010",
  15648=>"011001001",
  15649=>"000101000",
  15650=>"111111011",
  15651=>"000100000",
  15652=>"001011010",
  15653=>"000010101",
  15654=>"111111000",
  15655=>"011110011",
  15656=>"001001101",
  15657=>"100110010",
  15658=>"011010100",
  15659=>"010100000",
  15660=>"011110100",
  15661=>"111010010",
  15662=>"011111111",
  15663=>"010111111",
  15664=>"101110000",
  15665=>"100011011",
  15666=>"110110100",
  15667=>"110101111",
  15668=>"101000001",
  15669=>"100111101",
  15670=>"101111100",
  15671=>"010010010",
  15672=>"011010100",
  15673=>"100010010",
  15674=>"101111100",
  15675=>"001111111",
  15676=>"000010110",
  15677=>"111110110",
  15678=>"000110111",
  15679=>"001011000",
  15680=>"100101100",
  15681=>"111000011",
  15682=>"110111000",
  15683=>"001011000",
  15684=>"000110001",
  15685=>"001110010",
  15686=>"110011100",
  15687=>"000110000",
  15688=>"000011100",
  15689=>"010000101",
  15690=>"000001011",
  15691=>"000101110",
  15692=>"010011000",
  15693=>"011000000",
  15694=>"000010001",
  15695=>"101010110",
  15696=>"100100100",
  15697=>"011101101",
  15698=>"000101111",
  15699=>"011111011",
  15700=>"011110001",
  15701=>"011011011",
  15702=>"011110010",
  15703=>"100111010",
  15704=>"110000000",
  15705=>"000110100",
  15706=>"110010011",
  15707=>"111010100",
  15708=>"111011110",
  15709=>"100100001",
  15710=>"100001101",
  15711=>"001111110",
  15712=>"100100010",
  15713=>"101011011",
  15714=>"000100110",
  15715=>"001100110",
  15716=>"010100001",
  15717=>"111110111",
  15718=>"000001000",
  15719=>"111111111",
  15720=>"111101000",
  15721=>"110000100",
  15722=>"100110101",
  15723=>"010111110",
  15724=>"000010101",
  15725=>"011000001",
  15726=>"111111011",
  15727=>"100010110",
  15728=>"011111101",
  15729=>"110110000",
  15730=>"001000001",
  15731=>"101000100",
  15732=>"010000000",
  15733=>"110100101",
  15734=>"110100111",
  15735=>"101011110",
  15736=>"100111110",
  15737=>"000001010",
  15738=>"111100101",
  15739=>"001001100",
  15740=>"110101101",
  15741=>"100101111",
  15742=>"010111000",
  15743=>"100110110",
  15744=>"010101001",
  15745=>"001000101",
  15746=>"100000010",
  15747=>"001000101",
  15748=>"010001001",
  15749=>"000000000",
  15750=>"100111101",
  15751=>"010000110",
  15752=>"000001000",
  15753=>"011001000",
  15754=>"001001111",
  15755=>"001010110",
  15756=>"110000100",
  15757=>"100000110",
  15758=>"010011100",
  15759=>"001101000",
  15760=>"001011000",
  15761=>"000111001",
  15762=>"101100100",
  15763=>"100110010",
  15764=>"000101100",
  15765=>"110000001",
  15766=>"001010110",
  15767=>"100000011",
  15768=>"110001010",
  15769=>"110101111",
  15770=>"100000001",
  15771=>"111000010",
  15772=>"100100011",
  15773=>"101010110",
  15774=>"110001100",
  15775=>"101000111",
  15776=>"110011010",
  15777=>"001001101",
  15778=>"000010000",
  15779=>"010110110",
  15780=>"111100100",
  15781=>"001011101",
  15782=>"011101000",
  15783=>"100110110",
  15784=>"111000011",
  15785=>"101111010",
  15786=>"100010110",
  15787=>"101100100",
  15788=>"110001010",
  15789=>"001001101",
  15790=>"110110111",
  15791=>"000101110",
  15792=>"000100010",
  15793=>"001111110",
  15794=>"011110110",
  15795=>"000110001",
  15796=>"010100110",
  15797=>"010111101",
  15798=>"100111111",
  15799=>"010001111",
  15800=>"011000010",
  15801=>"000001001",
  15802=>"010110110",
  15803=>"100010000",
  15804=>"011001100",
  15805=>"110110011",
  15806=>"100001110",
  15807=>"111100111",
  15808=>"011001000",
  15809=>"000101100",
  15810=>"101011111",
  15811=>"000101000",
  15812=>"111110011",
  15813=>"010001110",
  15814=>"001000001",
  15815=>"010111010",
  15816=>"001001001",
  15817=>"110101000",
  15818=>"110111101",
  15819=>"001111011",
  15820=>"011111000",
  15821=>"110100101",
  15822=>"110110011",
  15823=>"000000001",
  15824=>"000011110",
  15825=>"100100100",
  15826=>"011101000",
  15827=>"100001011",
  15828=>"000101010",
  15829=>"000000000",
  15830=>"010101101",
  15831=>"110000100",
  15832=>"110001110",
  15833=>"111110000",
  15834=>"101101011",
  15835=>"100100000",
  15836=>"011010010",
  15837=>"110011111",
  15838=>"110011101",
  15839=>"110110100",
  15840=>"001001100",
  15841=>"011001100",
  15842=>"011010110",
  15843=>"100101101",
  15844=>"001111110",
  15845=>"001111100",
  15846=>"111110010",
  15847=>"111010100",
  15848=>"001110000",
  15849=>"011010010",
  15850=>"011100100",
  15851=>"100101011",
  15852=>"111111110",
  15853=>"101010111",
  15854=>"001000010",
  15855=>"100001010",
  15856=>"110111110",
  15857=>"011100010",
  15858=>"100010001",
  15859=>"011000100",
  15860=>"000101011",
  15861=>"110111111",
  15862=>"011000111",
  15863=>"110110110",
  15864=>"011001110",
  15865=>"011111110",
  15866=>"111100010",
  15867=>"011101101",
  15868=>"111110100",
  15869=>"100101010",
  15870=>"110001111",
  15871=>"000010010",
  15872=>"111111101",
  15873=>"111001000",
  15874=>"101010110",
  15875=>"100111110",
  15876=>"010001100",
  15877=>"001000111",
  15878=>"111011111",
  15879=>"111100101",
  15880=>"100010000",
  15881=>"010011100",
  15882=>"111101010",
  15883=>"010011010",
  15884=>"011001001",
  15885=>"101011010",
  15886=>"011001110",
  15887=>"000100000",
  15888=>"000100010",
  15889=>"011010001",
  15890=>"111001011",
  15891=>"000001111",
  15892=>"010000000",
  15893=>"100110010",
  15894=>"001000010",
  15895=>"111111001",
  15896=>"101111001",
  15897=>"111101100",
  15898=>"101100110",
  15899=>"011111001",
  15900=>"010000100",
  15901=>"110111101",
  15902=>"010100010",
  15903=>"100010010",
  15904=>"110000001",
  15905=>"010100000",
  15906=>"110100010",
  15907=>"000101010",
  15908=>"100001111",
  15909=>"100000011",
  15910=>"001110110",
  15911=>"000011110",
  15912=>"011000110",
  15913=>"110101010",
  15914=>"101111000",
  15915=>"010000001",
  15916=>"000111111",
  15917=>"010011010",
  15918=>"111101111",
  15919=>"101000000",
  15920=>"101101010",
  15921=>"111011100",
  15922=>"011101100",
  15923=>"111101000",
  15924=>"001011010",
  15925=>"110110110",
  15926=>"000101000",
  15927=>"000010111",
  15928=>"011010110",
  15929=>"011010111",
  15930=>"011000001",
  15931=>"011001011",
  15932=>"100011000",
  15933=>"001001010",
  15934=>"000100010",
  15935=>"001110111",
  15936=>"100101110",
  15937=>"110110101",
  15938=>"101000111",
  15939=>"011001000",
  15940=>"111000001",
  15941=>"100000000",
  15942=>"000010001",
  15943=>"101001000",
  15944=>"001010100",
  15945=>"010111010",
  15946=>"110011001",
  15947=>"100010110",
  15948=>"001100111",
  15949=>"011111011",
  15950=>"001110100",
  15951=>"000101001",
  15952=>"010011000",
  15953=>"010110100",
  15954=>"000010101",
  15955=>"001011100",
  15956=>"000110101",
  15957=>"100000000",
  15958=>"000111111",
  15959=>"111010101",
  15960=>"100100100",
  15961=>"011011010",
  15962=>"010111001",
  15963=>"000010001",
  15964=>"011101000",
  15965=>"010010110",
  15966=>"110000110",
  15967=>"011101111",
  15968=>"111011101",
  15969=>"100010101",
  15970=>"110000010",
  15971=>"101001011",
  15972=>"100100110",
  15973=>"100100100",
  15974=>"010010000",
  15975=>"100000111",
  15976=>"011001000",
  15977=>"100000010",
  15978=>"110011011",
  15979=>"110110001",
  15980=>"011010110",
  15981=>"001110111",
  15982=>"011111101",
  15983=>"001000110",
  15984=>"011000001",
  15985=>"101000000",
  15986=>"010101000",
  15987=>"101100100",
  15988=>"110110001",
  15989=>"011010100",
  15990=>"010001001",
  15991=>"100001110",
  15992=>"111001011",
  15993=>"110011100",
  15994=>"011011101",
  15995=>"001100011",
  15996=>"000011010",
  15997=>"011001000",
  15998=>"100111000",
  15999=>"110101110",
  16000=>"010111100",
  16001=>"101101010",
  16002=>"000010101",
  16003=>"010000111",
  16004=>"110110010",
  16005=>"110110100",
  16006=>"011010101",
  16007=>"101100100",
  16008=>"011100100",
  16009=>"010100000",
  16010=>"110011000",
  16011=>"001010101",
  16012=>"010001001",
  16013=>"110111111",
  16014=>"001100001",
  16015=>"101001011",
  16016=>"000001000",
  16017=>"010111101",
  16018=>"100110101",
  16019=>"000101011",
  16020=>"011101000",
  16021=>"101001011",
  16022=>"101000101",
  16023=>"100000010",
  16024=>"000010010",
  16025=>"101111101",
  16026=>"111011110",
  16027=>"010010001",
  16028=>"100000110",
  16029=>"000100010",
  16030=>"000000010",
  16031=>"001011101",
  16032=>"011011100",
  16033=>"111110111",
  16034=>"100000000",
  16035=>"010001101",
  16036=>"010111001",
  16037=>"010011001",
  16038=>"110100100",
  16039=>"110111100",
  16040=>"110000100",
  16041=>"000000110",
  16042=>"110010101",
  16043=>"011100010",
  16044=>"011011110",
  16045=>"001001100",
  16046=>"011100100",
  16047=>"001100011",
  16048=>"000011000",
  16049=>"110000011",
  16050=>"111111110",
  16051=>"110111010",
  16052=>"010010110",
  16053=>"110101001",
  16054=>"010111101",
  16055=>"010010101",
  16056=>"101101110",
  16057=>"101000010",
  16058=>"111011101",
  16059=>"110110110",
  16060=>"000100100",
  16061=>"010001001",
  16062=>"100000101",
  16063=>"110001011",
  16064=>"000100000",
  16065=>"011000000",
  16066=>"101111100",
  16067=>"100111111",
  16068=>"110001001",
  16069=>"100000110",
  16070=>"011100000",
  16071=>"010111000",
  16072=>"100110011",
  16073=>"010111001",
  16074=>"111111111",
  16075=>"111110011",
  16076=>"111000010",
  16077=>"001111110",
  16078=>"110010101",
  16079=>"100110100",
  16080=>"010110000",
  16081=>"001101100",
  16082=>"100101001",
  16083=>"111100111",
  16084=>"001001001",
  16085=>"100100001",
  16086=>"101001011",
  16087=>"110110001",
  16088=>"100110011",
  16089=>"111011000",
  16090=>"111101010",
  16091=>"011011011",
  16092=>"101001100",
  16093=>"100101000",
  16094=>"000110010",
  16095=>"111111001",
  16096=>"010101010",
  16097=>"000000011",
  16098=>"111011001",
  16099=>"010100011",
  16100=>"101101110",
  16101=>"000010101",
  16102=>"000011100",
  16103=>"010100111",
  16104=>"011111101",
  16105=>"001110001",
  16106=>"000001000",
  16107=>"011111011",
  16108=>"001100001",
  16109=>"010000010",
  16110=>"000001001",
  16111=>"111110111",
  16112=>"110000000",
  16113=>"110111001",
  16114=>"000001001",
  16115=>"011001101",
  16116=>"010100100",
  16117=>"010001101",
  16118=>"100110000",
  16119=>"111111001",
  16120=>"000010100",
  16121=>"011000111",
  16122=>"000011000",
  16123=>"011010001",
  16124=>"001001011",
  16125=>"011011011",
  16126=>"110011011",
  16127=>"000000011",
  16128=>"111100100",
  16129=>"111010010",
  16130=>"000110111",
  16131=>"101001011",
  16132=>"010101000",
  16133=>"010110100",
  16134=>"000110100",
  16135=>"010011001",
  16136=>"010101110",
  16137=>"111101101",
  16138=>"010001101",
  16139=>"010001011",
  16140=>"011001111",
  16141=>"110011001",
  16142=>"011101101",
  16143=>"111110101",
  16144=>"100110111",
  16145=>"000101101",
  16146=>"000001111",
  16147=>"011101010",
  16148=>"100111100",
  16149=>"001011101",
  16150=>"011110110",
  16151=>"101110001",
  16152=>"010100010",
  16153=>"000000100",
  16154=>"000010011",
  16155=>"110000111",
  16156=>"010001101",
  16157=>"000011100",
  16158=>"111101110",
  16159=>"001101011",
  16160=>"110110000",
  16161=>"010101101",
  16162=>"110111011",
  16163=>"011100000",
  16164=>"100110111",
  16165=>"101001111",
  16166=>"011010111",
  16167=>"011000111",
  16168=>"000111110",
  16169=>"001001000",
  16170=>"100101010",
  16171=>"111010110",
  16172=>"000111110",
  16173=>"100001010",
  16174=>"001001010",
  16175=>"100010011",
  16176=>"100111011",
  16177=>"001001110",
  16178=>"000000001",
  16179=>"110001100",
  16180=>"010010001",
  16181=>"100101100",
  16182=>"111100001",
  16183=>"000001001",
  16184=>"111110100",
  16185=>"111110100",
  16186=>"000001101",
  16187=>"010001010",
  16188=>"011101000",
  16189=>"011000000",
  16190=>"111000001",
  16191=>"001111111",
  16192=>"000111110",
  16193=>"101110100",
  16194=>"110111011",
  16195=>"100010010",
  16196=>"011000100",
  16197=>"110111111",
  16198=>"111000111",
  16199=>"001011001",
  16200=>"011011011",
  16201=>"000001110",
  16202=>"101100011",
  16203=>"111101000",
  16204=>"010100101",
  16205=>"110111100",
  16206=>"101101111",
  16207=>"010111110",
  16208=>"010100011",
  16209=>"110011000",
  16210=>"100001100",
  16211=>"000000111",
  16212=>"001111000",
  16213=>"001011000",
  16214=>"010101111",
  16215=>"011011111",
  16216=>"011011101",
  16217=>"111111000",
  16218=>"111111010",
  16219=>"000110100",
  16220=>"000010010",
  16221=>"100001000",
  16222=>"001100010",
  16223=>"100001111",
  16224=>"010011011",
  16225=>"110100011",
  16226=>"100100001",
  16227=>"111010110",
  16228=>"111011101",
  16229=>"111001011",
  16230=>"101110000",
  16231=>"101111000",
  16232=>"010000100",
  16233=>"111001101",
  16234=>"010000000",
  16235=>"110111101",
  16236=>"111110110",
  16237=>"011000011",
  16238=>"111111101",
  16239=>"111011110",
  16240=>"000110010",
  16241=>"110011001",
  16242=>"100110000",
  16243=>"110010001",
  16244=>"010000010",
  16245=>"010111100",
  16246=>"110010110",
  16247=>"101111010",
  16248=>"001001101",
  16249=>"000001111",
  16250=>"000101111",
  16251=>"001101011",
  16252=>"000100000",
  16253=>"011110000",
  16254=>"011100010",
  16255=>"110101101",
  16256=>"001101100",
  16257=>"101111101",
  16258=>"100000100",
  16259=>"001011100",
  16260=>"001110111",
  16261=>"101000110",
  16262=>"100011011",
  16263=>"011101011",
  16264=>"001100111",
  16265=>"010010100",
  16266=>"101001111",
  16267=>"111100010",
  16268=>"011110000",
  16269=>"110101101",
  16270=>"001001001",
  16271=>"011111010",
  16272=>"101110001",
  16273=>"110001010",
  16274=>"000110110",
  16275=>"011100001",
  16276=>"000111000",
  16277=>"110111011",
  16278=>"100011000",
  16279=>"001110100",
  16280=>"110100101",
  16281=>"101010011",
  16282=>"010101010",
  16283=>"111111000",
  16284=>"000010010",
  16285=>"000000000",
  16286=>"010001010",
  16287=>"001011001",
  16288=>"100100001",
  16289=>"011010000",
  16290=>"010111010",
  16291=>"000110010",
  16292=>"111010100",
  16293=>"101001100",
  16294=>"010000000",
  16295=>"111101100",
  16296=>"000001000",
  16297=>"100100110",
  16298=>"011110100",
  16299=>"000010110",
  16300=>"101001110",
  16301=>"000110011",
  16302=>"100100111",
  16303=>"011110010",
  16304=>"011000110",
  16305=>"111111100",
  16306=>"101101111",
  16307=>"101000101",
  16308=>"011011101",
  16309=>"110110101",
  16310=>"101001101",
  16311=>"001101011",
  16312=>"001011000",
  16313=>"101011111",
  16314=>"000100110",
  16315=>"101101101",
  16316=>"010000001",
  16317=>"100101101",
  16318=>"001011110",
  16319=>"100000010",
  16320=>"011011010",
  16321=>"110100010",
  16322=>"111101010",
  16323=>"000101100",
  16324=>"110011111",
  16325=>"001110001",
  16326=>"011101101",
  16327=>"000010100",
  16328=>"011001100",
  16329=>"011100011",
  16330=>"100000101",
  16331=>"010011111",
  16332=>"100000000",
  16333=>"100100101",
  16334=>"101101100",
  16335=>"100001110",
  16336=>"100001011",
  16337=>"001010000",
  16338=>"101010000",
  16339=>"011011111",
  16340=>"101010101",
  16341=>"000110000",
  16342=>"000110111",
  16343=>"011001001",
  16344=>"111101111",
  16345=>"001000101",
  16346=>"110100110",
  16347=>"111000101",
  16348=>"100000011",
  16349=>"010011101",
  16350=>"001110111",
  16351=>"100010101",
  16352=>"001000010",
  16353=>"110111000",
  16354=>"000000000",
  16355=>"000010110",
  16356=>"000000110",
  16357=>"111101101",
  16358=>"100011110",
  16359=>"110110100",
  16360=>"000011001",
  16361=>"010100011",
  16362=>"101000000",
  16363=>"111001101",
  16364=>"000001010",
  16365=>"001011000",
  16366=>"010110000",
  16367=>"011001001",
  16368=>"011001011",
  16369=>"010001111",
  16370=>"000011011",
  16371=>"010001110",
  16372=>"111110111",
  16373=>"000011000",
  16374=>"100010110",
  16375=>"011001010",
  16376=>"110000111",
  16377=>"101000001",
  16378=>"010011001",
  16379=>"111010100",
  16380=>"110111110",
  16381=>"011010000",
  16382=>"011100010",
  16383=>"100100101",
  16384=>"100111001",
  16385=>"110110011",
  16386=>"101111110",
  16387=>"001111100",
  16388=>"100110010",
  16389=>"101010100",
  16390=>"101000111",
  16391=>"010011111",
  16392=>"000010000",
  16393=>"111011010",
  16394=>"000010000",
  16395=>"011100001",
  16396=>"101011101",
  16397=>"111110001",
  16398=>"010010110",
  16399=>"010111111",
  16400=>"101000100",
  16401=>"101100100",
  16402=>"100101000",
  16403=>"000100001",
  16404=>"101101000",
  16405=>"110011010",
  16406=>"111011011",
  16407=>"110001001",
  16408=>"011101000",
  16409=>"110011111",
  16410=>"111111101",
  16411=>"010001010",
  16412=>"111010001",
  16413=>"000010100",
  16414=>"000000000",
  16415=>"000110110",
  16416=>"001001001",
  16417=>"101000100",
  16418=>"010110001",
  16419=>"111010111",
  16420=>"001000000",
  16421=>"101100100",
  16422=>"101111100",
  16423=>"111010011",
  16424=>"010000010",
  16425=>"001101011",
  16426=>"001001000",
  16427=>"110010000",
  16428=>"000010101",
  16429=>"110011001",
  16430=>"000101100",
  16431=>"111001001",
  16432=>"111001100",
  16433=>"111110010",
  16434=>"100000010",
  16435=>"110111001",
  16436=>"111110100",
  16437=>"101110011",
  16438=>"010011101",
  16439=>"001001100",
  16440=>"011000100",
  16441=>"010110100",
  16442=>"010001111",
  16443=>"111111011",
  16444=>"111011111",
  16445=>"101111010",
  16446=>"011101110",
  16447=>"000111111",
  16448=>"001101110",
  16449=>"011110110",
  16450=>"010110111",
  16451=>"001010100",
  16452=>"101011111",
  16453=>"001010000",
  16454=>"101110111",
  16455=>"110101100",
  16456=>"111010000",
  16457=>"110111000",
  16458=>"110011101",
  16459=>"000110100",
  16460=>"110000111",
  16461=>"000010101",
  16462=>"110110101",
  16463=>"110011111",
  16464=>"100111000",
  16465=>"000110100",
  16466=>"000100101",
  16467=>"001000101",
  16468=>"101001101",
  16469=>"101100000",
  16470=>"100111001",
  16471=>"010000111",
  16472=>"100101100",
  16473=>"111111111",
  16474=>"001011010",
  16475=>"100000100",
  16476=>"111101011",
  16477=>"011010001",
  16478=>"110001110",
  16479=>"100111110",
  16480=>"111110010",
  16481=>"110011100",
  16482=>"001110000",
  16483=>"011010101",
  16484=>"011001111",
  16485=>"101000000",
  16486=>"101000100",
  16487=>"111111001",
  16488=>"101001100",
  16489=>"000110010",
  16490=>"011000111",
  16491=>"100010110",
  16492=>"111001110",
  16493=>"000001010",
  16494=>"000010000",
  16495=>"100011000",
  16496=>"000100101",
  16497=>"100011011",
  16498=>"000110111",
  16499=>"100011110",
  16500=>"011100010",
  16501=>"100110110",
  16502=>"010101000",
  16503=>"100001010",
  16504=>"001111101",
  16505=>"000011000",
  16506=>"110001110",
  16507=>"110100101",
  16508=>"001101010",
  16509=>"110110101",
  16510=>"100110000",
  16511=>"010000011",
  16512=>"001000100",
  16513=>"011100001",
  16514=>"010100010",
  16515=>"100110010",
  16516=>"110000000",
  16517=>"000110001",
  16518=>"000001111",
  16519=>"100001101",
  16520=>"110110000",
  16521=>"110110000",
  16522=>"010111011",
  16523=>"010101100",
  16524=>"011010000",
  16525=>"110000111",
  16526=>"001000111",
  16527=>"111100100",
  16528=>"111010010",
  16529=>"111011111",
  16530=>"001111011",
  16531=>"001101110",
  16532=>"100011100",
  16533=>"000000110",
  16534=>"111010101",
  16535=>"011111110",
  16536=>"011101101",
  16537=>"100010010",
  16538=>"001011010",
  16539=>"100011001",
  16540=>"110110010",
  16541=>"011000010",
  16542=>"111110011",
  16543=>"101111001",
  16544=>"000100011",
  16545=>"111110110",
  16546=>"011010011",
  16547=>"010101001",
  16548=>"011111000",
  16549=>"110001111",
  16550=>"101001110",
  16551=>"110001001",
  16552=>"110001000",
  16553=>"000100011",
  16554=>"100100010",
  16555=>"111000000",
  16556=>"100110000",
  16557=>"010111001",
  16558=>"100000111",
  16559=>"101010010",
  16560=>"011000001",
  16561=>"110001100",
  16562=>"101010100",
  16563=>"110000100",
  16564=>"000100010",
  16565=>"111011001",
  16566=>"111110111",
  16567=>"001000000",
  16568=>"000001100",
  16569=>"100111110",
  16570=>"111011100",
  16571=>"000111111",
  16572=>"010111101",
  16573=>"011110100",
  16574=>"100100010",
  16575=>"100101011",
  16576=>"011001111",
  16577=>"001010010",
  16578=>"101100111",
  16579=>"100101100",
  16580=>"011100100",
  16581=>"101000000",
  16582=>"000110100",
  16583=>"110010010",
  16584=>"011110110",
  16585=>"101101110",
  16586=>"111011011",
  16587=>"000100010",
  16588=>"100010000",
  16589=>"110010011",
  16590=>"001001100",
  16591=>"000000000",
  16592=>"010110010",
  16593=>"001111010",
  16594=>"000111110",
  16595=>"000101100",
  16596=>"000000100",
  16597=>"111001010",
  16598=>"011001110",
  16599=>"111011100",
  16600=>"100110110",
  16601=>"111110101",
  16602=>"110111010",
  16603=>"101011111",
  16604=>"111000011",
  16605=>"001001010",
  16606=>"001101001",
  16607=>"010110001",
  16608=>"001010010",
  16609=>"100000110",
  16610=>"100100011",
  16611=>"100111110",
  16612=>"010110110",
  16613=>"111011101",
  16614=>"111101001",
  16615=>"110100001",
  16616=>"001001000",
  16617=>"101100111",
  16618=>"101011111",
  16619=>"111111101",
  16620=>"001100001",
  16621=>"111011110",
  16622=>"100011001",
  16623=>"101100010",
  16624=>"100010111",
  16625=>"010111101",
  16626=>"110000100",
  16627=>"110001110",
  16628=>"110100011",
  16629=>"100010010",
  16630=>"011110011",
  16631=>"011100111",
  16632=>"110101110",
  16633=>"000000001",
  16634=>"011010101",
  16635=>"001100011",
  16636=>"111001110",
  16637=>"110000001",
  16638=>"000010111",
  16639=>"111110011",
  16640=>"110100010",
  16641=>"010001101",
  16642=>"010101111",
  16643=>"100011110",
  16644=>"011101011",
  16645=>"100111010",
  16646=>"010010000",
  16647=>"011001000",
  16648=>"101100010",
  16649=>"011110110",
  16650=>"010111010",
  16651=>"110011101",
  16652=>"011011101",
  16653=>"010001111",
  16654=>"010010011",
  16655=>"010100111",
  16656=>"001111011",
  16657=>"000000111",
  16658=>"010110011",
  16659=>"100011110",
  16660=>"111010000",
  16661=>"101101001",
  16662=>"011001001",
  16663=>"010100011",
  16664=>"100011011",
  16665=>"110101001",
  16666=>"001111100",
  16667=>"111110010",
  16668=>"010010000",
  16669=>"010001000",
  16670=>"001011100",
  16671=>"101101000",
  16672=>"101100110",
  16673=>"001101100",
  16674=>"001100100",
  16675=>"011101100",
  16676=>"111011110",
  16677=>"001011010",
  16678=>"000111010",
  16679=>"101000001",
  16680=>"011111101",
  16681=>"100111000",
  16682=>"010000110",
  16683=>"111111001",
  16684=>"001100101",
  16685=>"000001100",
  16686=>"000110010",
  16687=>"001000000",
  16688=>"010001100",
  16689=>"100100101",
  16690=>"010101110",
  16691=>"110010101",
  16692=>"111001100",
  16693=>"010110111",
  16694=>"000001011",
  16695=>"001111010",
  16696=>"110011111",
  16697=>"000101000",
  16698=>"101000001",
  16699=>"001001101",
  16700=>"000100111",
  16701=>"101010101",
  16702=>"111110100",
  16703=>"011111011",
  16704=>"101001100",
  16705=>"111111000",
  16706=>"000100000",
  16707=>"101010010",
  16708=>"110000001",
  16709=>"110000011",
  16710=>"001000011",
  16711=>"011110101",
  16712=>"001100010",
  16713=>"010010100",
  16714=>"110101000",
  16715=>"001000000",
  16716=>"101010010",
  16717=>"011110110",
  16718=>"101010101",
  16719=>"010001101",
  16720=>"001000100",
  16721=>"001011011",
  16722=>"110111001",
  16723=>"110000100",
  16724=>"001011001",
  16725=>"001000000",
  16726=>"111010010",
  16727=>"111000010",
  16728=>"100000001",
  16729=>"111110000",
  16730=>"010110010",
  16731=>"111111000",
  16732=>"110101011",
  16733=>"000101111",
  16734=>"100000000",
  16735=>"000110010",
  16736=>"110110111",
  16737=>"100001111",
  16738=>"111010100",
  16739=>"101100000",
  16740=>"101000010",
  16741=>"000100101",
  16742=>"110101100",
  16743=>"110101101",
  16744=>"110010111",
  16745=>"101000100",
  16746=>"111100100",
  16747=>"000110101",
  16748=>"010101111",
  16749=>"111100010",
  16750=>"111101111",
  16751=>"111101110",
  16752=>"101011010",
  16753=>"110101001",
  16754=>"111011001",
  16755=>"100111111",
  16756=>"100101110",
  16757=>"110011000",
  16758=>"000010111",
  16759=>"011000110",
  16760=>"010001010",
  16761=>"010001110",
  16762=>"000001110",
  16763=>"000011000",
  16764=>"010101010",
  16765=>"100000111",
  16766=>"000110110",
  16767=>"000100110",
  16768=>"111010001",
  16769=>"001110001",
  16770=>"110100000",
  16771=>"110101101",
  16772=>"000000100",
  16773=>"100000101",
  16774=>"011100101",
  16775=>"111000101",
  16776=>"111000011",
  16777=>"100001010",
  16778=>"110110100",
  16779=>"111010010",
  16780=>"100000001",
  16781=>"011110110",
  16782=>"101000000",
  16783=>"010111111",
  16784=>"101110101",
  16785=>"011011111",
  16786=>"001000111",
  16787=>"010110101",
  16788=>"100101001",
  16789=>"001001101",
  16790=>"011000111",
  16791=>"111100100",
  16792=>"110001010",
  16793=>"100100110",
  16794=>"110101110",
  16795=>"010110001",
  16796=>"101000001",
  16797=>"111111100",
  16798=>"010011000",
  16799=>"011111111",
  16800=>"000011100",
  16801=>"100111101",
  16802=>"111010111",
  16803=>"000011010",
  16804=>"111000000",
  16805=>"001011011",
  16806=>"100101111",
  16807=>"110001010",
  16808=>"010000000",
  16809=>"011100010",
  16810=>"001100101",
  16811=>"100110000",
  16812=>"101001000",
  16813=>"000100110",
  16814=>"011111110",
  16815=>"110011010",
  16816=>"011101110",
  16817=>"100001000",
  16818=>"101101110",
  16819=>"010100010",
  16820=>"001000101",
  16821=>"011100101",
  16822=>"010100000",
  16823=>"010000010",
  16824=>"101011101",
  16825=>"010101000",
  16826=>"100101111",
  16827=>"001111110",
  16828=>"111110101",
  16829=>"111101010",
  16830=>"111100011",
  16831=>"111011100",
  16832=>"111111010",
  16833=>"111111110",
  16834=>"011010111",
  16835=>"011011110",
  16836=>"100010111",
  16837=>"110111001",
  16838=>"111000101",
  16839=>"001011011",
  16840=>"001110000",
  16841=>"110100011",
  16842=>"110010100",
  16843=>"111110011",
  16844=>"110011101",
  16845=>"110001001",
  16846=>"100111100",
  16847=>"101100111",
  16848=>"110001111",
  16849=>"000010010",
  16850=>"011000011",
  16851=>"100100100",
  16852=>"110100101",
  16853=>"011110000",
  16854=>"010111001",
  16855=>"111001010",
  16856=>"001010110",
  16857=>"111011000",
  16858=>"101100100",
  16859=>"000111110",
  16860=>"010111101",
  16861=>"000101111",
  16862=>"011110010",
  16863=>"110101101",
  16864=>"011000000",
  16865=>"110111001",
  16866=>"100000010",
  16867=>"000111110",
  16868=>"111010101",
  16869=>"110011100",
  16870=>"101100101",
  16871=>"101010000",
  16872=>"011001000",
  16873=>"000011110",
  16874=>"001000001",
  16875=>"010111011",
  16876=>"100000100",
  16877=>"101010010",
  16878=>"001000010",
  16879=>"100100100",
  16880=>"011001111",
  16881=>"111110111",
  16882=>"001001011",
  16883=>"110110010",
  16884=>"111001000",
  16885=>"011101001",
  16886=>"010000101",
  16887=>"111010011",
  16888=>"111011011",
  16889=>"110001000",
  16890=>"011001010",
  16891=>"011100000",
  16892=>"010110010",
  16893=>"100010100",
  16894=>"100101000",
  16895=>"111010001",
  16896=>"110100110",
  16897=>"010001110",
  16898=>"000001011",
  16899=>"000111000",
  16900=>"100001111",
  16901=>"000001100",
  16902=>"101001000",
  16903=>"011101110",
  16904=>"101110011",
  16905=>"011001000",
  16906=>"111001010",
  16907=>"001000011",
  16908=>"111010001",
  16909=>"000101100",
  16910=>"001010010",
  16911=>"000011001",
  16912=>"101001011",
  16913=>"000011100",
  16914=>"010101110",
  16915=>"110000101",
  16916=>"101000111",
  16917=>"000111011",
  16918=>"101100010",
  16919=>"101000111",
  16920=>"000111001",
  16921=>"110101010",
  16922=>"001101000",
  16923=>"001000101",
  16924=>"000000100",
  16925=>"000110000",
  16926=>"010001100",
  16927=>"111110011",
  16928=>"011101111",
  16929=>"111101101",
  16930=>"000100001",
  16931=>"100001101",
  16932=>"011111101",
  16933=>"000011011",
  16934=>"010110001",
  16935=>"001001100",
  16936=>"000001100",
  16937=>"011001010",
  16938=>"101001000",
  16939=>"101001111",
  16940=>"010111000",
  16941=>"001010000",
  16942=>"010000010",
  16943=>"000000100",
  16944=>"111111101",
  16945=>"110011100",
  16946=>"001000011",
  16947=>"011101000",
  16948=>"011110010",
  16949=>"100111111",
  16950=>"101101011",
  16951=>"000001000",
  16952=>"100010111",
  16953=>"101011101",
  16954=>"110110101",
  16955=>"011100010",
  16956=>"011001100",
  16957=>"111011101",
  16958=>"000011001",
  16959=>"011000100",
  16960=>"000011110",
  16961=>"111101100",
  16962=>"000001011",
  16963=>"100000100",
  16964=>"101011001",
  16965=>"001110001",
  16966=>"100111011",
  16967=>"101101101",
  16968=>"010010010",
  16969=>"010110010",
  16970=>"010111101",
  16971=>"100111111",
  16972=>"011000010",
  16973=>"101001100",
  16974=>"101011000",
  16975=>"001000111",
  16976=>"010010001",
  16977=>"110100111",
  16978=>"000010001",
  16979=>"000000010",
  16980=>"110101100",
  16981=>"111000100",
  16982=>"001111010",
  16983=>"111001001",
  16984=>"010010000",
  16985=>"000101101",
  16986=>"101110100",
  16987=>"110000101",
  16988=>"100110011",
  16989=>"011000100",
  16990=>"100110000",
  16991=>"011011011",
  16992=>"101000100",
  16993=>"101011010",
  16994=>"101010110",
  16995=>"100110011",
  16996=>"010110010",
  16997=>"101010101",
  16998=>"011111101",
  16999=>"001100000",
  17000=>"000000010",
  17001=>"111010101",
  17002=>"101100011",
  17003=>"011101110",
  17004=>"001110101",
  17005=>"010010000",
  17006=>"000110010",
  17007=>"010101011",
  17008=>"001011110",
  17009=>"111001111",
  17010=>"101101101",
  17011=>"110000110",
  17012=>"101101111",
  17013=>"011011000",
  17014=>"110111011",
  17015=>"000001000",
  17016=>"010111100",
  17017=>"000001110",
  17018=>"010001101",
  17019=>"111110110",
  17020=>"101001001",
  17021=>"000100110",
  17022=>"001010110",
  17023=>"001011101",
  17024=>"111101001",
  17025=>"000110010",
  17026=>"101110000",
  17027=>"000100001",
  17028=>"111001110",
  17029=>"010011001",
  17030=>"011111111",
  17031=>"000001111",
  17032=>"111111000",
  17033=>"110010001",
  17034=>"101101100",
  17035=>"100010010",
  17036=>"110111000",
  17037=>"001001010",
  17038=>"001000110",
  17039=>"111101010",
  17040=>"000111111",
  17041=>"010111001",
  17042=>"000100000",
  17043=>"010010011",
  17044=>"100001011",
  17045=>"000001110",
  17046=>"101000000",
  17047=>"101111100",
  17048=>"110100100",
  17049=>"100100111",
  17050=>"010110100",
  17051=>"100110100",
  17052=>"001110110",
  17053=>"001111000",
  17054=>"101111111",
  17055=>"000100010",
  17056=>"100010111",
  17057=>"110101100",
  17058=>"001010111",
  17059=>"100001000",
  17060=>"001000001",
  17061=>"101110110",
  17062=>"001100000",
  17063=>"111101000",
  17064=>"101101111",
  17065=>"010001001",
  17066=>"001110111",
  17067=>"001101011",
  17068=>"010110111",
  17069=>"111000000",
  17070=>"001001011",
  17071=>"101100110",
  17072=>"010100001",
  17073=>"011011000",
  17074=>"010101111",
  17075=>"111010101",
  17076=>"100011100",
  17077=>"101000101",
  17078=>"101111101",
  17079=>"111111100",
  17080=>"001110010",
  17081=>"001101110",
  17082=>"011101110",
  17083=>"001101111",
  17084=>"100011101",
  17085=>"001000100",
  17086=>"000000100",
  17087=>"111010101",
  17088=>"011101000",
  17089=>"001111010",
  17090=>"111000100",
  17091=>"110010110",
  17092=>"100001100",
  17093=>"111111111",
  17094=>"010001001",
  17095=>"000101000",
  17096=>"001011000",
  17097=>"000100010",
  17098=>"111101010",
  17099=>"000000010",
  17100=>"101001100",
  17101=>"100100010",
  17102=>"000001111",
  17103=>"010000111",
  17104=>"000011010",
  17105=>"000101110",
  17106=>"011111000",
  17107=>"101010110",
  17108=>"010000111",
  17109=>"100111000",
  17110=>"111101110",
  17111=>"010000000",
  17112=>"111001110",
  17113=>"101110011",
  17114=>"100010011",
  17115=>"000010010",
  17116=>"000010100",
  17117=>"010011110",
  17118=>"110000011",
  17119=>"111010000",
  17120=>"001010011",
  17121=>"100000011",
  17122=>"000000100",
  17123=>"001011010",
  17124=>"100010111",
  17125=>"101110110",
  17126=>"011111000",
  17127=>"000010100",
  17128=>"000010011",
  17129=>"000010000",
  17130=>"110001111",
  17131=>"010101000",
  17132=>"010000000",
  17133=>"111101011",
  17134=>"110001011",
  17135=>"100010010",
  17136=>"000100111",
  17137=>"010110000",
  17138=>"010010011",
  17139=>"111100110",
  17140=>"000000101",
  17141=>"101010110",
  17142=>"101110011",
  17143=>"111101010",
  17144=>"001100101",
  17145=>"111100000",
  17146=>"111101000",
  17147=>"001001101",
  17148=>"000011100",
  17149=>"010001010",
  17150=>"110001101",
  17151=>"100110101",
  17152=>"001110111",
  17153=>"101000000",
  17154=>"011010011",
  17155=>"110111110",
  17156=>"100100000",
  17157=>"111011000",
  17158=>"101010100",
  17159=>"011110010",
  17160=>"101011001",
  17161=>"111101111",
  17162=>"110000101",
  17163=>"101011100",
  17164=>"001101011",
  17165=>"010111010",
  17166=>"010000110",
  17167=>"011100110",
  17168=>"000101001",
  17169=>"000001100",
  17170=>"001101001",
  17171=>"101101000",
  17172=>"000111100",
  17173=>"110111100",
  17174=>"111011010",
  17175=>"011000111",
  17176=>"010101001",
  17177=>"100010101",
  17178=>"100001111",
  17179=>"111100110",
  17180=>"110111111",
  17181=>"100001100",
  17182=>"010011011",
  17183=>"111000011",
  17184=>"111101111",
  17185=>"110110001",
  17186=>"001010111",
  17187=>"111110101",
  17188=>"001110111",
  17189=>"111110010",
  17190=>"101000000",
  17191=>"011101110",
  17192=>"100111100",
  17193=>"111011111",
  17194=>"011111111",
  17195=>"000101111",
  17196=>"111101000",
  17197=>"000000110",
  17198=>"000010001",
  17199=>"011111100",
  17200=>"011101000",
  17201=>"011000001",
  17202=>"111111001",
  17203=>"011000111",
  17204=>"000101010",
  17205=>"000001011",
  17206=>"111011001",
  17207=>"101100001",
  17208=>"101011000",
  17209=>"101000011",
  17210=>"101100111",
  17211=>"011010101",
  17212=>"110110001",
  17213=>"101101111",
  17214=>"111011001",
  17215=>"011000000",
  17216=>"101001101",
  17217=>"001000011",
  17218=>"111110010",
  17219=>"111111110",
  17220=>"000011101",
  17221=>"100010101",
  17222=>"010000101",
  17223=>"011011111",
  17224=>"011001011",
  17225=>"100001111",
  17226=>"000111011",
  17227=>"001110011",
  17228=>"101001100",
  17229=>"011010011",
  17230=>"111101011",
  17231=>"101000100",
  17232=>"110000000",
  17233=>"001001111",
  17234=>"111000110",
  17235=>"001000111",
  17236=>"111110100",
  17237=>"110100111",
  17238=>"110011110",
  17239=>"001100100",
  17240=>"100010111",
  17241=>"000100111",
  17242=>"011000000",
  17243=>"010010000",
  17244=>"110111111",
  17245=>"100111001",
  17246=>"001001100",
  17247=>"010000000",
  17248=>"010000101",
  17249=>"001011000",
  17250=>"100000101",
  17251=>"000100101",
  17252=>"011100101",
  17253=>"110100000",
  17254=>"100110111",
  17255=>"000111100",
  17256=>"111101101",
  17257=>"100001010",
  17258=>"110111111",
  17259=>"101000111",
  17260=>"011110110",
  17261=>"100111100",
  17262=>"100011011",
  17263=>"110111010",
  17264=>"111001011",
  17265=>"111000010",
  17266=>"110011001",
  17267=>"010011010",
  17268=>"001110110",
  17269=>"101110010",
  17270=>"110000100",
  17271=>"111101010",
  17272=>"011101000",
  17273=>"001001111",
  17274=>"010000000",
  17275=>"110101010",
  17276=>"111100110",
  17277=>"010011101",
  17278=>"110001111",
  17279=>"010010010",
  17280=>"000111101",
  17281=>"011010000",
  17282=>"011110001",
  17283=>"000111001",
  17284=>"101100110",
  17285=>"110001001",
  17286=>"111011110",
  17287=>"001011111",
  17288=>"000010110",
  17289=>"001111001",
  17290=>"011011111",
  17291=>"010001100",
  17292=>"010101010",
  17293=>"110110001",
  17294=>"000110000",
  17295=>"101101001",
  17296=>"000110010",
  17297=>"010110011",
  17298=>"000000000",
  17299=>"001011110",
  17300=>"010000110",
  17301=>"111101111",
  17302=>"001110010",
  17303=>"010101010",
  17304=>"001001101",
  17305=>"001000000",
  17306=>"111111000",
  17307=>"001000110",
  17308=>"111001000",
  17309=>"010001000",
  17310=>"001000101",
  17311=>"000100010",
  17312=>"010001010",
  17313=>"001100011",
  17314=>"100010101",
  17315=>"101110111",
  17316=>"011100011",
  17317=>"100011111",
  17318=>"110011100",
  17319=>"000010001",
  17320=>"001011100",
  17321=>"101000111",
  17322=>"011110000",
  17323=>"110010100",
  17324=>"010101000",
  17325=>"011100110",
  17326=>"100110111",
  17327=>"001011111",
  17328=>"101101000",
  17329=>"110100000",
  17330=>"011010100",
  17331=>"111010000",
  17332=>"011000011",
  17333=>"100001101",
  17334=>"101011010",
  17335=>"000001101",
  17336=>"011111110",
  17337=>"101001011",
  17338=>"100111011",
  17339=>"010110111",
  17340=>"010101010",
  17341=>"111010000",
  17342=>"011101001",
  17343=>"110011100",
  17344=>"000100101",
  17345=>"101000001",
  17346=>"101000010",
  17347=>"100101010",
  17348=>"000001010",
  17349=>"110110001",
  17350=>"110111111",
  17351=>"101000100",
  17352=>"110110110",
  17353=>"110100001",
  17354=>"100110001",
  17355=>"110011100",
  17356=>"100110001",
  17357=>"011010100",
  17358=>"010100001",
  17359=>"011000001",
  17360=>"001010001",
  17361=>"101001101",
  17362=>"111011101",
  17363=>"110111101",
  17364=>"100001010",
  17365=>"000001111",
  17366=>"000000000",
  17367=>"000111000",
  17368=>"000000101",
  17369=>"100001000",
  17370=>"011111101",
  17371=>"110110111",
  17372=>"010100001",
  17373=>"111011110",
  17374=>"101000000",
  17375=>"111000011",
  17376=>"111010010",
  17377=>"111001101",
  17378=>"011001000",
  17379=>"111001101",
  17380=>"110111001",
  17381=>"010011011",
  17382=>"010011011",
  17383=>"110000111",
  17384=>"111111101",
  17385=>"101001001",
  17386=>"000100110",
  17387=>"001101111",
  17388=>"111101011",
  17389=>"100100101",
  17390=>"011000000",
  17391=>"010111100",
  17392=>"001010000",
  17393=>"010100100",
  17394=>"011110111",
  17395=>"101010111",
  17396=>"101011011",
  17397=>"101100011",
  17398=>"111011000",
  17399=>"010010101",
  17400=>"110101100",
  17401=>"101101000",
  17402=>"011000000",
  17403=>"001000111",
  17404=>"110101101",
  17405=>"010010011",
  17406=>"000111011",
  17407=>"101100011",
  17408=>"101111010",
  17409=>"100101111",
  17410=>"000100010",
  17411=>"010111100",
  17412=>"110100010",
  17413=>"110010011",
  17414=>"100010100",
  17415=>"001111101",
  17416=>"111000110",
  17417=>"100010101",
  17418=>"000011000",
  17419=>"000011001",
  17420=>"110010010",
  17421=>"010000011",
  17422=>"010000010",
  17423=>"000010101",
  17424=>"001000011",
  17425=>"010001010",
  17426=>"100100010",
  17427=>"000000111",
  17428=>"000110011",
  17429=>"100010010",
  17430=>"100110111",
  17431=>"100010101",
  17432=>"111000000",
  17433=>"111000011",
  17434=>"010001010",
  17435=>"110101000",
  17436=>"111101101",
  17437=>"111111111",
  17438=>"001011001",
  17439=>"110101101",
  17440=>"110101010",
  17441=>"110101101",
  17442=>"100100100",
  17443=>"111010001",
  17444=>"001100000",
  17445=>"111110011",
  17446=>"000110111",
  17447=>"001111111",
  17448=>"100001000",
  17449=>"000101010",
  17450=>"000011110",
  17451=>"001011000",
  17452=>"100000101",
  17453=>"111110010",
  17454=>"111000001",
  17455=>"100100011",
  17456=>"101010110",
  17457=>"010010010",
  17458=>"011010000",
  17459=>"000100110",
  17460=>"010011100",
  17461=>"000100001",
  17462=>"010110110",
  17463=>"011010100",
  17464=>"010101111",
  17465=>"000101001",
  17466=>"011110110",
  17467=>"000111111",
  17468=>"011000001",
  17469=>"111001011",
  17470=>"000110100",
  17471=>"101110011",
  17472=>"101111111",
  17473=>"011000010",
  17474=>"111101010",
  17475=>"001110111",
  17476=>"001010111",
  17477=>"101110001",
  17478=>"000011001",
  17479=>"000001110",
  17480=>"011111011",
  17481=>"111010100",
  17482=>"010001000",
  17483=>"111110110",
  17484=>"111000000",
  17485=>"111110000",
  17486=>"111110110",
  17487=>"000001010",
  17488=>"110100011",
  17489=>"000110011",
  17490=>"000100111",
  17491=>"110101000",
  17492=>"100010100",
  17493=>"001010011",
  17494=>"111111111",
  17495=>"001000001",
  17496=>"100111110",
  17497=>"000010001",
  17498=>"100110110",
  17499=>"001010111",
  17500=>"011111110",
  17501=>"111001101",
  17502=>"111001011",
  17503=>"000011100",
  17504=>"000001010",
  17505=>"011110011",
  17506=>"100011110",
  17507=>"001010000",
  17508=>"011011000",
  17509=>"100000111",
  17510=>"101000011",
  17511=>"000011010",
  17512=>"101000010",
  17513=>"011000011",
  17514=>"010001000",
  17515=>"010111110",
  17516=>"110101101",
  17517=>"011110100",
  17518=>"111011110",
  17519=>"000100110",
  17520=>"111110000",
  17521=>"000101100",
  17522=>"000011001",
  17523=>"000110011",
  17524=>"101110100",
  17525=>"101111010",
  17526=>"100111010",
  17527=>"100110100",
  17528=>"100111010",
  17529=>"110110001",
  17530=>"111101010",
  17531=>"101100011",
  17532=>"101010110",
  17533=>"001110110",
  17534=>"111011001",
  17535=>"000001110",
  17536=>"000000100",
  17537=>"110101110",
  17538=>"111101001",
  17539=>"111011100",
  17540=>"001010010",
  17541=>"011100001",
  17542=>"101101011",
  17543=>"001001101",
  17544=>"111101101",
  17545=>"110101001",
  17546=>"110011000",
  17547=>"011001100",
  17548=>"000001110",
  17549=>"110111100",
  17550=>"100000111",
  17551=>"001110101",
  17552=>"110101111",
  17553=>"011100001",
  17554=>"000011101",
  17555=>"100111110",
  17556=>"000010010",
  17557=>"011001100",
  17558=>"101101011",
  17559=>"000111001",
  17560=>"011110011",
  17561=>"001110100",
  17562=>"110011110",
  17563=>"011011111",
  17564=>"110001000",
  17565=>"111000010",
  17566=>"101011110",
  17567=>"100001110",
  17568=>"001110011",
  17569=>"000111101",
  17570=>"101010000",
  17571=>"000110001",
  17572=>"110001110",
  17573=>"001001101",
  17574=>"110000011",
  17575=>"010000000",
  17576=>"001111111",
  17577=>"000110010",
  17578=>"000000100",
  17579=>"000100001",
  17580=>"110110110",
  17581=>"111000011",
  17582=>"011111110",
  17583=>"010101111",
  17584=>"000000000",
  17585=>"001111001",
  17586=>"000001100",
  17587=>"001000110",
  17588=>"100111100",
  17589=>"011110001",
  17590=>"110100100",
  17591=>"101110001",
  17592=>"010111011",
  17593=>"101001011",
  17594=>"100100100",
  17595=>"110110100",
  17596=>"101110100",
  17597=>"000101011",
  17598=>"110001001",
  17599=>"101100110",
  17600=>"100101111",
  17601=>"010001000",
  17602=>"110011101",
  17603=>"010101101",
  17604=>"010001110",
  17605=>"001111010",
  17606=>"110101110",
  17607=>"010000001",
  17608=>"010000000",
  17609=>"110110100",
  17610=>"101110010",
  17611=>"101001010",
  17612=>"110000111",
  17613=>"010100001",
  17614=>"001111001",
  17615=>"100100010",
  17616=>"000000100",
  17617=>"100111001",
  17618=>"101100010",
  17619=>"101010101",
  17620=>"110001000",
  17621=>"001100000",
  17622=>"000101010",
  17623=>"101101000",
  17624=>"100001101",
  17625=>"001010101",
  17626=>"010110000",
  17627=>"000001110",
  17628=>"010010011",
  17629=>"010101110",
  17630=>"011110101",
  17631=>"100111110",
  17632=>"010001001",
  17633=>"000000000",
  17634=>"101111110",
  17635=>"111101001",
  17636=>"010010101",
  17637=>"011101011",
  17638=>"110101101",
  17639=>"000001101",
  17640=>"100001010",
  17641=>"110001001",
  17642=>"001110000",
  17643=>"111101111",
  17644=>"011110111",
  17645=>"010011010",
  17646=>"011110001",
  17647=>"000000101",
  17648=>"011000100",
  17649=>"001110000",
  17650=>"111000110",
  17651=>"010001001",
  17652=>"100111000",
  17653=>"111111110",
  17654=>"001010010",
  17655=>"011001010",
  17656=>"110010011",
  17657=>"110111101",
  17658=>"011110011",
  17659=>"101001100",
  17660=>"010100000",
  17661=>"100101010",
  17662=>"010110110",
  17663=>"111001111",
  17664=>"000110111",
  17665=>"000111100",
  17666=>"100010000",
  17667=>"110100110",
  17668=>"001111100",
  17669=>"011101011",
  17670=>"011000000",
  17671=>"100100000",
  17672=>"100000101",
  17673=>"100000001",
  17674=>"011101010",
  17675=>"000101000",
  17676=>"000111000",
  17677=>"000011110",
  17678=>"110010100",
  17679=>"001111111",
  17680=>"101000010",
  17681=>"011001010",
  17682=>"101010100",
  17683=>"100110101",
  17684=>"100001110",
  17685=>"100011101",
  17686=>"001011000",
  17687=>"001000100",
  17688=>"100010000",
  17689=>"110010100",
  17690=>"111000010",
  17691=>"011101100",
  17692=>"011011110",
  17693=>"111011110",
  17694=>"100001101",
  17695=>"010011100",
  17696=>"010101110",
  17697=>"000000011",
  17698=>"100100000",
  17699=>"110001010",
  17700=>"001001100",
  17701=>"101000100",
  17702=>"000000010",
  17703=>"000000110",
  17704=>"011000111",
  17705=>"001000011",
  17706=>"100000000",
  17707=>"011100000",
  17708=>"101100111",
  17709=>"100010011",
  17710=>"100111000",
  17711=>"000011110",
  17712=>"001111110",
  17713=>"000111000",
  17714=>"011001101",
  17715=>"100110101",
  17716=>"111110011",
  17717=>"100000101",
  17718=>"011001110",
  17719=>"101100010",
  17720=>"100110000",
  17721=>"111001010",
  17722=>"101010110",
  17723=>"111111011",
  17724=>"011110001",
  17725=>"001001001",
  17726=>"000111000",
  17727=>"011111111",
  17728=>"111101001",
  17729=>"111111110",
  17730=>"101000010",
  17731=>"101000011",
  17732=>"001110000",
  17733=>"111010110",
  17734=>"000010101",
  17735=>"011111111",
  17736=>"011011011",
  17737=>"010111110",
  17738=>"000011001",
  17739=>"100000101",
  17740=>"110011111",
  17741=>"000111110",
  17742=>"111011011",
  17743=>"000010101",
  17744=>"100011011",
  17745=>"010000010",
  17746=>"111100010",
  17747=>"000111100",
  17748=>"101010110",
  17749=>"001011010",
  17750=>"100001110",
  17751=>"010001110",
  17752=>"100000010",
  17753=>"100010001",
  17754=>"111000101",
  17755=>"100000001",
  17756=>"101100001",
  17757=>"001001110",
  17758=>"001111101",
  17759=>"000010110",
  17760=>"111100110",
  17761=>"111110000",
  17762=>"110010011",
  17763=>"010110011",
  17764=>"100111110",
  17765=>"100001010",
  17766=>"110000101",
  17767=>"100011010",
  17768=>"000100111",
  17769=>"000100100",
  17770=>"000101001",
  17771=>"011100100",
  17772=>"011000001",
  17773=>"100101001",
  17774=>"010111000",
  17775=>"000110110",
  17776=>"000000001",
  17777=>"001100100",
  17778=>"111000001",
  17779=>"001110010",
  17780=>"000101000",
  17781=>"101011100",
  17782=>"101010010",
  17783=>"100001001",
  17784=>"110110010",
  17785=>"000001001",
  17786=>"010001000",
  17787=>"110101111",
  17788=>"001001101",
  17789=>"000111010",
  17790=>"101011011",
  17791=>"001110011",
  17792=>"011110001",
  17793=>"101000000",
  17794=>"111100101",
  17795=>"111101101",
  17796=>"100001010",
  17797=>"010110010",
  17798=>"000001110",
  17799=>"100001100",
  17800=>"101101000",
  17801=>"001110010",
  17802=>"101000111",
  17803=>"101100101",
  17804=>"110110111",
  17805=>"110010010",
  17806=>"000111111",
  17807=>"100111101",
  17808=>"100100011",
  17809=>"010100110",
  17810=>"011001010",
  17811=>"011111001",
  17812=>"010101111",
  17813=>"011000101",
  17814=>"111110111",
  17815=>"010110100",
  17816=>"000001001",
  17817=>"110110000",
  17818=>"111111000",
  17819=>"001111100",
  17820=>"101100111",
  17821=>"000011010",
  17822=>"111001110",
  17823=>"111101010",
  17824=>"111111000",
  17825=>"000010000",
  17826=>"010000001",
  17827=>"011000000",
  17828=>"100010100",
  17829=>"100000111",
  17830=>"001100000",
  17831=>"111110111",
  17832=>"011001110",
  17833=>"010110101",
  17834=>"110011101",
  17835=>"110001000",
  17836=>"010011000",
  17837=>"111010111",
  17838=>"110000010",
  17839=>"011000100",
  17840=>"010110010",
  17841=>"100001100",
  17842=>"100110100",
  17843=>"011000011",
  17844=>"101010010",
  17845=>"000001101",
  17846=>"111011111",
  17847=>"111101110",
  17848=>"111000110",
  17849=>"100110100",
  17850=>"010011101",
  17851=>"111011111",
  17852=>"010100000",
  17853=>"010101100",
  17854=>"101011000",
  17855=>"111000010",
  17856=>"110011000",
  17857=>"001111101",
  17858=>"001111000",
  17859=>"111101101",
  17860=>"111101000",
  17861=>"000011011",
  17862=>"111010001",
  17863=>"111001000",
  17864=>"111101000",
  17865=>"101000001",
  17866=>"001101010",
  17867=>"011111101",
  17868=>"000000011",
  17869=>"010010001",
  17870=>"100000010",
  17871=>"111000011",
  17872=>"110101111",
  17873=>"110100011",
  17874=>"111000011",
  17875=>"000110111",
  17876=>"110111010",
  17877=>"011001011",
  17878=>"111001111",
  17879=>"110010101",
  17880=>"000110100",
  17881=>"000011111",
  17882=>"101100110",
  17883=>"000011000",
  17884=>"111001001",
  17885=>"000000010",
  17886=>"000110011",
  17887=>"100011010",
  17888=>"100011001",
  17889=>"001110111",
  17890=>"010111100",
  17891=>"101001100",
  17892=>"101001101",
  17893=>"011111010",
  17894=>"010101001",
  17895=>"000011011",
  17896=>"111011011",
  17897=>"101001110",
  17898=>"001000111",
  17899=>"011011010",
  17900=>"100110100",
  17901=>"100010010",
  17902=>"000001110",
  17903=>"000000000",
  17904=>"110011100",
  17905=>"011110101",
  17906=>"100111111",
  17907=>"000010100",
  17908=>"010101011",
  17909=>"101001100",
  17910=>"000100000",
  17911=>"111000010",
  17912=>"001110001",
  17913=>"011001100",
  17914=>"010010111",
  17915=>"100101110",
  17916=>"001101111",
  17917=>"100000111",
  17918=>"010101101",
  17919=>"010111101",
  17920=>"100010111",
  17921=>"110111000",
  17922=>"100011011",
  17923=>"000010001",
  17924=>"011100000",
  17925=>"001000011",
  17926=>"111000100",
  17927=>"000010111",
  17928=>"011100000",
  17929=>"111100001",
  17930=>"101000100",
  17931=>"001001100",
  17932=>"000100010",
  17933=>"011111110",
  17934=>"000000011",
  17935=>"010011110",
  17936=>"111000011",
  17937=>"010010100",
  17938=>"111111010",
  17939=>"010001100",
  17940=>"100101011",
  17941=>"101100011",
  17942=>"001101101",
  17943=>"110111100",
  17944=>"001001100",
  17945=>"011111100",
  17946=>"000011110",
  17947=>"011000111",
  17948=>"111110010",
  17949=>"000000000",
  17950=>"010101010",
  17951=>"101010001",
  17952=>"101010101",
  17953=>"010100110",
  17954=>"100011100",
  17955=>"000001101",
  17956=>"000011101",
  17957=>"100001101",
  17958=>"001000000",
  17959=>"001010011",
  17960=>"010000000",
  17961=>"011101000",
  17962=>"111000000",
  17963=>"100000101",
  17964=>"010110000",
  17965=>"010010001",
  17966=>"100110100",
  17967=>"011110100",
  17968=>"011010100",
  17969=>"100011010",
  17970=>"101000100",
  17971=>"101100101",
  17972=>"100110000",
  17973=>"111101000",
  17974=>"100110010",
  17975=>"101101101",
  17976=>"100010110",
  17977=>"100110011",
  17978=>"101110111",
  17979=>"111110100",
  17980=>"001110110",
  17981=>"100110000",
  17982=>"111011001",
  17983=>"001001011",
  17984=>"001111110",
  17985=>"001111000",
  17986=>"100011001",
  17987=>"011101111",
  17988=>"010100011",
  17989=>"110010100",
  17990=>"010011110",
  17991=>"101111011",
  17992=>"100100110",
  17993=>"100000111",
  17994=>"101100110",
  17995=>"011000110",
  17996=>"001001100",
  17997=>"101010000",
  17998=>"011101010",
  17999=>"011110100",
  18000=>"111101010",
  18001=>"101001010",
  18002=>"100111111",
  18003=>"101110101",
  18004=>"101001000",
  18005=>"001010011",
  18006=>"001111011",
  18007=>"100001111",
  18008=>"111111101",
  18009=>"110111010",
  18010=>"010111010",
  18011=>"111000111",
  18012=>"100101010",
  18013=>"010000101",
  18014=>"100100000",
  18015=>"100101101",
  18016=>"000110101",
  18017=>"011110000",
  18018=>"111110000",
  18019=>"110100001",
  18020=>"001001110",
  18021=>"101001100",
  18022=>"111001100",
  18023=>"100111110",
  18024=>"000100101",
  18025=>"011110111",
  18026=>"001001111",
  18027=>"100101100",
  18028=>"111000000",
  18029=>"111000111",
  18030=>"100010101",
  18031=>"001101011",
  18032=>"010101000",
  18033=>"101011101",
  18034=>"010000110",
  18035=>"111101011",
  18036=>"010000110",
  18037=>"110010110",
  18038=>"010101110",
  18039=>"010001001",
  18040=>"101110000",
  18041=>"110011010",
  18042=>"001011110",
  18043=>"110100100",
  18044=>"110001001",
  18045=>"011111011",
  18046=>"011000001",
  18047=>"110111110",
  18048=>"110101000",
  18049=>"000111010",
  18050=>"100000100",
  18051=>"001011101",
  18052=>"110111001",
  18053=>"000001110",
  18054=>"010000010",
  18055=>"100000000",
  18056=>"111001110",
  18057=>"001111001",
  18058=>"000110011",
  18059=>"000111010",
  18060=>"100110111",
  18061=>"111001111",
  18062=>"111101111",
  18063=>"110111011",
  18064=>"111011101",
  18065=>"110110101",
  18066=>"000111011",
  18067=>"010001101",
  18068=>"001001000",
  18069=>"111111011",
  18070=>"010100001",
  18071=>"110110111",
  18072=>"011100101",
  18073=>"101101011",
  18074=>"101001011",
  18075=>"110111010",
  18076=>"100100000",
  18077=>"100010000",
  18078=>"110111100",
  18079=>"000001110",
  18080=>"110011111",
  18081=>"011111100",
  18082=>"011100011",
  18083=>"100000101",
  18084=>"010100111",
  18085=>"001110011",
  18086=>"110011001",
  18087=>"010010000",
  18088=>"101110000",
  18089=>"101111000",
  18090=>"101000100",
  18091=>"110100000",
  18092=>"000100101",
  18093=>"000111101",
  18094=>"111001010",
  18095=>"100011110",
  18096=>"100100100",
  18097=>"011110110",
  18098=>"010110010",
  18099=>"101101010",
  18100=>"100100001",
  18101=>"001110000",
  18102=>"110101100",
  18103=>"110101110",
  18104=>"101101000",
  18105=>"101010011",
  18106=>"110001101",
  18107=>"011011100",
  18108=>"101001011",
  18109=>"111010011",
  18110=>"010010110",
  18111=>"111111011",
  18112=>"010000011",
  18113=>"101011011",
  18114=>"111000001",
  18115=>"111101111",
  18116=>"111000011",
  18117=>"101010100",
  18118=>"001010100",
  18119=>"100001010",
  18120=>"011011101",
  18121=>"111011111",
  18122=>"010101100",
  18123=>"110110010",
  18124=>"111001111",
  18125=>"101110000",
  18126=>"011110100",
  18127=>"010000101",
  18128=>"000111010",
  18129=>"110000011",
  18130=>"110011010",
  18131=>"100010110",
  18132=>"100100100",
  18133=>"010010010",
  18134=>"001010001",
  18135=>"100011001",
  18136=>"000101000",
  18137=>"010010010",
  18138=>"000000111",
  18139=>"110010001",
  18140=>"000100011",
  18141=>"001010101",
  18142=>"011011011",
  18143=>"100110101",
  18144=>"101111100",
  18145=>"101001000",
  18146=>"110110101",
  18147=>"000101111",
  18148=>"001100111",
  18149=>"011111110",
  18150=>"001101001",
  18151=>"101011000",
  18152=>"001101101",
  18153=>"010010011",
  18154=>"111010110",
  18155=>"101001100",
  18156=>"000000000",
  18157=>"100000011",
  18158=>"111011010",
  18159=>"101010111",
  18160=>"101110000",
  18161=>"010101110",
  18162=>"111100010",
  18163=>"111010001",
  18164=>"001100101",
  18165=>"110101100",
  18166=>"110100100",
  18167=>"101010010",
  18168=>"101010011",
  18169=>"001001011",
  18170=>"111100011",
  18171=>"010101000",
  18172=>"110010000",
  18173=>"010011100",
  18174=>"101111100",
  18175=>"000010000",
  18176=>"100010110",
  18177=>"000000001",
  18178=>"110101011",
  18179=>"101101101",
  18180=>"100101110",
  18181=>"010010000",
  18182=>"111000110",
  18183=>"000001001",
  18184=>"001001100",
  18185=>"100001001",
  18186=>"011010111",
  18187=>"011011000",
  18188=>"100011001",
  18189=>"110011010",
  18190=>"101010000",
  18191=>"101111111",
  18192=>"101110101",
  18193=>"100101110",
  18194=>"010101001",
  18195=>"001000011",
  18196=>"011010001",
  18197=>"000101101",
  18198=>"110001100",
  18199=>"110101100",
  18200=>"111101111",
  18201=>"011000101",
  18202=>"100010100",
  18203=>"001111100",
  18204=>"110101101",
  18205=>"000010100",
  18206=>"110000000",
  18207=>"111001001",
  18208=>"110100111",
  18209=>"101101110",
  18210=>"110101011",
  18211=>"111111100",
  18212=>"111111010",
  18213=>"001000010",
  18214=>"111110100",
  18215=>"010000010",
  18216=>"001000011",
  18217=>"010110101",
  18218=>"000001110",
  18219=>"100000001",
  18220=>"000110011",
  18221=>"010010001",
  18222=>"001001001",
  18223=>"100001000",
  18224=>"101100010",
  18225=>"111011011",
  18226=>"000010010",
  18227=>"101111110",
  18228=>"011100011",
  18229=>"011000001",
  18230=>"000101001",
  18231=>"010001110",
  18232=>"001011011",
  18233=>"000111011",
  18234=>"111111100",
  18235=>"111101100",
  18236=>"000001111",
  18237=>"011000001",
  18238=>"011011110",
  18239=>"100000011",
  18240=>"000001100",
  18241=>"011011000",
  18242=>"001010111",
  18243=>"011111100",
  18244=>"101000100",
  18245=>"010010101",
  18246=>"001000110",
  18247=>"010110011",
  18248=>"010001101",
  18249=>"001001100",
  18250=>"011101011",
  18251=>"101110100",
  18252=>"101101101",
  18253=>"100100000",
  18254=>"000100010",
  18255=>"110010111",
  18256=>"001001000",
  18257=>"000011110",
  18258=>"001001100",
  18259=>"011001000",
  18260=>"111110011",
  18261=>"011000110",
  18262=>"100100110",
  18263=>"110011000",
  18264=>"110111010",
  18265=>"011001100",
  18266=>"011101100",
  18267=>"110101011",
  18268=>"000101011",
  18269=>"011111100",
  18270=>"101110101",
  18271=>"100010000",
  18272=>"111000001",
  18273=>"001011101",
  18274=>"001110001",
  18275=>"010000010",
  18276=>"001011011",
  18277=>"111101011",
  18278=>"111001110",
  18279=>"010101010",
  18280=>"010110000",
  18281=>"000011000",
  18282=>"100001010",
  18283=>"000111100",
  18284=>"111001011",
  18285=>"001000010",
  18286=>"001111110",
  18287=>"010010010",
  18288=>"100001011",
  18289=>"111100000",
  18290=>"111000100",
  18291=>"101111100",
  18292=>"011000101",
  18293=>"101001101",
  18294=>"001001111",
  18295=>"100101000",
  18296=>"100011001",
  18297=>"110110010",
  18298=>"111010110",
  18299=>"101111101",
  18300=>"000000010",
  18301=>"110100111",
  18302=>"101011101",
  18303=>"111000101",
  18304=>"001000111",
  18305=>"110110011",
  18306=>"110010010",
  18307=>"101000010",
  18308=>"110100011",
  18309=>"011001010",
  18310=>"010100110",
  18311=>"111000000",
  18312=>"101010011",
  18313=>"101010011",
  18314=>"101101101",
  18315=>"111000101",
  18316=>"011001011",
  18317=>"110000000",
  18318=>"111010011",
  18319=>"011101101",
  18320=>"010110001",
  18321=>"111101010",
  18322=>"001000111",
  18323=>"001001100",
  18324=>"000000111",
  18325=>"000000100",
  18326=>"111010001",
  18327=>"111111111",
  18328=>"101011111",
  18329=>"010101101",
  18330=>"001001000",
  18331=>"110101010",
  18332=>"110111001",
  18333=>"100111111",
  18334=>"010011101",
  18335=>"101110010",
  18336=>"100011100",
  18337=>"001010011",
  18338=>"011100100",
  18339=>"000000000",
  18340=>"001010010",
  18341=>"100001000",
  18342=>"010100001",
  18343=>"010100000",
  18344=>"010100011",
  18345=>"011001011",
  18346=>"000001110",
  18347=>"101010011",
  18348=>"000000000",
  18349=>"100110111",
  18350=>"101100100",
  18351=>"101100000",
  18352=>"011101000",
  18353=>"111011011",
  18354=>"000001111",
  18355=>"110111001",
  18356=>"100010001",
  18357=>"110110110",
  18358=>"000010001",
  18359=>"111111111",
  18360=>"110111100",
  18361=>"000110111",
  18362=>"011000011",
  18363=>"010100111",
  18364=>"010110011",
  18365=>"000101110",
  18366=>"100101010",
  18367=>"010101101",
  18368=>"000100101",
  18369=>"111101101",
  18370=>"001000101",
  18371=>"100000001",
  18372=>"100011110",
  18373=>"110010111",
  18374=>"010110011",
  18375=>"001011001",
  18376=>"100001000",
  18377=>"100101100",
  18378=>"000010000",
  18379=>"000100011",
  18380=>"100011010",
  18381=>"011100100",
  18382=>"010111010",
  18383=>"010001111",
  18384=>"100100110",
  18385=>"011010110",
  18386=>"011000110",
  18387=>"000100000",
  18388=>"011100100",
  18389=>"010001110",
  18390=>"001110110",
  18391=>"000000000",
  18392=>"111011001",
  18393=>"000001101",
  18394=>"101011010",
  18395=>"111111011",
  18396=>"101100111",
  18397=>"110101011",
  18398=>"111010100",
  18399=>"111000100",
  18400=>"100111100",
  18401=>"111111010",
  18402=>"110100101",
  18403=>"101011001",
  18404=>"011010110",
  18405=>"001011111",
  18406=>"111111011",
  18407=>"100000000",
  18408=>"100000010",
  18409=>"110101000",
  18410=>"000000101",
  18411=>"110000011",
  18412=>"011000111",
  18413=>"001010110",
  18414=>"100101000",
  18415=>"101011000",
  18416=>"010010100",
  18417=>"111010000",
  18418=>"001110100",
  18419=>"000011010",
  18420=>"111110111",
  18421=>"000100100",
  18422=>"110001010",
  18423=>"000101010",
  18424=>"111111111",
  18425=>"100000000",
  18426=>"000100110",
  18427=>"100110101",
  18428=>"111101111",
  18429=>"101001000",
  18430=>"010111000",
  18431=>"001010111",
  18432=>"000110010",
  18433=>"011100101",
  18434=>"100110011",
  18435=>"001111101",
  18436=>"111010111",
  18437=>"011101110",
  18438=>"000001100",
  18439=>"100101101",
  18440=>"000100100",
  18441=>"110000101",
  18442=>"110011011",
  18443=>"010001100",
  18444=>"010100100",
  18445=>"110110010",
  18446=>"100010001",
  18447=>"010110000",
  18448=>"011001100",
  18449=>"000001110",
  18450=>"010100000",
  18451=>"100010001",
  18452=>"110000100",
  18453=>"000100001",
  18454=>"011000110",
  18455=>"010001000",
  18456=>"110111000",
  18457=>"000110101",
  18458=>"010010001",
  18459=>"001000100",
  18460=>"101100100",
  18461=>"110010110",
  18462=>"100101100",
  18463=>"001111010",
  18464=>"100101001",
  18465=>"101101110",
  18466=>"001101001",
  18467=>"011001001",
  18468=>"010011101",
  18469=>"100111110",
  18470=>"000001100",
  18471=>"001010011",
  18472=>"111000001",
  18473=>"001111010",
  18474=>"000011111",
  18475=>"001110101",
  18476=>"110111100",
  18477=>"011000111",
  18478=>"111001101",
  18479=>"001011110",
  18480=>"011111000",
  18481=>"111111011",
  18482=>"110100100",
  18483=>"010101110",
  18484=>"110100111",
  18485=>"101111101",
  18486=>"101001000",
  18487=>"100101111",
  18488=>"010000010",
  18489=>"111001010",
  18490=>"111001111",
  18491=>"111101001",
  18492=>"001100101",
  18493=>"111110000",
  18494=>"110101001",
  18495=>"100101011",
  18496=>"100000111",
  18497=>"011011001",
  18498=>"010110000",
  18499=>"110101110",
  18500=>"011011000",
  18501=>"101111111",
  18502=>"111000101",
  18503=>"111111111",
  18504=>"000001110",
  18505=>"000101110",
  18506=>"010010000",
  18507=>"111010000",
  18508=>"011101101",
  18509=>"100101000",
  18510=>"000100001",
  18511=>"110100010",
  18512=>"111011100",
  18513=>"010011010",
  18514=>"100111101",
  18515=>"101001010",
  18516=>"001010111",
  18517=>"100110010",
  18518=>"100101010",
  18519=>"010101100",
  18520=>"101011011",
  18521=>"111110011",
  18522=>"010000010",
  18523=>"101011001",
  18524=>"011101010",
  18525=>"000100001",
  18526=>"000100110",
  18527=>"010011111",
  18528=>"001011101",
  18529=>"010101000",
  18530=>"011001100",
  18531=>"010110001",
  18532=>"010100100",
  18533=>"100010010",
  18534=>"100000100",
  18535=>"110110100",
  18536=>"101010101",
  18537=>"010010111",
  18538=>"001000110",
  18539=>"011111111",
  18540=>"110011100",
  18541=>"111000010",
  18542=>"010011010",
  18543=>"000111100",
  18544=>"011001111",
  18545=>"111101111",
  18546=>"010111011",
  18547=>"111101000",
  18548=>"110111000",
  18549=>"010001101",
  18550=>"101101111",
  18551=>"010011010",
  18552=>"001110111",
  18553=>"101101000",
  18554=>"011101010",
  18555=>"100010111",
  18556=>"000101000",
  18557=>"000011101",
  18558=>"010101001",
  18559=>"001000110",
  18560=>"000111110",
  18561=>"011100001",
  18562=>"001110000",
  18563=>"010100011",
  18564=>"111000001",
  18565=>"001011111",
  18566=>"011001101",
  18567=>"101000101",
  18568=>"011101100",
  18569=>"001000100",
  18570=>"000010001",
  18571=>"101000010",
  18572=>"110100001",
  18573=>"010000010",
  18574=>"110110001",
  18575=>"001100101",
  18576=>"010001100",
  18577=>"010110001",
  18578=>"101010100",
  18579=>"001010001",
  18580=>"010001100",
  18581=>"100101100",
  18582=>"001001111",
  18583=>"111100010",
  18584=>"010101101",
  18585=>"011010001",
  18586=>"111000101",
  18587=>"001001100",
  18588=>"010100110",
  18589=>"010111110",
  18590=>"011001110",
  18591=>"100100000",
  18592=>"011011010",
  18593=>"000110110",
  18594=>"000010000",
  18595=>"110110100",
  18596=>"100011011",
  18597=>"011111101",
  18598=>"110111101",
  18599=>"001010111",
  18600=>"100010010",
  18601=>"010101110",
  18602=>"111011110",
  18603=>"101111001",
  18604=>"110100010",
  18605=>"011011111",
  18606=>"110001101",
  18607=>"101100110",
  18608=>"100000011",
  18609=>"111110100",
  18610=>"000100010",
  18611=>"010110001",
  18612=>"001100011",
  18613=>"010110011",
  18614=>"101110110",
  18615=>"010011101",
  18616=>"001010010",
  18617=>"011111101",
  18618=>"101000110",
  18619=>"000010100",
  18620=>"101100100",
  18621=>"110010100",
  18622=>"011001100",
  18623=>"110110001",
  18624=>"110000000",
  18625=>"100100100",
  18626=>"101000011",
  18627=>"100100001",
  18628=>"111111110",
  18629=>"101011101",
  18630=>"001100101",
  18631=>"001110100",
  18632=>"101111001",
  18633=>"011000110",
  18634=>"011001011",
  18635=>"010000100",
  18636=>"010010110",
  18637=>"110010000",
  18638=>"010101010",
  18639=>"100101101",
  18640=>"110010000",
  18641=>"000100110",
  18642=>"000010110",
  18643=>"101010110",
  18644=>"000010000",
  18645=>"100000010",
  18646=>"010100010",
  18647=>"001100011",
  18648=>"001101001",
  18649=>"111001011",
  18650=>"011000101",
  18651=>"100101011",
  18652=>"101111100",
  18653=>"000011100",
  18654=>"010010000",
  18655=>"110100100",
  18656=>"000111111",
  18657=>"010000101",
  18658=>"010000011",
  18659=>"111000100",
  18660=>"000110100",
  18661=>"110111100",
  18662=>"110101000",
  18663=>"110010110",
  18664=>"010111100",
  18665=>"110111100",
  18666=>"110110000",
  18667=>"111101110",
  18668=>"101110010",
  18669=>"111001000",
  18670=>"011001000",
  18671=>"001101001",
  18672=>"000100101",
  18673=>"000101111",
  18674=>"101101011",
  18675=>"011101000",
  18676=>"010001001",
  18677=>"000011001",
  18678=>"011110010",
  18679=>"010000001",
  18680=>"100000111",
  18681=>"001010000",
  18682=>"111001111",
  18683=>"000001001",
  18684=>"001111111",
  18685=>"001010100",
  18686=>"101100101",
  18687=>"110011110",
  18688=>"101101101",
  18689=>"111000010",
  18690=>"000111000",
  18691=>"111100110",
  18692=>"011110100",
  18693=>"101110110",
  18694=>"010100101",
  18695=>"110110010",
  18696=>"000110000",
  18697=>"111110011",
  18698=>"101110010",
  18699=>"001010110",
  18700=>"101110010",
  18701=>"001110000",
  18702=>"101110100",
  18703=>"001111001",
  18704=>"110100100",
  18705=>"011001000",
  18706=>"101100110",
  18707=>"101010110",
  18708=>"010001010",
  18709=>"010110000",
  18710=>"000111010",
  18711=>"010110000",
  18712=>"001011110",
  18713=>"111111100",
  18714=>"000011100",
  18715=>"001010001",
  18716=>"010000001",
  18717=>"010001110",
  18718=>"101000010",
  18719=>"000001010",
  18720=>"100101110",
  18721=>"001000011",
  18722=>"100001000",
  18723=>"010010001",
  18724=>"000011110",
  18725=>"010010110",
  18726=>"101111110",
  18727=>"000101010",
  18728=>"111011001",
  18729=>"001110011",
  18730=>"110010111",
  18731=>"111010010",
  18732=>"000111100",
  18733=>"010111101",
  18734=>"110000101",
  18735=>"101000001",
  18736=>"000101101",
  18737=>"101000001",
  18738=>"000001001",
  18739=>"011011010",
  18740=>"010000111",
  18741=>"000010111",
  18742=>"111101001",
  18743=>"000011111",
  18744=>"000011001",
  18745=>"100001001",
  18746=>"110010011",
  18747=>"100111000",
  18748=>"111110111",
  18749=>"101110111",
  18750=>"011101001",
  18751=>"001101000",
  18752=>"000110011",
  18753=>"011010110",
  18754=>"010001010",
  18755=>"110000110",
  18756=>"000111010",
  18757=>"000010100",
  18758=>"001001011",
  18759=>"111111100",
  18760=>"101100100",
  18761=>"110011100",
  18762=>"010000111",
  18763=>"000100111",
  18764=>"011010000",
  18765=>"011100101",
  18766=>"101111111",
  18767=>"101000100",
  18768=>"000110010",
  18769=>"000100100",
  18770=>"001111100",
  18771=>"010101111",
  18772=>"011011110",
  18773=>"010011000",
  18774=>"101011001",
  18775=>"001100110",
  18776=>"000101100",
  18777=>"100001010",
  18778=>"100000101",
  18779=>"010100110",
  18780=>"001001100",
  18781=>"001000111",
  18782=>"001111101",
  18783=>"011100000",
  18784=>"001000000",
  18785=>"111000100",
  18786=>"001100110",
  18787=>"101001111",
  18788=>"001100101",
  18789=>"111011110",
  18790=>"100010111",
  18791=>"111111100",
  18792=>"111110010",
  18793=>"000001000",
  18794=>"100011111",
  18795=>"101110010",
  18796=>"111110101",
  18797=>"011101010",
  18798=>"110100001",
  18799=>"100101111",
  18800=>"001110001",
  18801=>"000000011",
  18802=>"011010110",
  18803=>"110010010",
  18804=>"111011000",
  18805=>"010101111",
  18806=>"100111001",
  18807=>"100110001",
  18808=>"010011010",
  18809=>"001011011",
  18810=>"011100011",
  18811=>"000000011",
  18812=>"001001000",
  18813=>"110000001",
  18814=>"000011011",
  18815=>"010000101",
  18816=>"110110010",
  18817=>"000000001",
  18818=>"011100000",
  18819=>"111001000",
  18820=>"101110110",
  18821=>"001001101",
  18822=>"011100000",
  18823=>"011011010",
  18824=>"001001000",
  18825=>"111100000",
  18826=>"111111001",
  18827=>"101111110",
  18828=>"000100110",
  18829=>"101000100",
  18830=>"011001000",
  18831=>"110010111",
  18832=>"010100111",
  18833=>"000000011",
  18834=>"000000101",
  18835=>"100001000",
  18836=>"001010001",
  18837=>"111111001",
  18838=>"010110111",
  18839=>"111000100",
  18840=>"011110011",
  18841=>"010101101",
  18842=>"000110000",
  18843=>"100100011",
  18844=>"101101111",
  18845=>"111000011",
  18846=>"101011010",
  18847=>"001010110",
  18848=>"100000010",
  18849=>"001010010",
  18850=>"111110010",
  18851=>"011100110",
  18852=>"111001011",
  18853=>"011000110",
  18854=>"111101001",
  18855=>"110000111",
  18856=>"110110101",
  18857=>"100001100",
  18858=>"010010111",
  18859=>"010110000",
  18860=>"101001000",
  18861=>"010111011",
  18862=>"111110111",
  18863=>"110100010",
  18864=>"000100111",
  18865=>"100010010",
  18866=>"001111111",
  18867=>"000000001",
  18868=>"111001011",
  18869=>"000000000",
  18870=>"010000101",
  18871=>"011111100",
  18872=>"111010110",
  18873=>"010100110",
  18874=>"001111110",
  18875=>"101110110",
  18876=>"111011110",
  18877=>"001111110",
  18878=>"111110111",
  18879=>"001111101",
  18880=>"010011001",
  18881=>"000101101",
  18882=>"100000100",
  18883=>"101010100",
  18884=>"000011000",
  18885=>"001010000",
  18886=>"011110011",
  18887=>"000000010",
  18888=>"001001000",
  18889=>"110000111",
  18890=>"011000001",
  18891=>"001011110",
  18892=>"101111101",
  18893=>"000101000",
  18894=>"000001111",
  18895=>"110100010",
  18896=>"010110100",
  18897=>"111010010",
  18898=>"011110100",
  18899=>"011000010",
  18900=>"011011110",
  18901=>"000000111",
  18902=>"110010110",
  18903=>"010101110",
  18904=>"100100000",
  18905=>"011001000",
  18906=>"101101011",
  18907=>"110000001",
  18908=>"001001000",
  18909=>"111010110",
  18910=>"110101100",
  18911=>"100100011",
  18912=>"000010011",
  18913=>"111110100",
  18914=>"101110001",
  18915=>"101101111",
  18916=>"011100010",
  18917=>"111111000",
  18918=>"011001110",
  18919=>"001110011",
  18920=>"101100001",
  18921=>"010100001",
  18922=>"001100000",
  18923=>"001101100",
  18924=>"000010000",
  18925=>"000101001",
  18926=>"110111110",
  18927=>"100101011",
  18928=>"010001100",
  18929=>"100100101",
  18930=>"011001111",
  18931=>"101001111",
  18932=>"010010101",
  18933=>"101110111",
  18934=>"011001010",
  18935=>"101110100",
  18936=>"101001110",
  18937=>"000111110",
  18938=>"011010010",
  18939=>"011011101",
  18940=>"111101111",
  18941=>"001010000",
  18942=>"101000011",
  18943=>"111100000",
  18944=>"000001011",
  18945=>"101001000",
  18946=>"111001101",
  18947=>"011100101",
  18948=>"111001110",
  18949=>"010010010",
  18950=>"111100110",
  18951=>"111110101",
  18952=>"101101010",
  18953=>"000100110",
  18954=>"101001100",
  18955=>"110100001",
  18956=>"011010110",
  18957=>"100110111",
  18958=>"001011000",
  18959=>"110111101",
  18960=>"100010010",
  18961=>"111100111",
  18962=>"010011111",
  18963=>"100100110",
  18964=>"011001011",
  18965=>"100011011",
  18966=>"110010111",
  18967=>"010001000",
  18968=>"110010110",
  18969=>"001011010",
  18970=>"100001000",
  18971=>"000000011",
  18972=>"001010011",
  18973=>"111101000",
  18974=>"111111100",
  18975=>"111110111",
  18976=>"010011111",
  18977=>"011100001",
  18978=>"010001101",
  18979=>"111000100",
  18980=>"001010001",
  18981=>"110100110",
  18982=>"111000011",
  18983=>"001010111",
  18984=>"011001110",
  18985=>"110001100",
  18986=>"010010001",
  18987=>"010110100",
  18988=>"010111110",
  18989=>"110101100",
  18990=>"001100010",
  18991=>"000011100",
  18992=>"100111001",
  18993=>"101100000",
  18994=>"001000111",
  18995=>"010100101",
  18996=>"100110101",
  18997=>"111110101",
  18998=>"100110101",
  18999=>"001011011",
  19000=>"100111111",
  19001=>"111000101",
  19002=>"000100010",
  19003=>"001010010",
  19004=>"001100011",
  19005=>"001000000",
  19006=>"111111111",
  19007=>"100101101",
  19008=>"001011110",
  19009=>"010001001",
  19010=>"010100011",
  19011=>"001000111",
  19012=>"000000111",
  19013=>"001101000",
  19014=>"111110111",
  19015=>"100101110",
  19016=>"001110110",
  19017=>"011100101",
  19018=>"011111100",
  19019=>"001110101",
  19020=>"100110011",
  19021=>"001001000",
  19022=>"101010011",
  19023=>"011000101",
  19024=>"110100011",
  19025=>"011111010",
  19026=>"100001010",
  19027=>"000001101",
  19028=>"110000011",
  19029=>"000001101",
  19030=>"110111101",
  19031=>"010010000",
  19032=>"100000111",
  19033=>"110101011",
  19034=>"111101011",
  19035=>"100111100",
  19036=>"001011001",
  19037=>"101101001",
  19038=>"000101011",
  19039=>"111000101",
  19040=>"110111001",
  19041=>"010001111",
  19042=>"011011111",
  19043=>"011111011",
  19044=>"100001111",
  19045=>"000010110",
  19046=>"010010011",
  19047=>"111000011",
  19048=>"000000111",
  19049=>"111110011",
  19050=>"110001110",
  19051=>"010101000",
  19052=>"100111011",
  19053=>"011101110",
  19054=>"100011001",
  19055=>"100010000",
  19056=>"111110000",
  19057=>"100000000",
  19058=>"100101101",
  19059=>"010001100",
  19060=>"001101100",
  19061=>"010010100",
  19062=>"101100111",
  19063=>"001100011",
  19064=>"010011110",
  19065=>"110000111",
  19066=>"000110111",
  19067=>"011100101",
  19068=>"101110011",
  19069=>"110011111",
  19070=>"100111000",
  19071=>"000010010",
  19072=>"110111101",
  19073=>"010011001",
  19074=>"001010101",
  19075=>"101000010",
  19076=>"100101100",
  19077=>"000100100",
  19078=>"111110110",
  19079=>"000011111",
  19080=>"001110011",
  19081=>"110000100",
  19082=>"110010010",
  19083=>"100111000",
  19084=>"111111111",
  19085=>"001000001",
  19086=>"001101011",
  19087=>"100001010",
  19088=>"110011111",
  19089=>"001111001",
  19090=>"001011000",
  19091=>"000111101",
  19092=>"011110011",
  19093=>"001111111",
  19094=>"111110100",
  19095=>"100101001",
  19096=>"000001100",
  19097=>"101010100",
  19098=>"000011000",
  19099=>"000011110",
  19100=>"001111010",
  19101=>"111111001",
  19102=>"000011010",
  19103=>"111000101",
  19104=>"111100110",
  19105=>"000001101",
  19106=>"000000110",
  19107=>"101110011",
  19108=>"011111110",
  19109=>"100000101",
  19110=>"001001011",
  19111=>"110011100",
  19112=>"101001100",
  19113=>"000101001",
  19114=>"010100000",
  19115=>"011101011",
  19116=>"100001001",
  19117=>"010001011",
  19118=>"100111000",
  19119=>"101101000",
  19120=>"100000100",
  19121=>"010000000",
  19122=>"000001110",
  19123=>"101111000",
  19124=>"111101000",
  19125=>"100110001",
  19126=>"100010010",
  19127=>"001100001",
  19128=>"001010110",
  19129=>"110010100",
  19130=>"001000100",
  19131=>"011111110",
  19132=>"110111010",
  19133=>"010111000",
  19134=>"010111000",
  19135=>"110011011",
  19136=>"010101100",
  19137=>"111101001",
  19138=>"000110000",
  19139=>"001101011",
  19140=>"010101001",
  19141=>"110100110",
  19142=>"001001000",
  19143=>"100110101",
  19144=>"000010010",
  19145=>"110111011",
  19146=>"010010101",
  19147=>"101010101",
  19148=>"000010111",
  19149=>"010010000",
  19150=>"110001001",
  19151=>"001000010",
  19152=>"001101011",
  19153=>"101001001",
  19154=>"011100110",
  19155=>"111011010",
  19156=>"100001101",
  19157=>"000000001",
  19158=>"010010110",
  19159=>"111000000",
  19160=>"010111100",
  19161=>"100001101",
  19162=>"100111111",
  19163=>"100101011",
  19164=>"110110110",
  19165=>"101001101",
  19166=>"110001100",
  19167=>"000011010",
  19168=>"100111100",
  19169=>"000100000",
  19170=>"111001011",
  19171=>"001010110",
  19172=>"100111010",
  19173=>"011111011",
  19174=>"011010100",
  19175=>"000001000",
  19176=>"001111000",
  19177=>"111111110",
  19178=>"101000000",
  19179=>"111000110",
  19180=>"010101001",
  19181=>"100001100",
  19182=>"001101000",
  19183=>"101010101",
  19184=>"111011111",
  19185=>"000101000",
  19186=>"111000000",
  19187=>"101000010",
  19188=>"101111100",
  19189=>"110001010",
  19190=>"011101010",
  19191=>"100111110",
  19192=>"011000100",
  19193=>"110111100",
  19194=>"110110111",
  19195=>"000101100",
  19196=>"001010110",
  19197=>"001110111",
  19198=>"111001100",
  19199=>"000110000",
  19200=>"011000110",
  19201=>"011001000",
  19202=>"000111001",
  19203=>"111101111",
  19204=>"001010010",
  19205=>"110000110",
  19206=>"000101100",
  19207=>"111110001",
  19208=>"101110110",
  19209=>"100100101",
  19210=>"100110000",
  19211=>"111101000",
  19212=>"001011000",
  19213=>"101001100",
  19214=>"011000101",
  19215=>"001010011",
  19216=>"010011110",
  19217=>"110111000",
  19218=>"100000111",
  19219=>"101100101",
  19220=>"101111101",
  19221=>"110110101",
  19222=>"011001111",
  19223=>"010010010",
  19224=>"101101110",
  19225=>"110010011",
  19226=>"000000110",
  19227=>"111000010",
  19228=>"101000110",
  19229=>"110100010",
  19230=>"100011100",
  19231=>"010011011",
  19232=>"000000010",
  19233=>"111010010",
  19234=>"001000010",
  19235=>"100001010",
  19236=>"000010100",
  19237=>"001001010",
  19238=>"100000111",
  19239=>"001101111",
  19240=>"101100111",
  19241=>"101101101",
  19242=>"101111001",
  19243=>"010010001",
  19244=>"100001101",
  19245=>"010011110",
  19246=>"000000011",
  19247=>"100001110",
  19248=>"000010101",
  19249=>"010100001",
  19250=>"001001100",
  19251=>"111100110",
  19252=>"001111001",
  19253=>"010001010",
  19254=>"010100111",
  19255=>"011010111",
  19256=>"010010000",
  19257=>"010001111",
  19258=>"011001111",
  19259=>"100111011",
  19260=>"000011001",
  19261=>"010101110",
  19262=>"001110001",
  19263=>"011001001",
  19264=>"111110010",
  19265=>"000010010",
  19266=>"111110011",
  19267=>"010011100",
  19268=>"010111100",
  19269=>"000100011",
  19270=>"111111100",
  19271=>"000100100",
  19272=>"010001011",
  19273=>"000010100",
  19274=>"110110000",
  19275=>"101101101",
  19276=>"111001100",
  19277=>"000010111",
  19278=>"100010101",
  19279=>"100010101",
  19280=>"101100010",
  19281=>"101101101",
  19282=>"001011101",
  19283=>"101011010",
  19284=>"101000110",
  19285=>"111010011",
  19286=>"111101010",
  19287=>"111001011",
  19288=>"001010001",
  19289=>"011000010",
  19290=>"110011101",
  19291=>"000001111",
  19292=>"011100101",
  19293=>"110000111",
  19294=>"011100011",
  19295=>"000100000",
  19296=>"101010011",
  19297=>"001010001",
  19298=>"110000101",
  19299=>"010110011",
  19300=>"101110111",
  19301=>"010100100",
  19302=>"011011000",
  19303=>"000000111",
  19304=>"001000101",
  19305=>"001101001",
  19306=>"000010110",
  19307=>"000010001",
  19308=>"110010001",
  19309=>"111011101",
  19310=>"101011010",
  19311=>"100100010",
  19312=>"011110000",
  19313=>"011100011",
  19314=>"110111011",
  19315=>"010010100",
  19316=>"000111110",
  19317=>"101001111",
  19318=>"100101111",
  19319=>"011000110",
  19320=>"000100111",
  19321=>"000100001",
  19322=>"101000010",
  19323=>"100011001",
  19324=>"010000000",
  19325=>"101111000",
  19326=>"100010000",
  19327=>"000010110",
  19328=>"000000000",
  19329=>"011110010",
  19330=>"100001000",
  19331=>"000111101",
  19332=>"000110111",
  19333=>"111110110",
  19334=>"100010010",
  19335=>"101111010",
  19336=>"001011101",
  19337=>"101101111",
  19338=>"110000101",
  19339=>"111011000",
  19340=>"110110001",
  19341=>"111111110",
  19342=>"001001101",
  19343=>"101001010",
  19344=>"010011000",
  19345=>"111001011",
  19346=>"100001101",
  19347=>"111100110",
  19348=>"011100110",
  19349=>"011000010",
  19350=>"111100011",
  19351=>"100111000",
  19352=>"100101110",
  19353=>"011111001",
  19354=>"110001100",
  19355=>"110100101",
  19356=>"100100111",
  19357=>"111111100",
  19358=>"110000001",
  19359=>"000100010",
  19360=>"000100111",
  19361=>"111111110",
  19362=>"011111000",
  19363=>"001100000",
  19364=>"000010001",
  19365=>"111011110",
  19366=>"110101100",
  19367=>"100001010",
  19368=>"110110001",
  19369=>"011001101",
  19370=>"010010111",
  19371=>"001001110",
  19372=>"111110011",
  19373=>"000101100",
  19374=>"000010101",
  19375=>"010001110",
  19376=>"001100100",
  19377=>"101000011",
  19378=>"101100001",
  19379=>"001001001",
  19380=>"100110011",
  19381=>"000000000",
  19382=>"111001010",
  19383=>"111101111",
  19384=>"011111100",
  19385=>"101101000",
  19386=>"011111001",
  19387=>"101000010",
  19388=>"000001011",
  19389=>"000011100",
  19390=>"000011111",
  19391=>"001001111",
  19392=>"011000001",
  19393=>"000101011",
  19394=>"001000111",
  19395=>"100100000",
  19396=>"111111110",
  19397=>"111001110",
  19398=>"101000011",
  19399=>"000101011",
  19400=>"110100110",
  19401=>"001001001",
  19402=>"000011110",
  19403=>"110111110",
  19404=>"100011000",
  19405=>"101000100",
  19406=>"111101011",
  19407=>"110011001",
  19408=>"100110110",
  19409=>"100001100",
  19410=>"101100101",
  19411=>"111000100",
  19412=>"000001000",
  19413=>"100110001",
  19414=>"000001000",
  19415=>"001001101",
  19416=>"101111111",
  19417=>"010100011",
  19418=>"011111001",
  19419=>"001110110",
  19420=>"101101100",
  19421=>"001100111",
  19422=>"111111111",
  19423=>"111111111",
  19424=>"001000000",
  19425=>"001001111",
  19426=>"111110001",
  19427=>"000100101",
  19428=>"101011100",
  19429=>"101001101",
  19430=>"101101100",
  19431=>"000010010",
  19432=>"111010111",
  19433=>"001101111",
  19434=>"010000000",
  19435=>"100000001",
  19436=>"100011101",
  19437=>"111111000",
  19438=>"111010010",
  19439=>"000001000",
  19440=>"001011011",
  19441=>"110011110",
  19442=>"101111011",
  19443=>"100000001",
  19444=>"100101100",
  19445=>"000000100",
  19446=>"001001101",
  19447=>"110110000",
  19448=>"100000001",
  19449=>"100111101",
  19450=>"110001100",
  19451=>"101000100",
  19452=>"111001000",
  19453=>"010101010",
  19454=>"000001111",
  19455=>"100101110",
  19456=>"000000000",
  19457=>"111011000",
  19458=>"010100001",
  19459=>"110100011",
  19460=>"010111010",
  19461=>"001100101",
  19462=>"001101111",
  19463=>"100010011",
  19464=>"111001100",
  19465=>"001100100",
  19466=>"111000111",
  19467=>"101101000",
  19468=>"010100000",
  19469=>"100110001",
  19470=>"010110110",
  19471=>"101111101",
  19472=>"110000111",
  19473=>"001111111",
  19474=>"111101110",
  19475=>"000001010",
  19476=>"111111010",
  19477=>"011000000",
  19478=>"010001011",
  19479=>"101110000",
  19480=>"100010001",
  19481=>"111011010",
  19482=>"001010001",
  19483=>"000111101",
  19484=>"001110110",
  19485=>"001110010",
  19486=>"110000110",
  19487=>"011001111",
  19488=>"001011000",
  19489=>"110100110",
  19490=>"000110010",
  19491=>"110110110",
  19492=>"010101000",
  19493=>"010100000",
  19494=>"011110101",
  19495=>"001001000",
  19496=>"000011011",
  19497=>"000010101",
  19498=>"000000101",
  19499=>"110111111",
  19500=>"100000101",
  19501=>"110110100",
  19502=>"001110100",
  19503=>"111100010",
  19504=>"101100000",
  19505=>"110000111",
  19506=>"011001001",
  19507=>"100001111",
  19508=>"001001001",
  19509=>"001100100",
  19510=>"011000000",
  19511=>"001000100",
  19512=>"101110011",
  19513=>"101001010",
  19514=>"000100001",
  19515=>"100111011",
  19516=>"000001010",
  19517=>"101100000",
  19518=>"110000110",
  19519=>"001010010",
  19520=>"010000001",
  19521=>"001000110",
  19522=>"100011000",
  19523=>"001110100",
  19524=>"000111101",
  19525=>"110011011",
  19526=>"011000010",
  19527=>"110110101",
  19528=>"000111000",
  19529=>"110011001",
  19530=>"001010000",
  19531=>"010101101",
  19532=>"001100100",
  19533=>"110100101",
  19534=>"110101000",
  19535=>"001101000",
  19536=>"001000110",
  19537=>"101101100",
  19538=>"111011110",
  19539=>"101100100",
  19540=>"000101001",
  19541=>"000001101",
  19542=>"110110111",
  19543=>"000100011",
  19544=>"100100010",
  19545=>"111010011",
  19546=>"001011110",
  19547=>"010010011",
  19548=>"010001111",
  19549=>"010011110",
  19550=>"000000111",
  19551=>"010110000",
  19552=>"000101110",
  19553=>"000011100",
  19554=>"011000010",
  19555=>"001100000",
  19556=>"111000001",
  19557=>"011011101",
  19558=>"011100000",
  19559=>"111101111",
  19560=>"100100011",
  19561=>"010011000",
  19562=>"001110111",
  19563=>"000100111",
  19564=>"000100111",
  19565=>"110000110",
  19566=>"100010000",
  19567=>"000001100",
  19568=>"000101011",
  19569=>"111100100",
  19570=>"001000111",
  19571=>"010110110",
  19572=>"100101001",
  19573=>"011101101",
  19574=>"111100111",
  19575=>"111101111",
  19576=>"111010011",
  19577=>"100100111",
  19578=>"110100000",
  19579=>"100100000",
  19580=>"011101010",
  19581=>"000001100",
  19582=>"101000110",
  19583=>"001000000",
  19584=>"010101100",
  19585=>"111110101",
  19586=>"010100011",
  19587=>"001101000",
  19588=>"111000001",
  19589=>"001011101",
  19590=>"111111010",
  19591=>"110010001",
  19592=>"000011010",
  19593=>"100000010",
  19594=>"000100011",
  19595=>"110000110",
  19596=>"110001110",
  19597=>"000001010",
  19598=>"001011000",
  19599=>"101011000",
  19600=>"110010001",
  19601=>"100111100",
  19602=>"100100110",
  19603=>"010010110",
  19604=>"100001101",
  19605=>"011000100",
  19606=>"000100111",
  19607=>"001010100",
  19608=>"010101010",
  19609=>"111011000",
  19610=>"001010011",
  19611=>"001001001",
  19612=>"010101100",
  19613=>"111101110",
  19614=>"101100111",
  19615=>"101111111",
  19616=>"000111011",
  19617=>"010000001",
  19618=>"000000111",
  19619=>"100011101",
  19620=>"110010100",
  19621=>"000111010",
  19622=>"110101110",
  19623=>"111100110",
  19624=>"000100000",
  19625=>"100010001",
  19626=>"000011100",
  19627=>"001000010",
  19628=>"111011011",
  19629=>"000111011",
  19630=>"011010110",
  19631=>"001111010",
  19632=>"000100000",
  19633=>"010111110",
  19634=>"110000100",
  19635=>"110111011",
  19636=>"100101100",
  19637=>"000010010",
  19638=>"111001101",
  19639=>"010000101",
  19640=>"001111111",
  19641=>"001110001",
  19642=>"011110101",
  19643=>"101001001",
  19644=>"010100010",
  19645=>"111000000",
  19646=>"000101110",
  19647=>"100000101",
  19648=>"100000110",
  19649=>"001100011",
  19650=>"010101001",
  19651=>"001110010",
  19652=>"110110111",
  19653=>"011100010",
  19654=>"101000001",
  19655=>"101111010",
  19656=>"100100100",
  19657=>"000101001",
  19658=>"010011000",
  19659=>"111100010",
  19660=>"000011001",
  19661=>"010100011",
  19662=>"110101101",
  19663=>"101000101",
  19664=>"100100001",
  19665=>"000010110",
  19666=>"001110010",
  19667=>"100100100",
  19668=>"010101100",
  19669=>"111011110",
  19670=>"000000101",
  19671=>"100101000",
  19672=>"110110110",
  19673=>"011110100",
  19674=>"011000011",
  19675=>"011001100",
  19676=>"101001000",
  19677=>"111110011",
  19678=>"000000011",
  19679=>"100100101",
  19680=>"000111000",
  19681=>"001001100",
  19682=>"101001000",
  19683=>"100011110",
  19684=>"110101111",
  19685=>"100111110",
  19686=>"010101010",
  19687=>"111011111",
  19688=>"000010110",
  19689=>"101110000",
  19690=>"100000101",
  19691=>"100010110",
  19692=>"010000001",
  19693=>"000001000",
  19694=>"001010101",
  19695=>"011010001",
  19696=>"101111110",
  19697=>"100001101",
  19698=>"011111000",
  19699=>"111000010",
  19700=>"011001100",
  19701=>"001011001",
  19702=>"110001010",
  19703=>"001000011",
  19704=>"000111000",
  19705=>"011011010",
  19706=>"010000110",
  19707=>"100000110",
  19708=>"001000111",
  19709=>"111110001",
  19710=>"000100011",
  19711=>"111110001",
  19712=>"111111111",
  19713=>"110001100",
  19714=>"101000000",
  19715=>"000000111",
  19716=>"000101101",
  19717=>"001110101",
  19718=>"001000101",
  19719=>"010111111",
  19720=>"100110100",
  19721=>"100100111",
  19722=>"001101011",
  19723=>"011110100",
  19724=>"011001011",
  19725=>"100010000",
  19726=>"110010001",
  19727=>"000101100",
  19728=>"011010011",
  19729=>"010101110",
  19730=>"000110101",
  19731=>"100111110",
  19732=>"000001000",
  19733=>"100100101",
  19734=>"100011010",
  19735=>"011111110",
  19736=>"101011000",
  19737=>"100110100",
  19738=>"000011000",
  19739=>"100100000",
  19740=>"011011011",
  19741=>"111000001",
  19742=>"110001011",
  19743=>"100001010",
  19744=>"100100001",
  19745=>"101110000",
  19746=>"110001110",
  19747=>"111010000",
  19748=>"010100010",
  19749=>"110011000",
  19750=>"110011011",
  19751=>"001011011",
  19752=>"001111110",
  19753=>"101001000",
  19754=>"101001001",
  19755=>"111111001",
  19756=>"000001001",
  19757=>"100100001",
  19758=>"110111101",
  19759=>"100011001",
  19760=>"101111111",
  19761=>"000110011",
  19762=>"110101100",
  19763=>"101001011",
  19764=>"100110010",
  19765=>"010011000",
  19766=>"100011111",
  19767=>"100001111",
  19768=>"000101010",
  19769=>"010001010",
  19770=>"010100010",
  19771=>"000100111",
  19772=>"110100001",
  19773=>"011110111",
  19774=>"110010111",
  19775=>"100010110",
  19776=>"100110010",
  19777=>"001100010",
  19778=>"001010100",
  19779=>"110011100",
  19780=>"000010011",
  19781=>"111011011",
  19782=>"001101100",
  19783=>"011000001",
  19784=>"010000010",
  19785=>"100001001",
  19786=>"100010001",
  19787=>"000111011",
  19788=>"011001000",
  19789=>"111111010",
  19790=>"010000101",
  19791=>"111110111",
  19792=>"000111010",
  19793=>"100010010",
  19794=>"000011111",
  19795=>"000110001",
  19796=>"100000001",
  19797=>"101110111",
  19798=>"010111010",
  19799=>"100001001",
  19800=>"111110011",
  19801=>"110100000",
  19802=>"111011101",
  19803=>"010000101",
  19804=>"111101111",
  19805=>"011011100",
  19806=>"110100011",
  19807=>"000001110",
  19808=>"101011010",
  19809=>"010100000",
  19810=>"110011011",
  19811=>"000001111",
  19812=>"000111110",
  19813=>"011101110",
  19814=>"010111101",
  19815=>"011000011",
  19816=>"011011101",
  19817=>"001001111",
  19818=>"110100011",
  19819=>"010011110",
  19820=>"001011100",
  19821=>"100011100",
  19822=>"111111010",
  19823=>"100001000",
  19824=>"001011111",
  19825=>"001111111",
  19826=>"000000000",
  19827=>"001101110",
  19828=>"000000000",
  19829=>"110011001",
  19830=>"110111110",
  19831=>"110010001",
  19832=>"101100011",
  19833=>"101111011",
  19834=>"000101101",
  19835=>"101011000",
  19836=>"101001000",
  19837=>"100001101",
  19838=>"010011001",
  19839=>"111000101",
  19840=>"111010000",
  19841=>"111111010",
  19842=>"100000000",
  19843=>"101111010",
  19844=>"000100111",
  19845=>"111011100",
  19846=>"110110100",
  19847=>"000110011",
  19848=>"010011011",
  19849=>"001000100",
  19850=>"110111100",
  19851=>"000100111",
  19852=>"101110010",
  19853=>"111101010",
  19854=>"100100001",
  19855=>"001001110",
  19856=>"000011010",
  19857=>"111101100",
  19858=>"001000110",
  19859=>"101001111",
  19860=>"111110011",
  19861=>"011111110",
  19862=>"111101110",
  19863=>"101011111",
  19864=>"010101101",
  19865=>"111110011",
  19866=>"011000011",
  19867=>"100011000",
  19868=>"001111000",
  19869=>"111010000",
  19870=>"001100110",
  19871=>"101111011",
  19872=>"100011111",
  19873=>"110001111",
  19874=>"001000010",
  19875=>"000111110",
  19876=>"100100100",
  19877=>"001000010",
  19878=>"100100101",
  19879=>"010011111",
  19880=>"101100111",
  19881=>"111001011",
  19882=>"111111001",
  19883=>"010110111",
  19884=>"110101010",
  19885=>"111111111",
  19886=>"101001101",
  19887=>"110111101",
  19888=>"100100110",
  19889=>"011110100",
  19890=>"000100111",
  19891=>"001000010",
  19892=>"100101101",
  19893=>"111000111",
  19894=>"111110110",
  19895=>"101011010",
  19896=>"000101111",
  19897=>"101110000",
  19898=>"010011011",
  19899=>"000001000",
  19900=>"001110100",
  19901=>"101011110",
  19902=>"011110000",
  19903=>"011011010",
  19904=>"001000000",
  19905=>"111001010",
  19906=>"001100011",
  19907=>"010100010",
  19908=>"001001001",
  19909=>"111110000",
  19910=>"011010001",
  19911=>"101000000",
  19912=>"011000110",
  19913=>"111010101",
  19914=>"110010010",
  19915=>"000101011",
  19916=>"101100100",
  19917=>"100110101",
  19918=>"101111000",
  19919=>"001010100",
  19920=>"011011111",
  19921=>"101010001",
  19922=>"001001000",
  19923=>"000110010",
  19924=>"000100010",
  19925=>"100000101",
  19926=>"000111000",
  19927=>"100001001",
  19928=>"110100100",
  19929=>"001010110",
  19930=>"000100001",
  19931=>"010101010",
  19932=>"111100110",
  19933=>"000011011",
  19934=>"110100111",
  19935=>"000011011",
  19936=>"101101101",
  19937=>"110000101",
  19938=>"111001000",
  19939=>"011001111",
  19940=>"110000110",
  19941=>"011110101",
  19942=>"000010110",
  19943=>"111111100",
  19944=>"110000100",
  19945=>"010111000",
  19946=>"000001000",
  19947=>"101001001",
  19948=>"101001000",
  19949=>"101101100",
  19950=>"110011111",
  19951=>"000010011",
  19952=>"101010010",
  19953=>"101001100",
  19954=>"100000111",
  19955=>"001000001",
  19956=>"011100100",
  19957=>"111111100",
  19958=>"010000110",
  19959=>"101110000",
  19960=>"000110001",
  19961=>"101001000",
  19962=>"001001010",
  19963=>"101110111",
  19964=>"110011011",
  19965=>"110111111",
  19966=>"111000111",
  19967=>"011100011",
  19968=>"110111001",
  19969=>"100010110",
  19970=>"110110010",
  19971=>"010011000",
  19972=>"001001001",
  19973=>"110110010",
  19974=>"011101111",
  19975=>"111000101",
  19976=>"111001100",
  19977=>"001011110",
  19978=>"111001101",
  19979=>"000101000",
  19980=>"000101001",
  19981=>"000110011",
  19982=>"110100011",
  19983=>"100010000",
  19984=>"001111001",
  19985=>"110010100",
  19986=>"000101100",
  19987=>"110000101",
  19988=>"111000011",
  19989=>"000101010",
  19990=>"011111011",
  19991=>"011010111",
  19992=>"110100100",
  19993=>"000111010",
  19994=>"011101100",
  19995=>"100010100",
  19996=>"100000010",
  19997=>"001001001",
  19998=>"010010000",
  19999=>"011110010",
  20000=>"000100111",
  20001=>"001000001",
  20002=>"111111010",
  20003=>"100010010",
  20004=>"100010111",
  20005=>"001010110",
  20006=>"110100011",
  20007=>"011101110",
  20008=>"011101001",
  20009=>"101010010",
  20010=>"011011010",
  20011=>"100111101",
  20012=>"001001001",
  20013=>"011110110",
  20014=>"001000001",
  20015=>"010101111",
  20016=>"100000011",
  20017=>"001000110",
  20018=>"000000001",
  20019=>"100110011",
  20020=>"000011110",
  20021=>"010100000",
  20022=>"000110010",
  20023=>"110000101",
  20024=>"101000011",
  20025=>"011001111",
  20026=>"101000110",
  20027=>"111011111",
  20028=>"010100001",
  20029=>"000011100",
  20030=>"100001110",
  20031=>"110000000",
  20032=>"111011111",
  20033=>"011000011",
  20034=>"011101011",
  20035=>"011100001",
  20036=>"011110101",
  20037=>"001010001",
  20038=>"101111101",
  20039=>"000010101",
  20040=>"000110011",
  20041=>"111000000",
  20042=>"111111110",
  20043=>"101110110",
  20044=>"000010000",
  20045=>"010111000",
  20046=>"000101000",
  20047=>"100100110",
  20048=>"111000111",
  20049=>"000110110",
  20050=>"100000111",
  20051=>"011010010",
  20052=>"000011001",
  20053=>"100001011",
  20054=>"011110111",
  20055=>"111010101",
  20056=>"000100101",
  20057=>"111010100",
  20058=>"001110011",
  20059=>"000000000",
  20060=>"101110001",
  20061=>"000000110",
  20062=>"000011010",
  20063=>"101011111",
  20064=>"111111001",
  20065=>"001101001",
  20066=>"100000100",
  20067=>"011101100",
  20068=>"101011000",
  20069=>"100001101",
  20070=>"011000001",
  20071=>"111000111",
  20072=>"000101000",
  20073=>"010110101",
  20074=>"100001010",
  20075=>"001010010",
  20076=>"110111011",
  20077=>"111000010",
  20078=>"100110000",
  20079=>"011011011",
  20080=>"010111101",
  20081=>"101011000",
  20082=>"101001000",
  20083=>"101011000",
  20084=>"010011111",
  20085=>"000010010",
  20086=>"011010011",
  20087=>"100001010",
  20088=>"000110100",
  20089=>"001011000",
  20090=>"110010111",
  20091=>"100100010",
  20092=>"010111111",
  20093=>"011100000",
  20094=>"000010010",
  20095=>"110101111",
  20096=>"100001101",
  20097=>"100010011",
  20098=>"000011101",
  20099=>"101011010",
  20100=>"110101111",
  20101=>"001001000",
  20102=>"011001111",
  20103=>"111111111",
  20104=>"101011110",
  20105=>"000100111",
  20106=>"100010011",
  20107=>"000001010",
  20108=>"110000100",
  20109=>"010001111",
  20110=>"110101111",
  20111=>"111110100",
  20112=>"100011010",
  20113=>"010101100",
  20114=>"111001011",
  20115=>"111110011",
  20116=>"011111101",
  20117=>"001011000",
  20118=>"111011110",
  20119=>"011010101",
  20120=>"011000111",
  20121=>"100111110",
  20122=>"000010011",
  20123=>"100010010",
  20124=>"011000000",
  20125=>"100011001",
  20126=>"010001111",
  20127=>"101001110",
  20128=>"111111110",
  20129=>"101010000",
  20130=>"000010111",
  20131=>"011111100",
  20132=>"000110010",
  20133=>"011111110",
  20134=>"010000101",
  20135=>"010100101",
  20136=>"011010011",
  20137=>"111011101",
  20138=>"111101111",
  20139=>"000101101",
  20140=>"000010001",
  20141=>"111011001",
  20142=>"111101101",
  20143=>"010001010",
  20144=>"011101110",
  20145=>"111000111",
  20146=>"111111000",
  20147=>"000110111",
  20148=>"000100110",
  20149=>"100010011",
  20150=>"000101000",
  20151=>"011100000",
  20152=>"011111001",
  20153=>"000111010",
  20154=>"110010111",
  20155=>"011001010",
  20156=>"000100000",
  20157=>"101000000",
  20158=>"101011110",
  20159=>"010110011",
  20160=>"111111111",
  20161=>"101110100",
  20162=>"110011000",
  20163=>"100011001",
  20164=>"011111111",
  20165=>"110010010",
  20166=>"001111100",
  20167=>"101111010",
  20168=>"110001100",
  20169=>"010010110",
  20170=>"110100111",
  20171=>"010011101",
  20172=>"110000000",
  20173=>"101011000",
  20174=>"110000111",
  20175=>"111111011",
  20176=>"000000001",
  20177=>"001010000",
  20178=>"001010000",
  20179=>"010111001",
  20180=>"001000100",
  20181=>"010001011",
  20182=>"110111011",
  20183=>"111100010",
  20184=>"110111010",
  20185=>"101011111",
  20186=>"100010111",
  20187=>"000111100",
  20188=>"110110111",
  20189=>"111101101",
  20190=>"000100111",
  20191=>"000101100",
  20192=>"101111001",
  20193=>"101001110",
  20194=>"000111001",
  20195=>"100000010",
  20196=>"101001011",
  20197=>"100101011",
  20198=>"110111111",
  20199=>"001000100",
  20200=>"111110001",
  20201=>"001100010",
  20202=>"101100111",
  20203=>"110101010",
  20204=>"110111110",
  20205=>"101000110",
  20206=>"000011010",
  20207=>"000000110",
  20208=>"101100100",
  20209=>"110100000",
  20210=>"010011111",
  20211=>"111101101",
  20212=>"110011000",
  20213=>"111010001",
  20214=>"111111000",
  20215=>"010010011",
  20216=>"000011110",
  20217=>"000100100",
  20218=>"011000100",
  20219=>"000110101",
  20220=>"101100001",
  20221=>"011101001",
  20222=>"011100011",
  20223=>"110100000",
  20224=>"100000000",
  20225=>"101011001",
  20226=>"101110100",
  20227=>"100001110",
  20228=>"110010000",
  20229=>"100000110",
  20230=>"001100000",
  20231=>"111010010",
  20232=>"110111001",
  20233=>"110000010",
  20234=>"010010111",
  20235=>"101111110",
  20236=>"010110110",
  20237=>"010110000",
  20238=>"000000010",
  20239=>"101011100",
  20240=>"001101101",
  20241=>"001011000",
  20242=>"100001010",
  20243=>"101101110",
  20244=>"010001101",
  20245=>"111110101",
  20246=>"100011100",
  20247=>"100011111",
  20248=>"000101110",
  20249=>"010100011",
  20250=>"100101110",
  20251=>"111111011",
  20252=>"101100001",
  20253=>"001000101",
  20254=>"001111011",
  20255=>"001010111",
  20256=>"010011101",
  20257=>"111101001",
  20258=>"101111011",
  20259=>"000110010",
  20260=>"100010000",
  20261=>"100111101",
  20262=>"010011100",
  20263=>"111100010",
  20264=>"010110001",
  20265=>"111100001",
  20266=>"111010011",
  20267=>"010001110",
  20268=>"111010011",
  20269=>"111101011",
  20270=>"000010000",
  20271=>"000100010",
  20272=>"111110001",
  20273=>"100011001",
  20274=>"110110000",
  20275=>"111111000",
  20276=>"100001000",
  20277=>"111000101",
  20278=>"110000001",
  20279=>"011010110",
  20280=>"101011000",
  20281=>"011010101",
  20282=>"001001011",
  20283=>"011100010",
  20284=>"010000000",
  20285=>"100101010",
  20286=>"000100101",
  20287=>"110100110",
  20288=>"100011100",
  20289=>"100100001",
  20290=>"010110010",
  20291=>"000000100",
  20292=>"110100000",
  20293=>"010010111",
  20294=>"111101111",
  20295=>"001011010",
  20296=>"011100110",
  20297=>"001001100",
  20298=>"000011011",
  20299=>"100010100",
  20300=>"101100100",
  20301=>"001100010",
  20302=>"010100101",
  20303=>"100010011",
  20304=>"001101110",
  20305=>"011000111",
  20306=>"000001010",
  20307=>"010101111",
  20308=>"100000100",
  20309=>"100001110",
  20310=>"001111111",
  20311=>"111101010",
  20312=>"101010110",
  20313=>"101100110",
  20314=>"111001111",
  20315=>"110101110",
  20316=>"010101001",
  20317=>"111101110",
  20318=>"010000101",
  20319=>"000100110",
  20320=>"000010001",
  20321=>"000010010",
  20322=>"001111000",
  20323=>"101111011",
  20324=>"000101010",
  20325=>"101010101",
  20326=>"100011110",
  20327=>"110111010",
  20328=>"101010010",
  20329=>"010010111",
  20330=>"110111111",
  20331=>"111111101",
  20332=>"101000000",
  20333=>"100010101",
  20334=>"010111011",
  20335=>"101000100",
  20336=>"000110110",
  20337=>"101110001",
  20338=>"010111011",
  20339=>"110000110",
  20340=>"011010110",
  20341=>"010010110",
  20342=>"000010101",
  20343=>"010010010",
  20344=>"011001101",
  20345=>"100101111",
  20346=>"001101000",
  20347=>"100010000",
  20348=>"101101010",
  20349=>"111011010",
  20350=>"110011001",
  20351=>"000100111",
  20352=>"000111000",
  20353=>"000101101",
  20354=>"111100100",
  20355=>"110000001",
  20356=>"010110101",
  20357=>"101100001",
  20358=>"101101100",
  20359=>"010001000",
  20360=>"111010100",
  20361=>"011001101",
  20362=>"110100000",
  20363=>"110000001",
  20364=>"000011110",
  20365=>"110100100",
  20366=>"100000110",
  20367=>"100101010",
  20368=>"111000010",
  20369=>"011110010",
  20370=>"010000100",
  20371=>"110111010",
  20372=>"110011101",
  20373=>"010111111",
  20374=>"111000111",
  20375=>"001110111",
  20376=>"111010100",
  20377=>"011010100",
  20378=>"010010101",
  20379=>"001010010",
  20380=>"010110100",
  20381=>"010100111",
  20382=>"001101110",
  20383=>"011001001",
  20384=>"101101110",
  20385=>"011110111",
  20386=>"001100000",
  20387=>"011000001",
  20388=>"001101101",
  20389=>"110111011",
  20390=>"100000101",
  20391=>"000010011",
  20392=>"101010110",
  20393=>"101111110",
  20394=>"101111101",
  20395=>"000010100",
  20396=>"001001000",
  20397=>"110111101",
  20398=>"001111100",
  20399=>"001010111",
  20400=>"100001010",
  20401=>"101000101",
  20402=>"101001110",
  20403=>"000100101",
  20404=>"111011011",
  20405=>"011010101",
  20406=>"110001010",
  20407=>"111000011",
  20408=>"000001001",
  20409=>"010111110",
  20410=>"101001111",
  20411=>"010110000",
  20412=>"100000000",
  20413=>"010010010",
  20414=>"001010100",
  20415=>"000100011",
  20416=>"100101111",
  20417=>"000110001",
  20418=>"100110001",
  20419=>"101011010",
  20420=>"010011100",
  20421=>"111010110",
  20422=>"011100000",
  20423=>"011101111",
  20424=>"000101111",
  20425=>"110010001",
  20426=>"011001010",
  20427=>"111100101",
  20428=>"111000111",
  20429=>"110000010",
  20430=>"001010001",
  20431=>"001010100",
  20432=>"011111000",
  20433=>"111110111",
  20434=>"011101110",
  20435=>"101101100",
  20436=>"101111011",
  20437=>"000100000",
  20438=>"001100000",
  20439=>"111001111",
  20440=>"100001101",
  20441=>"111010001",
  20442=>"010110010",
  20443=>"010100011",
  20444=>"101000001",
  20445=>"010111011",
  20446=>"110000100",
  20447=>"100100110",
  20448=>"111101001",
  20449=>"100010110",
  20450=>"100001010",
  20451=>"101001001",
  20452=>"001100000",
  20453=>"001000101",
  20454=>"111100000",
  20455=>"100101111",
  20456=>"100100110",
  20457=>"101010001",
  20458=>"010010010",
  20459=>"101001011",
  20460=>"110011101",
  20461=>"000000010",
  20462=>"101010000",
  20463=>"110101010",
  20464=>"011111010",
  20465=>"000100010",
  20466=>"010001100",
  20467=>"001100000",
  20468=>"011011101",
  20469=>"100011010",
  20470=>"000111100",
  20471=>"100001011",
  20472=>"001100100",
  20473=>"111111100",
  20474=>"110110011",
  20475=>"100101011",
  20476=>"010101010",
  20477=>"001110011",
  20478=>"111111100",
  20479=>"001011011",
  20480=>"100001001",
  20481=>"000011000",
  20482=>"100111111",
  20483=>"110010001",
  20484=>"000100100",
  20485=>"111001100",
  20486=>"000010010",
  20487=>"100101111",
  20488=>"010101010",
  20489=>"000101100",
  20490=>"100100010",
  20491=>"010010101",
  20492=>"111100010",
  20493=>"000001111",
  20494=>"111000101",
  20495=>"110101011",
  20496=>"001000110",
  20497=>"011001110",
  20498=>"100111101",
  20499=>"111111000",
  20500=>"010001001",
  20501=>"110001110",
  20502=>"011000110",
  20503=>"101100010",
  20504=>"100000010",
  20505=>"110111110",
  20506=>"011101000",
  20507=>"000100111",
  20508=>"111000101",
  20509=>"001100111",
  20510=>"010101111",
  20511=>"011110001",
  20512=>"111010101",
  20513=>"010100001",
  20514=>"110100010",
  20515=>"001110101",
  20516=>"111101101",
  20517=>"101111001",
  20518=>"101101001",
  20519=>"101101111",
  20520=>"001001110",
  20521=>"111111000",
  20522=>"001100100",
  20523=>"010100111",
  20524=>"101101000",
  20525=>"011110000",
  20526=>"111111011",
  20527=>"100111111",
  20528=>"000111000",
  20529=>"001101011",
  20530=>"000100001",
  20531=>"111011110",
  20532=>"111001100",
  20533=>"110010011",
  20534=>"111100010",
  20535=>"101111011",
  20536=>"010011110",
  20537=>"101010001",
  20538=>"000000010",
  20539=>"100100011",
  20540=>"100000000",
  20541=>"001011001",
  20542=>"001100111",
  20543=>"111100000",
  20544=>"100010000",
  20545=>"010011100",
  20546=>"111111010",
  20547=>"011010110",
  20548=>"000101000",
  20549=>"000000010",
  20550=>"111101110",
  20551=>"101110010",
  20552=>"001000100",
  20553=>"010011010",
  20554=>"101110110",
  20555=>"101001010",
  20556=>"000110101",
  20557=>"100011110",
  20558=>"100000111",
  20559=>"110101000",
  20560=>"000001100",
  20561=>"101100000",
  20562=>"101111111",
  20563=>"011100010",
  20564=>"100110100",
  20565=>"100000001",
  20566=>"110010001",
  20567=>"011101000",
  20568=>"110011101",
  20569=>"001111000",
  20570=>"011000110",
  20571=>"000011011",
  20572=>"001011101",
  20573=>"101011111",
  20574=>"101010011",
  20575=>"001100111",
  20576=>"100000000",
  20577=>"001100100",
  20578=>"110110011",
  20579=>"000001010",
  20580=>"101100001",
  20581=>"101101110",
  20582=>"000111011",
  20583=>"111111100",
  20584=>"111001101",
  20585=>"111111010",
  20586=>"110111011",
  20587=>"001110011",
  20588=>"011100000",
  20589=>"000101101",
  20590=>"110100010",
  20591=>"100001010",
  20592=>"101001000",
  20593=>"000011001",
  20594=>"101111101",
  20595=>"111100001",
  20596=>"011101100",
  20597=>"111101101",
  20598=>"010011000",
  20599=>"011101010",
  20600=>"010110000",
  20601=>"010000001",
  20602=>"101110001",
  20603=>"010010001",
  20604=>"011101011",
  20605=>"101010101",
  20606=>"001101001",
  20607=>"010101100",
  20608=>"101011011",
  20609=>"000101100",
  20610=>"100000000",
  20611=>"011101000",
  20612=>"011011110",
  20613=>"010101110",
  20614=>"010100010",
  20615=>"111000010",
  20616=>"010011100",
  20617=>"101111101",
  20618=>"100000010",
  20619=>"111010000",
  20620=>"011101010",
  20621=>"110110111",
  20622=>"010001000",
  20623=>"111101011",
  20624=>"011111000",
  20625=>"000001010",
  20626=>"110111101",
  20627=>"011011111",
  20628=>"111110111",
  20629=>"110001010",
  20630=>"001010111",
  20631=>"010101011",
  20632=>"011111111",
  20633=>"101000101",
  20634=>"101110101",
  20635=>"000010011",
  20636=>"111100001",
  20637=>"000000111",
  20638=>"001100000",
  20639=>"110011101",
  20640=>"101111111",
  20641=>"110011010",
  20642=>"101100101",
  20643=>"100100011",
  20644=>"101000110",
  20645=>"100010111",
  20646=>"010100011",
  20647=>"010011000",
  20648=>"101000001",
  20649=>"011010010",
  20650=>"000110011",
  20651=>"000010001",
  20652=>"001011011",
  20653=>"011111110",
  20654=>"010101011",
  20655=>"011001111",
  20656=>"111101010",
  20657=>"011011110",
  20658=>"011100001",
  20659=>"001100010",
  20660=>"000101111",
  20661=>"101110001",
  20662=>"000011111",
  20663=>"001101001",
  20664=>"000100011",
  20665=>"100101100",
  20666=>"101100001",
  20667=>"101100100",
  20668=>"011010100",
  20669=>"000111001",
  20670=>"111000000",
  20671=>"101011001",
  20672=>"110000110",
  20673=>"001110101",
  20674=>"011111110",
  20675=>"100100110",
  20676=>"001001001",
  20677=>"001101010",
  20678=>"000110001",
  20679=>"000000110",
  20680=>"110010010",
  20681=>"100110010",
  20682=>"111011000",
  20683=>"011110000",
  20684=>"110000000",
  20685=>"110001101",
  20686=>"011001000",
  20687=>"001010111",
  20688=>"000100100",
  20689=>"111000011",
  20690=>"001110110",
  20691=>"001000010",
  20692=>"111111001",
  20693=>"111011010",
  20694=>"000001001",
  20695=>"011110000",
  20696=>"110101000",
  20697=>"110110011",
  20698=>"110000001",
  20699=>"111111101",
  20700=>"110001000",
  20701=>"001111100",
  20702=>"001100111",
  20703=>"010101100",
  20704=>"000110000",
  20705=>"011100000",
  20706=>"010011110",
  20707=>"110111100",
  20708=>"111100011",
  20709=>"111111011",
  20710=>"010001110",
  20711=>"001100010",
  20712=>"110100101",
  20713=>"001100110",
  20714=>"011101000",
  20715=>"011111011",
  20716=>"001110000",
  20717=>"011011011",
  20718=>"011000101",
  20719=>"001011100",
  20720=>"111010100",
  20721=>"000001010",
  20722=>"111101000",
  20723=>"101100100",
  20724=>"011100111",
  20725=>"110000010",
  20726=>"000111111",
  20727=>"011111111",
  20728=>"100001100",
  20729=>"011001111",
  20730=>"010111111",
  20731=>"000011100",
  20732=>"100100110",
  20733=>"010011001",
  20734=>"101011110",
  20735=>"001101101",
  20736=>"110001000",
  20737=>"001111100",
  20738=>"010000011",
  20739=>"111010111",
  20740=>"011110010",
  20741=>"010010100",
  20742=>"000101010",
  20743=>"000111001",
  20744=>"111000010",
  20745=>"111111100",
  20746=>"110001010",
  20747=>"001001110",
  20748=>"001010101",
  20749=>"100100000",
  20750=>"101011011",
  20751=>"000110110",
  20752=>"010101001",
  20753=>"000110000",
  20754=>"000100011",
  20755=>"111111011",
  20756=>"111100110",
  20757=>"000100100",
  20758=>"110100100",
  20759=>"111110100",
  20760=>"100010001",
  20761=>"100011110",
  20762=>"101111010",
  20763=>"101100101",
  20764=>"011001001",
  20765=>"010100000",
  20766=>"011110111",
  20767=>"101110000",
  20768=>"011011010",
  20769=>"101101101",
  20770=>"010101010",
  20771=>"001100000",
  20772=>"010100001",
  20773=>"000000010",
  20774=>"000010001",
  20775=>"100000000",
  20776=>"000111011",
  20777=>"001101011",
  20778=>"110100101",
  20779=>"011010111",
  20780=>"111000000",
  20781=>"111001101",
  20782=>"100101011",
  20783=>"000100011",
  20784=>"010111100",
  20785=>"010111001",
  20786=>"100100100",
  20787=>"010100111",
  20788=>"000100001",
  20789=>"000011111",
  20790=>"110100010",
  20791=>"111011100",
  20792=>"010101001",
  20793=>"101011111",
  20794=>"100010111",
  20795=>"101000001",
  20796=>"000100100",
  20797=>"101000101",
  20798=>"100101100",
  20799=>"011010010",
  20800=>"111101100",
  20801=>"100001111",
  20802=>"111110111",
  20803=>"111100001",
  20804=>"010000111",
  20805=>"000111001",
  20806=>"011011111",
  20807=>"011011001",
  20808=>"110011110",
  20809=>"001001000",
  20810=>"011100100",
  20811=>"011000110",
  20812=>"000000001",
  20813=>"010011011",
  20814=>"100111000",
  20815=>"111001110",
  20816=>"010110011",
  20817=>"001000100",
  20818=>"010010010",
  20819=>"011011100",
  20820=>"111100001",
  20821=>"011111111",
  20822=>"111010111",
  20823=>"000101011",
  20824=>"000111001",
  20825=>"100101000",
  20826=>"110000011",
  20827=>"000001110",
  20828=>"001000110",
  20829=>"001001101",
  20830=>"011101000",
  20831=>"110011011",
  20832=>"001111010",
  20833=>"011010110",
  20834=>"100100101",
  20835=>"000001101",
  20836=>"110111011",
  20837=>"100000010",
  20838=>"011101000",
  20839=>"010111100",
  20840=>"000100100",
  20841=>"010110010",
  20842=>"001001110",
  20843=>"001110100",
  20844=>"000101101",
  20845=>"001000100",
  20846=>"101110010",
  20847=>"011100011",
  20848=>"011011101",
  20849=>"100011011",
  20850=>"100110100",
  20851=>"110001111",
  20852=>"100100110",
  20853=>"111010101",
  20854=>"110011010",
  20855=>"011100111",
  20856=>"011010011",
  20857=>"010000011",
  20858=>"011110010",
  20859=>"110010100",
  20860=>"001100101",
  20861=>"110101011",
  20862=>"001100010",
  20863=>"010110001",
  20864=>"000000000",
  20865=>"000010101",
  20866=>"100101100",
  20867=>"001010011",
  20868=>"001111110",
  20869=>"001111110",
  20870=>"010001001",
  20871=>"000111100",
  20872=>"001101001",
  20873=>"111011001",
  20874=>"011110011",
  20875=>"110010111",
  20876=>"110111111",
  20877=>"000001011",
  20878=>"111010011",
  20879=>"111100100",
  20880=>"111010100",
  20881=>"010100010",
  20882=>"001011011",
  20883=>"110101111",
  20884=>"101011000",
  20885=>"111101110",
  20886=>"010001001",
  20887=>"000100000",
  20888=>"010000001",
  20889=>"110000111",
  20890=>"011100011",
  20891=>"100011100",
  20892=>"101001101",
  20893=>"010100000",
  20894=>"100100110",
  20895=>"100110100",
  20896=>"011011010",
  20897=>"000101110",
  20898=>"001111010",
  20899=>"000110110",
  20900=>"100100110",
  20901=>"111100010",
  20902=>"000001000",
  20903=>"011100000",
  20904=>"000111000",
  20905=>"110010101",
  20906=>"111011111",
  20907=>"010000011",
  20908=>"101101110",
  20909=>"010101011",
  20910=>"000000011",
  20911=>"000111101",
  20912=>"011011110",
  20913=>"001100111",
  20914=>"010101000",
  20915=>"110001011",
  20916=>"001011011",
  20917=>"010000010",
  20918=>"010010110",
  20919=>"001111010",
  20920=>"101101011",
  20921=>"001011110",
  20922=>"100110001",
  20923=>"011001011",
  20924=>"010101110",
  20925=>"010000000",
  20926=>"101010001",
  20927=>"011101001",
  20928=>"110010001",
  20929=>"111110101",
  20930=>"001110101",
  20931=>"010011011",
  20932=>"011000100",
  20933=>"110101010",
  20934=>"101000011",
  20935=>"000110101",
  20936=>"001001111",
  20937=>"101010011",
  20938=>"101100100",
  20939=>"010010001",
  20940=>"011011011",
  20941=>"010001111",
  20942=>"011111101",
  20943=>"001011100",
  20944=>"101001110",
  20945=>"011110011",
  20946=>"111010101",
  20947=>"110100101",
  20948=>"010011011",
  20949=>"000111101",
  20950=>"101011101",
  20951=>"110000010",
  20952=>"011111111",
  20953=>"100110100",
  20954=>"010010101",
  20955=>"010011001",
  20956=>"010011010",
  20957=>"101101010",
  20958=>"110011011",
  20959=>"001101001",
  20960=>"110000111",
  20961=>"010101101",
  20962=>"110111111",
  20963=>"000101100",
  20964=>"101001100",
  20965=>"100010110",
  20966=>"011110000",
  20967=>"110110101",
  20968=>"011111001",
  20969=>"010010011",
  20970=>"110010110",
  20971=>"110100111",
  20972=>"011001101",
  20973=>"110010000",
  20974=>"000001011",
  20975=>"000010011",
  20976=>"101110000",
  20977=>"101101100",
  20978=>"001010011",
  20979=>"101100011",
  20980=>"110000100",
  20981=>"100111110",
  20982=>"010000110",
  20983=>"100101101",
  20984=>"000001100",
  20985=>"010101101",
  20986=>"001010111",
  20987=>"010110101",
  20988=>"111101111",
  20989=>"001001011",
  20990=>"100010000",
  20991=>"010111111",
  20992=>"001111100",
  20993=>"001010101",
  20994=>"010010010",
  20995=>"001000101",
  20996=>"101100111",
  20997=>"100011101",
  20998=>"100011010",
  20999=>"010000000",
  21000=>"011000000",
  21001=>"100001110",
  21002=>"010011100",
  21003=>"000111011",
  21004=>"111110010",
  21005=>"110011101",
  21006=>"011001110",
  21007=>"011101000",
  21008=>"010111110",
  21009=>"111010000",
  21010=>"111100101",
  21011=>"000011011",
  21012=>"010001111",
  21013=>"011011011",
  21014=>"100101110",
  21015=>"110011101",
  21016=>"101000011",
  21017=>"110100101",
  21018=>"000100110",
  21019=>"000001101",
  21020=>"110110111",
  21021=>"111111111",
  21022=>"100111011",
  21023=>"110101001",
  21024=>"010111101",
  21025=>"101010111",
  21026=>"001010111",
  21027=>"111001000",
  21028=>"110000010",
  21029=>"000000000",
  21030=>"001011111",
  21031=>"000101010",
  21032=>"010111111",
  21033=>"000010010",
  21034=>"100110100",
  21035=>"110010111",
  21036=>"011011000",
  21037=>"001000000",
  21038=>"001010000",
  21039=>"010001100",
  21040=>"111111100",
  21041=>"000110110",
  21042=>"111000000",
  21043=>"000110011",
  21044=>"011011111",
  21045=>"010110101",
  21046=>"101010101",
  21047=>"101010111",
  21048=>"000000000",
  21049=>"000001110",
  21050=>"000001100",
  21051=>"101111011",
  21052=>"110101000",
  21053=>"001110110",
  21054=>"000100010",
  21055=>"001010010",
  21056=>"100000011",
  21057=>"010001101",
  21058=>"011011101",
  21059=>"010011011",
  21060=>"111110101",
  21061=>"011100000",
  21062=>"000111010",
  21063=>"000111001",
  21064=>"010011110",
  21065=>"011010001",
  21066=>"101001001",
  21067=>"011101101",
  21068=>"101001111",
  21069=>"101101100",
  21070=>"000001100",
  21071=>"010111110",
  21072=>"111010101",
  21073=>"110111011",
  21074=>"010001111",
  21075=>"001010001",
  21076=>"001110010",
  21077=>"111111111",
  21078=>"100111001",
  21079=>"101011110",
  21080=>"110111111",
  21081=>"100001111",
  21082=>"001110110",
  21083=>"101001000",
  21084=>"101000011",
  21085=>"111011110",
  21086=>"000011111",
  21087=>"010100111",
  21088=>"000101010",
  21089=>"001011111",
  21090=>"010101000",
  21091=>"001101000",
  21092=>"110011110",
  21093=>"101000001",
  21094=>"101100101",
  21095=>"101001001",
  21096=>"100110111",
  21097=>"111011010",
  21098=>"100011111",
  21099=>"100100010",
  21100=>"001111000",
  21101=>"011101000",
  21102=>"100111011",
  21103=>"011010000",
  21104=>"111100011",
  21105=>"000110010",
  21106=>"111000010",
  21107=>"111001100",
  21108=>"010000010",
  21109=>"101101111",
  21110=>"101010001",
  21111=>"101001011",
  21112=>"011010010",
  21113=>"101100001",
  21114=>"111001000",
  21115=>"101111101",
  21116=>"100001011",
  21117=>"000101110",
  21118=>"011100101",
  21119=>"011010110",
  21120=>"000100001",
  21121=>"011010101",
  21122=>"011100110",
  21123=>"000000001",
  21124=>"011011110",
  21125=>"111010111",
  21126=>"111111111",
  21127=>"001101110",
  21128=>"010111011",
  21129=>"110100010",
  21130=>"111011010",
  21131=>"111100101",
  21132=>"101010011",
  21133=>"010100001",
  21134=>"010001100",
  21135=>"000011101",
  21136=>"000111001",
  21137=>"000001000",
  21138=>"000011110",
  21139=>"010001100",
  21140=>"011011011",
  21141=>"000001100",
  21142=>"001001111",
  21143=>"000100000",
  21144=>"110110001",
  21145=>"111101110",
  21146=>"101111100",
  21147=>"001100111",
  21148=>"010010110",
  21149=>"001001011",
  21150=>"111000111",
  21151=>"100100001",
  21152=>"010011111",
  21153=>"111011010",
  21154=>"110111110",
  21155=>"010011101",
  21156=>"000001110",
  21157=>"100011010",
  21158=>"100111110",
  21159=>"001111111",
  21160=>"111010010",
  21161=>"011111110",
  21162=>"101010010",
  21163=>"110101000",
  21164=>"110000000",
  21165=>"111001001",
  21166=>"000001000",
  21167=>"011111001",
  21168=>"000101000",
  21169=>"100011100",
  21170=>"100011110",
  21171=>"111000111",
  21172=>"111110000",
  21173=>"000011000",
  21174=>"001111001",
  21175=>"011110110",
  21176=>"110110000",
  21177=>"111111110",
  21178=>"111110111",
  21179=>"000101111",
  21180=>"011010110",
  21181=>"000101000",
  21182=>"001011000",
  21183=>"010011001",
  21184=>"000111101",
  21185=>"110111110",
  21186=>"000110110",
  21187=>"110001000",
  21188=>"101110101",
  21189=>"011000111",
  21190=>"101110011",
  21191=>"101100111",
  21192=>"001001011",
  21193=>"001111011",
  21194=>"111001001",
  21195=>"001110101",
  21196=>"001001011",
  21197=>"100011000",
  21198=>"100110110",
  21199=>"101101011",
  21200=>"011110001",
  21201=>"111100100",
  21202=>"011110010",
  21203=>"011010011",
  21204=>"000001010",
  21205=>"000000000",
  21206=>"001110000",
  21207=>"100110111",
  21208=>"010000101",
  21209=>"010000011",
  21210=>"111100100",
  21211=>"101000000",
  21212=>"110101111",
  21213=>"110100111",
  21214=>"010001100",
  21215=>"010110100",
  21216=>"011010111",
  21217=>"000001001",
  21218=>"110101010",
  21219=>"011001010",
  21220=>"001011000",
  21221=>"100100000",
  21222=>"110011100",
  21223=>"101011110",
  21224=>"100001010",
  21225=>"110010101",
  21226=>"000111111",
  21227=>"110010111",
  21228=>"000110000",
  21229=>"010000010",
  21230=>"100001000",
  21231=>"100010101",
  21232=>"100111011",
  21233=>"101011011",
  21234=>"100010011",
  21235=>"101000001",
  21236=>"000101000",
  21237=>"000000011",
  21238=>"111100010",
  21239=>"100001101",
  21240=>"010110011",
  21241=>"010000001",
  21242=>"010100010",
  21243=>"111101111",
  21244=>"001100111",
  21245=>"111000011",
  21246=>"111010110",
  21247=>"100000001",
  21248=>"011111101",
  21249=>"110111111",
  21250=>"101010111",
  21251=>"011001111",
  21252=>"001100001",
  21253=>"010100111",
  21254=>"011111010",
  21255=>"010100101",
  21256=>"000111001",
  21257=>"000001010",
  21258=>"000010010",
  21259=>"100100001",
  21260=>"000000111",
  21261=>"000101110",
  21262=>"111000010",
  21263=>"100100110",
  21264=>"011111000",
  21265=>"000000010",
  21266=>"010001000",
  21267=>"110001110",
  21268=>"101101110",
  21269=>"101010111",
  21270=>"001001001",
  21271=>"111011011",
  21272=>"100110101",
  21273=>"011001111",
  21274=>"101101001",
  21275=>"010110010",
  21276=>"001011101",
  21277=>"100100110",
  21278=>"101001101",
  21279=>"000000001",
  21280=>"110001111",
  21281=>"001111000",
  21282=>"010110001",
  21283=>"111000111",
  21284=>"000011001",
  21285=>"011000110",
  21286=>"000010100",
  21287=>"000110000",
  21288=>"100110000",
  21289=>"000100010",
  21290=>"110011010",
  21291=>"110111001",
  21292=>"111100001",
  21293=>"010000100",
  21294=>"001001101",
  21295=>"110000001",
  21296=>"001111001",
  21297=>"010101000",
  21298=>"000110000",
  21299=>"011111111",
  21300=>"111111111",
  21301=>"011110010",
  21302=>"010011011",
  21303=>"011000001",
  21304=>"100111000",
  21305=>"000011101",
  21306=>"110111000",
  21307=>"111011100",
  21308=>"001100111",
  21309=>"110011101",
  21310=>"110101000",
  21311=>"100000101",
  21312=>"100110001",
  21313=>"111100110",
  21314=>"101111001",
  21315=>"111110111",
  21316=>"110011000",
  21317=>"001101111",
  21318=>"111001101",
  21319=>"100111100",
  21320=>"101111110",
  21321=>"111001011",
  21322=>"111110110",
  21323=>"000101000",
  21324=>"010011010",
  21325=>"101000011",
  21326=>"000010110",
  21327=>"000000011",
  21328=>"011010110",
  21329=>"010001101",
  21330=>"110000001",
  21331=>"101111111",
  21332=>"001110000",
  21333=>"111011111",
  21334=>"111001111",
  21335=>"000000100",
  21336=>"000110101",
  21337=>"001010110",
  21338=>"100011001",
  21339=>"001001101",
  21340=>"000011100",
  21341=>"001000101",
  21342=>"100001011",
  21343=>"111110011",
  21344=>"111011001",
  21345=>"011001000",
  21346=>"011111110",
  21347=>"010010011",
  21348=>"010101000",
  21349=>"111100111",
  21350=>"001101010",
  21351=>"011010000",
  21352=>"011000000",
  21353=>"010100101",
  21354=>"000010010",
  21355=>"101000011",
  21356=>"110101010",
  21357=>"010001110",
  21358=>"010010000",
  21359=>"100010010",
  21360=>"010101101",
  21361=>"100100101",
  21362=>"011001100",
  21363=>"111011011",
  21364=>"101101110",
  21365=>"010110100",
  21366=>"101000000",
  21367=>"101000010",
  21368=>"110010000",
  21369=>"101111010",
  21370=>"100111111",
  21371=>"110011010",
  21372=>"001001111",
  21373=>"101011000",
  21374=>"100110111",
  21375=>"101010110",
  21376=>"111110111",
  21377=>"001100111",
  21378=>"000100101",
  21379=>"001001010",
  21380=>"001110100",
  21381=>"111101001",
  21382=>"101001101",
  21383=>"011001010",
  21384=>"011110001",
  21385=>"011110010",
  21386=>"111110010",
  21387=>"110000011",
  21388=>"000100101",
  21389=>"111000011",
  21390=>"001110101",
  21391=>"100111110",
  21392=>"011110111",
  21393=>"111111111",
  21394=>"001110100",
  21395=>"001101000",
  21396=>"111010001",
  21397=>"111000100",
  21398=>"010001111",
  21399=>"000111001",
  21400=>"001101101",
  21401=>"001000000",
  21402=>"010111111",
  21403=>"101100000",
  21404=>"100100101",
  21405=>"001100100",
  21406=>"001100011",
  21407=>"101100011",
  21408=>"111010101",
  21409=>"011001010",
  21410=>"001101111",
  21411=>"111000001",
  21412=>"001110111",
  21413=>"011100000",
  21414=>"111011010",
  21415=>"001111000",
  21416=>"110100011",
  21417=>"000010011",
  21418=>"111101010",
  21419=>"101011000",
  21420=>"000110110",
  21421=>"010010000",
  21422=>"111000001",
  21423=>"010011000",
  21424=>"111111110",
  21425=>"111010100",
  21426=>"011110010",
  21427=>"101010011",
  21428=>"101000100",
  21429=>"100001001",
  21430=>"000100000",
  21431=>"101000001",
  21432=>"101110000",
  21433=>"001110000",
  21434=>"111100110",
  21435=>"111001011",
  21436=>"100000111",
  21437=>"110010001",
  21438=>"001100111",
  21439=>"111001001",
  21440=>"101101010",
  21441=>"000111001",
  21442=>"110100011",
  21443=>"101111001",
  21444=>"110011110",
  21445=>"111001011",
  21446=>"111111001",
  21447=>"011011111",
  21448=>"011101100",
  21449=>"010011011",
  21450=>"001111110",
  21451=>"001111011",
  21452=>"001101101",
  21453=>"110001010",
  21454=>"100101111",
  21455=>"000110100",
  21456=>"101001110",
  21457=>"011001001",
  21458=>"000111111",
  21459=>"110111111",
  21460=>"000011100",
  21461=>"001000111",
  21462=>"111001111",
  21463=>"001100100",
  21464=>"100111011",
  21465=>"111000111",
  21466=>"100110000",
  21467=>"001010101",
  21468=>"111111011",
  21469=>"011111011",
  21470=>"001000011",
  21471=>"000110111",
  21472=>"101111011",
  21473=>"010100101",
  21474=>"100100000",
  21475=>"011111101",
  21476=>"010101111",
  21477=>"010011101",
  21478=>"000011010",
  21479=>"101010000",
  21480=>"000000001",
  21481=>"110111100",
  21482=>"110111100",
  21483=>"011110010",
  21484=>"001101010",
  21485=>"111001100",
  21486=>"010001011",
  21487=>"111011110",
  21488=>"101111101",
  21489=>"000100010",
  21490=>"001110110",
  21491=>"100110011",
  21492=>"000110011",
  21493=>"010010000",
  21494=>"101110101",
  21495=>"111110110",
  21496=>"111000110",
  21497=>"011011100",
  21498=>"000011110",
  21499=>"011010100",
  21500=>"011101000",
  21501=>"001010111",
  21502=>"000111011",
  21503=>"111001111",
  21504=>"101100110",
  21505=>"110100111",
  21506=>"000110110",
  21507=>"010101100",
  21508=>"010101011",
  21509=>"000110010",
  21510=>"100000101",
  21511=>"000101100",
  21512=>"001000001",
  21513=>"011001000",
  21514=>"001010001",
  21515=>"101111110",
  21516=>"101100000",
  21517=>"011111100",
  21518=>"101011011",
  21519=>"100000101",
  21520=>"000100000",
  21521=>"010110110",
  21522=>"010011001",
  21523=>"100100101",
  21524=>"011010001",
  21525=>"101011011",
  21526=>"101100111",
  21527=>"011110000",
  21528=>"101101000",
  21529=>"101000000",
  21530=>"111111011",
  21531=>"101110111",
  21532=>"011011000",
  21533=>"010010000",
  21534=>"111001001",
  21535=>"010111000",
  21536=>"001000100",
  21537=>"110110101",
  21538=>"100010000",
  21539=>"011111010",
  21540=>"111100100",
  21541=>"110100011",
  21542=>"110110100",
  21543=>"010101011",
  21544=>"101101110",
  21545=>"010000000",
  21546=>"000111101",
  21547=>"001000010",
  21548=>"111111100",
  21549=>"100111011",
  21550=>"000001011",
  21551=>"011100100",
  21552=>"000001110",
  21553=>"010000001",
  21554=>"101010001",
  21555=>"111100000",
  21556=>"110001000",
  21557=>"110000011",
  21558=>"110111101",
  21559=>"000000110",
  21560=>"101100100",
  21561=>"000011010",
  21562=>"010100101",
  21563=>"001111001",
  21564=>"010010001",
  21565=>"001001001",
  21566=>"100100011",
  21567=>"111101100",
  21568=>"011010100",
  21569=>"111011101",
  21570=>"111100001",
  21571=>"000101101",
  21572=>"100011111",
  21573=>"111000111",
  21574=>"001101101",
  21575=>"110000001",
  21576=>"111000111",
  21577=>"000100100",
  21578=>"011000111",
  21579=>"101111110",
  21580=>"011110011",
  21581=>"010110101",
  21582=>"011111011",
  21583=>"000000000",
  21584=>"010001000",
  21585=>"111001111",
  21586=>"100011110",
  21587=>"011000111",
  21588=>"101000010",
  21589=>"100110110",
  21590=>"111111010",
  21591=>"101001110",
  21592=>"010110100",
  21593=>"000011011",
  21594=>"101011100",
  21595=>"101001010",
  21596=>"111111111",
  21597=>"100110000",
  21598=>"111011011",
  21599=>"011111000",
  21600=>"000100010",
  21601=>"010110011",
  21602=>"001001010",
  21603=>"000111011",
  21604=>"011000111",
  21605=>"001100010",
  21606=>"010011100",
  21607=>"010001111",
  21608=>"110110110",
  21609=>"100001111",
  21610=>"000101000",
  21611=>"001001100",
  21612=>"110011011",
  21613=>"100110101",
  21614=>"110111111",
  21615=>"000001000",
  21616=>"100101111",
  21617=>"010000001",
  21618=>"011011001",
  21619=>"001000110",
  21620=>"011011111",
  21621=>"100101101",
  21622=>"111110100",
  21623=>"111110101",
  21624=>"010000011",
  21625=>"110101000",
  21626=>"010100000",
  21627=>"110111010",
  21628=>"101000011",
  21629=>"001011001",
  21630=>"111111001",
  21631=>"000001010",
  21632=>"000000000",
  21633=>"010010011",
  21634=>"111011111",
  21635=>"010100110",
  21636=>"011001111",
  21637=>"110110101",
  21638=>"011101000",
  21639=>"011101100",
  21640=>"111101101",
  21641=>"111100011",
  21642=>"000000000",
  21643=>"000001010",
  21644=>"100101010",
  21645=>"100100111",
  21646=>"111010000",
  21647=>"001001110",
  21648=>"111110111",
  21649=>"110010110",
  21650=>"000001110",
  21651=>"101101110",
  21652=>"000001000",
  21653=>"100100001",
  21654=>"100111111",
  21655=>"010111001",
  21656=>"110011101",
  21657=>"101010001",
  21658=>"001110000",
  21659=>"100100101",
  21660=>"001110110",
  21661=>"111101100",
  21662=>"100001001",
  21663=>"010100100",
  21664=>"100000101",
  21665=>"010110011",
  21666=>"111101000",
  21667=>"000100100",
  21668=>"010000011",
  21669=>"110111001",
  21670=>"100100001",
  21671=>"100010000",
  21672=>"100001011",
  21673=>"101101111",
  21674=>"101110110",
  21675=>"000101111",
  21676=>"111001011",
  21677=>"001100111",
  21678=>"100111001",
  21679=>"100101110",
  21680=>"010011001",
  21681=>"000010011",
  21682=>"000010111",
  21683=>"000010000",
  21684=>"110110000",
  21685=>"000010000",
  21686=>"011100011",
  21687=>"110111011",
  21688=>"101111000",
  21689=>"011110000",
  21690=>"110111101",
  21691=>"100111000",
  21692=>"100011100",
  21693=>"000111100",
  21694=>"101101110",
  21695=>"011110100",
  21696=>"101001001",
  21697=>"001110000",
  21698=>"001011001",
  21699=>"011001110",
  21700=>"000000101",
  21701=>"011010101",
  21702=>"100001000",
  21703=>"101001100",
  21704=>"100001101",
  21705=>"101101101",
  21706=>"110101101",
  21707=>"011000000",
  21708=>"001000110",
  21709=>"010001101",
  21710=>"010111100",
  21711=>"011001001",
  21712=>"011000001",
  21713=>"111110110",
  21714=>"111011001",
  21715=>"001001101",
  21716=>"001100110",
  21717=>"100101011",
  21718=>"111110010",
  21719=>"011110100",
  21720=>"111000001",
  21721=>"011110100",
  21722=>"010010011",
  21723=>"100100111",
  21724=>"110111010",
  21725=>"100010100",
  21726=>"110101001",
  21727=>"010110000",
  21728=>"111000110",
  21729=>"001001101",
  21730=>"101111100",
  21731=>"111101000",
  21732=>"101000101",
  21733=>"011110101",
  21734=>"111110100",
  21735=>"110110111",
  21736=>"001011001",
  21737=>"001101000",
  21738=>"111100010",
  21739=>"111000001",
  21740=>"000111101",
  21741=>"010100001",
  21742=>"101101111",
  21743=>"111000111",
  21744=>"011001111",
  21745=>"000010111",
  21746=>"100000011",
  21747=>"110001001",
  21748=>"111000001",
  21749=>"101110000",
  21750=>"010101111",
  21751=>"111101111",
  21752=>"100110010",
  21753=>"011101110",
  21754=>"011110111",
  21755=>"100110100",
  21756=>"011101111",
  21757=>"011011010",
  21758=>"011001101",
  21759=>"100011010",
  21760=>"101111100",
  21761=>"100011110",
  21762=>"111101101",
  21763=>"000001010",
  21764=>"100001000",
  21765=>"010111000",
  21766=>"110101001",
  21767=>"111011001",
  21768=>"010000111",
  21769=>"101100010",
  21770=>"111011111",
  21771=>"101100100",
  21772=>"100000010",
  21773=>"000110100",
  21774=>"101110100",
  21775=>"101010000",
  21776=>"100011110",
  21777=>"000011011",
  21778=>"001001001",
  21779=>"111101111",
  21780=>"100001100",
  21781=>"001110110",
  21782=>"110001101",
  21783=>"110000110",
  21784=>"011110011",
  21785=>"001001101",
  21786=>"000000011",
  21787=>"110000011",
  21788=>"101010000",
  21789=>"111101101",
  21790=>"111100010",
  21791=>"011010111",
  21792=>"110001001",
  21793=>"100110000",
  21794=>"010110101",
  21795=>"101011010",
  21796=>"100100010",
  21797=>"001100000",
  21798=>"001111000",
  21799=>"111101000",
  21800=>"011010011",
  21801=>"011110110",
  21802=>"000100011",
  21803=>"001010000",
  21804=>"000111111",
  21805=>"100000000",
  21806=>"001101110",
  21807=>"010000010",
  21808=>"010001100",
  21809=>"000111000",
  21810=>"000001111",
  21811=>"001010111",
  21812=>"001000101",
  21813=>"100100011",
  21814=>"100101110",
  21815=>"111010000",
  21816=>"111001101",
  21817=>"110101100",
  21818=>"010111000",
  21819=>"001110000",
  21820=>"111100000",
  21821=>"101011010",
  21822=>"110100001",
  21823=>"011001100",
  21824=>"100001111",
  21825=>"100000111",
  21826=>"110111100",
  21827=>"010010011",
  21828=>"111111111",
  21829=>"100010011",
  21830=>"000001010",
  21831=>"111011000",
  21832=>"101010100",
  21833=>"101111100",
  21834=>"100010100",
  21835=>"000010000",
  21836=>"100111010",
  21837=>"010001111",
  21838=>"101100010",
  21839=>"000011101",
  21840=>"111110111",
  21841=>"100001001",
  21842=>"111111101",
  21843=>"110001100",
  21844=>"111000001",
  21845=>"011001110",
  21846=>"111100100",
  21847=>"011011001",
  21848=>"101010011",
  21849=>"010011101",
  21850=>"101111011",
  21851=>"101110000",
  21852=>"110011101",
  21853=>"011110101",
  21854=>"010000000",
  21855=>"011000010",
  21856=>"111101101",
  21857=>"111000111",
  21858=>"011001011",
  21859=>"101101000",
  21860=>"100001111",
  21861=>"000100110",
  21862=>"010001100",
  21863=>"111111111",
  21864=>"011010111",
  21865=>"110000101",
  21866=>"010101010",
  21867=>"011011010",
  21868=>"000100000",
  21869=>"000010001",
  21870=>"110011100",
  21871=>"111000001",
  21872=>"001111010",
  21873=>"111100000",
  21874=>"101010001",
  21875=>"001101101",
  21876=>"010111000",
  21877=>"111010010",
  21878=>"010001110",
  21879=>"100001101",
  21880=>"011111100",
  21881=>"101011111",
  21882=>"010000010",
  21883=>"011100100",
  21884=>"010111010",
  21885=>"100011110",
  21886=>"000011111",
  21887=>"000101011",
  21888=>"100011000",
  21889=>"000001110",
  21890=>"110111111",
  21891=>"010101101",
  21892=>"011011110",
  21893=>"001010010",
  21894=>"001011101",
  21895=>"010100001",
  21896=>"000110001",
  21897=>"100000110",
  21898=>"001011110",
  21899=>"001000100",
  21900=>"000001000",
  21901=>"000111110",
  21902=>"001111000",
  21903=>"100011010",
  21904=>"111011010",
  21905=>"110100010",
  21906=>"001001100",
  21907=>"110100001",
  21908=>"110000000",
  21909=>"010001110",
  21910=>"100000100",
  21911=>"101101010",
  21912=>"010100110",
  21913=>"000001000",
  21914=>"010111111",
  21915=>"010011100",
  21916=>"100011011",
  21917=>"100010110",
  21918=>"101110001",
  21919=>"110010110",
  21920=>"111110100",
  21921=>"111100101",
  21922=>"100101110",
  21923=>"000010110",
  21924=>"100100110",
  21925=>"101001110",
  21926=>"111110011",
  21927=>"001000110",
  21928=>"100001111",
  21929=>"100011110",
  21930=>"011001111",
  21931=>"111011011",
  21932=>"111011011",
  21933=>"001001111",
  21934=>"101100100",
  21935=>"000101000",
  21936=>"111010111",
  21937=>"110101011",
  21938=>"010011001",
  21939=>"010001011",
  21940=>"111100111",
  21941=>"101100101",
  21942=>"010010000",
  21943=>"000000110",
  21944=>"100000000",
  21945=>"001110000",
  21946=>"111000001",
  21947=>"010011001",
  21948=>"111010101",
  21949=>"010101101",
  21950=>"100000100",
  21951=>"111101011",
  21952=>"001011010",
  21953=>"001000001",
  21954=>"101111110",
  21955=>"101000001",
  21956=>"010010011",
  21957=>"111100111",
  21958=>"110100111",
  21959=>"101101110",
  21960=>"010000001",
  21961=>"010011010",
  21962=>"100000010",
  21963=>"101111001",
  21964=>"101001110",
  21965=>"110101001",
  21966=>"010101101",
  21967=>"001101001",
  21968=>"000110111",
  21969=>"011110101",
  21970=>"011000110",
  21971=>"001001110",
  21972=>"010011001",
  21973=>"001011111",
  21974=>"001011000",
  21975=>"010101101",
  21976=>"001011000",
  21977=>"101100010",
  21978=>"010100010",
  21979=>"111100110",
  21980=>"010110110",
  21981=>"100100000",
  21982=>"001101010",
  21983=>"001001101",
  21984=>"110110111",
  21985=>"110100111",
  21986=>"101101100",
  21987=>"110010101",
  21988=>"110110110",
  21989=>"010000101",
  21990=>"001111000",
  21991=>"011011100",
  21992=>"000111100",
  21993=>"011100111",
  21994=>"110001100",
  21995=>"011100111",
  21996=>"101011001",
  21997=>"000000000",
  21998=>"011000000",
  21999=>"000010001",
  22000=>"100001111",
  22001=>"010111100",
  22002=>"000000110",
  22003=>"100101000",
  22004=>"000010011",
  22005=>"001000110",
  22006=>"101000101",
  22007=>"000001001",
  22008=>"110111000",
  22009=>"110110101",
  22010=>"011110101",
  22011=>"101000110",
  22012=>"000010111",
  22013=>"100101111",
  22014=>"111100101",
  22015=>"110100010",
  22016=>"101001010",
  22017=>"010101000",
  22018=>"111010011",
  22019=>"100101011",
  22020=>"001000011",
  22021=>"000010011",
  22022=>"101011110",
  22023=>"010000100",
  22024=>"010110111",
  22025=>"011101110",
  22026=>"010100100",
  22027=>"010010000",
  22028=>"101101000",
  22029=>"000111100",
  22030=>"101100011",
  22031=>"000001110",
  22032=>"001101110",
  22033=>"111110101",
  22034=>"110100101",
  22035=>"111101010",
  22036=>"100011110",
  22037=>"100010010",
  22038=>"101010101",
  22039=>"100101101",
  22040=>"100100100",
  22041=>"110011111",
  22042=>"011010100",
  22043=>"001000100",
  22044=>"011001010",
  22045=>"111001011",
  22046=>"101100110",
  22047=>"100001100",
  22048=>"001000011",
  22049=>"110000001",
  22050=>"010000110",
  22051=>"101000001",
  22052=>"111011101",
  22053=>"101011100",
  22054=>"100011100",
  22055=>"000000101",
  22056=>"011000011",
  22057=>"011010110",
  22058=>"000010110",
  22059=>"010101110",
  22060=>"101011010",
  22061=>"000011100",
  22062=>"100100000",
  22063=>"110011101",
  22064=>"100010001",
  22065=>"110011111",
  22066=>"110000110",
  22067=>"110001101",
  22068=>"110110011",
  22069=>"110100011",
  22070=>"000011101",
  22071=>"000101010",
  22072=>"000011110",
  22073=>"111001101",
  22074=>"010100100",
  22075=>"100001001",
  22076=>"010011001",
  22077=>"010100000",
  22078=>"110010111",
  22079=>"001101010",
  22080=>"110110011",
  22081=>"110100010",
  22082=>"001011100",
  22083=>"001101000",
  22084=>"001110001",
  22085=>"111111100",
  22086=>"001001000",
  22087=>"100111101",
  22088=>"001000100",
  22089=>"110100010",
  22090=>"001000001",
  22091=>"100000001",
  22092=>"101010111",
  22093=>"011001101",
  22094=>"011111111",
  22095=>"100010001",
  22096=>"110111001",
  22097=>"001001000",
  22098=>"100110010",
  22099=>"100101011",
  22100=>"101110110",
  22101=>"011111010",
  22102=>"110100000",
  22103=>"111111101",
  22104=>"110001100",
  22105=>"101111100",
  22106=>"000101000",
  22107=>"011111111",
  22108=>"110000110",
  22109=>"111100000",
  22110=>"001011001",
  22111=>"111000101",
  22112=>"101110011",
  22113=>"101011111",
  22114=>"100010011",
  22115=>"100010111",
  22116=>"101001010",
  22117=>"100000011",
  22118=>"110000001",
  22119=>"110110000",
  22120=>"111110110",
  22121=>"000100011",
  22122=>"101011101",
  22123=>"000011110",
  22124=>"010110010",
  22125=>"010100111",
  22126=>"001011111",
  22127=>"010110111",
  22128=>"000110101",
  22129=>"111101010",
  22130=>"000101011",
  22131=>"010011110",
  22132=>"101111001",
  22133=>"101011100",
  22134=>"000111111",
  22135=>"000001010",
  22136=>"010011000",
  22137=>"111010011",
  22138=>"011100011",
  22139=>"000000001",
  22140=>"000001001",
  22141=>"011000010",
  22142=>"101100010",
  22143=>"001100010",
  22144=>"101101011",
  22145=>"101110100",
  22146=>"110010011",
  22147=>"010000001",
  22148=>"011111111",
  22149=>"101000011",
  22150=>"011110111",
  22151=>"001100000",
  22152=>"001110101",
  22153=>"100010000",
  22154=>"001001100",
  22155=>"010010000",
  22156=>"110000000",
  22157=>"101010010",
  22158=>"111110000",
  22159=>"101010100",
  22160=>"010101010",
  22161=>"010111011",
  22162=>"111110010",
  22163=>"110111101",
  22164=>"110010001",
  22165=>"110010001",
  22166=>"011001100",
  22167=>"001110000",
  22168=>"011001111",
  22169=>"100111111",
  22170=>"010111110",
  22171=>"011100111",
  22172=>"111011010",
  22173=>"000011110",
  22174=>"001101010",
  22175=>"110101010",
  22176=>"001001001",
  22177=>"000010010",
  22178=>"010011010",
  22179=>"111001110",
  22180=>"011110001",
  22181=>"001000010",
  22182=>"001001001",
  22183=>"110010110",
  22184=>"010101010",
  22185=>"111001001",
  22186=>"101100000",
  22187=>"101100101",
  22188=>"110110010",
  22189=>"100001010",
  22190=>"000011000",
  22191=>"101110100",
  22192=>"000000110",
  22193=>"111101010",
  22194=>"101001100",
  22195=>"000001001",
  22196=>"000110000",
  22197=>"001101000",
  22198=>"110110000",
  22199=>"111110011",
  22200=>"010100010",
  22201=>"011011100",
  22202=>"111010000",
  22203=>"001011001",
  22204=>"111101100",
  22205=>"001011000",
  22206=>"001000011",
  22207=>"110101000",
  22208=>"011111101",
  22209=>"001110011",
  22210=>"000110011",
  22211=>"001001110",
  22212=>"000111000",
  22213=>"100010110",
  22214=>"111011010",
  22215=>"111100011",
  22216=>"110001000",
  22217=>"111111100",
  22218=>"110101101",
  22219=>"001000000",
  22220=>"101000110",
  22221=>"011111100",
  22222=>"100001011",
  22223=>"111110010",
  22224=>"000010111",
  22225=>"101100011",
  22226=>"000100101",
  22227=>"011100100",
  22228=>"111111111",
  22229=>"110010111",
  22230=>"110110100",
  22231=>"001010010",
  22232=>"110011000",
  22233=>"110111111",
  22234=>"001101011",
  22235=>"110110010",
  22236=>"000101101",
  22237=>"100000000",
  22238=>"001001000",
  22239=>"100101000",
  22240=>"000010100",
  22241=>"100000111",
  22242=>"101101010",
  22243=>"101001111",
  22244=>"011010111",
  22245=>"111101001",
  22246=>"001101000",
  22247=>"011100100",
  22248=>"000111000",
  22249=>"010111111",
  22250=>"011001011",
  22251=>"111111111",
  22252=>"111000010",
  22253=>"100010010",
  22254=>"101110011",
  22255=>"111110111",
  22256=>"000111100",
  22257=>"100100111",
  22258=>"001110001",
  22259=>"001101101",
  22260=>"001010110",
  22261=>"110110000",
  22262=>"101111000",
  22263=>"000010100",
  22264=>"000011100",
  22265=>"011010101",
  22266=>"110011101",
  22267=>"001101111",
  22268=>"110110001",
  22269=>"000011101",
  22270=>"111001010",
  22271=>"011000010",
  22272=>"111011011",
  22273=>"101001011",
  22274=>"010001101",
  22275=>"111110100",
  22276=>"100101010",
  22277=>"111010110",
  22278=>"010001011",
  22279=>"001100010",
  22280=>"011011110",
  22281=>"000010010",
  22282=>"100100100",
  22283=>"001111010",
  22284=>"110011000",
  22285=>"000000111",
  22286=>"010000001",
  22287=>"011101110",
  22288=>"010100000",
  22289=>"100100100",
  22290=>"000001110",
  22291=>"000010110",
  22292=>"101111111",
  22293=>"001010111",
  22294=>"010011101",
  22295=>"111011101",
  22296=>"000000110",
  22297=>"000100011",
  22298=>"100100001",
  22299=>"000010111",
  22300=>"110010101",
  22301=>"111110001",
  22302=>"010101001",
  22303=>"000011001",
  22304=>"100101010",
  22305=>"111010110",
  22306=>"011101001",
  22307=>"110000101",
  22308=>"111100010",
  22309=>"100010010",
  22310=>"010011001",
  22311=>"101001101",
  22312=>"011110010",
  22313=>"000101111",
  22314=>"110010011",
  22315=>"111001010",
  22316=>"010100111",
  22317=>"000000000",
  22318=>"111000011",
  22319=>"110000011",
  22320=>"111100111",
  22321=>"110000110",
  22322=>"101001000",
  22323=>"111101111",
  22324=>"001100001",
  22325=>"010010011",
  22326=>"001000011",
  22327=>"111110110",
  22328=>"001101010",
  22329=>"100001010",
  22330=>"110111001",
  22331=>"011111111",
  22332=>"011110101",
  22333=>"110100101",
  22334=>"110011101",
  22335=>"101100010",
  22336=>"111000110",
  22337=>"111111110",
  22338=>"111101000",
  22339=>"011100000",
  22340=>"010011000",
  22341=>"100001111",
  22342=>"110101110",
  22343=>"111010000",
  22344=>"010101100",
  22345=>"001010010",
  22346=>"000110001",
  22347=>"110111010",
  22348=>"101111101",
  22349=>"011111001",
  22350=>"001010000",
  22351=>"001001001",
  22352=>"110100001",
  22353=>"001100101",
  22354=>"110000111",
  22355=>"011011011",
  22356=>"111100111",
  22357=>"110111110",
  22358=>"001111011",
  22359=>"001011011",
  22360=>"001101110",
  22361=>"110110101",
  22362=>"111010010",
  22363=>"111110000",
  22364=>"000111110",
  22365=>"101111101",
  22366=>"001010110",
  22367=>"000011000",
  22368=>"100101101",
  22369=>"011001101",
  22370=>"000000010",
  22371=>"101011110",
  22372=>"010010110",
  22373=>"101011111",
  22374=>"100011101",
  22375=>"001110111",
  22376=>"111000100",
  22377=>"100001001",
  22378=>"100110000",
  22379=>"010011110",
  22380=>"111000101",
  22381=>"011111101",
  22382=>"001111111",
  22383=>"100001100",
  22384=>"100011110",
  22385=>"100010010",
  22386=>"101000100",
  22387=>"001010101",
  22388=>"110011110",
  22389=>"110110011",
  22390=>"000110000",
  22391=>"000010011",
  22392=>"011111110",
  22393=>"001010000",
  22394=>"100110001",
  22395=>"011011111",
  22396=>"001010010",
  22397=>"100101101",
  22398=>"011011010",
  22399=>"111011000",
  22400=>"111101010",
  22401=>"111111010",
  22402=>"100111100",
  22403=>"001000010",
  22404=>"010110101",
  22405=>"111001000",
  22406=>"001101011",
  22407=>"101101011",
  22408=>"000101011",
  22409=>"110111111",
  22410=>"000111011",
  22411=>"000111110",
  22412=>"110111110",
  22413=>"001010111",
  22414=>"011001110",
  22415=>"010101110",
  22416=>"001110010",
  22417=>"111101101",
  22418=>"100101000",
  22419=>"110011111",
  22420=>"000011110",
  22421=>"001001101",
  22422=>"111101100",
  22423=>"101101011",
  22424=>"000100111",
  22425=>"001000010",
  22426=>"011100000",
  22427=>"000110101",
  22428=>"010111111",
  22429=>"101001011",
  22430=>"000001010",
  22431=>"100110011",
  22432=>"001101110",
  22433=>"011011000",
  22434=>"101010010",
  22435=>"111110011",
  22436=>"000011011",
  22437=>"000010100",
  22438=>"001101111",
  22439=>"110010101",
  22440=>"001000100",
  22441=>"000000000",
  22442=>"010101011",
  22443=>"001000010",
  22444=>"000000011",
  22445=>"101011011",
  22446=>"011100110",
  22447=>"110011100",
  22448=>"110001001",
  22449=>"100110011",
  22450=>"100010010",
  22451=>"010011001",
  22452=>"000011110",
  22453=>"000101010",
  22454=>"011011100",
  22455=>"000010000",
  22456=>"000110100",
  22457=>"011011001",
  22458=>"011110101",
  22459=>"000100111",
  22460=>"010011000",
  22461=>"101110010",
  22462=>"010001110",
  22463=>"010001010",
  22464=>"010110100",
  22465=>"010001011",
  22466=>"011011011",
  22467=>"101000000",
  22468=>"001101100",
  22469=>"110111000",
  22470=>"100100101",
  22471=>"000110001",
  22472=>"011011000",
  22473=>"011111101",
  22474=>"001111000",
  22475=>"010010001",
  22476=>"101111000",
  22477=>"111110111",
  22478=>"010001101",
  22479=>"111100111",
  22480=>"001111101",
  22481=>"100101110",
  22482=>"100101001",
  22483=>"011000011",
  22484=>"110010000",
  22485=>"100110001",
  22486=>"011000101",
  22487=>"110101100",
  22488=>"011101111",
  22489=>"010111001",
  22490=>"110011010",
  22491=>"011110001",
  22492=>"010111101",
  22493=>"111001111",
  22494=>"100101000",
  22495=>"000110100",
  22496=>"101111100",
  22497=>"010101110",
  22498=>"000001001",
  22499=>"000110010",
  22500=>"110100010",
  22501=>"010011110",
  22502=>"000011001",
  22503=>"100100010",
  22504=>"001000110",
  22505=>"001000101",
  22506=>"011000000",
  22507=>"000000011",
  22508=>"110110001",
  22509=>"101010110",
  22510=>"000011100",
  22511=>"100010011",
  22512=>"001100001",
  22513=>"001100011",
  22514=>"001010010",
  22515=>"101000010",
  22516=>"111110001",
  22517=>"010010001",
  22518=>"001100111",
  22519=>"110010101",
  22520=>"000101101",
  22521=>"000011100",
  22522=>"001010000",
  22523=>"101100110",
  22524=>"111100101",
  22525=>"000011011",
  22526=>"101011111",
  22527=>"011101011",
  22528=>"011000111",
  22529=>"001001101",
  22530=>"100101011",
  22531=>"101001011",
  22532=>"100011011",
  22533=>"100100110",
  22534=>"010000001",
  22535=>"111101010",
  22536=>"100101111",
  22537=>"110000111",
  22538=>"001001111",
  22539=>"101011011",
  22540=>"001101001",
  22541=>"001110110",
  22542=>"000000100",
  22543=>"111111011",
  22544=>"111011010",
  22545=>"011110110",
  22546=>"111000110",
  22547=>"011000110",
  22548=>"111101010",
  22549=>"000001000",
  22550=>"101111001",
  22551=>"101110100",
  22552=>"001110001",
  22553=>"000010001",
  22554=>"111111000",
  22555=>"000101100",
  22556=>"101100110",
  22557=>"111001010",
  22558=>"110000111",
  22559=>"111110001",
  22560=>"011000110",
  22561=>"010111100",
  22562=>"000111100",
  22563=>"100001110",
  22564=>"000101101",
  22565=>"111111011",
  22566=>"111100100",
  22567=>"101000000",
  22568=>"000111110",
  22569=>"110011001",
  22570=>"100100101",
  22571=>"000110010",
  22572=>"000000011",
  22573=>"001010010",
  22574=>"101110100",
  22575=>"011101101",
  22576=>"110010010",
  22577=>"000011110",
  22578=>"011010101",
  22579=>"011100010",
  22580=>"110100000",
  22581=>"000001000",
  22582=>"110011011",
  22583=>"110010000",
  22584=>"110011001",
  22585=>"000100101",
  22586=>"100010000",
  22587=>"110111010",
  22588=>"101101101",
  22589=>"010000110",
  22590=>"110111100",
  22591=>"100001110",
  22592=>"111110101",
  22593=>"110001010",
  22594=>"010000110",
  22595=>"111110111",
  22596=>"111111010",
  22597=>"101100101",
  22598=>"001100001",
  22599=>"001100111",
  22600=>"111111100",
  22601=>"010000110",
  22602=>"011011111",
  22603=>"010010110",
  22604=>"100101011",
  22605=>"110110110",
  22606=>"110010101",
  22607=>"010001001",
  22608=>"000010101",
  22609=>"001111011",
  22610=>"011110000",
  22611=>"100010000",
  22612=>"000110101",
  22613=>"011111001",
  22614=>"011110011",
  22615=>"110110011",
  22616=>"110011000",
  22617=>"100111110",
  22618=>"010000000",
  22619=>"001000010",
  22620=>"000011101",
  22621=>"100101101",
  22622=>"110100100",
  22623=>"010010100",
  22624=>"111001100",
  22625=>"111010010",
  22626=>"010010101",
  22627=>"100110001",
  22628=>"100100010",
  22629=>"000011111",
  22630=>"110110110",
  22631=>"100101111",
  22632=>"111111000",
  22633=>"101100111",
  22634=>"110010000",
  22635=>"001011111",
  22636=>"011111000",
  22637=>"000001001",
  22638=>"111010111",
  22639=>"000000011",
  22640=>"000000111",
  22641=>"001101110",
  22642=>"010001111",
  22643=>"101101010",
  22644=>"000001000",
  22645=>"101101000",
  22646=>"110010011",
  22647=>"011001001",
  22648=>"010000000",
  22649=>"101111000",
  22650=>"111011101",
  22651=>"000001001",
  22652=>"011110001",
  22653=>"100010000",
  22654=>"010000010",
  22655=>"011000011",
  22656=>"001010010",
  22657=>"000010011",
  22658=>"000110000",
  22659=>"110000001",
  22660=>"111011100",
  22661=>"101010100",
  22662=>"110110110",
  22663=>"101111101",
  22664=>"011010101",
  22665=>"001101010",
  22666=>"011110100",
  22667=>"100001011",
  22668=>"001100100",
  22669=>"100111111",
  22670=>"101111111",
  22671=>"101100101",
  22672=>"110011010",
  22673=>"000100101",
  22674=>"101111100",
  22675=>"110010010",
  22676=>"001110100",
  22677=>"111101101",
  22678=>"100110111",
  22679=>"001000001",
  22680=>"010110011",
  22681=>"000110110",
  22682=>"111010001",
  22683=>"011101010",
  22684=>"000101011",
  22685=>"110101111",
  22686=>"101010000",
  22687=>"101001101",
  22688=>"100011111",
  22689=>"100000001",
  22690=>"110111011",
  22691=>"011001111",
  22692=>"100100110",
  22693=>"001010001",
  22694=>"001111001",
  22695=>"000100100",
  22696=>"001101100",
  22697=>"011010001",
  22698=>"110110011",
  22699=>"011010010",
  22700=>"111010111",
  22701=>"000110101",
  22702=>"100000000",
  22703=>"101100000",
  22704=>"000000100",
  22705=>"110111000",
  22706=>"010001011",
  22707=>"001001110",
  22708=>"000001001",
  22709=>"000111111",
  22710=>"001101000",
  22711=>"101101111",
  22712=>"111010000",
  22713=>"100010101",
  22714=>"110110101",
  22715=>"011001111",
  22716=>"000000001",
  22717=>"100011111",
  22718=>"000010011",
  22719=>"110110101",
  22720=>"010110001",
  22721=>"001010101",
  22722=>"000101011",
  22723=>"110111111",
  22724=>"111110001",
  22725=>"000000000",
  22726=>"110011000",
  22727=>"111011010",
  22728=>"001011011",
  22729=>"010100111",
  22730=>"101111101",
  22731=>"110111010",
  22732=>"111100001",
  22733=>"001111111",
  22734=>"110001110",
  22735=>"000000100",
  22736=>"001001111",
  22737=>"100011001",
  22738=>"111000000",
  22739=>"001100011",
  22740=>"010101001",
  22741=>"011011011",
  22742=>"010100011",
  22743=>"101010100",
  22744=>"011110111",
  22745=>"010000011",
  22746=>"000110011",
  22747=>"110111001",
  22748=>"111101001",
  22749=>"111010111",
  22750=>"001010001",
  22751=>"010010100",
  22752=>"111000000",
  22753=>"110011010",
  22754=>"000010011",
  22755=>"010001011",
  22756=>"110001011",
  22757=>"011100101",
  22758=>"101111111",
  22759=>"000110110",
  22760=>"100100010",
  22761=>"111100000",
  22762=>"110101110",
  22763=>"110010001",
  22764=>"011100100",
  22765=>"111011111",
  22766=>"001000100",
  22767=>"010100001",
  22768=>"101110101",
  22769=>"011010101",
  22770=>"010010011",
  22771=>"100010010",
  22772=>"000011010",
  22773=>"111011101",
  22774=>"110000010",
  22775=>"111000011",
  22776=>"100000100",
  22777=>"111010110",
  22778=>"110000011",
  22779=>"010111001",
  22780=>"111001010",
  22781=>"100001010",
  22782=>"111010010",
  22783=>"101101101",
  22784=>"011101101",
  22785=>"100101101",
  22786=>"100001011",
  22787=>"101101001",
  22788=>"011000111",
  22789=>"001000100",
  22790=>"000101101",
  22791=>"011010010",
  22792=>"001011010",
  22793=>"111011111",
  22794=>"110011101",
  22795=>"101111011",
  22796=>"100011110",
  22797=>"100101101",
  22798=>"101010111",
  22799=>"001001000",
  22800=>"000111111",
  22801=>"100011001",
  22802=>"000011100",
  22803=>"111011001",
  22804=>"100101011",
  22805=>"011100001",
  22806=>"100011110",
  22807=>"101101100",
  22808=>"000010010",
  22809=>"101001100",
  22810=>"101111101",
  22811=>"011110000",
  22812=>"101110010",
  22813=>"001111100",
  22814=>"010010110",
  22815=>"100010110",
  22816=>"001000110",
  22817=>"111111111",
  22818=>"111100110",
  22819=>"001110000",
  22820=>"101111110",
  22821=>"010011100",
  22822=>"101100111",
  22823=>"111111110",
  22824=>"001111100",
  22825=>"111111000",
  22826=>"010000100",
  22827=>"110001110",
  22828=>"100111000",
  22829=>"110101000",
  22830=>"010100110",
  22831=>"011100110",
  22832=>"100100000",
  22833=>"100010011",
  22834=>"101110100",
  22835=>"100100001",
  22836=>"111110011",
  22837=>"100111100",
  22838=>"011001111",
  22839=>"001010000",
  22840=>"101011101",
  22841=>"001000010",
  22842=>"100010011",
  22843=>"100101000",
  22844=>"010010100",
  22845=>"110001110",
  22846=>"010010001",
  22847=>"100011111",
  22848=>"000101010",
  22849=>"110011011",
  22850=>"100000111",
  22851=>"001000001",
  22852=>"001110110",
  22853=>"000011001",
  22854=>"000010011",
  22855=>"000100010",
  22856=>"100011010",
  22857=>"101111100",
  22858=>"000000000",
  22859=>"110011010",
  22860=>"100111000",
  22861=>"010101100",
  22862=>"000100101",
  22863=>"001011111",
  22864=>"000110000",
  22865=>"100101011",
  22866=>"001011101",
  22867=>"111100011",
  22868=>"111110010",
  22869=>"110011010",
  22870=>"010100101",
  22871=>"110100001",
  22872=>"100001000",
  22873=>"101000101",
  22874=>"000101010",
  22875=>"100101001",
  22876=>"100011010",
  22877=>"110101101",
  22878=>"011100000",
  22879=>"001110011",
  22880=>"101110000",
  22881=>"010101000",
  22882=>"100100100",
  22883=>"100010101",
  22884=>"000100000",
  22885=>"010011001",
  22886=>"110010001",
  22887=>"111110110",
  22888=>"111001110",
  22889=>"101101101",
  22890=>"000100111",
  22891=>"000000100",
  22892=>"001111000",
  22893=>"100101000",
  22894=>"000100110",
  22895=>"011001011",
  22896=>"010010100",
  22897=>"111101010",
  22898=>"111111001",
  22899=>"100010001",
  22900=>"110010010",
  22901=>"010111000",
  22902=>"100001011",
  22903=>"101010001",
  22904=>"000101111",
  22905=>"110011011",
  22906=>"110010100",
  22907=>"100101010",
  22908=>"011101110",
  22909=>"000011010",
  22910=>"100001110",
  22911=>"101101110",
  22912=>"011011100",
  22913=>"000101110",
  22914=>"101111111",
  22915=>"101111101",
  22916=>"010101010",
  22917=>"111101001",
  22918=>"101111111",
  22919=>"111001101",
  22920=>"100111010",
  22921=>"000000111",
  22922=>"100000100",
  22923=>"000010010",
  22924=>"011100100",
  22925=>"000101101",
  22926=>"101101011",
  22927=>"000100110",
  22928=>"101010000",
  22929=>"110000110",
  22930=>"101111100",
  22931=>"111110111",
  22932=>"101101001",
  22933=>"101101000",
  22934=>"101110011",
  22935=>"111111011",
  22936=>"111111001",
  22937=>"000000100",
  22938=>"101110101",
  22939=>"000001110",
  22940=>"001001010",
  22941=>"000001110",
  22942=>"101100101",
  22943=>"101010100",
  22944=>"100000010",
  22945=>"000111101",
  22946=>"010010101",
  22947=>"100011001",
  22948=>"111011110",
  22949=>"101000001",
  22950=>"100000110",
  22951=>"000011101",
  22952=>"100111001",
  22953=>"111001011",
  22954=>"100101010",
  22955=>"101011010",
  22956=>"001110011",
  22957=>"100111100",
  22958=>"000110100",
  22959=>"110010011",
  22960=>"111011111",
  22961=>"011110111",
  22962=>"101000010",
  22963=>"111111000",
  22964=>"100000110",
  22965=>"000101111",
  22966=>"000111101",
  22967=>"001100001",
  22968=>"111010010",
  22969=>"110010111",
  22970=>"101010011",
  22971=>"110010010",
  22972=>"010110101",
  22973=>"110111111",
  22974=>"100010010",
  22975=>"111011011",
  22976=>"111111100",
  22977=>"100010101",
  22978=>"010010111",
  22979=>"101010011",
  22980=>"111101111",
  22981=>"111001100",
  22982=>"110110011",
  22983=>"010000000",
  22984=>"100110101",
  22985=>"101100110",
  22986=>"100110001",
  22987=>"100100110",
  22988=>"001001111",
  22989=>"111010010",
  22990=>"110110000",
  22991=>"001001011",
  22992=>"111100111",
  22993=>"110110101",
  22994=>"101010001",
  22995=>"100011110",
  22996=>"001110011",
  22997=>"110000000",
  22998=>"010100010",
  22999=>"101101001",
  23000=>"110001000",
  23001=>"100110001",
  23002=>"010001000",
  23003=>"111100000",
  23004=>"111100101",
  23005=>"111011000",
  23006=>"101000110",
  23007=>"110010001",
  23008=>"100011100",
  23009=>"011111010",
  23010=>"001101010",
  23011=>"010101000",
  23012=>"111000111",
  23013=>"100101100",
  23014=>"001111101",
  23015=>"001101001",
  23016=>"001111001",
  23017=>"011000011",
  23018=>"110110101",
  23019=>"100010000",
  23020=>"110100110",
  23021=>"111010000",
  23022=>"000101000",
  23023=>"011011010",
  23024=>"011100010",
  23025=>"011111110",
  23026=>"111011101",
  23027=>"111110001",
  23028=>"101000111",
  23029=>"000100000",
  23030=>"000001111",
  23031=>"100001001",
  23032=>"111010100",
  23033=>"011001101",
  23034=>"011000110",
  23035=>"010000101",
  23036=>"000001011",
  23037=>"101110101",
  23038=>"000000101",
  23039=>"001011110",
  23040=>"111011010",
  23041=>"110110100",
  23042=>"101100010",
  23043=>"000010100",
  23044=>"100001000",
  23045=>"110010111",
  23046=>"101010011",
  23047=>"111010011",
  23048=>"101000101",
  23049=>"110111101",
  23050=>"110110011",
  23051=>"110010010",
  23052=>"111011100",
  23053=>"110000011",
  23054=>"101001110",
  23055=>"000001010",
  23056=>"110100010",
  23057=>"000001100",
  23058=>"101001101",
  23059=>"000011110",
  23060=>"110000100",
  23061=>"100100101",
  23062=>"111011001",
  23063=>"100010000",
  23064=>"111010000",
  23065=>"001001000",
  23066=>"101111011",
  23067=>"001111110",
  23068=>"011100110",
  23069=>"011110101",
  23070=>"001001110",
  23071=>"111101010",
  23072=>"011110100",
  23073=>"101110010",
  23074=>"010100100",
  23075=>"010001001",
  23076=>"110011100",
  23077=>"001111100",
  23078=>"010111110",
  23079=>"110110111",
  23080=>"001000011",
  23081=>"111100000",
  23082=>"001000111",
  23083=>"000101111",
  23084=>"111001001",
  23085=>"100001111",
  23086=>"010110000",
  23087=>"110101110",
  23088=>"101010110",
  23089=>"110011010",
  23090=>"111111100",
  23091=>"100010100",
  23092=>"100011011",
  23093=>"000100010",
  23094=>"001101101",
  23095=>"001000011",
  23096=>"101100011",
  23097=>"101110000",
  23098=>"011111111",
  23099=>"100000011",
  23100=>"111101110",
  23101=>"110010101",
  23102=>"001011100",
  23103=>"111101001",
  23104=>"011011101",
  23105=>"110100101",
  23106=>"010111000",
  23107=>"010110000",
  23108=>"111010000",
  23109=>"011000010",
  23110=>"111101100",
  23111=>"000000101",
  23112=>"110001110",
  23113=>"000111100",
  23114=>"010101111",
  23115=>"100100000",
  23116=>"101111000",
  23117=>"100100010",
  23118=>"101100110",
  23119=>"001011110",
  23120=>"111111001",
  23121=>"100101111",
  23122=>"111111011",
  23123=>"010000000",
  23124=>"110101101",
  23125=>"111101000",
  23126=>"010111100",
  23127=>"101111000",
  23128=>"001000110",
  23129=>"000001001",
  23130=>"011110110",
  23131=>"000101100",
  23132=>"100100011",
  23133=>"101010000",
  23134=>"010000101",
  23135=>"110110001",
  23136=>"001111100",
  23137=>"001101010",
  23138=>"000011010",
  23139=>"110000001",
  23140=>"110110011",
  23141=>"101110010",
  23142=>"101111001",
  23143=>"001001010",
  23144=>"010111111",
  23145=>"011001000",
  23146=>"110110111",
  23147=>"110101000",
  23148=>"001011111",
  23149=>"010011110",
  23150=>"010101100",
  23151=>"111000001",
  23152=>"100100000",
  23153=>"110001010",
  23154=>"010010000",
  23155=>"000000111",
  23156=>"011111111",
  23157=>"001101110",
  23158=>"110101001",
  23159=>"110000000",
  23160=>"000110110",
  23161=>"011111110",
  23162=>"011011100",
  23163=>"110110011",
  23164=>"001100111",
  23165=>"111100001",
  23166=>"100111110",
  23167=>"101010000",
  23168=>"100111110",
  23169=>"001001111",
  23170=>"001101111",
  23171=>"101000001",
  23172=>"001010010",
  23173=>"000100111",
  23174=>"100100111",
  23175=>"110101010",
  23176=>"110111110",
  23177=>"100011111",
  23178=>"110010000",
  23179=>"000010110",
  23180=>"010010010",
  23181=>"110100111",
  23182=>"100000011",
  23183=>"100100111",
  23184=>"001101111",
  23185=>"111011010",
  23186=>"100110011",
  23187=>"011000010",
  23188=>"001010011",
  23189=>"000001011",
  23190=>"110100100",
  23191=>"110110000",
  23192=>"100100000",
  23193=>"100000110",
  23194=>"001000110",
  23195=>"000001011",
  23196=>"111010000",
  23197=>"010111101",
  23198=>"110110001",
  23199=>"010010011",
  23200=>"001101101",
  23201=>"111111011",
  23202=>"111111001",
  23203=>"111111100",
  23204=>"000000111",
  23205=>"110010011",
  23206=>"111111100",
  23207=>"000010110",
  23208=>"111111110",
  23209=>"101111000",
  23210=>"010111101",
  23211=>"111011110",
  23212=>"100100110",
  23213=>"000010110",
  23214=>"101101100",
  23215=>"001100001",
  23216=>"101111010",
  23217=>"110010100",
  23218=>"011101001",
  23219=>"100011100",
  23220=>"101011010",
  23221=>"111011001",
  23222=>"010110010",
  23223=>"111101110",
  23224=>"000111001",
  23225=>"110111110",
  23226=>"010101000",
  23227=>"011000100",
  23228=>"001000001",
  23229=>"000100001",
  23230=>"111011001",
  23231=>"011000111",
  23232=>"111101110",
  23233=>"110011000",
  23234=>"101110100",
  23235=>"001101011",
  23236=>"011111111",
  23237=>"101000110",
  23238=>"011010000",
  23239=>"101111110",
  23240=>"010000000",
  23241=>"100001010",
  23242=>"001010011",
  23243=>"101110110",
  23244=>"001111110",
  23245=>"010000000",
  23246=>"011110111",
  23247=>"111011001",
  23248=>"011000110",
  23249=>"011011010",
  23250=>"100101000",
  23251=>"011111001",
  23252=>"101000010",
  23253=>"000111101",
  23254=>"010100010",
  23255=>"100100101",
  23256=>"010110000",
  23257=>"000000010",
  23258=>"100100001",
  23259=>"110001011",
  23260=>"100100000",
  23261=>"100110100",
  23262=>"010110100",
  23263=>"100111110",
  23264=>"011101111",
  23265=>"000000101",
  23266=>"000101110",
  23267=>"111111111",
  23268=>"111101000",
  23269=>"010010001",
  23270=>"101000000",
  23271=>"110101011",
  23272=>"011001100",
  23273=>"000000000",
  23274=>"100000010",
  23275=>"010111110",
  23276=>"101001011",
  23277=>"111000000",
  23278=>"111111010",
  23279=>"111011010",
  23280=>"110000010",
  23281=>"001010010",
  23282=>"110011110",
  23283=>"001111000",
  23284=>"001011001",
  23285=>"101101001",
  23286=>"110001011",
  23287=>"100101110",
  23288=>"010000011",
  23289=>"111011000",
  23290=>"100110110",
  23291=>"000111111",
  23292=>"111111101",
  23293=>"001000000",
  23294=>"101110101",
  23295=>"101110000",
  23296=>"100001011",
  23297=>"001110011",
  23298=>"111011111",
  23299=>"011010011",
  23300=>"000101110",
  23301=>"000001000",
  23302=>"001101100",
  23303=>"111101100",
  23304=>"000100111",
  23305=>"101111101",
  23306=>"101000000",
  23307=>"001011001",
  23308=>"000010110",
  23309=>"000010111",
  23310=>"000110010",
  23311=>"101111010",
  23312=>"101110110",
  23313=>"110010010",
  23314=>"111111000",
  23315=>"110000000",
  23316=>"010001011",
  23317=>"110100100",
  23318=>"110101010",
  23319=>"110100111",
  23320=>"110011110",
  23321=>"011000000",
  23322=>"100011001",
  23323=>"100010000",
  23324=>"010101010",
  23325=>"000101110",
  23326=>"101011101",
  23327=>"001011101",
  23328=>"000000101",
  23329=>"011000110",
  23330=>"110101010",
  23331=>"101111100",
  23332=>"011010111",
  23333=>"001001111",
  23334=>"000011000",
  23335=>"000000111",
  23336=>"110110011",
  23337=>"100100100",
  23338=>"111111111",
  23339=>"000110101",
  23340=>"110001110",
  23341=>"111101110",
  23342=>"111000111",
  23343=>"110011111",
  23344=>"010000110",
  23345=>"010100000",
  23346=>"111101100",
  23347=>"111010100",
  23348=>"100111111",
  23349=>"101110100",
  23350=>"010011001",
  23351=>"100000111",
  23352=>"111001110",
  23353=>"011011000",
  23354=>"001001000",
  23355=>"111000111",
  23356=>"100000101",
  23357=>"001010110",
  23358=>"101010100",
  23359=>"110111111",
  23360=>"011111111",
  23361=>"011101101",
  23362=>"000000000",
  23363=>"110110101",
  23364=>"001100111",
  23365=>"111011101",
  23366=>"010001000",
  23367=>"011101001",
  23368=>"110001110",
  23369=>"000000001",
  23370=>"011101001",
  23371=>"110101110",
  23372=>"001101010",
  23373=>"101101110",
  23374=>"110110100",
  23375=>"011101000",
  23376=>"011100000",
  23377=>"000110111",
  23378=>"101011100",
  23379=>"101100111",
  23380=>"000110001",
  23381=>"110010011",
  23382=>"101010100",
  23383=>"010001000",
  23384=>"011010010",
  23385=>"010010100",
  23386=>"101011110",
  23387=>"101110011",
  23388=>"111011010",
  23389=>"000100000",
  23390=>"110101100",
  23391=>"011011010",
  23392=>"101011111",
  23393=>"010110000",
  23394=>"110000001",
  23395=>"111100111",
  23396=>"001010100",
  23397=>"100000111",
  23398=>"011111111",
  23399=>"111111010",
  23400=>"001100111",
  23401=>"101101101",
  23402=>"111011111",
  23403=>"010000110",
  23404=>"101001000",
  23405=>"000110001",
  23406=>"110100101",
  23407=>"110011100",
  23408=>"101110110",
  23409=>"110100000",
  23410=>"011100000",
  23411=>"110001100",
  23412=>"110011001",
  23413=>"000101000",
  23414=>"100000000",
  23415=>"011110010",
  23416=>"101000101",
  23417=>"101100000",
  23418=>"011101001",
  23419=>"100101000",
  23420=>"100001011",
  23421=>"011110111",
  23422=>"011111001",
  23423=>"010001001",
  23424=>"101110010",
  23425=>"111001110",
  23426=>"011001101",
  23427=>"010101001",
  23428=>"100101100",
  23429=>"111011001",
  23430=>"100100001",
  23431=>"100001101",
  23432=>"001110000",
  23433=>"010110010",
  23434=>"110111100",
  23435=>"000110010",
  23436=>"010110110",
  23437=>"010101011",
  23438=>"000001000",
  23439=>"110111111",
  23440=>"001110101",
  23441=>"100001000",
  23442=>"110101101",
  23443=>"010100001",
  23444=>"000000111",
  23445=>"000101110",
  23446=>"100001001",
  23447=>"111101110",
  23448=>"010100100",
  23449=>"110101010",
  23450=>"111011001",
  23451=>"000000000",
  23452=>"101001010",
  23453=>"001100001",
  23454=>"111111111",
  23455=>"100011011",
  23456=>"101100111",
  23457=>"011100010",
  23458=>"011011000",
  23459=>"100000101",
  23460=>"111000110",
  23461=>"000000001",
  23462=>"011110100",
  23463=>"000110110",
  23464=>"111111100",
  23465=>"101111110",
  23466=>"100001000",
  23467=>"011110010",
  23468=>"100110001",
  23469=>"110011010",
  23470=>"100111100",
  23471=>"010000100",
  23472=>"100110100",
  23473=>"111101100",
  23474=>"100001001",
  23475=>"110010100",
  23476=>"000011010",
  23477=>"101111101",
  23478=>"100000010",
  23479=>"000111101",
  23480=>"100101011",
  23481=>"001110000",
  23482=>"011100010",
  23483=>"010100010",
  23484=>"101000000",
  23485=>"000011011",
  23486=>"010110010",
  23487=>"100010101",
  23488=>"001010010",
  23489=>"001001001",
  23490=>"011001001",
  23491=>"110011000",
  23492=>"110000011",
  23493=>"011101110",
  23494=>"001011011",
  23495=>"111010111",
  23496=>"100000010",
  23497=>"101111010",
  23498=>"000101011",
  23499=>"110001101",
  23500=>"101110110",
  23501=>"111111101",
  23502=>"101111010",
  23503=>"100111011",
  23504=>"100101100",
  23505=>"100001010",
  23506=>"111011001",
  23507=>"010100001",
  23508=>"111001111",
  23509=>"011001000",
  23510=>"111101110",
  23511=>"101110101",
  23512=>"010011110",
  23513=>"110011001",
  23514=>"100010100",
  23515=>"101010111",
  23516=>"011001110",
  23517=>"000111001",
  23518=>"110010101",
  23519=>"111111100",
  23520=>"011100000",
  23521=>"000000111",
  23522=>"110111011",
  23523=>"101011111",
  23524=>"010100100",
  23525=>"111111011",
  23526=>"100001001",
  23527=>"110000010",
  23528=>"001100000",
  23529=>"000100000",
  23530=>"000100000",
  23531=>"011110011",
  23532=>"001000100",
  23533=>"100100000",
  23534=>"000010010",
  23535=>"011111100",
  23536=>"110100000",
  23537=>"000101011",
  23538=>"000110011",
  23539=>"000001000",
  23540=>"000010110",
  23541=>"011001010",
  23542=>"000000111",
  23543=>"100101001",
  23544=>"000000110",
  23545=>"100010000",
  23546=>"101010110",
  23547=>"100000101",
  23548=>"100011100",
  23549=>"011011011",
  23550=>"010111101",
  23551=>"100000100",
  23552=>"000000011",
  23553=>"111011100",
  23554=>"001011001",
  23555=>"000000101",
  23556=>"001110000",
  23557=>"100000100",
  23558=>"111110101",
  23559=>"101001101",
  23560=>"111110011",
  23561=>"110001111",
  23562=>"010100111",
  23563=>"111110101",
  23564=>"111010101",
  23565=>"000100000",
  23566=>"110011001",
  23567=>"111111001",
  23568=>"111011111",
  23569=>"010111010",
  23570=>"000100111",
  23571=>"001000100",
  23572=>"000010101",
  23573=>"011101010",
  23574=>"111100101",
  23575=>"111000010",
  23576=>"011110010",
  23577=>"011110010",
  23578=>"000100000",
  23579=>"001000000",
  23580=>"111011010",
  23581=>"010000110",
  23582=>"110011010",
  23583=>"000001110",
  23584=>"110100000",
  23585=>"010111000",
  23586=>"100100000",
  23587=>"010100100",
  23588=>"001111000",
  23589=>"000011010",
  23590=>"111010000",
  23591=>"001010101",
  23592=>"001111011",
  23593=>"101101101",
  23594=>"001110101",
  23595=>"000011100",
  23596=>"100001101",
  23597=>"011100110",
  23598=>"001001101",
  23599=>"000110111",
  23600=>"101111011",
  23601=>"111110000",
  23602=>"010100000",
  23603=>"001010001",
  23604=>"011100010",
  23605=>"100100110",
  23606=>"000110000",
  23607=>"000001100",
  23608=>"010000101",
  23609=>"100011100",
  23610=>"111101100",
  23611=>"101101111",
  23612=>"000100000",
  23613=>"101011111",
  23614=>"101001110",
  23615=>"000011011",
  23616=>"010000101",
  23617=>"000100000",
  23618=>"000101000",
  23619=>"010011100",
  23620=>"111001000",
  23621=>"100111011",
  23622=>"100001001",
  23623=>"011011110",
  23624=>"100111011",
  23625=>"110010011",
  23626=>"100110011",
  23627=>"010011110",
  23628=>"010101100",
  23629=>"010111000",
  23630=>"010111011",
  23631=>"110010010",
  23632=>"111011111",
  23633=>"010011011",
  23634=>"101010100",
  23635=>"001100110",
  23636=>"100111111",
  23637=>"010000100",
  23638=>"111101100",
  23639=>"001011010",
  23640=>"010101100",
  23641=>"101011111",
  23642=>"011011001",
  23643=>"011010111",
  23644=>"110100000",
  23645=>"101100010",
  23646=>"001100100",
  23647=>"000101011",
  23648=>"000000010",
  23649=>"101111011",
  23650=>"100110000",
  23651=>"010011100",
  23652=>"101110010",
  23653=>"110011010",
  23654=>"110111001",
  23655=>"110110101",
  23656=>"000000010",
  23657=>"001011110",
  23658=>"111100000",
  23659=>"111110000",
  23660=>"110110001",
  23661=>"010001110",
  23662=>"000001011",
  23663=>"010111101",
  23664=>"111101111",
  23665=>"111101110",
  23666=>"111011100",
  23667=>"100011000",
  23668=>"101111011",
  23669=>"000001111",
  23670=>"110100100",
  23671=>"001010001",
  23672=>"101110110",
  23673=>"110001011",
  23674=>"111010100",
  23675=>"100110001",
  23676=>"101010001",
  23677=>"101000000",
  23678=>"000101000",
  23679=>"010010011",
  23680=>"111010101",
  23681=>"010000101",
  23682=>"001010000",
  23683=>"101010000",
  23684=>"111010000",
  23685=>"100111001",
  23686=>"101111001",
  23687=>"110000010",
  23688=>"100100010",
  23689=>"110011101",
  23690=>"110101110",
  23691=>"100111010",
  23692=>"011111111",
  23693=>"010001000",
  23694=>"110010110",
  23695=>"111101111",
  23696=>"110001000",
  23697=>"100001111",
  23698=>"011000011",
  23699=>"000010110",
  23700=>"111111111",
  23701=>"111011110",
  23702=>"000100111",
  23703=>"100000010",
  23704=>"010110110",
  23705=>"110100110",
  23706=>"000001101",
  23707=>"000010001",
  23708=>"111000010",
  23709=>"010101111",
  23710=>"001010111",
  23711=>"100001000",
  23712=>"001110001",
  23713=>"101101000",
  23714=>"100101111",
  23715=>"111110111",
  23716=>"010011101",
  23717=>"011111001",
  23718=>"100001001",
  23719=>"110100100",
  23720=>"011000100",
  23721=>"111001001",
  23722=>"010001010",
  23723=>"110000001",
  23724=>"100111101",
  23725=>"011011011",
  23726=>"001001101",
  23727=>"110110110",
  23728=>"000000111",
  23729=>"000001000",
  23730=>"001111010",
  23731=>"100010001",
  23732=>"010101111",
  23733=>"110110110",
  23734=>"101010111",
  23735=>"001000100",
  23736=>"100010000",
  23737=>"110110111",
  23738=>"000010000",
  23739=>"101101010",
  23740=>"101111111",
  23741=>"101011100",
  23742=>"011111000",
  23743=>"011110100",
  23744=>"001110001",
  23745=>"000100011",
  23746=>"010000011",
  23747=>"000111011",
  23748=>"101000000",
  23749=>"110011110",
  23750=>"100101000",
  23751=>"101011100",
  23752=>"010001011",
  23753=>"010010001",
  23754=>"111100000",
  23755=>"000001110",
  23756=>"100000111",
  23757=>"110111111",
  23758=>"100000011",
  23759=>"000100111",
  23760=>"101000110",
  23761=>"010010010",
  23762=>"100101001",
  23763=>"000101011",
  23764=>"100110111",
  23765=>"011101110",
  23766=>"000011100",
  23767=>"010100000",
  23768=>"010111011",
  23769=>"001011110",
  23770=>"000100110",
  23771=>"010000010",
  23772=>"101010111",
  23773=>"110111111",
  23774=>"100000110",
  23775=>"010101110",
  23776=>"111000000",
  23777=>"010011110",
  23778=>"111000111",
  23779=>"011011010",
  23780=>"001101001",
  23781=>"100000110",
  23782=>"000011010",
  23783=>"110000111",
  23784=>"100000000",
  23785=>"011111100",
  23786=>"000010000",
  23787=>"110011111",
  23788=>"111101100",
  23789=>"001011011",
  23790=>"011011100",
  23791=>"100010010",
  23792=>"011101111",
  23793=>"010010010",
  23794=>"110101100",
  23795=>"111111000",
  23796=>"001111001",
  23797=>"110111110",
  23798=>"011110000",
  23799=>"000000010",
  23800=>"100101111",
  23801=>"011100100",
  23802=>"010011110",
  23803=>"011010110",
  23804=>"100001100",
  23805=>"010011101",
  23806=>"111100010",
  23807=>"000111101",
  23808=>"101111011",
  23809=>"111101011",
  23810=>"000001101",
  23811=>"011000100",
  23812=>"000011001",
  23813=>"101111000",
  23814=>"000000111",
  23815=>"100101101",
  23816=>"100101101",
  23817=>"001011110",
  23818=>"011110100",
  23819=>"110101101",
  23820=>"001110110",
  23821=>"011111010",
  23822=>"001010100",
  23823=>"001000000",
  23824=>"100110101",
  23825=>"000101011",
  23826=>"110001000",
  23827=>"011100111",
  23828=>"101110001",
  23829=>"111100000",
  23830=>"001000010",
  23831=>"010010010",
  23832=>"011100000",
  23833=>"100010001",
  23834=>"011100010",
  23835=>"111111011",
  23836=>"110100010",
  23837=>"010000101",
  23838=>"001110110",
  23839=>"010000001",
  23840=>"111110010",
  23841=>"111100011",
  23842=>"010110101",
  23843=>"011000110",
  23844=>"011111101",
  23845=>"101110000",
  23846=>"010100110",
  23847=>"001011000",
  23848=>"110111000",
  23849=>"100110011",
  23850=>"000010111",
  23851=>"100100011",
  23852=>"111010111",
  23853=>"010001000",
  23854=>"101001111",
  23855=>"101000011",
  23856=>"100110011",
  23857=>"000111001",
  23858=>"101111011",
  23859=>"010111101",
  23860=>"000111101",
  23861=>"001001011",
  23862=>"000010101",
  23863=>"110000111",
  23864=>"011100100",
  23865=>"110010101",
  23866=>"000111110",
  23867=>"011111111",
  23868=>"111000010",
  23869=>"110111111",
  23870=>"001010010",
  23871=>"101100001",
  23872=>"010100010",
  23873=>"111101010",
  23874=>"001000010",
  23875=>"111000101",
  23876=>"001010111",
  23877=>"110000010",
  23878=>"101110101",
  23879=>"010010010",
  23880=>"111001001",
  23881=>"110110010",
  23882=>"000110100",
  23883=>"000011111",
  23884=>"000011001",
  23885=>"110011010",
  23886=>"000111111",
  23887=>"110101100",
  23888=>"010111111",
  23889=>"010111000",
  23890=>"000110000",
  23891=>"011000111",
  23892=>"010100001",
  23893=>"010110111",
  23894=>"000001000",
  23895=>"111001100",
  23896=>"001000010",
  23897=>"111110100",
  23898=>"111111101",
  23899=>"011010011",
  23900=>"001011000",
  23901=>"011111101",
  23902=>"110110001",
  23903=>"100001110",
  23904=>"010100110",
  23905=>"010011111",
  23906=>"010101110",
  23907=>"000010110",
  23908=>"001001111",
  23909=>"010001011",
  23910=>"000010110",
  23911=>"010001010",
  23912=>"010110110",
  23913=>"000101110",
  23914=>"000001110",
  23915=>"001100000",
  23916=>"010010001",
  23917=>"100100101",
  23918=>"100101010",
  23919=>"000101101",
  23920=>"110111011",
  23921=>"111001101",
  23922=>"001101110",
  23923=>"101000011",
  23924=>"100000111",
  23925=>"101111000",
  23926=>"011001111",
  23927=>"101111000",
  23928=>"100110100",
  23929=>"110110010",
  23930=>"000000110",
  23931=>"101011010",
  23932=>"101100011",
  23933=>"001111111",
  23934=>"011010111",
  23935=>"101001110",
  23936=>"011100111",
  23937=>"010010000",
  23938=>"000011110",
  23939=>"100100100",
  23940=>"111010100",
  23941=>"000011011",
  23942=>"000111000",
  23943=>"010000111",
  23944=>"111010011",
  23945=>"111101001",
  23946=>"000000010",
  23947=>"110101000",
  23948=>"110111110",
  23949=>"010011100",
  23950=>"110101101",
  23951=>"100010001",
  23952=>"001010110",
  23953=>"000101101",
  23954=>"011001010",
  23955=>"000010110",
  23956=>"011001010",
  23957=>"000010101",
  23958=>"100010001",
  23959=>"011111101",
  23960=>"110111111",
  23961=>"111100001",
  23962=>"001011011",
  23963=>"100010100",
  23964=>"101010110",
  23965=>"100111111",
  23966=>"101101111",
  23967=>"011011010",
  23968=>"010110000",
  23969=>"100101110",
  23970=>"001111000",
  23971=>"111111100",
  23972=>"101100000",
  23973=>"011001001",
  23974=>"001010001",
  23975=>"100000011",
  23976=>"100000000",
  23977=>"010111101",
  23978=>"111110110",
  23979=>"000010010",
  23980=>"011011110",
  23981=>"001000011",
  23982=>"000111100",
  23983=>"100101010",
  23984=>"000001001",
  23985=>"010011101",
  23986=>"010100001",
  23987=>"110101011",
  23988=>"110001111",
  23989=>"101011110",
  23990=>"110111111",
  23991=>"010010101",
  23992=>"100011011",
  23993=>"110010110",
  23994=>"111111110",
  23995=>"100010010",
  23996=>"010111110",
  23997=>"000100111",
  23998=>"001010101",
  23999=>"001111100",
  24000=>"000000111",
  24001=>"010100110",
  24002=>"100111100",
  24003=>"111100011",
  24004=>"111011000",
  24005=>"100101000",
  24006=>"111100000",
  24007=>"000111000",
  24008=>"001110010",
  24009=>"010110000",
  24010=>"000001000",
  24011=>"000101100",
  24012=>"111011001",
  24013=>"101101100",
  24014=>"111011100",
  24015=>"000111110",
  24016=>"101110010",
  24017=>"001111010",
  24018=>"010010010",
  24019=>"000101010",
  24020=>"000110001",
  24021=>"011011110",
  24022=>"000000110",
  24023=>"000111110",
  24024=>"001010011",
  24025=>"101001010",
  24026=>"110101100",
  24027=>"000000000",
  24028=>"110001010",
  24029=>"010001100",
  24030=>"010101110",
  24031=>"111110101",
  24032=>"100100010",
  24033=>"101010001",
  24034=>"011011000",
  24035=>"100010000",
  24036=>"010110011",
  24037=>"110011111",
  24038=>"100010100",
  24039=>"001001000",
  24040=>"100111110",
  24041=>"110111111",
  24042=>"100011010",
  24043=>"110010001",
  24044=>"010101110",
  24045=>"111111010",
  24046=>"110111111",
  24047=>"110011100",
  24048=>"100101111",
  24049=>"100111100",
  24050=>"111111001",
  24051=>"000010110",
  24052=>"100000001",
  24053=>"010110101",
  24054=>"100100100",
  24055=>"111001100",
  24056=>"111100001",
  24057=>"011001010",
  24058=>"111101010",
  24059=>"110000001",
  24060=>"101000111",
  24061=>"111100011",
  24062=>"000001001",
  24063=>"101011101",
  24064=>"011100010",
  24065=>"000000000",
  24066=>"111110100",
  24067=>"110101010",
  24068=>"100110001",
  24069=>"001101011",
  24070=>"001001001",
  24071=>"001110000",
  24072=>"110110100",
  24073=>"110110100",
  24074=>"011101000",
  24075=>"001000000",
  24076=>"111011101",
  24077=>"111111101",
  24078=>"110000001",
  24079=>"100011010",
  24080=>"110010001",
  24081=>"100100110",
  24082=>"011111101",
  24083=>"111000111",
  24084=>"100000101",
  24085=>"111001110",
  24086=>"111111111",
  24087=>"000011001",
  24088=>"100000000",
  24089=>"011011000",
  24090=>"011001101",
  24091=>"100100110",
  24092=>"111101110",
  24093=>"111110010",
  24094=>"011000010",
  24095=>"110010110",
  24096=>"000110000",
  24097=>"111110011",
  24098=>"101110001",
  24099=>"000001101",
  24100=>"101010100",
  24101=>"011100011",
  24102=>"110100001",
  24103=>"111110010",
  24104=>"111110100",
  24105=>"110110100",
  24106=>"011110111",
  24107=>"110111000",
  24108=>"111111000",
  24109=>"001100001",
  24110=>"001101010",
  24111=>"110010111",
  24112=>"110110011",
  24113=>"110110011",
  24114=>"100001110",
  24115=>"111011110",
  24116=>"100011101",
  24117=>"111011011",
  24118=>"000111010",
  24119=>"000100111",
  24120=>"000110110",
  24121=>"000000001",
  24122=>"001100100",
  24123=>"101111111",
  24124=>"101111110",
  24125=>"000011000",
  24126=>"000111011",
  24127=>"001101001",
  24128=>"010001000",
  24129=>"101011101",
  24130=>"010001111",
  24131=>"001101001",
  24132=>"010111010",
  24133=>"111101001",
  24134=>"111101010",
  24135=>"000000011",
  24136=>"001100010",
  24137=>"011011101",
  24138=>"110111010",
  24139=>"001001010",
  24140=>"001101001",
  24141=>"100011111",
  24142=>"110101111",
  24143=>"000110001",
  24144=>"010010111",
  24145=>"010100000",
  24146=>"110101111",
  24147=>"111001011",
  24148=>"010000101",
  24149=>"101100011",
  24150=>"010111101",
  24151=>"000111001",
  24152=>"011000000",
  24153=>"011110000",
  24154=>"111001001",
  24155=>"101001000",
  24156=>"000010011",
  24157=>"110011110",
  24158=>"100111001",
  24159=>"011010100",
  24160=>"001101101",
  24161=>"111101101",
  24162=>"110011101",
  24163=>"001001000",
  24164=>"010110001",
  24165=>"101110010",
  24166=>"110010101",
  24167=>"101101000",
  24168=>"011100100",
  24169=>"001011000",
  24170=>"111110111",
  24171=>"010011010",
  24172=>"010010000",
  24173=>"111001100",
  24174=>"111000000",
  24175=>"110100101",
  24176=>"011110011",
  24177=>"110000101",
  24178=>"010110000",
  24179=>"001010011",
  24180=>"111111110",
  24181=>"100011010",
  24182=>"011000001",
  24183=>"000000110",
  24184=>"101000110",
  24185=>"111101111",
  24186=>"101110000",
  24187=>"111000001",
  24188=>"000110010",
  24189=>"001110000",
  24190=>"100111000",
  24191=>"111000000",
  24192=>"111101001",
  24193=>"110101100",
  24194=>"111100110",
  24195=>"111101101",
  24196=>"001001011",
  24197=>"101001110",
  24198=>"011111010",
  24199=>"101011100",
  24200=>"011000110",
  24201=>"111110101",
  24202=>"110101001",
  24203=>"001011010",
  24204=>"110001100",
  24205=>"101010110",
  24206=>"011100101",
  24207=>"001100101",
  24208=>"110011001",
  24209=>"000000010",
  24210=>"000010110",
  24211=>"011001110",
  24212=>"011111000",
  24213=>"011101001",
  24214=>"101110010",
  24215=>"100001100",
  24216=>"001010001",
  24217=>"101100001",
  24218=>"001100111",
  24219=>"010100110",
  24220=>"110000000",
  24221=>"110011010",
  24222=>"011010011",
  24223=>"000110101",
  24224=>"000001111",
  24225=>"111011111",
  24226=>"011001101",
  24227=>"101110001",
  24228=>"110101110",
  24229=>"100000001",
  24230=>"110110101",
  24231=>"011000110",
  24232=>"111010001",
  24233=>"001001000",
  24234=>"011001010",
  24235=>"100001101",
  24236=>"000101111",
  24237=>"011101011",
  24238=>"000001001",
  24239=>"010000010",
  24240=>"101011000",
  24241=>"111101001",
  24242=>"011101000",
  24243=>"101100110",
  24244=>"011001001",
  24245=>"000101101",
  24246=>"100110100",
  24247=>"010101010",
  24248=>"110010010",
  24249=>"011011001",
  24250=>"111011001",
  24251=>"101101011",
  24252=>"011101100",
  24253=>"011100100",
  24254=>"010011110",
  24255=>"111011011",
  24256=>"101001101",
  24257=>"110111010",
  24258=>"101000100",
  24259=>"010101100",
  24260=>"110011011",
  24261=>"110010010",
  24262=>"111010010",
  24263=>"000011010",
  24264=>"001000100",
  24265=>"011100101",
  24266=>"110011100",
  24267=>"000000011",
  24268=>"110111010",
  24269=>"101000000",
  24270=>"000101110",
  24271=>"000111011",
  24272=>"110100000",
  24273=>"011110100",
  24274=>"100101100",
  24275=>"001101010",
  24276=>"101010000",
  24277=>"000101110",
  24278=>"000111010",
  24279=>"010000101",
  24280=>"100001001",
  24281=>"001010101",
  24282=>"110110101",
  24283=>"010101010",
  24284=>"010011111",
  24285=>"001101011",
  24286=>"101010110",
  24287=>"010101011",
  24288=>"010100100",
  24289=>"110001010",
  24290=>"101111100",
  24291=>"101010001",
  24292=>"000111100",
  24293=>"001101111",
  24294=>"111000001",
  24295=>"000010110",
  24296=>"011100010",
  24297=>"010101010",
  24298=>"111000001",
  24299=>"111000110",
  24300=>"000011011",
  24301=>"000010010",
  24302=>"001001111",
  24303=>"001000011",
  24304=>"001011100",
  24305=>"100011111",
  24306=>"010011010",
  24307=>"001000110",
  24308=>"101010010",
  24309=>"010011001",
  24310=>"000001000",
  24311=>"000110110",
  24312=>"101001001",
  24313=>"111000010",
  24314=>"000100101",
  24315=>"001011000",
  24316=>"110000000",
  24317=>"010000010",
  24318=>"101101011",
  24319=>"010011110",
  24320=>"100000011",
  24321=>"010111111",
  24322=>"110100101",
  24323=>"000111000",
  24324=>"111000000",
  24325=>"011111001",
  24326=>"100010110",
  24327=>"110110110",
  24328=>"000010010",
  24329=>"101110111",
  24330=>"111000101",
  24331=>"111010100",
  24332=>"000000011",
  24333=>"111010110",
  24334=>"100100100",
  24335=>"010111100",
  24336=>"000111010",
  24337=>"101100000",
  24338=>"111100111",
  24339=>"101100101",
  24340=>"000110110",
  24341=>"100010100",
  24342=>"111100000",
  24343=>"101000010",
  24344=>"101101011",
  24345=>"111101100",
  24346=>"111010100",
  24347=>"111100001",
  24348=>"101011100",
  24349=>"000110001",
  24350=>"011010010",
  24351=>"110101011",
  24352=>"010100110",
  24353=>"100110000",
  24354=>"011110111",
  24355=>"110001011",
  24356=>"111111100",
  24357=>"101100000",
  24358=>"011111110",
  24359=>"011001011",
  24360=>"001101010",
  24361=>"110110100",
  24362=>"000010000",
  24363=>"101000100",
  24364=>"100101010",
  24365=>"001001111",
  24366=>"011110111",
  24367=>"111000000",
  24368=>"000111111",
  24369=>"000001000",
  24370=>"011000000",
  24371=>"011010100",
  24372=>"011010111",
  24373=>"001010001",
  24374=>"000001011",
  24375=>"010100010",
  24376=>"001110010",
  24377=>"100000100",
  24378=>"101010001",
  24379=>"100010010",
  24380=>"100001111",
  24381=>"110111100",
  24382=>"110111111",
  24383=>"000110110",
  24384=>"111101110",
  24385=>"010110101",
  24386=>"101101011",
  24387=>"000001011",
  24388=>"010000100",
  24389=>"101011110",
  24390=>"011100001",
  24391=>"000000010",
  24392=>"101010100",
  24393=>"101111110",
  24394=>"111011010",
  24395=>"000101011",
  24396=>"111100111",
  24397=>"011000000",
  24398=>"100001101",
  24399=>"000011001",
  24400=>"001011111",
  24401=>"101100101",
  24402=>"111010010",
  24403=>"011001000",
  24404=>"111100100",
  24405=>"100110011",
  24406=>"010010100",
  24407=>"010101111",
  24408=>"111110001",
  24409=>"101011100",
  24410=>"000111101",
  24411=>"101001000",
  24412=>"000010101",
  24413=>"010000100",
  24414=>"010011100",
  24415=>"100100010",
  24416=>"000000111",
  24417=>"011011011",
  24418=>"010101100",
  24419=>"011100111",
  24420=>"101100100",
  24421=>"010101100",
  24422=>"111000000",
  24423=>"010010011",
  24424=>"100111100",
  24425=>"100010111",
  24426=>"110101111",
  24427=>"100111110",
  24428=>"111111010",
  24429=>"101001011",
  24430=>"001001010",
  24431=>"100111001",
  24432=>"110000010",
  24433=>"100100100",
  24434=>"010110111",
  24435=>"110010010",
  24436=>"100110111",
  24437=>"000101100",
  24438=>"111011011",
  24439=>"000100010",
  24440=>"000001011",
  24441=>"001001000",
  24442=>"110001111",
  24443=>"000111111",
  24444=>"001100110",
  24445=>"111011001",
  24446=>"111111110",
  24447=>"001101000",
  24448=>"101110110",
  24449=>"100000010",
  24450=>"111001001",
  24451=>"010000111",
  24452=>"011000110",
  24453=>"110001100",
  24454=>"111011001",
  24455=>"101111111",
  24456=>"111001010",
  24457=>"001010101",
  24458=>"111101111",
  24459=>"000001000",
  24460=>"001000000",
  24461=>"110011110",
  24462=>"100011101",
  24463=>"001110011",
  24464=>"111101100",
  24465=>"100011000",
  24466=>"101011011",
  24467=>"000011111",
  24468=>"110110110",
  24469=>"000101010",
  24470=>"100010110",
  24471=>"111110100",
  24472=>"101101100",
  24473=>"000001010",
  24474=>"111110011",
  24475=>"110101100",
  24476=>"110111111",
  24477=>"001100101",
  24478=>"111010000",
  24479=>"010000111",
  24480=>"000101101",
  24481=>"111000100",
  24482=>"110110101",
  24483=>"010100001",
  24484=>"110000111",
  24485=>"111111111",
  24486=>"011010100",
  24487=>"010001100",
  24488=>"001010100",
  24489=>"001100010",
  24490=>"101001101",
  24491=>"100101110",
  24492=>"011001000",
  24493=>"111010010",
  24494=>"101111110",
  24495=>"001111000",
  24496=>"111101000",
  24497=>"100111111",
  24498=>"110001101",
  24499=>"111100010",
  24500=>"110001001",
  24501=>"110011110",
  24502=>"110001000",
  24503=>"000000111",
  24504=>"011111101",
  24505=>"110101100",
  24506=>"100101010",
  24507=>"101001000",
  24508=>"000100110",
  24509=>"110010000",
  24510=>"010000001",
  24511=>"110010110",
  24512=>"010010011",
  24513=>"100100011",
  24514=>"101010101",
  24515=>"110110011",
  24516=>"000101000",
  24517=>"001001001",
  24518=>"011001100",
  24519=>"100110010",
  24520=>"110110100",
  24521=>"101010010",
  24522=>"111000100",
  24523=>"000010100",
  24524=>"110111111",
  24525=>"100000000",
  24526=>"000010010",
  24527=>"001001100",
  24528=>"110010111",
  24529=>"100001000",
  24530=>"000001100",
  24531=>"110100100",
  24532=>"000010111",
  24533=>"101011110",
  24534=>"010100001",
  24535=>"100111111",
  24536=>"111110011",
  24537=>"011100011",
  24538=>"000000110",
  24539=>"111011001",
  24540=>"010110011",
  24541=>"101011101",
  24542=>"001011001",
  24543=>"111101101",
  24544=>"010111111",
  24545=>"011010101",
  24546=>"000000011",
  24547=>"111100111",
  24548=>"000000000",
  24549=>"000010000",
  24550=>"100100010",
  24551=>"111100000",
  24552=>"111010000",
  24553=>"110000100",
  24554=>"110001000",
  24555=>"000100111",
  24556=>"000110110",
  24557=>"000101000",
  24558=>"000011110",
  24559=>"000001110",
  24560=>"101111111",
  24561=>"110010101",
  24562=>"111101000",
  24563=>"100100100",
  24564=>"001000101",
  24565=>"100111001",
  24566=>"110011011",
  24567=>"100101001",
  24568=>"000000011",
  24569=>"010010111",
  24570=>"101111110",
  24571=>"111110110",
  24572=>"010111101",
  24573=>"101011001",
  24574=>"000110101",
  24575=>"110010011",
  24576=>"010000010",
  24577=>"001100010",
  24578=>"000101100",
  24579=>"000001110",
  24580=>"001111010",
  24581=>"111000000",
  24582=>"010100111",
  24583=>"011011000",
  24584=>"001001000",
  24585=>"000110000",
  24586=>"100010000",
  24587=>"100001011",
  24588=>"111100010",
  24589=>"011111111",
  24590=>"011111110",
  24591=>"011011110",
  24592=>"011010111",
  24593=>"100000011",
  24594=>"110011110",
  24595=>"111100000",
  24596=>"101111000",
  24597=>"001000000",
  24598=>"100010110",
  24599=>"101111000",
  24600=>"000001101",
  24601=>"111000100",
  24602=>"001001110",
  24603=>"001001111",
  24604=>"001000010",
  24605=>"001101101",
  24606=>"001101101",
  24607=>"000011111",
  24608=>"110000100",
  24609=>"100000101",
  24610=>"000001110",
  24611=>"001000001",
  24612=>"100010111",
  24613=>"110010001",
  24614=>"111100110",
  24615=>"001010001",
  24616=>"101000111",
  24617=>"100000011",
  24618=>"001111110",
  24619=>"101100011",
  24620=>"101001100",
  24621=>"010001110",
  24622=>"010010000",
  24623=>"110111001",
  24624=>"011100000",
  24625=>"011111100",
  24626=>"011100010",
  24627=>"100000001",
  24628=>"000010010",
  24629=>"110110010",
  24630=>"110111100",
  24631=>"111011101",
  24632=>"011000100",
  24633=>"111001000",
  24634=>"011000100",
  24635=>"101110111",
  24636=>"000010110",
  24637=>"100100110",
  24638=>"010011000",
  24639=>"000101000",
  24640=>"100110011",
  24641=>"001000100",
  24642=>"000000111",
  24643=>"000100100",
  24644=>"011100111",
  24645=>"001000110",
  24646=>"100010001",
  24647=>"101110101",
  24648=>"100100101",
  24649=>"110011111",
  24650=>"110111110",
  24651=>"001100001",
  24652=>"000100001",
  24653=>"110010101",
  24654=>"010011110",
  24655=>"111101101",
  24656=>"101101110",
  24657=>"111111000",
  24658=>"100011111",
  24659=>"010100111",
  24660=>"010101001",
  24661=>"100001010",
  24662=>"000011001",
  24663=>"001011010",
  24664=>"100110000",
  24665=>"011111110",
  24666=>"101110111",
  24667=>"000011001",
  24668=>"001100101",
  24669=>"001101101",
  24670=>"111011010",
  24671=>"000011100",
  24672=>"010011110",
  24673=>"100110001",
  24674=>"111101011",
  24675=>"001001100",
  24676=>"001011011",
  24677=>"010011011",
  24678=>"100000011",
  24679=>"000100110",
  24680=>"111000000",
  24681=>"000001000",
  24682=>"110100000",
  24683=>"011101111",
  24684=>"000101110",
  24685=>"010111111",
  24686=>"011001111",
  24687=>"001011001",
  24688=>"000111101",
  24689=>"111010000",
  24690=>"011100111",
  24691=>"011101010",
  24692=>"011110000",
  24693=>"000010011",
  24694=>"000000110",
  24695=>"101000101",
  24696=>"100010000",
  24697=>"111101111",
  24698=>"111100100",
  24699=>"111111111",
  24700=>"000000111",
  24701=>"000111111",
  24702=>"000000000",
  24703=>"100001101",
  24704=>"100100111",
  24705=>"000100101",
  24706=>"111101111",
  24707=>"000100111",
  24708=>"001101011",
  24709=>"000001100",
  24710=>"101110011",
  24711=>"101100101",
  24712=>"000100011",
  24713=>"011010001",
  24714=>"000001010",
  24715=>"100110110",
  24716=>"010111110",
  24717=>"101101111",
  24718=>"111110000",
  24719=>"101100100",
  24720=>"110010110",
  24721=>"101101011",
  24722=>"111100101",
  24723=>"101110000",
  24724=>"000000010",
  24725=>"000011110",
  24726=>"010010010",
  24727=>"110100111",
  24728=>"001011011",
  24729=>"010010010",
  24730=>"111101011",
  24731=>"010011000",
  24732=>"010011011",
  24733=>"100011100",
  24734=>"111001101",
  24735=>"010001000",
  24736=>"000000001",
  24737=>"111100001",
  24738=>"110010101",
  24739=>"110110000",
  24740=>"100100011",
  24741=>"000000101",
  24742=>"110011111",
  24743=>"011100010",
  24744=>"011000010",
  24745=>"000011001",
  24746=>"111111110",
  24747=>"111101110",
  24748=>"111101011",
  24749=>"110111101",
  24750=>"010000011",
  24751=>"100110110",
  24752=>"011010010",
  24753=>"100100001",
  24754=>"110001100",
  24755=>"100111101",
  24756=>"100100001",
  24757=>"111101111",
  24758=>"001110011",
  24759=>"001000100",
  24760=>"010111101",
  24761=>"011111100",
  24762=>"101010011",
  24763=>"000111001",
  24764=>"111110010",
  24765=>"001011011",
  24766=>"100101100",
  24767=>"101100110",
  24768=>"001101111",
  24769=>"111011110",
  24770=>"000000000",
  24771=>"000111001",
  24772=>"101001110",
  24773=>"110101111",
  24774=>"100011111",
  24775=>"101110000",
  24776=>"111101110",
  24777=>"111110011",
  24778=>"000100000",
  24779=>"111101001",
  24780=>"011010001",
  24781=>"001100000",
  24782=>"001110100",
  24783=>"010010111",
  24784=>"011110010",
  24785=>"111101001",
  24786=>"010011101",
  24787=>"111100000",
  24788=>"100010000",
  24789=>"111010000",
  24790=>"010110000",
  24791=>"110001101",
  24792=>"100111010",
  24793=>"101111111",
  24794=>"001001100",
  24795=>"101011010",
  24796=>"010100000",
  24797=>"101101111",
  24798=>"010000011",
  24799=>"001110111",
  24800=>"000011111",
  24801=>"111001100",
  24802=>"110101000",
  24803=>"100000100",
  24804=>"011001011",
  24805=>"110110000",
  24806=>"111010111",
  24807=>"101100101",
  24808=>"001001110",
  24809=>"100101111",
  24810=>"100110010",
  24811=>"111010100",
  24812=>"010100011",
  24813=>"111111101",
  24814=>"010101101",
  24815=>"101110001",
  24816=>"000000111",
  24817=>"110011111",
  24818=>"001100100",
  24819=>"001011111",
  24820=>"001010011",
  24821=>"000100111",
  24822=>"111111101",
  24823=>"011010110",
  24824=>"100101000",
  24825=>"111000110",
  24826=>"000110101",
  24827=>"011010110",
  24828=>"000000000",
  24829=>"110100000",
  24830=>"000000010",
  24831=>"001110100",
  24832=>"100000001",
  24833=>"101001110",
  24834=>"111000111",
  24835=>"011011010",
  24836=>"100010001",
  24837=>"011111011",
  24838=>"011110011",
  24839=>"101111000",
  24840=>"100110011",
  24841=>"100101001",
  24842=>"010101011",
  24843=>"000000011",
  24844=>"101011110",
  24845=>"010010010",
  24846=>"100101011",
  24847=>"000001111",
  24848=>"000110011",
  24849=>"001100111",
  24850=>"010001100",
  24851=>"101110001",
  24852=>"001010100",
  24853=>"100010110",
  24854=>"111111111",
  24855=>"010011000",
  24856=>"010111000",
  24857=>"010100111",
  24858=>"100110100",
  24859=>"000110011",
  24860=>"010101111",
  24861=>"001101100",
  24862=>"110100000",
  24863=>"000010011",
  24864=>"010010110",
  24865=>"000011111",
  24866=>"010111111",
  24867=>"000100001",
  24868=>"010101111",
  24869=>"110100111",
  24870=>"001001001",
  24871=>"010000110",
  24872=>"110001111",
  24873=>"000111010",
  24874=>"100111101",
  24875=>"110000010",
  24876=>"101100000",
  24877=>"000000010",
  24878=>"111010001",
  24879=>"010011010",
  24880=>"010110000",
  24881=>"111101011",
  24882=>"110010101",
  24883=>"100100111",
  24884=>"100101111",
  24885=>"011000010",
  24886=>"100001111",
  24887=>"111110010",
  24888=>"100111010",
  24889=>"100011101",
  24890=>"001010110",
  24891=>"111010011",
  24892=>"000110100",
  24893=>"111101001",
  24894=>"101001100",
  24895=>"111001011",
  24896=>"111001111",
  24897=>"010101001",
  24898=>"110101111",
  24899=>"000010010",
  24900=>"100100100",
  24901=>"011101100",
  24902=>"110101010",
  24903=>"001001010",
  24904=>"011100011",
  24905=>"010111100",
  24906=>"011000011",
  24907=>"000000000",
  24908=>"100110100",
  24909=>"111101111",
  24910=>"111010001",
  24911=>"010110001",
  24912=>"011011010",
  24913=>"101101110",
  24914=>"110111111",
  24915=>"000001000",
  24916=>"001000010",
  24917=>"101010101",
  24918=>"010101000",
  24919=>"111110100",
  24920=>"100001001",
  24921=>"011100011",
  24922=>"001000110",
  24923=>"001001100",
  24924=>"010100100",
  24925=>"100010011",
  24926=>"000100011",
  24927=>"001010100",
  24928=>"001111111",
  24929=>"100001111",
  24930=>"101000001",
  24931=>"010011111",
  24932=>"001011100",
  24933=>"111110011",
  24934=>"011101000",
  24935=>"111100010",
  24936=>"000010010",
  24937=>"011011010",
  24938=>"101011111",
  24939=>"010000101",
  24940=>"111110110",
  24941=>"110110010",
  24942=>"110110110",
  24943=>"001000101",
  24944=>"011001101",
  24945=>"010010110",
  24946=>"110011111",
  24947=>"011011100",
  24948=>"010010101",
  24949=>"000011000",
  24950=>"101000001",
  24951=>"001011111",
  24952=>"001010100",
  24953=>"000100011",
  24954=>"001001111",
  24955=>"111010000",
  24956=>"010000111",
  24957=>"011111101",
  24958=>"010110010",
  24959=>"101111111",
  24960=>"010111101",
  24961=>"001111111",
  24962=>"000011101",
  24963=>"001100011",
  24964=>"111100110",
  24965=>"110010100",
  24966=>"000000001",
  24967=>"111101101",
  24968=>"001100010",
  24969=>"001011100",
  24970=>"111100011",
  24971=>"111101001",
  24972=>"100001111",
  24973=>"100110110",
  24974=>"001101101",
  24975=>"000100001",
  24976=>"001110010",
  24977=>"111110111",
  24978=>"011100001",
  24979=>"010011011",
  24980=>"000101000",
  24981=>"011110111",
  24982=>"010001000",
  24983=>"110000000",
  24984=>"111010010",
  24985=>"010110111",
  24986=>"000010000",
  24987=>"100000000",
  24988=>"000011110",
  24989=>"110000100",
  24990=>"111110011",
  24991=>"110010010",
  24992=>"101010100",
  24993=>"011101000",
  24994=>"010111011",
  24995=>"110111000",
  24996=>"110011001",
  24997=>"110010001",
  24998=>"010100010",
  24999=>"100001001",
  25000=>"110111110",
  25001=>"011010100",
  25002=>"000101000",
  25003=>"100000001",
  25004=>"010101011",
  25005=>"010110111",
  25006=>"111101010",
  25007=>"001011100",
  25008=>"101001000",
  25009=>"111101111",
  25010=>"010011010",
  25011=>"011001100",
  25012=>"110010001",
  25013=>"010010001",
  25014=>"101010101",
  25015=>"100010100",
  25016=>"110111011",
  25017=>"000000100",
  25018=>"000100000",
  25019=>"110111100",
  25020=>"100100101",
  25021=>"001000000",
  25022=>"011101011",
  25023=>"010100000",
  25024=>"111100110",
  25025=>"111000101",
  25026=>"010000111",
  25027=>"011001000",
  25028=>"011101110",
  25029=>"111100100",
  25030=>"110111110",
  25031=>"010001010",
  25032=>"100001001",
  25033=>"000011100",
  25034=>"010100011",
  25035=>"010010010",
  25036=>"001111101",
  25037=>"011011001",
  25038=>"000100111",
  25039=>"001101001",
  25040=>"010110111",
  25041=>"111000111",
  25042=>"111010101",
  25043=>"111001110",
  25044=>"111001001",
  25045=>"111000010",
  25046=>"111111100",
  25047=>"011100000",
  25048=>"000110010",
  25049=>"110111000",
  25050=>"000000000",
  25051=>"010000010",
  25052=>"010110000",
  25053=>"101001110",
  25054=>"110000101",
  25055=>"100110000",
  25056=>"111111111",
  25057=>"100100000",
  25058=>"101111011",
  25059=>"101100011",
  25060=>"010100101",
  25061=>"111001111",
  25062=>"111011000",
  25063=>"011110010",
  25064=>"101010000",
  25065=>"010100111",
  25066=>"011100000",
  25067=>"100010100",
  25068=>"101001000",
  25069=>"111001110",
  25070=>"100001100",
  25071=>"100010101",
  25072=>"001001001",
  25073=>"111111010",
  25074=>"100000100",
  25075=>"010111111",
  25076=>"010011100",
  25077=>"111101001",
  25078=>"011111110",
  25079=>"000011011",
  25080=>"010101110",
  25081=>"010000110",
  25082=>"010111000",
  25083=>"000101011",
  25084=>"110110000",
  25085=>"111000010",
  25086=>"100011011",
  25087=>"110001001",
  25088=>"011001001",
  25089=>"111111111",
  25090=>"010101000",
  25091=>"100111100",
  25092=>"001010101",
  25093=>"110011001",
  25094=>"111000101",
  25095=>"111000111",
  25096=>"001011001",
  25097=>"000011000",
  25098=>"111000001",
  25099=>"000110010",
  25100=>"000111110",
  25101=>"101100011",
  25102=>"100001100",
  25103=>"010001111",
  25104=>"011111001",
  25105=>"111010001",
  25106=>"000100010",
  25107=>"100010101",
  25108=>"000011101",
  25109=>"010010010",
  25110=>"111000011",
  25111=>"110000010",
  25112=>"111110110",
  25113=>"101010111",
  25114=>"001011011",
  25115=>"110111111",
  25116=>"000101100",
  25117=>"000000001",
  25118=>"011101000",
  25119=>"111000100",
  25120=>"000000101",
  25121=>"010010101",
  25122=>"000000010",
  25123=>"111100011",
  25124=>"110110010",
  25125=>"011110000",
  25126=>"010000100",
  25127=>"111001101",
  25128=>"101000001",
  25129=>"110010111",
  25130=>"110100101",
  25131=>"000010101",
  25132=>"010001011",
  25133=>"101110110",
  25134=>"001010010",
  25135=>"111000101",
  25136=>"110001111",
  25137=>"110010010",
  25138=>"000001111",
  25139=>"010001001",
  25140=>"010110111",
  25141=>"111000010",
  25142=>"010011011",
  25143=>"100101100",
  25144=>"010111110",
  25145=>"101101111",
  25146=>"010011010",
  25147=>"000010001",
  25148=>"001101010",
  25149=>"010000100",
  25150=>"111010001",
  25151=>"110111011",
  25152=>"000000100",
  25153=>"011101000",
  25154=>"111101011",
  25155=>"101001001",
  25156=>"100011001",
  25157=>"101110011",
  25158=>"001011110",
  25159=>"001100100",
  25160=>"000000110",
  25161=>"001011111",
  25162=>"111011110",
  25163=>"111111000",
  25164=>"000010011",
  25165=>"011110011",
  25166=>"010001111",
  25167=>"110100111",
  25168=>"010000111",
  25169=>"100100010",
  25170=>"001001011",
  25171=>"111100000",
  25172=>"000110011",
  25173=>"010101101",
  25174=>"001011111",
  25175=>"010000100",
  25176=>"011111001",
  25177=>"000011101",
  25178=>"000000110",
  25179=>"010001000",
  25180=>"000110010",
  25181=>"000100101",
  25182=>"011000111",
  25183=>"001100101",
  25184=>"110111001",
  25185=>"100000011",
  25186=>"100001011",
  25187=>"001000001",
  25188=>"101110100",
  25189=>"001001011",
  25190=>"101100100",
  25191=>"010111101",
  25192=>"000001100",
  25193=>"100100011",
  25194=>"010110011",
  25195=>"011010111",
  25196=>"011100110",
  25197=>"001100001",
  25198=>"000110111",
  25199=>"101110111",
  25200=>"101001100",
  25201=>"100101000",
  25202=>"000001110",
  25203=>"000110001",
  25204=>"010110001",
  25205=>"000010110",
  25206=>"111111101",
  25207=>"111001110",
  25208=>"111000011",
  25209=>"111110101",
  25210=>"100010010",
  25211=>"001011101",
  25212=>"010000101",
  25213=>"010010001",
  25214=>"001001011",
  25215=>"011011110",
  25216=>"111011100",
  25217=>"000111100",
  25218=>"001011010",
  25219=>"111010100",
  25220=>"100100000",
  25221=>"110101101",
  25222=>"001100001",
  25223=>"111011010",
  25224=>"110001010",
  25225=>"011000101",
  25226=>"101110000",
  25227=>"001011111",
  25228=>"111101001",
  25229=>"010010000",
  25230=>"110000011",
  25231=>"100010100",
  25232=>"000010110",
  25233=>"111110111",
  25234=>"111011000",
  25235=>"011100101",
  25236=>"010010000",
  25237=>"111100001",
  25238=>"110011101",
  25239=>"100110101",
  25240=>"100101110",
  25241=>"011010010",
  25242=>"100101010",
  25243=>"011011001",
  25244=>"001000001",
  25245=>"000001110",
  25246=>"010101000",
  25247=>"001011110",
  25248=>"000010111",
  25249=>"110101101",
  25250=>"011110101",
  25251=>"011101101",
  25252=>"011111100",
  25253=>"011000000",
  25254=>"011101011",
  25255=>"000011000",
  25256=>"011100011",
  25257=>"000110000",
  25258=>"010100110",
  25259=>"110110000",
  25260=>"010100000",
  25261=>"111000001",
  25262=>"110101010",
  25263=>"011100110",
  25264=>"100101001",
  25265=>"110001101",
  25266=>"011111011",
  25267=>"111010010",
  25268=>"001001010",
  25269=>"101110110",
  25270=>"011010010",
  25271=>"000100001",
  25272=>"010001001",
  25273=>"000110101",
  25274=>"101010100",
  25275=>"011110001",
  25276=>"000001010",
  25277=>"100000011",
  25278=>"000101001",
  25279=>"011101000",
  25280=>"111111100",
  25281=>"011010010",
  25282=>"001101111",
  25283=>"111110000",
  25284=>"010000100",
  25285=>"101000001",
  25286=>"100111001",
  25287=>"010111010",
  25288=>"110100110",
  25289=>"011100010",
  25290=>"101010110",
  25291=>"000000100",
  25292=>"010000011",
  25293=>"111111001",
  25294=>"011010100",
  25295=>"010100000",
  25296=>"000010100",
  25297=>"100011001",
  25298=>"010100000",
  25299=>"100001000",
  25300=>"101111100",
  25301=>"101011111",
  25302=>"110101101",
  25303=>"111011000",
  25304=>"101000101",
  25305=>"000000010",
  25306=>"111101000",
  25307=>"101001000",
  25308=>"001011111",
  25309=>"001100100",
  25310=>"101101010",
  25311=>"011001100",
  25312=>"110100001",
  25313=>"100011010",
  25314=>"101111010",
  25315=>"110010010",
  25316=>"110100000",
  25317=>"100100101",
  25318=>"001001100",
  25319=>"011010101",
  25320=>"110011000",
  25321=>"100010001",
  25322=>"100001111",
  25323=>"010001101",
  25324=>"001001111",
  25325=>"111111111",
  25326=>"000111011",
  25327=>"010111000",
  25328=>"111111100",
  25329=>"111000100",
  25330=>"000001111",
  25331=>"000001011",
  25332=>"000010011",
  25333=>"111100100",
  25334=>"000011011",
  25335=>"010101000",
  25336=>"000000110",
  25337=>"011101101",
  25338=>"100010110",
  25339=>"011100000",
  25340=>"001001011",
  25341=>"010111110",
  25342=>"011011111",
  25343=>"100001110",
  25344=>"100000011",
  25345=>"111110100",
  25346=>"001011100",
  25347=>"010000110",
  25348=>"111011011",
  25349=>"001001111",
  25350=>"111001010",
  25351=>"001001011",
  25352=>"110111011",
  25353=>"111100000",
  25354=>"010010010",
  25355=>"000011100",
  25356=>"010011100",
  25357=>"111001010",
  25358=>"110010000",
  25359=>"101010011",
  25360=>"101000001",
  25361=>"111000110",
  25362=>"110010110",
  25363=>"111010001",
  25364=>"101011100",
  25365=>"011001101",
  25366=>"000010110",
  25367=>"010111110",
  25368=>"000011000",
  25369=>"000000110",
  25370=>"001010101",
  25371=>"000110001",
  25372=>"011011100",
  25373=>"000111011",
  25374=>"101111011",
  25375=>"000011110",
  25376=>"110111000",
  25377=>"110110110",
  25378=>"010000001",
  25379=>"001110111",
  25380=>"111110100",
  25381=>"101001011",
  25382=>"001011100",
  25383=>"111001010",
  25384=>"111100101",
  25385=>"111011011",
  25386=>"101111100",
  25387=>"010101101",
  25388=>"110100010",
  25389=>"100101001",
  25390=>"101110101",
  25391=>"101001010",
  25392=>"110100000",
  25393=>"110100101",
  25394=>"000110100",
  25395=>"010101100",
  25396=>"111101101",
  25397=>"010000110",
  25398=>"110001010",
  25399=>"111111011",
  25400=>"111101111",
  25401=>"001010000",
  25402=>"000000000",
  25403=>"110010011",
  25404=>"000011101",
  25405=>"000010001",
  25406=>"000101001",
  25407=>"111101001",
  25408=>"101000011",
  25409=>"100001001",
  25410=>"011011111",
  25411=>"111011100",
  25412=>"000010011",
  25413=>"100111110",
  25414=>"100110101",
  25415=>"101100001",
  25416=>"001001011",
  25417=>"100101110",
  25418=>"010100100",
  25419=>"101100110",
  25420=>"010100001",
  25421=>"101000101",
  25422=>"111010000",
  25423=>"010101100",
  25424=>"010111011",
  25425=>"100000101",
  25426=>"111000111",
  25427=>"100001110",
  25428=>"001010010",
  25429=>"011001001",
  25430=>"100111111",
  25431=>"101101011",
  25432=>"110111101",
  25433=>"011011101",
  25434=>"101010001",
  25435=>"110001111",
  25436=>"111011000",
  25437=>"010100110",
  25438=>"000000010",
  25439=>"110001011",
  25440=>"111111011",
  25441=>"101010110",
  25442=>"100101110",
  25443=>"111011011",
  25444=>"010111000",
  25445=>"010110001",
  25446=>"011011000",
  25447=>"001101001",
  25448=>"011000100",
  25449=>"000111101",
  25450=>"010100100",
  25451=>"001110101",
  25452=>"110011010",
  25453=>"001111001",
  25454=>"011100001",
  25455=>"011011011",
  25456=>"111010010",
  25457=>"011001011",
  25458=>"000101100",
  25459=>"110111101",
  25460=>"100011011",
  25461=>"100101100",
  25462=>"101011000",
  25463=>"001101001",
  25464=>"001001101",
  25465=>"101110111",
  25466=>"101001101",
  25467=>"110010111",
  25468=>"101011001",
  25469=>"001101111",
  25470=>"110010011",
  25471=>"110000011",
  25472=>"110000100",
  25473=>"001000010",
  25474=>"000011000",
  25475=>"101010000",
  25476=>"111001001",
  25477=>"100011001",
  25478=>"111010000",
  25479=>"010110010",
  25480=>"110011111",
  25481=>"100111001",
  25482=>"000011100",
  25483=>"100110011",
  25484=>"011001010",
  25485=>"100011000",
  25486=>"010010110",
  25487=>"001111110",
  25488=>"000110000",
  25489=>"100000100",
  25490=>"001001010",
  25491=>"111101101",
  25492=>"000001001",
  25493=>"101101001",
  25494=>"001000000",
  25495=>"000011000",
  25496=>"001111100",
  25497=>"111101010",
  25498=>"110100101",
  25499=>"011011001",
  25500=>"001011001",
  25501=>"000011110",
  25502=>"100001010",
  25503=>"000100101",
  25504=>"011000111",
  25505=>"001101110",
  25506=>"110110110",
  25507=>"101110011",
  25508=>"100010000",
  25509=>"101100110",
  25510=>"010111111",
  25511=>"110001001",
  25512=>"000111111",
  25513=>"111010111",
  25514=>"010011100",
  25515=>"110000010",
  25516=>"000101101",
  25517=>"000110110",
  25518=>"000011001",
  25519=>"111010001",
  25520=>"001001101",
  25521=>"111101001",
  25522=>"011110111",
  25523=>"000111111",
  25524=>"111011110",
  25525=>"101000000",
  25526=>"111110110",
  25527=>"001011001",
  25528=>"110100110",
  25529=>"101110100",
  25530=>"000010001",
  25531=>"000101000",
  25532=>"110010100",
  25533=>"000111100",
  25534=>"000100110",
  25535=>"101000000",
  25536=>"111110101",
  25537=>"101100001",
  25538=>"101110110",
  25539=>"000011000",
  25540=>"001111011",
  25541=>"011011001",
  25542=>"011001111",
  25543=>"011010111",
  25544=>"110000000",
  25545=>"011011110",
  25546=>"101000000",
  25547=>"010000010",
  25548=>"110001000",
  25549=>"001010001",
  25550=>"100011110",
  25551=>"001011111",
  25552=>"001101001",
  25553=>"110001010",
  25554=>"110011111",
  25555=>"010100110",
  25556=>"101101001",
  25557=>"011111100",
  25558=>"001100001",
  25559=>"110010000",
  25560=>"110110101",
  25561=>"000110011",
  25562=>"111111000",
  25563=>"001000010",
  25564=>"100111100",
  25565=>"000110000",
  25566=>"100011111",
  25567=>"001110101",
  25568=>"010110000",
  25569=>"111010010",
  25570=>"011001111",
  25571=>"001010001",
  25572=>"111000101",
  25573=>"011011011",
  25574=>"010111001",
  25575=>"000001001",
  25576=>"000001011",
  25577=>"011110010",
  25578=>"000111110",
  25579=>"001001110",
  25580=>"000001101",
  25581=>"010111100",
  25582=>"100000111",
  25583=>"001010001",
  25584=>"111001100",
  25585=>"111101010",
  25586=>"001010010",
  25587=>"100010000",
  25588=>"100011100",
  25589=>"010001111",
  25590=>"111001101",
  25591=>"110010011",
  25592=>"100110001",
  25593=>"001010100",
  25594=>"101000001",
  25595=>"111110100",
  25596=>"001111111",
  25597=>"011100011",
  25598=>"110001010",
  25599=>"010111011",
  25600=>"100000000",
  25601=>"011111001",
  25602=>"111000110",
  25603=>"110010111",
  25604=>"110000100",
  25605=>"101001101",
  25606=>"010100101",
  25607=>"000110111",
  25608=>"011010000",
  25609=>"010100010",
  25610=>"011011000",
  25611=>"010110111",
  25612=>"100101000",
  25613=>"000100001",
  25614=>"001100001",
  25615=>"010000001",
  25616=>"010011101",
  25617=>"110110010",
  25618=>"011110001",
  25619=>"000011101",
  25620=>"010000110",
  25621=>"101001101",
  25622=>"001110001",
  25623=>"011100011",
  25624=>"001111001",
  25625=>"001100001",
  25626=>"110011000",
  25627=>"111001011",
  25628=>"100110111",
  25629=>"110001110",
  25630=>"110100010",
  25631=>"011000001",
  25632=>"110011010",
  25633=>"110011110",
  25634=>"101110111",
  25635=>"011010011",
  25636=>"000000000",
  25637=>"000010001",
  25638=>"010100111",
  25639=>"111100110",
  25640=>"101111010",
  25641=>"011000000",
  25642=>"100110111",
  25643=>"111000101",
  25644=>"101101010",
  25645=>"100000100",
  25646=>"010010010",
  25647=>"010011010",
  25648=>"101100010",
  25649=>"001111010",
  25650=>"011100100",
  25651=>"110010011",
  25652=>"110101110",
  25653=>"000000010",
  25654=>"111111101",
  25655=>"000011001",
  25656=>"011101110",
  25657=>"111010111",
  25658=>"001001000",
  25659=>"111111000",
  25660=>"011010010",
  25661=>"000101000",
  25662=>"001010011",
  25663=>"000010101",
  25664=>"100001101",
  25665=>"011100000",
  25666=>"100001110",
  25667=>"000101001",
  25668=>"100111110",
  25669=>"101000001",
  25670=>"100101000",
  25671=>"101011001",
  25672=>"111001110",
  25673=>"011111011",
  25674=>"010010101",
  25675=>"110111000",
  25676=>"000111111",
  25677=>"111111100",
  25678=>"100110101",
  25679=>"010110111",
  25680=>"110100010",
  25681=>"111101111",
  25682=>"101010000",
  25683=>"100111100",
  25684=>"000010101",
  25685=>"011101001",
  25686=>"110001010",
  25687=>"010001000",
  25688=>"110000110",
  25689=>"101100100",
  25690=>"010010100",
  25691=>"110010100",
  25692=>"111110010",
  25693=>"010011101",
  25694=>"101110000",
  25695=>"001110011",
  25696=>"101111010",
  25697=>"000100100",
  25698=>"101001111",
  25699=>"000111000",
  25700=>"111010000",
  25701=>"110011010",
  25702=>"011110000",
  25703=>"001001100",
  25704=>"111010011",
  25705=>"001001001",
  25706=>"010011101",
  25707=>"110011111",
  25708=>"100100011",
  25709=>"110011100",
  25710=>"001001000",
  25711=>"010111001",
  25712=>"111100100",
  25713=>"010100001",
  25714=>"010001111",
  25715=>"110111000",
  25716=>"001111010",
  25717=>"101101111",
  25718=>"010010011",
  25719=>"100011101",
  25720=>"000100011",
  25721=>"000011001",
  25722=>"111001101",
  25723=>"100111001",
  25724=>"111011011",
  25725=>"011100000",
  25726=>"111010010",
  25727=>"010000000",
  25728=>"010010011",
  25729=>"111001000",
  25730=>"000110001",
  25731=>"001110000",
  25732=>"000111001",
  25733=>"110010100",
  25734=>"110110010",
  25735=>"110001011",
  25736=>"000000000",
  25737=>"001000110",
  25738=>"000110010",
  25739=>"001110010",
  25740=>"110110111",
  25741=>"000001100",
  25742=>"100100101",
  25743=>"010111111",
  25744=>"110010001",
  25745=>"011000001",
  25746=>"100101101",
  25747=>"110011010",
  25748=>"100110011",
  25749=>"100101101",
  25750=>"011111000",
  25751=>"000000111",
  25752=>"001100010",
  25753=>"010000010",
  25754=>"101001001",
  25755=>"010110010",
  25756=>"010101011",
  25757=>"001100000",
  25758=>"001110100",
  25759=>"111111010",
  25760=>"010000000",
  25761=>"001010000",
  25762=>"111101101",
  25763=>"001110111",
  25764=>"011110100",
  25765=>"101111000",
  25766=>"011101111",
  25767=>"001100111",
  25768=>"110000100",
  25769=>"100100000",
  25770=>"111110111",
  25771=>"101111010",
  25772=>"110111101",
  25773=>"111001101",
  25774=>"100000000",
  25775=>"100010011",
  25776=>"100100000",
  25777=>"000101001",
  25778=>"010110010",
  25779=>"000111000",
  25780=>"001001101",
  25781=>"011000000",
  25782=>"111110010",
  25783=>"011001000",
  25784=>"001001110",
  25785=>"100001101",
  25786=>"010000111",
  25787=>"110100101",
  25788=>"011011111",
  25789=>"110010111",
  25790=>"110000010",
  25791=>"110110011",
  25792=>"001011000",
  25793=>"110010000",
  25794=>"011011100",
  25795=>"100110000",
  25796=>"011000011",
  25797=>"011010001",
  25798=>"111110101",
  25799=>"010000001",
  25800=>"111110110",
  25801=>"110110101",
  25802=>"100011111",
  25803=>"001000011",
  25804=>"001001110",
  25805=>"111101111",
  25806=>"111110010",
  25807=>"111010010",
  25808=>"110101001",
  25809=>"110011001",
  25810=>"000111000",
  25811=>"100101110",
  25812=>"110000110",
  25813=>"010111010",
  25814=>"100001001",
  25815=>"011000110",
  25816=>"000011010",
  25817=>"011101000",
  25818=>"010010111",
  25819=>"011000011",
  25820=>"110000110",
  25821=>"101000101",
  25822=>"001000100",
  25823=>"101111110",
  25824=>"110110011",
  25825=>"100101101",
  25826=>"001100100",
  25827=>"110111111",
  25828=>"000011000",
  25829=>"011001010",
  25830=>"000001011",
  25831=>"010100100",
  25832=>"011111011",
  25833=>"010001111",
  25834=>"101001101",
  25835=>"111010111",
  25836=>"011101010",
  25837=>"101110100",
  25838=>"011001011",
  25839=>"000010000",
  25840=>"111011111",
  25841=>"111110001",
  25842=>"001110001",
  25843=>"000000101",
  25844=>"101111001",
  25845=>"110110110",
  25846=>"100110011",
  25847=>"111001001",
  25848=>"001101100",
  25849=>"010011010",
  25850=>"110010100",
  25851=>"000101100",
  25852=>"001101100",
  25853=>"100010001",
  25854=>"111101110",
  25855=>"100010110",
  25856=>"010100001",
  25857=>"011001110",
  25858=>"110101010",
  25859=>"000111100",
  25860=>"111100101",
  25861=>"110110011",
  25862=>"101010011",
  25863=>"010111011",
  25864=>"001101010",
  25865=>"000011101",
  25866=>"011110101",
  25867=>"100111111",
  25868=>"001011011",
  25869=>"010111001",
  25870=>"100110100",
  25871=>"000000001",
  25872=>"111111110",
  25873=>"101011001",
  25874=>"100010001",
  25875=>"000011011",
  25876=>"000100000",
  25877=>"001000000",
  25878=>"101111111",
  25879=>"000010100",
  25880=>"011101000",
  25881=>"111011001",
  25882=>"011100010",
  25883=>"011001111",
  25884=>"110000001",
  25885=>"011011110",
  25886=>"000110010",
  25887=>"110111111",
  25888=>"000110110",
  25889=>"101010100",
  25890=>"101001110",
  25891=>"001011111",
  25892=>"100100111",
  25893=>"001000010",
  25894=>"101001100",
  25895=>"111110011",
  25896=>"000101111",
  25897=>"000010001",
  25898=>"110010101",
  25899=>"001111111",
  25900=>"101011111",
  25901=>"000000000",
  25902=>"011000110",
  25903=>"011000011",
  25904=>"110001001",
  25905=>"010101111",
  25906=>"101100011",
  25907=>"110010100",
  25908=>"011000011",
  25909=>"001000100",
  25910=>"001101000",
  25911=>"011100101",
  25912=>"110000010",
  25913=>"010111001",
  25914=>"011111011",
  25915=>"000100010",
  25916=>"001000010",
  25917=>"101110000",
  25918=>"001110101",
  25919=>"010010001",
  25920=>"101000011",
  25921=>"001000000",
  25922=>"101110010",
  25923=>"000011011",
  25924=>"011101111",
  25925=>"101001100",
  25926=>"100010000",
  25927=>"101101100",
  25928=>"011110110",
  25929=>"011001101",
  25930=>"111110101",
  25931=>"011000000",
  25932=>"100001111",
  25933=>"000010100",
  25934=>"001111001",
  25935=>"111010011",
  25936=>"110100100",
  25937=>"100101010",
  25938=>"101101000",
  25939=>"110001001",
  25940=>"100110000",
  25941=>"010011001",
  25942=>"110110011",
  25943=>"111111101",
  25944=>"011010100",
  25945=>"011001100",
  25946=>"111010000",
  25947=>"000100110",
  25948=>"000011100",
  25949=>"111110001",
  25950=>"110000110",
  25951=>"000110010",
  25952=>"011111000",
  25953=>"111011011",
  25954=>"101111111",
  25955=>"000100011",
  25956=>"001111000",
  25957=>"001000000",
  25958=>"011001100",
  25959=>"100010010",
  25960=>"101001001",
  25961=>"111111101",
  25962=>"000111100",
  25963=>"011011010",
  25964=>"000001000",
  25965=>"001111011",
  25966=>"000101100",
  25967=>"110100011",
  25968=>"101010100",
  25969=>"101011111",
  25970=>"000100001",
  25971=>"001001000",
  25972=>"100111111",
  25973=>"010001010",
  25974=>"101011111",
  25975=>"000110010",
  25976=>"101001001",
  25977=>"011001100",
  25978=>"100010100",
  25979=>"100001110",
  25980=>"001010100",
  25981=>"111001011",
  25982=>"001010011",
  25983=>"111011110",
  25984=>"111010001",
  25985=>"111100110",
  25986=>"010111111",
  25987=>"000100001",
  25988=>"110101000",
  25989=>"111111110",
  25990=>"001010100",
  25991=>"111111110",
  25992=>"010110000",
  25993=>"101011110",
  25994=>"101001101",
  25995=>"100100011",
  25996=>"010110110",
  25997=>"011110110",
  25998=>"111010010",
  25999=>"110010010",
  26000=>"100101100",
  26001=>"011010011",
  26002=>"000011001",
  26003=>"100000000",
  26004=>"000101001",
  26005=>"111110110",
  26006=>"110111111",
  26007=>"000000101",
  26008=>"001000111",
  26009=>"010000101",
  26010=>"011011001",
  26011=>"010100101",
  26012=>"000011100",
  26013=>"000010010",
  26014=>"000010011",
  26015=>"100010011",
  26016=>"010111000",
  26017=>"110111000",
  26018=>"111100010",
  26019=>"100101100",
  26020=>"101011111",
  26021=>"100000101",
  26022=>"010000001",
  26023=>"001010110",
  26024=>"001010011",
  26025=>"110111000",
  26026=>"010010100",
  26027=>"001011011",
  26028=>"000011011",
  26029=>"111111011",
  26030=>"111000001",
  26031=>"101111111",
  26032=>"010011011",
  26033=>"101100101",
  26034=>"101000011",
  26035=>"011101111",
  26036=>"100000110",
  26037=>"000101011",
  26038=>"101100001",
  26039=>"110001011",
  26040=>"101100010",
  26041=>"100000001",
  26042=>"001001110",
  26043=>"001000111",
  26044=>"001011001",
  26045=>"111100001",
  26046=>"010001001",
  26047=>"001001001",
  26048=>"010110001",
  26049=>"111011101",
  26050=>"010110000",
  26051=>"100100100",
  26052=>"011000100",
  26053=>"111011011",
  26054=>"101101011",
  26055=>"011110111",
  26056=>"011011111",
  26057=>"100110101",
  26058=>"000111000",
  26059=>"101101010",
  26060=>"010100000",
  26061=>"111011011",
  26062=>"001111100",
  26063=>"011111111",
  26064=>"000111101",
  26065=>"111001110",
  26066=>"111100110",
  26067=>"101111001",
  26068=>"101111101",
  26069=>"011110010",
  26070=>"110111010",
  26071=>"111011001",
  26072=>"101111000",
  26073=>"110000101",
  26074=>"111000001",
  26075=>"000011010",
  26076=>"111110011",
  26077=>"001110000",
  26078=>"111011111",
  26079=>"000000000",
  26080=>"001011001",
  26081=>"110001100",
  26082=>"100001111",
  26083=>"110111110",
  26084=>"111100100",
  26085=>"000010001",
  26086=>"110010111",
  26087=>"010010011",
  26088=>"010101011",
  26089=>"000100110",
  26090=>"001111001",
  26091=>"001010010",
  26092=>"010110011",
  26093=>"100111100",
  26094=>"101011111",
  26095=>"000110001",
  26096=>"101100001",
  26097=>"001000011",
  26098=>"011100001",
  26099=>"000001111",
  26100=>"100000011",
  26101=>"001000010",
  26102=>"101001000",
  26103=>"111110101",
  26104=>"110101011",
  26105=>"111001101",
  26106=>"110100100",
  26107=>"010111010",
  26108=>"101110101",
  26109=>"000010111",
  26110=>"101101001",
  26111=>"010000111",
  26112=>"101010101",
  26113=>"110011110",
  26114=>"010100101",
  26115=>"101111100",
  26116=>"110100010",
  26117=>"101011011",
  26118=>"000111100",
  26119=>"110010100",
  26120=>"000000010",
  26121=>"110111010",
  26122=>"001101000",
  26123=>"000101111",
  26124=>"010000101",
  26125=>"100011100",
  26126=>"010000111",
  26127=>"001100011",
  26128=>"010000111",
  26129=>"001010010",
  26130=>"010110111",
  26131=>"011000001",
  26132=>"011000101",
  26133=>"000110101",
  26134=>"000100011",
  26135=>"010111100",
  26136=>"101011101",
  26137=>"100110001",
  26138=>"110011101",
  26139=>"101110101",
  26140=>"010010101",
  26141=>"100000110",
  26142=>"101011010",
  26143=>"101010011",
  26144=>"101101111",
  26145=>"010000110",
  26146=>"001110011",
  26147=>"000101110",
  26148=>"110101100",
  26149=>"000110001",
  26150=>"000011111",
  26151=>"101101001",
  26152=>"000010001",
  26153=>"110101100",
  26154=>"110111011",
  26155=>"011110100",
  26156=>"110110100",
  26157=>"000000101",
  26158=>"111110000",
  26159=>"000110011",
  26160=>"001101000",
  26161=>"001001011",
  26162=>"001010111",
  26163=>"001110100",
  26164=>"010101110",
  26165=>"111010001",
  26166=>"001001110",
  26167=>"110111111",
  26168=>"110111111",
  26169=>"111110100",
  26170=>"010101111",
  26171=>"000000010",
  26172=>"001100110",
  26173=>"101111001",
  26174=>"100011111",
  26175=>"001001010",
  26176=>"110000101",
  26177=>"000101100",
  26178=>"111010000",
  26179=>"100111100",
  26180=>"010000000",
  26181=>"011000001",
  26182=>"001110111",
  26183=>"110011001",
  26184=>"011110100",
  26185=>"000110100",
  26186=>"011000010",
  26187=>"001100100",
  26188=>"111010111",
  26189=>"011001001",
  26190=>"100001100",
  26191=>"110000110",
  26192=>"101100010",
  26193=>"100011101",
  26194=>"011011110",
  26195=>"111110000",
  26196=>"010001000",
  26197=>"101000011",
  26198=>"111010001",
  26199=>"010110100",
  26200=>"101101110",
  26201=>"011110011",
  26202=>"110010111",
  26203=>"001100111",
  26204=>"010011100",
  26205=>"010011101",
  26206=>"111111110",
  26207=>"011100111",
  26208=>"110001000",
  26209=>"100010010",
  26210=>"001010101",
  26211=>"101001001",
  26212=>"010001100",
  26213=>"000001100",
  26214=>"100111001",
  26215=>"011000111",
  26216=>"110010111",
  26217=>"011001011",
  26218=>"100101001",
  26219=>"111110101",
  26220=>"011100100",
  26221=>"111001011",
  26222=>"011000110",
  26223=>"110011101",
  26224=>"010101011",
  26225=>"000101000",
  26226=>"011010011",
  26227=>"111101011",
  26228=>"011101001",
  26229=>"010100001",
  26230=>"101100101",
  26231=>"000000001",
  26232=>"110101010",
  26233=>"000000101",
  26234=>"011110011",
  26235=>"111111101",
  26236=>"001011110",
  26237=>"010101100",
  26238=>"100001010",
  26239=>"001110001",
  26240=>"010010000",
  26241=>"001111000",
  26242=>"001100000",
  26243=>"011000000",
  26244=>"111000110",
  26245=>"100101101",
  26246=>"111001011",
  26247=>"101000010",
  26248=>"001010101",
  26249=>"000111000",
  26250=>"000000101",
  26251=>"000010010",
  26252=>"101011000",
  26253=>"000101111",
  26254=>"001010001",
  26255=>"111101000",
  26256=>"101011000",
  26257=>"110101101",
  26258=>"111000100",
  26259=>"001100111",
  26260=>"010100110",
  26261=>"000101100",
  26262=>"100011010",
  26263=>"000011000",
  26264=>"010100000",
  26265=>"110010100",
  26266=>"001110111",
  26267=>"100010001",
  26268=>"101001001",
  26269=>"101010001",
  26270=>"000011000",
  26271=>"000101110",
  26272=>"001111100",
  26273=>"100000000",
  26274=>"111111010",
  26275=>"101111111",
  26276=>"001101110",
  26277=>"110110001",
  26278=>"010001101",
  26279=>"110100011",
  26280=>"000011110",
  26281=>"101101011",
  26282=>"010000110",
  26283=>"010001100",
  26284=>"100110101",
  26285=>"110101101",
  26286=>"001010011",
  26287=>"110100010",
  26288=>"011000000",
  26289=>"000000100",
  26290=>"010011001",
  26291=>"101111100",
  26292=>"010110110",
  26293=>"011101100",
  26294=>"011000010",
  26295=>"100101011",
  26296=>"010100100",
  26297=>"101100100",
  26298=>"110110101",
  26299=>"100010100",
  26300=>"001111110",
  26301=>"001010011",
  26302=>"010000011",
  26303=>"111111011",
  26304=>"000001110",
  26305=>"010111100",
  26306=>"001011100",
  26307=>"100111011",
  26308=>"101000001",
  26309=>"101100111",
  26310=>"010111100",
  26311=>"001010011",
  26312=>"000011011",
  26313=>"011011001",
  26314=>"011001001",
  26315=>"001011010",
  26316=>"010011000",
  26317=>"010001000",
  26318=>"000011010",
  26319=>"001100010",
  26320=>"111100111",
  26321=>"111110000",
  26322=>"100000110",
  26323=>"000110111",
  26324=>"101101100",
  26325=>"011010110",
  26326=>"000110011",
  26327=>"111011110",
  26328=>"101000011",
  26329=>"000111101",
  26330=>"011100111",
  26331=>"010011001",
  26332=>"001101010",
  26333=>"000100000",
  26334=>"110001100",
  26335=>"010010011",
  26336=>"110000010",
  26337=>"000000010",
  26338=>"101110010",
  26339=>"111011001",
  26340=>"001011011",
  26341=>"110011110",
  26342=>"010000100",
  26343=>"111111010",
  26344=>"011000000",
  26345=>"101001011",
  26346=>"000001010",
  26347=>"100101001",
  26348=>"000110110",
  26349=>"100111101",
  26350=>"101001110",
  26351=>"011111101",
  26352=>"000111110",
  26353=>"011111111",
  26354=>"001100001",
  26355=>"101010111",
  26356=>"101111010",
  26357=>"100111101",
  26358=>"101110011",
  26359=>"010001010",
  26360=>"101100011",
  26361=>"010001011",
  26362=>"000100000",
  26363=>"110000100",
  26364=>"100111010",
  26365=>"000101001",
  26366=>"000111110",
  26367=>"110101101",
  26368=>"111101110",
  26369=>"010100010",
  26370=>"110011101",
  26371=>"001111001",
  26372=>"001010011",
  26373=>"110111000",
  26374=>"011101110",
  26375=>"001100010",
  26376=>"100110111",
  26377=>"101101111",
  26378=>"011100101",
  26379=>"011111111",
  26380=>"111101101",
  26381=>"011001110",
  26382=>"010111100",
  26383=>"110011001",
  26384=>"100101111",
  26385=>"011000001",
  26386=>"001001010",
  26387=>"001100101",
  26388=>"111000111",
  26389=>"100100111",
  26390=>"001101000",
  26391=>"100111010",
  26392=>"011111010",
  26393=>"010010111",
  26394=>"001111100",
  26395=>"100010111",
  26396=>"110001101",
  26397=>"100011101",
  26398=>"100101001",
  26399=>"000010001",
  26400=>"011000000",
  26401=>"001100000",
  26402=>"111010010",
  26403=>"100001110",
  26404=>"101100101",
  26405=>"111100111",
  26406=>"000101000",
  26407=>"101011100",
  26408=>"010101010",
  26409=>"001010010",
  26410=>"001000001",
  26411=>"101100010",
  26412=>"000001101",
  26413=>"000001010",
  26414=>"011010000",
  26415=>"000011011",
  26416=>"000011001",
  26417=>"000110010",
  26418=>"110011010",
  26419=>"101111010",
  26420=>"100101011",
  26421=>"000100101",
  26422=>"111111101",
  26423=>"110000010",
  26424=>"011100010",
  26425=>"110001110",
  26426=>"110111110",
  26427=>"001111101",
  26428=>"100110111",
  26429=>"010001010",
  26430=>"001001000",
  26431=>"110001011",
  26432=>"010010101",
  26433=>"111110101",
  26434=>"100100111",
  26435=>"011100000",
  26436=>"010011101",
  26437=>"101110010",
  26438=>"100101111",
  26439=>"110000000",
  26440=>"011110111",
  26441=>"011111101",
  26442=>"111110110",
  26443=>"101011110",
  26444=>"000010000",
  26445=>"100100010",
  26446=>"000101011",
  26447=>"110101110",
  26448=>"010011101",
  26449=>"011010100",
  26450=>"001111001",
  26451=>"100101000",
  26452=>"010001111",
  26453=>"011000001",
  26454=>"110000011",
  26455=>"001111110",
  26456=>"111010001",
  26457=>"000011001",
  26458=>"111100000",
  26459=>"000001011",
  26460=>"101001001",
  26461=>"011011101",
  26462=>"000111100",
  26463=>"110000111",
  26464=>"101011011",
  26465=>"110010100",
  26466=>"000100110",
  26467=>"100000001",
  26468=>"011001110",
  26469=>"111100010",
  26470=>"111110010",
  26471=>"000000010",
  26472=>"110010110",
  26473=>"000011011",
  26474=>"010001110",
  26475=>"000101000",
  26476=>"000000101",
  26477=>"000010110",
  26478=>"111010010",
  26479=>"110000010",
  26480=>"111100001",
  26481=>"001111111",
  26482=>"101001111",
  26483=>"001011001",
  26484=>"011110000",
  26485=>"101000000",
  26486=>"101111001",
  26487=>"010111110",
  26488=>"101100100",
  26489=>"101001111",
  26490=>"010011011",
  26491=>"001100010",
  26492=>"000100000",
  26493=>"111011010",
  26494=>"000001111",
  26495=>"100000001",
  26496=>"111110001",
  26497=>"011111111",
  26498=>"011000000",
  26499=>"110101001",
  26500=>"100001000",
  26501=>"010011010",
  26502=>"000010111",
  26503=>"100100111",
  26504=>"001001110",
  26505=>"011010100",
  26506=>"100111111",
  26507=>"110101011",
  26508=>"100110001",
  26509=>"110000000",
  26510=>"111011000",
  26511=>"000011100",
  26512=>"111111010",
  26513=>"000001111",
  26514=>"111000101",
  26515=>"101001110",
  26516=>"010110101",
  26517=>"100010010",
  26518=>"001100100",
  26519=>"011110100",
  26520=>"100010111",
  26521=>"111001101",
  26522=>"011010000",
  26523=>"100111000",
  26524=>"100000001",
  26525=>"101101000",
  26526=>"011001101",
  26527=>"000010001",
  26528=>"111001100",
  26529=>"111110001",
  26530=>"001010000",
  26531=>"001000101",
  26532=>"101000011",
  26533=>"000111101",
  26534=>"010110001",
  26535=>"101010111",
  26536=>"111111111",
  26537=>"011111101",
  26538=>"000000000",
  26539=>"011111011",
  26540=>"010011011",
  26541=>"101110101",
  26542=>"101111000",
  26543=>"011111101",
  26544=>"110101011",
  26545=>"111001100",
  26546=>"010111101",
  26547=>"100001010",
  26548=>"100010100",
  26549=>"110000001",
  26550=>"000001101",
  26551=>"110100010",
  26552=>"011111111",
  26553=>"101111111",
  26554=>"010001100",
  26555=>"001100001",
  26556=>"001011110",
  26557=>"100111100",
  26558=>"110000110",
  26559=>"010000110",
  26560=>"101000000",
  26561=>"000010010",
  26562=>"110001000",
  26563=>"000001000",
  26564=>"111111010",
  26565=>"000000010",
  26566=>"001000010",
  26567=>"001100011",
  26568=>"001000110",
  26569=>"111000010",
  26570=>"000110000",
  26571=>"000010011",
  26572=>"000100100",
  26573=>"101100001",
  26574=>"011100010",
  26575=>"101110101",
  26576=>"011000001",
  26577=>"001101101",
  26578=>"111110101",
  26579=>"000101000",
  26580=>"110010011",
  26581=>"101100011",
  26582=>"011001011",
  26583=>"010011011",
  26584=>"001110110",
  26585=>"010111011",
  26586=>"001100110",
  26587=>"111010001",
  26588=>"100100111",
  26589=>"100111000",
  26590=>"001011000",
  26591=>"111011001",
  26592=>"101001111",
  26593=>"100111101",
  26594=>"101010100",
  26595=>"111001110",
  26596=>"111110111",
  26597=>"000100010",
  26598=>"011000111",
  26599=>"001000000",
  26600=>"011000001",
  26601=>"001100111",
  26602=>"111001011",
  26603=>"011111000",
  26604=>"001101000",
  26605=>"110100100",
  26606=>"110001011",
  26607=>"001101100",
  26608=>"111000000",
  26609=>"000000000",
  26610=>"001110110",
  26611=>"100011011",
  26612=>"111101011",
  26613=>"001100100",
  26614=>"111100001",
  26615=>"100000010",
  26616=>"000000000",
  26617=>"011000001",
  26618=>"001000000",
  26619=>"010010000",
  26620=>"101000001",
  26621=>"100011011",
  26622=>"000010010",
  26623=>"101100100",
  26624=>"010101000",
  26625=>"111101011",
  26626=>"001000100",
  26627=>"011111111",
  26628=>"010000000",
  26629=>"011110100",
  26630=>"110101110",
  26631=>"001111101",
  26632=>"101000101",
  26633=>"111111011",
  26634=>"011111111",
  26635=>"110001010",
  26636=>"101001000",
  26637=>"110111000",
  26638=>"110101011",
  26639=>"001111010",
  26640=>"100001010",
  26641=>"110011000",
  26642=>"011111011",
  26643=>"110111010",
  26644=>"111011111",
  26645=>"001101000",
  26646=>"001101000",
  26647=>"001010000",
  26648=>"110000101",
  26649=>"100001011",
  26650=>"101001001",
  26651=>"111000011",
  26652=>"100100100",
  26653=>"001000101",
  26654=>"111110101",
  26655=>"011000010",
  26656=>"111000100",
  26657=>"101111111",
  26658=>"001110000",
  26659=>"110010100",
  26660=>"100011110",
  26661=>"001000110",
  26662=>"100010111",
  26663=>"110010011",
  26664=>"110001001",
  26665=>"001111100",
  26666=>"011110010",
  26667=>"010001010",
  26668=>"111101010",
  26669=>"110000100",
  26670=>"000000011",
  26671=>"111100000",
  26672=>"111001111",
  26673=>"001111100",
  26674=>"011001100",
  26675=>"101001110",
  26676=>"111010110",
  26677=>"000100010",
  26678=>"010001100",
  26679=>"001010010",
  26680=>"111100111",
  26681=>"001110011",
  26682=>"100101010",
  26683=>"110100000",
  26684=>"111101010",
  26685=>"000011111",
  26686=>"100000001",
  26687=>"110111011",
  26688=>"111001101",
  26689=>"000001100",
  26690=>"010010000",
  26691=>"101100000",
  26692=>"000010010",
  26693=>"111001000",
  26694=>"100100010",
  26695=>"101101010",
  26696=>"000110100",
  26697=>"000001011",
  26698=>"000111100",
  26699=>"110100010",
  26700=>"010100111",
  26701=>"001111000",
  26702=>"001111101",
  26703=>"011000110",
  26704=>"001010010",
  26705=>"000010000",
  26706=>"111100110",
  26707=>"100011111",
  26708=>"111111100",
  26709=>"010011111",
  26710=>"110010110",
  26711=>"110011101",
  26712=>"100101101",
  26713=>"111111100",
  26714=>"010000111",
  26715=>"110000111",
  26716=>"000100000",
  26717=>"000100011",
  26718=>"001010000",
  26719=>"110011011",
  26720=>"000000101",
  26721=>"000111110",
  26722=>"100001011",
  26723=>"110001111",
  26724=>"010110000",
  26725=>"100011101",
  26726=>"111010111",
  26727=>"110101000",
  26728=>"100100100",
  26729=>"000011111",
  26730=>"001101100",
  26731=>"001111111",
  26732=>"111000101",
  26733=>"001001111",
  26734=>"000100000",
  26735=>"001011011",
  26736=>"111011101",
  26737=>"001000111",
  26738=>"101110100",
  26739=>"010100111",
  26740=>"000010111",
  26741=>"111011011",
  26742=>"100110101",
  26743=>"000001010",
  26744=>"000100111",
  26745=>"110001001",
  26746=>"011110111",
  26747=>"001101010",
  26748=>"010110001",
  26749=>"111110101",
  26750=>"111000010",
  26751=>"000000101",
  26752=>"001110101",
  26753=>"111001110",
  26754=>"100000000",
  26755=>"000000110",
  26756=>"001100000",
  26757=>"011110111",
  26758=>"101011001",
  26759=>"101101011",
  26760=>"110000011",
  26761=>"001101001",
  26762=>"011001101",
  26763=>"111111111",
  26764=>"010011111",
  26765=>"100001101",
  26766=>"000010000",
  26767=>"100000000",
  26768=>"001010101",
  26769=>"011001011",
  26770=>"010010011",
  26771=>"100111110",
  26772=>"100010111",
  26773=>"100110111",
  26774=>"001100010",
  26775=>"111001001",
  26776=>"100001010",
  26777=>"110011011",
  26778=>"001110111",
  26779=>"000111011",
  26780=>"111000110",
  26781=>"101000101",
  26782=>"010000010",
  26783=>"001101100",
  26784=>"010101001",
  26785=>"000011101",
  26786=>"011110110",
  26787=>"111011111",
  26788=>"010000000",
  26789=>"100111100",
  26790=>"100101000",
  26791=>"111101101",
  26792=>"001000111",
  26793=>"011111001",
  26794=>"010011001",
  26795=>"000000000",
  26796=>"010001110",
  26797=>"011001111",
  26798=>"010100110",
  26799=>"110100010",
  26800=>"010000011",
  26801=>"010101110",
  26802=>"011010101",
  26803=>"010010000",
  26804=>"111111101",
  26805=>"100101111",
  26806=>"101100011",
  26807=>"001100011",
  26808=>"001110010",
  26809=>"111111010",
  26810=>"001011010",
  26811=>"000111111",
  26812=>"010010100",
  26813=>"100111010",
  26814=>"011000100",
  26815=>"111111000",
  26816=>"000011110",
  26817=>"001101111",
  26818=>"111111101",
  26819=>"101010010",
  26820=>"111011100",
  26821=>"010011010",
  26822=>"100101100",
  26823=>"100100100",
  26824=>"101111001",
  26825=>"100000100",
  26826=>"111111111",
  26827=>"000110010",
  26828=>"010110101",
  26829=>"011000100",
  26830=>"101110100",
  26831=>"011001111",
  26832=>"111000000",
  26833=>"101010111",
  26834=>"100000100",
  26835=>"100001110",
  26836=>"111111111",
  26837=>"011011110",
  26838=>"010000100",
  26839=>"000110001",
  26840=>"100010001",
  26841=>"000100010",
  26842=>"001101010",
  26843=>"001110000",
  26844=>"000110100",
  26845=>"001111000",
  26846=>"110010110",
  26847=>"100110001",
  26848=>"010101100",
  26849=>"111111111",
  26850=>"001000001",
  26851=>"100010011",
  26852=>"101001000",
  26853=>"100100001",
  26854=>"010010100",
  26855=>"011100111",
  26856=>"011111001",
  26857=>"100101111",
  26858=>"000011000",
  26859=>"101111010",
  26860=>"110110011",
  26861=>"000011010",
  26862=>"111011011",
  26863=>"010110111",
  26864=>"010101000",
  26865=>"101101100",
  26866=>"001011100",
  26867=>"100101101",
  26868=>"001111010",
  26869=>"100001010",
  26870=>"111110000",
  26871=>"110000110",
  26872=>"100110011",
  26873=>"110011100",
  26874=>"000000001",
  26875=>"100010110",
  26876=>"110000100",
  26877=>"110010100",
  26878=>"101110000",
  26879=>"110111000",
  26880=>"110111010",
  26881=>"000101011",
  26882=>"101011001",
  26883=>"011101111",
  26884=>"010101010",
  26885=>"110000011",
  26886=>"000111110",
  26887=>"001011111",
  26888=>"011000011",
  26889=>"010000011",
  26890=>"010011111",
  26891=>"111110111",
  26892=>"100110110",
  26893=>"100101001",
  26894=>"101111000",
  26895=>"000111010",
  26896=>"100100010",
  26897=>"111001101",
  26898=>"110011110",
  26899=>"011110100",
  26900=>"001000000",
  26901=>"110001110",
  26902=>"010000001",
  26903=>"010111001",
  26904=>"011010110",
  26905=>"010111001",
  26906=>"010001011",
  26907=>"100100001",
  26908=>"101011011",
  26909=>"111111110",
  26910=>"100101001",
  26911=>"010000101",
  26912=>"000000000",
  26913=>"110011111",
  26914=>"111100000",
  26915=>"011000010",
  26916=>"110010010",
  26917=>"100001111",
  26918=>"011101001",
  26919=>"001000100",
  26920=>"001100110",
  26921=>"110010000",
  26922=>"011111011",
  26923=>"100111110",
  26924=>"011110101",
  26925=>"001100000",
  26926=>"000001000",
  26927=>"100101111",
  26928=>"111100011",
  26929=>"101111011",
  26930=>"010111010",
  26931=>"110101110",
  26932=>"011100011",
  26933=>"101000010",
  26934=>"110011011",
  26935=>"011011100",
  26936=>"010100000",
  26937=>"010110110",
  26938=>"110011010",
  26939=>"010110111",
  26940=>"101001100",
  26941=>"011000010",
  26942=>"111001000",
  26943=>"110010101",
  26944=>"110110101",
  26945=>"010010011",
  26946=>"111001001",
  26947=>"111101111",
  26948=>"001000111",
  26949=>"111010111",
  26950=>"110001011",
  26951=>"111000011",
  26952=>"100110101",
  26953=>"100110011",
  26954=>"100110000",
  26955=>"110010110",
  26956=>"100010011",
  26957=>"111011111",
  26958=>"100010010",
  26959=>"101101101",
  26960=>"000010111",
  26961=>"100100000",
  26962=>"001000010",
  26963=>"010110011",
  26964=>"011010010",
  26965=>"111110100",
  26966=>"001110100",
  26967=>"010111011",
  26968=>"100101111",
  26969=>"111100100",
  26970=>"001001111",
  26971=>"111001110",
  26972=>"000101110",
  26973=>"110100110",
  26974=>"010101001",
  26975=>"000001001",
  26976=>"001000000",
  26977=>"011100100",
  26978=>"011111001",
  26979=>"100110111",
  26980=>"101011100",
  26981=>"100001001",
  26982=>"001000001",
  26983=>"000001010",
  26984=>"110010111",
  26985=>"001100100",
  26986=>"011000101",
  26987=>"100000001",
  26988=>"110101011",
  26989=>"010111000",
  26990=>"100110011",
  26991=>"000001001",
  26992=>"111001101",
  26993=>"101111011",
  26994=>"110100000",
  26995=>"001101110",
  26996=>"010111010",
  26997=>"110011100",
  26998=>"111111110",
  26999=>"001101100",
  27000=>"001011000",
  27001=>"010001000",
  27002=>"000110101",
  27003=>"100011110",
  27004=>"001100011",
  27005=>"100110111",
  27006=>"101110001",
  27007=>"011000000",
  27008=>"000100101",
  27009=>"011110100",
  27010=>"111111100",
  27011=>"100011001",
  27012=>"101001100",
  27013=>"011111110",
  27014=>"001101110",
  27015=>"001010000",
  27016=>"101000000",
  27017=>"111000100",
  27018=>"100010110",
  27019=>"111011110",
  27020=>"001011101",
  27021=>"110011110",
  27022=>"110000101",
  27023=>"001001001",
  27024=>"100000111",
  27025=>"100011100",
  27026=>"111000110",
  27027=>"011001100",
  27028=>"111011101",
  27029=>"001100001",
  27030=>"101111111",
  27031=>"100010001",
  27032=>"111100010",
  27033=>"101101101",
  27034=>"110101110",
  27035=>"000101110",
  27036=>"000101010",
  27037=>"000101010",
  27038=>"110010011",
  27039=>"100110100",
  27040=>"000000000",
  27041=>"111011000",
  27042=>"111000001",
  27043=>"010100011",
  27044=>"100001100",
  27045=>"001011001",
  27046=>"111100010",
  27047=>"101010101",
  27048=>"111001011",
  27049=>"000000010",
  27050=>"010000011",
  27051=>"010011110",
  27052=>"111001101",
  27053=>"101001010",
  27054=>"000010011",
  27055=>"101111110",
  27056=>"110000001",
  27057=>"101111001",
  27058=>"010101011",
  27059=>"100001011",
  27060=>"000001101",
  27061=>"001101001",
  27062=>"100101111",
  27063=>"110101001",
  27064=>"011000000",
  27065=>"100101010",
  27066=>"111010000",
  27067=>"001011010",
  27068=>"000010100",
  27069=>"110100010",
  27070=>"101000011",
  27071=>"001011100",
  27072=>"100011110",
  27073=>"001000101",
  27074=>"110101001",
  27075=>"011110100",
  27076=>"100001101",
  27077=>"001100010",
  27078=>"101100100",
  27079=>"101111001",
  27080=>"010001110",
  27081=>"010010001",
  27082=>"000000111",
  27083=>"111011001",
  27084=>"010111110",
  27085=>"011010000",
  27086=>"001000100",
  27087=>"010101011",
  27088=>"110111001",
  27089=>"101110101",
  27090=>"000001001",
  27091=>"000001011",
  27092=>"101101101",
  27093=>"110010011",
  27094=>"000101001",
  27095=>"101001011",
  27096=>"000111001",
  27097=>"101101100",
  27098=>"110101100",
  27099=>"000011011",
  27100=>"011100001",
  27101=>"001010101",
  27102=>"100111010",
  27103=>"000001000",
  27104=>"010101001",
  27105=>"000011110",
  27106=>"101100101",
  27107=>"011110100",
  27108=>"000100011",
  27109=>"010010000",
  27110=>"011000100",
  27111=>"011001010",
  27112=>"001011000",
  27113=>"000100111",
  27114=>"100111011",
  27115=>"011001101",
  27116=>"010111011",
  27117=>"100001010",
  27118=>"010010011",
  27119=>"001110000",
  27120=>"101011001",
  27121=>"011111110",
  27122=>"011100101",
  27123=>"101110100",
  27124=>"110010101",
  27125=>"110010101",
  27126=>"001110110",
  27127=>"110101010",
  27128=>"100000100",
  27129=>"110100111",
  27130=>"111100100",
  27131=>"101001101",
  27132=>"010010100",
  27133=>"111100001",
  27134=>"111111001",
  27135=>"101101111",
  27136=>"000000001",
  27137=>"001011000",
  27138=>"111001001",
  27139=>"001000000",
  27140=>"100011001",
  27141=>"001001101",
  27142=>"010000001",
  27143=>"010100010",
  27144=>"101000000",
  27145=>"101110100",
  27146=>"011010011",
  27147=>"110001101",
  27148=>"110011100",
  27149=>"001111011",
  27150=>"101000000",
  27151=>"100111000",
  27152=>"111001010",
  27153=>"100111111",
  27154=>"000100000",
  27155=>"100000101",
  27156=>"100000100",
  27157=>"011100101",
  27158=>"000000100",
  27159=>"011100110",
  27160=>"000010100",
  27161=>"001011110",
  27162=>"000000010",
  27163=>"010111110",
  27164=>"110100001",
  27165=>"110001110",
  27166=>"100011001",
  27167=>"111011001",
  27168=>"001001101",
  27169=>"110011010",
  27170=>"001100000",
  27171=>"000010000",
  27172=>"100110110",
  27173=>"101000100",
  27174=>"100011011",
  27175=>"010110000",
  27176=>"100110101",
  27177=>"111110011",
  27178=>"011101110",
  27179=>"001110110",
  27180=>"000101101",
  27181=>"100001000",
  27182=>"001111100",
  27183=>"101100110",
  27184=>"000101010",
  27185=>"101101101",
  27186=>"011001110",
  27187=>"110101000",
  27188=>"100101001",
  27189=>"010001001",
  27190=>"011010011",
  27191=>"011011000",
  27192=>"110100100",
  27193=>"000001000",
  27194=>"110111000",
  27195=>"000000110",
  27196=>"011001100",
  27197=>"011000010",
  27198=>"100001111",
  27199=>"101110000",
  27200=>"111100011",
  27201=>"110011010",
  27202=>"000100101",
  27203=>"110011000",
  27204=>"101111010",
  27205=>"110011011",
  27206=>"101110010",
  27207=>"000100000",
  27208=>"100001000",
  27209=>"111011001",
  27210=>"011000111",
  27211=>"001100000",
  27212=>"011111101",
  27213=>"000010000",
  27214=>"101101101",
  27215=>"110110000",
  27216=>"011010101",
  27217=>"100110001",
  27218=>"011100101",
  27219=>"001010010",
  27220=>"000011010",
  27221=>"010010011",
  27222=>"111011011",
  27223=>"010010110",
  27224=>"001111011",
  27225=>"000011111",
  27226=>"110101011",
  27227=>"101111000",
  27228=>"110110111",
  27229=>"111101101",
  27230=>"101111001",
  27231=>"111010000",
  27232=>"100111000",
  27233=>"110001100",
  27234=>"101001000",
  27235=>"111001010",
  27236=>"001011100",
  27237=>"000010000",
  27238=>"111010010",
  27239=>"111111010",
  27240=>"011101001",
  27241=>"001101000",
  27242=>"111010100",
  27243=>"111101100",
  27244=>"001101110",
  27245=>"111100100",
  27246=>"100111101",
  27247=>"110100001",
  27248=>"000010010",
  27249=>"001000100",
  27250=>"011010001",
  27251=>"111001111",
  27252=>"110010100",
  27253=>"011000110",
  27254=>"101111001",
  27255=>"010111111",
  27256=>"010010100",
  27257=>"000000010",
  27258=>"100100101",
  27259=>"110111100",
  27260=>"100011110",
  27261=>"100010101",
  27262=>"101111101",
  27263=>"101000001",
  27264=>"001001101",
  27265=>"001100110",
  27266=>"011001100",
  27267=>"010100111",
  27268=>"010110110",
  27269=>"111101100",
  27270=>"001001001",
  27271=>"101111110",
  27272=>"101000000",
  27273=>"110001111",
  27274=>"011010100",
  27275=>"001000001",
  27276=>"011100011",
  27277=>"000000111",
  27278=>"010000000",
  27279=>"000001100",
  27280=>"000111011",
  27281=>"011011001",
  27282=>"001010001",
  27283=>"010001110",
  27284=>"111100001",
  27285=>"100100010",
  27286=>"110100110",
  27287=>"010100110",
  27288=>"100101011",
  27289=>"010110100",
  27290=>"011000111",
  27291=>"000101001",
  27292=>"011011011",
  27293=>"110111001",
  27294=>"111010101",
  27295=>"101110010",
  27296=>"001010111",
  27297=>"011011110",
  27298=>"110111000",
  27299=>"000110000",
  27300=>"010010101",
  27301=>"101011100",
  27302=>"110101011",
  27303=>"100000111",
  27304=>"001111101",
  27305=>"100111011",
  27306=>"001101000",
  27307=>"101010011",
  27308=>"100110100",
  27309=>"111110111",
  27310=>"111001010",
  27311=>"011010100",
  27312=>"001000111",
  27313=>"100011000",
  27314=>"101111100",
  27315=>"001100000",
  27316=>"010011010",
  27317=>"010001001",
  27318=>"101001100",
  27319=>"000000111",
  27320=>"111101010",
  27321=>"010111110",
  27322=>"010111100",
  27323=>"000100000",
  27324=>"010011111",
  27325=>"110111111",
  27326=>"001001100",
  27327=>"011111101",
  27328=>"110010100",
  27329=>"011101001",
  27330=>"001011011",
  27331=>"111111110",
  27332=>"011011111",
  27333=>"100001010",
  27334=>"100111000",
  27335=>"101000111",
  27336=>"011101010",
  27337=>"101101111",
  27338=>"001011000",
  27339=>"010000101",
  27340=>"100100110",
  27341=>"100100010",
  27342=>"110000000",
  27343=>"000111010",
  27344=>"111100001",
  27345=>"000000000",
  27346=>"101111001",
  27347=>"011001000",
  27348=>"000101011",
  27349=>"101101000",
  27350=>"101000110",
  27351=>"111001110",
  27352=>"001110110",
  27353=>"110011000",
  27354=>"110111111",
  27355=>"011010001",
  27356=>"101110011",
  27357=>"010000111",
  27358=>"011100111",
  27359=>"111101011",
  27360=>"001000001",
  27361=>"000110110",
  27362=>"101110011",
  27363=>"010110011",
  27364=>"100101100",
  27365=>"011001001",
  27366=>"110010111",
  27367=>"011111000",
  27368=>"100000111",
  27369=>"101100000",
  27370=>"001011000",
  27371=>"000000011",
  27372=>"010011101",
  27373=>"110101100",
  27374=>"101100011",
  27375=>"010001100",
  27376=>"101110010",
  27377=>"001011110",
  27378=>"101001101",
  27379=>"000010110",
  27380=>"011111000",
  27381=>"011011111",
  27382=>"111010111",
  27383=>"010000010",
  27384=>"010111101",
  27385=>"001110111",
  27386=>"000001111",
  27387=>"001010000",
  27388=>"011111111",
  27389=>"101010101",
  27390=>"011011110",
  27391=>"001101000",
  27392=>"110101000",
  27393=>"111000011",
  27394=>"110010111",
  27395=>"100010000",
  27396=>"011010001",
  27397=>"010100110",
  27398=>"010110110",
  27399=>"000000010",
  27400=>"111000001",
  27401=>"111110101",
  27402=>"001001110",
  27403=>"010010110",
  27404=>"110100000",
  27405=>"010001100",
  27406=>"101101101",
  27407=>"000000011",
  27408=>"111111011",
  27409=>"110010100",
  27410=>"101001111",
  27411=>"001101010",
  27412=>"111111110",
  27413=>"110001010",
  27414=>"110110000",
  27415=>"011010000",
  27416=>"100000111",
  27417=>"111101001",
  27418=>"000110010",
  27419=>"111111101",
  27420=>"010100101",
  27421=>"101010110",
  27422=>"111001001",
  27423=>"111111111",
  27424=>"001010001",
  27425=>"000000011",
  27426=>"000101101",
  27427=>"000111111",
  27428=>"111101110",
  27429=>"100011000",
  27430=>"010000001",
  27431=>"011010001",
  27432=>"101101110",
  27433=>"001011111",
  27434=>"001001001",
  27435=>"100011110",
  27436=>"111010000",
  27437=>"101111110",
  27438=>"111100010",
  27439=>"110111100",
  27440=>"001001111",
  27441=>"100010101",
  27442=>"111011010",
  27443=>"000111011",
  27444=>"011011111",
  27445=>"110111010",
  27446=>"101100101",
  27447=>"001111111",
  27448=>"111100000",
  27449=>"101010001",
  27450=>"011100101",
  27451=>"001011010",
  27452=>"010000010",
  27453=>"101011001",
  27454=>"101101011",
  27455=>"011100011",
  27456=>"101011111",
  27457=>"111001000",
  27458=>"000001110",
  27459=>"101011000",
  27460=>"000110100",
  27461=>"000010011",
  27462=>"010000010",
  27463=>"111011110",
  27464=>"101000101",
  27465=>"011110101",
  27466=>"100010100",
  27467=>"001000000",
  27468=>"000011001",
  27469=>"011011001",
  27470=>"110111110",
  27471=>"111001101",
  27472=>"101000001",
  27473=>"011101101",
  27474=>"100100000",
  27475=>"001110000",
  27476=>"011111110",
  27477=>"001101011",
  27478=>"000100000",
  27479=>"110001011",
  27480=>"110101101",
  27481=>"001011000",
  27482=>"110111000",
  27483=>"000111111",
  27484=>"001010011",
  27485=>"100101011",
  27486=>"100001010",
  27487=>"010100100",
  27488=>"000101100",
  27489=>"100000101",
  27490=>"111000000",
  27491=>"110111011",
  27492=>"101000111",
  27493=>"110110010",
  27494=>"000010110",
  27495=>"111000010",
  27496=>"000101010",
  27497=>"111101111",
  27498=>"011000111",
  27499=>"001101101",
  27500=>"011011011",
  27501=>"110000110",
  27502=>"010011101",
  27503=>"000001011",
  27504=>"110111001",
  27505=>"000000000",
  27506=>"101111010",
  27507=>"101101110",
  27508=>"101001010",
  27509=>"000111100",
  27510=>"000010000",
  27511=>"000110011",
  27512=>"100111011",
  27513=>"100100010",
  27514=>"000101110",
  27515=>"000111010",
  27516=>"101111110",
  27517=>"001011100",
  27518=>"000100000",
  27519=>"011110101",
  27520=>"110111011",
  27521=>"010001010",
  27522=>"010001000",
  27523=>"111000111",
  27524=>"001011001",
  27525=>"101010011",
  27526=>"000110100",
  27527=>"010001100",
  27528=>"110011111",
  27529=>"100010001",
  27530=>"000111010",
  27531=>"100010010",
  27532=>"000101110",
  27533=>"011010011",
  27534=>"100011001",
  27535=>"101010000",
  27536=>"001000011",
  27537=>"010010010",
  27538=>"001101011",
  27539=>"001100111",
  27540=>"001111000",
  27541=>"110111111",
  27542=>"000011110",
  27543=>"001101001",
  27544=>"101110111",
  27545=>"000011010",
  27546=>"001011110",
  27547=>"110000100",
  27548=>"100111100",
  27549=>"001000011",
  27550=>"011001110",
  27551=>"111101000",
  27552=>"011001010",
  27553=>"001100111",
  27554=>"010011111",
  27555=>"000100001",
  27556=>"001101010",
  27557=>"011111111",
  27558=>"000011010",
  27559=>"100111111",
  27560=>"101110110",
  27561=>"011100110",
  27562=>"101100000",
  27563=>"110111111",
  27564=>"100111011",
  27565=>"111101101",
  27566=>"101001011",
  27567=>"001111001",
  27568=>"110110001",
  27569=>"111010011",
  27570=>"001111010",
  27571=>"011001100",
  27572=>"001100001",
  27573=>"111010110",
  27574=>"011101110",
  27575=>"111010100",
  27576=>"010000001",
  27577=>"011111111",
  27578=>"001110100",
  27579=>"110100000",
  27580=>"000010001",
  27581=>"111111111",
  27582=>"011001101",
  27583=>"101101001",
  27584=>"001011101",
  27585=>"100101000",
  27586=>"000001111",
  27587=>"001111111",
  27588=>"111011011",
  27589=>"000111111",
  27590=>"101011110",
  27591=>"001000101",
  27592=>"001000111",
  27593=>"010101000",
  27594=>"001000000",
  27595=>"101011011",
  27596=>"010110011",
  27597=>"100000010",
  27598=>"111011101",
  27599=>"000001101",
  27600=>"001111100",
  27601=>"001111010",
  27602=>"000110001",
  27603=>"000000100",
  27604=>"110000011",
  27605=>"101000100",
  27606=>"010001101",
  27607=>"101101101",
  27608=>"100101110",
  27609=>"101001001",
  27610=>"111110000",
  27611=>"010111011",
  27612=>"001100100",
  27613=>"011111110",
  27614=>"110010001",
  27615=>"110101010",
  27616=>"101110111",
  27617=>"001000001",
  27618=>"000000100",
  27619=>"110100101",
  27620=>"110011011",
  27621=>"000011000",
  27622=>"011100101",
  27623=>"011000001",
  27624=>"101010000",
  27625=>"000010101",
  27626=>"000101000",
  27627=>"110001101",
  27628=>"111111000",
  27629=>"101000000",
  27630=>"001001010",
  27631=>"000100111",
  27632=>"000110111",
  27633=>"000111011",
  27634=>"001011111",
  27635=>"101110100",
  27636=>"100011000",
  27637=>"010000000",
  27638=>"100111000",
  27639=>"100111011",
  27640=>"100010100",
  27641=>"000000010",
  27642=>"000000000",
  27643=>"010111000",
  27644=>"010100111",
  27645=>"011010101",
  27646=>"001011110",
  27647=>"000110010",
  27648=>"110011111",
  27649=>"000011100",
  27650=>"011101110",
  27651=>"011110111",
  27652=>"011000001",
  27653=>"001001111",
  27654=>"011111100",
  27655=>"010000100",
  27656=>"001101111",
  27657=>"000001010",
  27658=>"111011010",
  27659=>"010111010",
  27660=>"111001100",
  27661=>"001000101",
  27662=>"000100010",
  27663=>"010011111",
  27664=>"110101111",
  27665=>"010101011",
  27666=>"101100101",
  27667=>"101011110",
  27668=>"001000100",
  27669=>"000111001",
  27670=>"100111100",
  27671=>"000011100",
  27672=>"010100000",
  27673=>"110000100",
  27674=>"111111111",
  27675=>"010101010",
  27676=>"110011100",
  27677=>"010101000",
  27678=>"111010010",
  27679=>"010111111",
  27680=>"010010111",
  27681=>"001110010",
  27682=>"101111110",
  27683=>"101011000",
  27684=>"101001000",
  27685=>"111101100",
  27686=>"100100100",
  27687=>"111011100",
  27688=>"100010000",
  27689=>"001110110",
  27690=>"010000000",
  27691=>"100111001",
  27692=>"010010000",
  27693=>"000101111",
  27694=>"110100010",
  27695=>"100011111",
  27696=>"000100110",
  27697=>"101010111",
  27698=>"001011001",
  27699=>"010110101",
  27700=>"000010000",
  27701=>"100000101",
  27702=>"110011111",
  27703=>"110110100",
  27704=>"001001011",
  27705=>"111101000",
  27706=>"010111001",
  27707=>"101100111",
  27708=>"101011001",
  27709=>"000001001",
  27710=>"010011110",
  27711=>"010010010",
  27712=>"100100110",
  27713=>"111011111",
  27714=>"010110101",
  27715=>"001000001",
  27716=>"101110001",
  27717=>"011000110",
  27718=>"010111101",
  27719=>"010100000",
  27720=>"110011110",
  27721=>"110111011",
  27722=>"101010111",
  27723=>"001010000",
  27724=>"000001000",
  27725=>"010101111",
  27726=>"010110110",
  27727=>"000000011",
  27728=>"000101110",
  27729=>"100011100",
  27730=>"011110110",
  27731=>"000110100",
  27732=>"000011100",
  27733=>"001101100",
  27734=>"100001010",
  27735=>"000110010",
  27736=>"101111110",
  27737=>"000110111",
  27738=>"100111011",
  27739=>"110101101",
  27740=>"010100111",
  27741=>"111011101",
  27742=>"010110111",
  27743=>"100010000",
  27744=>"010000111",
  27745=>"100001111",
  27746=>"010001001",
  27747=>"001101001",
  27748=>"011011011",
  27749=>"011101001",
  27750=>"010100111",
  27751=>"011100001",
  27752=>"011011111",
  27753=>"100001111",
  27754=>"101001101",
  27755=>"110110100",
  27756=>"111100110",
  27757=>"110011011",
  27758=>"110111001",
  27759=>"111100100",
  27760=>"111000010",
  27761=>"000001000",
  27762=>"000111110",
  27763=>"110001010",
  27764=>"100010010",
  27765=>"110101011",
  27766=>"111110100",
  27767=>"110010010",
  27768=>"001010110",
  27769=>"110110111",
  27770=>"100000001",
  27771=>"001010100",
  27772=>"001111001",
  27773=>"000011100",
  27774=>"111110110",
  27775=>"110111011",
  27776=>"001101000",
  27777=>"101001111",
  27778=>"101000000",
  27779=>"011100000",
  27780=>"101000010",
  27781=>"101001101",
  27782=>"111111000",
  27783=>"100101111",
  27784=>"111011000",
  27785=>"100101110",
  27786=>"000011011",
  27787=>"100100100",
  27788=>"010101111",
  27789=>"001101111",
  27790=>"100011101",
  27791=>"010001000",
  27792=>"011001010",
  27793=>"111101101",
  27794=>"001000111",
  27795=>"010010000",
  27796=>"110011100",
  27797=>"001110100",
  27798=>"010000001",
  27799=>"000101000",
  27800=>"000101000",
  27801=>"100010011",
  27802=>"011110111",
  27803=>"110110011",
  27804=>"101011101",
  27805=>"100110011",
  27806=>"110000010",
  27807=>"011101011",
  27808=>"001100000",
  27809=>"000111001",
  27810=>"111011000",
  27811=>"101101110",
  27812=>"111101111",
  27813=>"110000110",
  27814=>"110010100",
  27815=>"010010110",
  27816=>"110100111",
  27817=>"010011011",
  27818=>"101111001",
  27819=>"111100111",
  27820=>"110011110",
  27821=>"111100100",
  27822=>"100011000",
  27823=>"000001011",
  27824=>"101111110",
  27825=>"110001010",
  27826=>"011001110",
  27827=>"101010111",
  27828=>"101000000",
  27829=>"111110000",
  27830=>"110110100",
  27831=>"101100000",
  27832=>"000111110",
  27833=>"101001000",
  27834=>"110010001",
  27835=>"000101011",
  27836=>"111011010",
  27837=>"001000101",
  27838=>"111010000",
  27839=>"100101001",
  27840=>"010110101",
  27841=>"111110100",
  27842=>"101001111",
  27843=>"111101000",
  27844=>"111000001",
  27845=>"100100010",
  27846=>"101111011",
  27847=>"011100011",
  27848=>"100110110",
  27849=>"110010101",
  27850=>"010111000",
  27851=>"110011000",
  27852=>"111011011",
  27853=>"011010010",
  27854=>"001110101",
  27855=>"110000011",
  27856=>"101101011",
  27857=>"101101110",
  27858=>"100101110",
  27859=>"110110101",
  27860=>"110010111",
  27861=>"101110011",
  27862=>"100000001",
  27863=>"000011100",
  27864=>"001110110",
  27865=>"001100011",
  27866=>"101000010",
  27867=>"101001001",
  27868=>"000001000",
  27869=>"000010111",
  27870=>"000101110",
  27871=>"110101111",
  27872=>"111101101",
  27873=>"001101011",
  27874=>"100100010",
  27875=>"101110111",
  27876=>"010100000",
  27877=>"000001111",
  27878=>"101100101",
  27879=>"111000001",
  27880=>"101010011",
  27881=>"101101101",
  27882=>"000110000",
  27883=>"011110111",
  27884=>"000001100",
  27885=>"000000100",
  27886=>"111011110",
  27887=>"110111001",
  27888=>"111100010",
  27889=>"001101011",
  27890=>"011100000",
  27891=>"101010100",
  27892=>"001000011",
  27893=>"100010111",
  27894=>"110100010",
  27895=>"101111111",
  27896=>"101110101",
  27897=>"001000011",
  27898=>"101101111",
  27899=>"010000100",
  27900=>"011001000",
  27901=>"000110000",
  27902=>"010111000",
  27903=>"000100001",
  27904=>"011110011",
  27905=>"000100001",
  27906=>"000010110",
  27907=>"011100010",
  27908=>"010000100",
  27909=>"011011101",
  27910=>"110000110",
  27911=>"100110011",
  27912=>"110100111",
  27913=>"000000010",
  27914=>"010100001",
  27915=>"001011011",
  27916=>"001010101",
  27917=>"100111100",
  27918=>"010001000",
  27919=>"110001111",
  27920=>"001110101",
  27921=>"101000000",
  27922=>"100010100",
  27923=>"101000111",
  27924=>"010110011",
  27925=>"101100010",
  27926=>"000111101",
  27927=>"111001111",
  27928=>"100010111",
  27929=>"010001010",
  27930=>"100100110",
  27931=>"000111010",
  27932=>"110111110",
  27933=>"001000011",
  27934=>"001111011",
  27935=>"001001111",
  27936=>"101101101",
  27937=>"111010010",
  27938=>"000100110",
  27939=>"010100000",
  27940=>"010011011",
  27941=>"000101100",
  27942=>"010111111",
  27943=>"111111000",
  27944=>"000100000",
  27945=>"011000010",
  27946=>"001111010",
  27947=>"000000011",
  27948=>"000000100",
  27949=>"100110011",
  27950=>"100001111",
  27951=>"011101111",
  27952=>"100001111",
  27953=>"001101001",
  27954=>"100000101",
  27955=>"100101101",
  27956=>"010001110",
  27957=>"001010110",
  27958=>"110001111",
  27959=>"001111001",
  27960=>"011011000",
  27961=>"010010111",
  27962=>"100000000",
  27963=>"100010101",
  27964=>"101101010",
  27965=>"010101110",
  27966=>"111100111",
  27967=>"011000000",
  27968=>"100000011",
  27969=>"000110001",
  27970=>"100110111",
  27971=>"111011110",
  27972=>"101101101",
  27973=>"000000010",
  27974=>"001101110",
  27975=>"000100010",
  27976=>"111100110",
  27977=>"010101000",
  27978=>"011110100",
  27979=>"000000010",
  27980=>"010100111",
  27981=>"101111100",
  27982=>"100001111",
  27983=>"011101111",
  27984=>"001000011",
  27985=>"100100000",
  27986=>"110101111",
  27987=>"011111101",
  27988=>"001000000",
  27989=>"101001011",
  27990=>"000001000",
  27991=>"101001000",
  27992=>"000100100",
  27993=>"010010111",
  27994=>"101011111",
  27995=>"100110011",
  27996=>"001110110",
  27997=>"001101111",
  27998=>"110101000",
  27999=>"101100000",
  28000=>"101111111",
  28001=>"001111010",
  28002=>"111101001",
  28003=>"000110011",
  28004=>"000010101",
  28005=>"101110000",
  28006=>"010010010",
  28007=>"111101111",
  28008=>"101001011",
  28009=>"010000101",
  28010=>"110110110",
  28011=>"101010101",
  28012=>"100001010",
  28013=>"100000000",
  28014=>"000111110",
  28015=>"011101110",
  28016=>"100101010",
  28017=>"010101000",
  28018=>"100100111",
  28019=>"011100110",
  28020=>"000100101",
  28021=>"001110000",
  28022=>"001110000",
  28023=>"000110001",
  28024=>"111001001",
  28025=>"000101100",
  28026=>"111111100",
  28027=>"010000100",
  28028=>"101111110",
  28029=>"000101011",
  28030=>"101010000",
  28031=>"011100010",
  28032=>"001010000",
  28033=>"000101101",
  28034=>"000100110",
  28035=>"101100111",
  28036=>"000111111",
  28037=>"000111010",
  28038=>"110111111",
  28039=>"100100100",
  28040=>"111011010",
  28041=>"100011000",
  28042=>"001001110",
  28043=>"010100111",
  28044=>"001011111",
  28045=>"010011100",
  28046=>"000100001",
  28047=>"010110100",
  28048=>"001011001",
  28049=>"111011000",
  28050=>"100001100",
  28051=>"001110111",
  28052=>"000110101",
  28053=>"010111100",
  28054=>"101000111",
  28055=>"000000000",
  28056=>"011000000",
  28057=>"110010000",
  28058=>"101001100",
  28059=>"011100001",
  28060=>"101001111",
  28061=>"111011000",
  28062=>"010010110",
  28063=>"111001100",
  28064=>"101110000",
  28065=>"111110011",
  28066=>"111101000",
  28067=>"000011011",
  28068=>"001100001",
  28069=>"011001001",
  28070=>"001000011",
  28071=>"110001000",
  28072=>"110010100",
  28073=>"101001000",
  28074=>"001100011",
  28075=>"101001111",
  28076=>"111100000",
  28077=>"001000101",
  28078=>"001101000",
  28079=>"011100100",
  28080=>"100001011",
  28081=>"110101010",
  28082=>"011001111",
  28083=>"111010001",
  28084=>"001001011",
  28085=>"000000010",
  28086=>"100101100",
  28087=>"010001100",
  28088=>"011001110",
  28089=>"110011011",
  28090=>"000101011",
  28091=>"111011101",
  28092=>"110100011",
  28093=>"001100111",
  28094=>"110011110",
  28095=>"010110111",
  28096=>"000000011",
  28097=>"111111111",
  28098=>"011101010",
  28099=>"011100010",
  28100=>"100001011",
  28101=>"101000011",
  28102=>"110000000",
  28103=>"001011000",
  28104=>"000010010",
  28105=>"000110000",
  28106=>"001010111",
  28107=>"101111111",
  28108=>"001101001",
  28109=>"001000001",
  28110=>"001110110",
  28111=>"110000111",
  28112=>"110000011",
  28113=>"010001010",
  28114=>"010100010",
  28115=>"101111101",
  28116=>"001110000",
  28117=>"111011100",
  28118=>"100001010",
  28119=>"110111010",
  28120=>"111001010",
  28121=>"001000100",
  28122=>"000101001",
  28123=>"110101100",
  28124=>"111010100",
  28125=>"101001000",
  28126=>"100000111",
  28127=>"111100101",
  28128=>"111111010",
  28129=>"111111100",
  28130=>"101011101",
  28131=>"111011011",
  28132=>"101001101",
  28133=>"111101100",
  28134=>"001111110",
  28135=>"011011010",
  28136=>"010100100",
  28137=>"000010110",
  28138=>"101010100",
  28139=>"100011110",
  28140=>"100001110",
  28141=>"010011110",
  28142=>"000101110",
  28143=>"111011111",
  28144=>"100000001",
  28145=>"010011010",
  28146=>"011000001",
  28147=>"100010101",
  28148=>"100000010",
  28149=>"000001011",
  28150=>"111010101",
  28151=>"111100100",
  28152=>"001111000",
  28153=>"011001000",
  28154=>"000000011",
  28155=>"101111111",
  28156=>"011110000",
  28157=>"111111011",
  28158=>"011011111",
  28159=>"100110011",
  28160=>"010010000",
  28161=>"110110101",
  28162=>"101101101",
  28163=>"000100111",
  28164=>"010101011",
  28165=>"010110101",
  28166=>"001100000",
  28167=>"110111110",
  28168=>"110110111",
  28169=>"000011110",
  28170=>"010111111",
  28171=>"110111001",
  28172=>"000110011",
  28173=>"111110000",
  28174=>"001111011",
  28175=>"111110011",
  28176=>"101010011",
  28177=>"100001000",
  28178=>"101101111",
  28179=>"110100010",
  28180=>"010000001",
  28181=>"000001101",
  28182=>"011000100",
  28183=>"101011011",
  28184=>"000111010",
  28185=>"000100011",
  28186=>"001101000",
  28187=>"000110000",
  28188=>"111111011",
  28189=>"011100111",
  28190=>"100101100",
  28191=>"001011111",
  28192=>"011000110",
  28193=>"000111011",
  28194=>"001001001",
  28195=>"000110110",
  28196=>"011011111",
  28197=>"010100100",
  28198=>"101100001",
  28199=>"100001111",
  28200=>"101011111",
  28201=>"101000011",
  28202=>"011011110",
  28203=>"001000101",
  28204=>"110111111",
  28205=>"110100011",
  28206=>"101111000",
  28207=>"111000011",
  28208=>"001111101",
  28209=>"110111001",
  28210=>"000000001",
  28211=>"000000100",
  28212=>"000000011",
  28213=>"010001100",
  28214=>"011101001",
  28215=>"111111010",
  28216=>"110000100",
  28217=>"110110110",
  28218=>"000010110",
  28219=>"110101011",
  28220=>"110100100",
  28221=>"011001000",
  28222=>"010000001",
  28223=>"001010000",
  28224=>"111100111",
  28225=>"111001110",
  28226=>"111111101",
  28227=>"000000111",
  28228=>"001111001",
  28229=>"001000100",
  28230=>"000001101",
  28231=>"001001101",
  28232=>"011111100",
  28233=>"000010010",
  28234=>"011111010",
  28235=>"000101101",
  28236=>"001000011",
  28237=>"101100100",
  28238=>"011110011",
  28239=>"000110111",
  28240=>"100111001",
  28241=>"100111101",
  28242=>"000001001",
  28243=>"001101011",
  28244=>"000111000",
  28245=>"111010100",
  28246=>"011000100",
  28247=>"111011111",
  28248=>"010111101",
  28249=>"111011101",
  28250=>"001010100",
  28251=>"101000110",
  28252=>"100111111",
  28253=>"010110110",
  28254=>"001010011",
  28255=>"000110111",
  28256=>"101110000",
  28257=>"001011000",
  28258=>"001010110",
  28259=>"001001101",
  28260=>"000001000",
  28261=>"111100101",
  28262=>"010011110",
  28263=>"110110000",
  28264=>"000101001",
  28265=>"010000110",
  28266=>"100001011",
  28267=>"101100011",
  28268=>"001011001",
  28269=>"101110010",
  28270=>"100101101",
  28271=>"100011110",
  28272=>"101010010",
  28273=>"010110101",
  28274=>"011111000",
  28275=>"101011111",
  28276=>"010010001",
  28277=>"110110111",
  28278=>"000010001",
  28279=>"111110100",
  28280=>"110110100",
  28281=>"010000000",
  28282=>"000100011",
  28283=>"111010111",
  28284=>"110010010",
  28285=>"011000101",
  28286=>"110010011",
  28287=>"100110111",
  28288=>"001000001",
  28289=>"000111111",
  28290=>"000010110",
  28291=>"111010111",
  28292=>"111011000",
  28293=>"000110110",
  28294=>"101100101",
  28295=>"000110000",
  28296=>"001000000",
  28297=>"101100110",
  28298=>"111100110",
  28299=>"010001010",
  28300=>"111101111",
  28301=>"111001011",
  28302=>"110100010",
  28303=>"100010111",
  28304=>"010001110",
  28305=>"010101000",
  28306=>"101111111",
  28307=>"011110101",
  28308=>"111000001",
  28309=>"001011011",
  28310=>"101101010",
  28311=>"111110000",
  28312=>"111110101",
  28313=>"101001010",
  28314=>"110000100",
  28315=>"010101001",
  28316=>"110000111",
  28317=>"110011100",
  28318=>"010001010",
  28319=>"001110100",
  28320=>"000001101",
  28321=>"111100001",
  28322=>"011110011",
  28323=>"111101111",
  28324=>"100001010",
  28325=>"111110000",
  28326=>"100011000",
  28327=>"001110100",
  28328=>"001100011",
  28329=>"101011010",
  28330=>"001000100",
  28331=>"111011100",
  28332=>"010000010",
  28333=>"100101110",
  28334=>"010100001",
  28335=>"010011100",
  28336=>"000010000",
  28337=>"110111001",
  28338=>"010011001",
  28339=>"111011001",
  28340=>"111101010",
  28341=>"011100001",
  28342=>"101101001",
  28343=>"011100101",
  28344=>"000010001",
  28345=>"011000011",
  28346=>"111111101",
  28347=>"111010110",
  28348=>"011000000",
  28349=>"001001111",
  28350=>"101011010",
  28351=>"101001101",
  28352=>"100011101",
  28353=>"011010101",
  28354=>"010110110",
  28355=>"000000100",
  28356=>"000010001",
  28357=>"010101011",
  28358=>"000010000",
  28359=>"011000010",
  28360=>"110000100",
  28361=>"001000101",
  28362=>"100001110",
  28363=>"001011101",
  28364=>"110100001",
  28365=>"101110110",
  28366=>"111001111",
  28367=>"001000010",
  28368=>"111001011",
  28369=>"011111111",
  28370=>"100011101",
  28371=>"101011110",
  28372=>"111001100",
  28373=>"011010010",
  28374=>"110100000",
  28375=>"001011011",
  28376=>"101000000",
  28377=>"000000010",
  28378=>"101001110",
  28379=>"110011001",
  28380=>"001010111",
  28381=>"100100001",
  28382=>"101011010",
  28383=>"010100111",
  28384=>"111000010",
  28385=>"011011011",
  28386=>"111111011",
  28387=>"010011010",
  28388=>"001000110",
  28389=>"101011011",
  28390=>"111100101",
  28391=>"111111110",
  28392=>"110100101",
  28393=>"001100111",
  28394=>"001001111",
  28395=>"111000011",
  28396=>"000011110",
  28397=>"001111101",
  28398=>"101001011",
  28399=>"011101010",
  28400=>"010010110",
  28401=>"011110000",
  28402=>"001011101",
  28403=>"000100100",
  28404=>"011101110",
  28405=>"000101001",
  28406=>"000010011",
  28407=>"011011100",
  28408=>"111100111",
  28409=>"000000010",
  28410=>"111000010",
  28411=>"101111101",
  28412=>"001110110",
  28413=>"000001000",
  28414=>"110101000",
  28415=>"101101101",
  28416=>"010101101",
  28417=>"000111000",
  28418=>"110011110",
  28419=>"000000100",
  28420=>"101110001",
  28421=>"100100101",
  28422=>"000110101",
  28423=>"010110000",
  28424=>"101001100",
  28425=>"011101010",
  28426=>"010010110",
  28427=>"110101011",
  28428=>"000001101",
  28429=>"111100001",
  28430=>"100110110",
  28431=>"101111101",
  28432=>"100111100",
  28433=>"101100010",
  28434=>"011100101",
  28435=>"011001010",
  28436=>"111110000",
  28437=>"110101010",
  28438=>"110010111",
  28439=>"000101000",
  28440=>"011001011",
  28441=>"010001101",
  28442=>"001110101",
  28443=>"101000000",
  28444=>"010110000",
  28445=>"000100111",
  28446=>"110110111",
  28447=>"011000110",
  28448=>"111011111",
  28449=>"110001010",
  28450=>"100110001",
  28451=>"010101010",
  28452=>"011101010",
  28453=>"101100010",
  28454=>"011010000",
  28455=>"101101011",
  28456=>"001010000",
  28457=>"100011110",
  28458=>"010111011",
  28459=>"100110101",
  28460=>"100001010",
  28461=>"100010001",
  28462=>"000111110",
  28463=>"100001100",
  28464=>"011110111",
  28465=>"000001100",
  28466=>"011111010",
  28467=>"100111100",
  28468=>"100111111",
  28469=>"010101011",
  28470=>"110111010",
  28471=>"000010110",
  28472=>"001001010",
  28473=>"110010011",
  28474=>"001011111",
  28475=>"011100000",
  28476=>"100000110",
  28477=>"111000110",
  28478=>"100010000",
  28479=>"000100001",
  28480=>"011011000",
  28481=>"010101000",
  28482=>"111100110",
  28483=>"011101110",
  28484=>"110100001",
  28485=>"011110110",
  28486=>"100111110",
  28487=>"111111100",
  28488=>"010111011",
  28489=>"101011011",
  28490=>"101011101",
  28491=>"000101101",
  28492=>"111110011",
  28493=>"011010111",
  28494=>"000010100",
  28495=>"001000100",
  28496=>"101110111",
  28497=>"000110010",
  28498=>"001111100",
  28499=>"010010110",
  28500=>"011110110",
  28501=>"010000000",
  28502=>"010000010",
  28503=>"010011010",
  28504=>"000001001",
  28505=>"000001010",
  28506=>"101101100",
  28507=>"101010001",
  28508=>"000001001",
  28509=>"011001001",
  28510=>"000010000",
  28511=>"001001001",
  28512=>"110101000",
  28513=>"011101111",
  28514=>"001110100",
  28515=>"110110000",
  28516=>"011011011",
  28517=>"000101100",
  28518=>"110011010",
  28519=>"000110000",
  28520=>"101000101",
  28521=>"001001111",
  28522=>"010101001",
  28523=>"101110101",
  28524=>"000101110",
  28525=>"011011000",
  28526=>"010101101",
  28527=>"010000101",
  28528=>"110000000",
  28529=>"011111011",
  28530=>"111101101",
  28531=>"011111110",
  28532=>"100110100",
  28533=>"111101101",
  28534=>"100001000",
  28535=>"011000101",
  28536=>"101100100",
  28537=>"110011001",
  28538=>"010011100",
  28539=>"011111011",
  28540=>"000011101",
  28541=>"011010011",
  28542=>"110011101",
  28543=>"100111111",
  28544=>"101010110",
  28545=>"110100010",
  28546=>"110110101",
  28547=>"010100011",
  28548=>"011110111",
  28549=>"111010001",
  28550=>"001011100",
  28551=>"010101111",
  28552=>"000011111",
  28553=>"011000001",
  28554=>"110000100",
  28555=>"111011111",
  28556=>"011111111",
  28557=>"101011001",
  28558=>"011000010",
  28559=>"101010000",
  28560=>"110010110",
  28561=>"101101010",
  28562=>"001101100",
  28563=>"001001100",
  28564=>"100011101",
  28565=>"011101011",
  28566=>"100101111",
  28567=>"001000110",
  28568=>"000111111",
  28569=>"111001100",
  28570=>"110001010",
  28571=>"011010110",
  28572=>"111101011",
  28573=>"000111000",
  28574=>"100111001",
  28575=>"100100000",
  28576=>"011011011",
  28577=>"010011000",
  28578=>"111110010",
  28579=>"000111011",
  28580=>"111010100",
  28581=>"101000110",
  28582=>"110000100",
  28583=>"011111111",
  28584=>"111001101",
  28585=>"001001001",
  28586=>"111101110",
  28587=>"011001101",
  28588=>"100101011",
  28589=>"111111000",
  28590=>"101010001",
  28591=>"100110100",
  28592=>"011100010",
  28593=>"111000100",
  28594=>"100100110",
  28595=>"001000001",
  28596=>"001100111",
  28597=>"100101010",
  28598=>"101010100",
  28599=>"010011011",
  28600=>"110010111",
  28601=>"010011010",
  28602=>"111100100",
  28603=>"111001010",
  28604=>"100101010",
  28605=>"101000111",
  28606=>"010100110",
  28607=>"110100100",
  28608=>"011110111",
  28609=>"010100101",
  28610=>"010110010",
  28611=>"101001110",
  28612=>"001101101",
  28613=>"001001110",
  28614=>"100011011",
  28615=>"111110110",
  28616=>"000000001",
  28617=>"010100110",
  28618=>"110111001",
  28619=>"100111111",
  28620=>"101101111",
  28621=>"011001010",
  28622=>"001111010",
  28623=>"000100010",
  28624=>"100101110",
  28625=>"100100101",
  28626=>"000101101",
  28627=>"110001000",
  28628=>"000100000",
  28629=>"110110000",
  28630=>"010110001",
  28631=>"110110101",
  28632=>"111000111",
  28633=>"000001101",
  28634=>"111000000",
  28635=>"110110000",
  28636=>"011001010",
  28637=>"000110100",
  28638=>"010000010",
  28639=>"101111111",
  28640=>"110000101",
  28641=>"101100111",
  28642=>"101101010",
  28643=>"111000011",
  28644=>"110010011",
  28645=>"100101011",
  28646=>"010101010",
  28647=>"001011000",
  28648=>"001101001",
  28649=>"110011101",
  28650=>"100101110",
  28651=>"001100101",
  28652=>"101111100",
  28653=>"000011110",
  28654=>"011111010",
  28655=>"000001011",
  28656=>"000100100",
  28657=>"110101011",
  28658=>"001010010",
  28659=>"110101111",
  28660=>"010100100",
  28661=>"111111001",
  28662=>"110100110",
  28663=>"011110000",
  28664=>"001010000",
  28665=>"000110001",
  28666=>"001111111",
  28667=>"100000110",
  28668=>"001000100",
  28669=>"001011000",
  28670=>"111000011",
  28671=>"111111110",
  28672=>"100111010",
  28673=>"101111100",
  28674=>"111100000",
  28675=>"011000101",
  28676=>"101010111",
  28677=>"100101010",
  28678=>"001000011",
  28679=>"011000000",
  28680=>"001001000",
  28681=>"011111000",
  28682=>"000011101",
  28683=>"010000101",
  28684=>"111001110",
  28685=>"101010010",
  28686=>"111110110",
  28687=>"011110111",
  28688=>"000100000",
  28689=>"001100000",
  28690=>"000101000",
  28691=>"100011100",
  28692=>"011010001",
  28693=>"111100100",
  28694=>"101000011",
  28695=>"010100011",
  28696=>"100111111",
  28697=>"110000001",
  28698=>"011000011",
  28699=>"101101101",
  28700=>"110111101",
  28701=>"010100100",
  28702=>"010111100",
  28703=>"000010000",
  28704=>"010001100",
  28705=>"110010101",
  28706=>"100000001",
  28707=>"110100010",
  28708=>"000001111",
  28709=>"000110010",
  28710=>"001101000",
  28711=>"111111100",
  28712=>"100001001",
  28713=>"001110010",
  28714=>"000010000",
  28715=>"001011101",
  28716=>"001001100",
  28717=>"100010101",
  28718=>"100100001",
  28719=>"111000001",
  28720=>"111010111",
  28721=>"111100100",
  28722=>"101010000",
  28723=>"101011101",
  28724=>"110100100",
  28725=>"111001111",
  28726=>"000100100",
  28727=>"101011110",
  28728=>"100001110",
  28729=>"110001101",
  28730=>"011111011",
  28731=>"111110001",
  28732=>"011010111",
  28733=>"001101110",
  28734=>"110100101",
  28735=>"001001010",
  28736=>"011110110",
  28737=>"001101001",
  28738=>"001100110",
  28739=>"000111110",
  28740=>"010011110",
  28741=>"110011111",
  28742=>"100011111",
  28743=>"011111110",
  28744=>"110101001",
  28745=>"100001110",
  28746=>"100010011",
  28747=>"101001011",
  28748=>"010001100",
  28749=>"011100001",
  28750=>"000100101",
  28751=>"000000011",
  28752=>"011001010",
  28753=>"000001001",
  28754=>"111000100",
  28755=>"110111101",
  28756=>"001100000",
  28757=>"110000010",
  28758=>"000100110",
  28759=>"100101110",
  28760=>"111111001",
  28761=>"000111011",
  28762=>"001101010",
  28763=>"000100010",
  28764=>"101110010",
  28765=>"011110110",
  28766=>"011110111",
  28767=>"110001111",
  28768=>"110010010",
  28769=>"000010001",
  28770=>"100000110",
  28771=>"001000000",
  28772=>"000111100",
  28773=>"011101010",
  28774=>"001011000",
  28775=>"000100101",
  28776=>"001100001",
  28777=>"000011001",
  28778=>"001010101",
  28779=>"101011000",
  28780=>"110000010",
  28781=>"000001000",
  28782=>"011011001",
  28783=>"001001110",
  28784=>"100000100",
  28785=>"010101000",
  28786=>"000101111",
  28787=>"001100100",
  28788=>"110001111",
  28789=>"010101111",
  28790=>"111101101",
  28791=>"111011011",
  28792=>"011101011",
  28793=>"111100001",
  28794=>"111000010",
  28795=>"010011111",
  28796=>"011100111",
  28797=>"011110000",
  28798=>"101010010",
  28799=>"001000111",
  28800=>"001100110",
  28801=>"000010110",
  28802=>"001000001",
  28803=>"010110110",
  28804=>"000010111",
  28805=>"011001111",
  28806=>"100001101",
  28807=>"110000011",
  28808=>"001000111",
  28809=>"100100110",
  28810=>"110001000",
  28811=>"010011101",
  28812=>"000111100",
  28813=>"100011100",
  28814=>"010111111",
  28815=>"001011111",
  28816=>"000100010",
  28817=>"100101000",
  28818=>"000011111",
  28819=>"110000101",
  28820=>"001001011",
  28821=>"001110011",
  28822=>"111011001",
  28823=>"111110000",
  28824=>"111100101",
  28825=>"100000101",
  28826=>"011100100",
  28827=>"101101111",
  28828=>"100110010",
  28829=>"000010011",
  28830=>"101010110",
  28831=>"001000011",
  28832=>"011100000",
  28833=>"101100011",
  28834=>"111011010",
  28835=>"000000000",
  28836=>"010111000",
  28837=>"011110010",
  28838=>"010100001",
  28839=>"111100111",
  28840=>"001011010",
  28841=>"111101100",
  28842=>"001010010",
  28843=>"100100010",
  28844=>"101010011",
  28845=>"110000100",
  28846=>"010110101",
  28847=>"111011111",
  28848=>"010010010",
  28849=>"110010011",
  28850=>"001001100",
  28851=>"101010110",
  28852=>"001001000",
  28853=>"110000010",
  28854=>"110101111",
  28855=>"110111111",
  28856=>"000100010",
  28857=>"000101000",
  28858=>"100000101",
  28859=>"111010111",
  28860=>"111111001",
  28861=>"111010010",
  28862=>"101110111",
  28863=>"001110110",
  28864=>"011011000",
  28865=>"110101100",
  28866=>"110101001",
  28867=>"111111100",
  28868=>"011100101",
  28869=>"010011100",
  28870=>"110101000",
  28871=>"111000110",
  28872=>"100110100",
  28873=>"101100111",
  28874=>"001101000",
  28875=>"010110100",
  28876=>"000011101",
  28877=>"000101111",
  28878=>"101001011",
  28879=>"110000000",
  28880=>"011111011",
  28881=>"111001010",
  28882=>"000100000",
  28883=>"011111010",
  28884=>"011000100",
  28885=>"101100000",
  28886=>"000111101",
  28887=>"100011000",
  28888=>"101111010",
  28889=>"111110001",
  28890=>"111110100",
  28891=>"100010001",
  28892=>"001110010",
  28893=>"011111101",
  28894=>"011011101",
  28895=>"101101011",
  28896=>"100101000",
  28897=>"100000010",
  28898=>"100101111",
  28899=>"000111110",
  28900=>"111101010",
  28901=>"010110100",
  28902=>"000000101",
  28903=>"100111010",
  28904=>"011101110",
  28905=>"010111110",
  28906=>"010000000",
  28907=>"101111101",
  28908=>"000001011",
  28909=>"000010010",
  28910=>"100000011",
  28911=>"110011101",
  28912=>"111010010",
  28913=>"001000100",
  28914=>"000101011",
  28915=>"111101010",
  28916=>"110101111",
  28917=>"111011010",
  28918=>"111111001",
  28919=>"111000101",
  28920=>"010010111",
  28921=>"111110101",
  28922=>"110011100",
  28923=>"000010100",
  28924=>"010010111",
  28925=>"110111100",
  28926=>"100111010",
  28927=>"000110110",
  28928=>"111000000",
  28929=>"010111000",
  28930=>"100110001",
  28931=>"001011000",
  28932=>"010100011",
  28933=>"100101111",
  28934=>"101111101",
  28935=>"001011101",
  28936=>"111110110",
  28937=>"110011010",
  28938=>"110101100",
  28939=>"001000101",
  28940=>"011000000",
  28941=>"111000000",
  28942=>"111011011",
  28943=>"001011100",
  28944=>"011111110",
  28945=>"100000001",
  28946=>"001110110",
  28947=>"010000011",
  28948=>"101101001",
  28949=>"000001100",
  28950=>"010000110",
  28951=>"100110010",
  28952=>"101110110",
  28953=>"000010111",
  28954=>"100000010",
  28955=>"100010111",
  28956=>"100000110",
  28957=>"010100010",
  28958=>"110000010",
  28959=>"111000111",
  28960=>"111110011",
  28961=>"010010010",
  28962=>"000010101",
  28963=>"001110011",
  28964=>"110110111",
  28965=>"100000000",
  28966=>"101100110",
  28967=>"001000111",
  28968=>"111010110",
  28969=>"001001000",
  28970=>"110000101",
  28971=>"010001110",
  28972=>"100101111",
  28973=>"000001000",
  28974=>"101000110",
  28975=>"111101010",
  28976=>"100111101",
  28977=>"110011100",
  28978=>"000011111",
  28979=>"111110001",
  28980=>"110100001",
  28981=>"100000111",
  28982=>"010000101",
  28983=>"100111111",
  28984=>"000100010",
  28985=>"000001111",
  28986=>"010011011",
  28987=>"110111100",
  28988=>"101001010",
  28989=>"000010011",
  28990=>"111111110",
  28991=>"011010010",
  28992=>"000100010",
  28993=>"010110001",
  28994=>"101001110",
  28995=>"000000100",
  28996=>"101001001",
  28997=>"101011110",
  28998=>"010000100",
  28999=>"010011011",
  29000=>"111001011",
  29001=>"011000010",
  29002=>"011111001",
  29003=>"100010001",
  29004=>"100000110",
  29005=>"001110100",
  29006=>"001100000",
  29007=>"010001111",
  29008=>"010100110",
  29009=>"001110111",
  29010=>"001010101",
  29011=>"011011101",
  29012=>"011100001",
  29013=>"010101101",
  29014=>"111100100",
  29015=>"011011100",
  29016=>"000111010",
  29017=>"010110111",
  29018=>"100010000",
  29019=>"001001100",
  29020=>"001101001",
  29021=>"011110100",
  29022=>"011111101",
  29023=>"000111110",
  29024=>"000011100",
  29025=>"001010110",
  29026=>"000001000",
  29027=>"101110001",
  29028=>"010010000",
  29029=>"101111010",
  29030=>"010111110",
  29031=>"011010000",
  29032=>"111111000",
  29033=>"001001101",
  29034=>"011111010",
  29035=>"101100001",
  29036=>"110100111",
  29037=>"000001001",
  29038=>"001010010",
  29039=>"001010010",
  29040=>"101111100",
  29041=>"010001010",
  29042=>"010100000",
  29043=>"010111001",
  29044=>"011111101",
  29045=>"000111101",
  29046=>"000010001",
  29047=>"110100011",
  29048=>"011100011",
  29049=>"011010010",
  29050=>"101001100",
  29051=>"110011011",
  29052=>"001100110",
  29053=>"000010000",
  29054=>"111011011",
  29055=>"101101000",
  29056=>"110100111",
  29057=>"010011010",
  29058=>"010110001",
  29059=>"010100000",
  29060=>"001001010",
  29061=>"010011010",
  29062=>"001111011",
  29063=>"110000000",
  29064=>"110010010",
  29065=>"011100011",
  29066=>"001000000",
  29067=>"001100000",
  29068=>"000011001",
  29069=>"001000110",
  29070=>"010101001",
  29071=>"101000010",
  29072=>"011101100",
  29073=>"101001101",
  29074=>"001001010",
  29075=>"001101000",
  29076=>"001111010",
  29077=>"100111010",
  29078=>"110000110",
  29079=>"101111101",
  29080=>"101101011",
  29081=>"000000010",
  29082=>"110010001",
  29083=>"111100000",
  29084=>"010110101",
  29085=>"011110111",
  29086=>"111111110",
  29087=>"110110010",
  29088=>"000011110",
  29089=>"110100100",
  29090=>"011111011",
  29091=>"000000010",
  29092=>"100011001",
  29093=>"000100011",
  29094=>"110101100",
  29095=>"000110111",
  29096=>"000010101",
  29097=>"101111101",
  29098=>"101001111",
  29099=>"110101011",
  29100=>"000000011",
  29101=>"111100010",
  29102=>"000011101",
  29103=>"011001011",
  29104=>"101000010",
  29105=>"000100110",
  29106=>"111111000",
  29107=>"000000010",
  29108=>"110000010",
  29109=>"010001011",
  29110=>"111110110",
  29111=>"011001001",
  29112=>"001111101",
  29113=>"001000110",
  29114=>"110011100",
  29115=>"111000010",
  29116=>"011011111",
  29117=>"011101100",
  29118=>"101100000",
  29119=>"110110011",
  29120=>"011010001",
  29121=>"101000001",
  29122=>"010001100",
  29123=>"111100000",
  29124=>"011101111",
  29125=>"111010101",
  29126=>"010110000",
  29127=>"111101011",
  29128=>"101100111",
  29129=>"010000111",
  29130=>"000010000",
  29131=>"111110010",
  29132=>"001111111",
  29133=>"101001111",
  29134=>"110010111",
  29135=>"010101010",
  29136=>"000101001",
  29137=>"001001000",
  29138=>"001011100",
  29139=>"010100010",
  29140=>"000011101",
  29141=>"110101100",
  29142=>"101011011",
  29143=>"101000010",
  29144=>"100101001",
  29145=>"000010010",
  29146=>"010010111",
  29147=>"000001101",
  29148=>"001000011",
  29149=>"101011010",
  29150=>"011010000",
  29151=>"010100101",
  29152=>"100100000",
  29153=>"010011001",
  29154=>"001001001",
  29155=>"100111011",
  29156=>"000101011",
  29157=>"111100100",
  29158=>"011011101",
  29159=>"010010011",
  29160=>"001010110",
  29161=>"001011000",
  29162=>"110010110",
  29163=>"101000100",
  29164=>"111111111",
  29165=>"001011100",
  29166=>"110100111",
  29167=>"110101010",
  29168=>"001011110",
  29169=>"010010111",
  29170=>"011111001",
  29171=>"001111011",
  29172=>"010010101",
  29173=>"010100111",
  29174=>"000111000",
  29175=>"001100010",
  29176=>"000011011",
  29177=>"001101010",
  29178=>"000011001",
  29179=>"111101000",
  29180=>"111011110",
  29181=>"000010101",
  29182=>"100010110",
  29183=>"110011111",
  29184=>"101110100",
  29185=>"000011001",
  29186=>"111101110",
  29187=>"011100101",
  29188=>"000010111",
  29189=>"101101010",
  29190=>"000010011",
  29191=>"000010000",
  29192=>"100010011",
  29193=>"000101011",
  29194=>"000110101",
  29195=>"010100010",
  29196=>"100010001",
  29197=>"010110000",
  29198=>"010001000",
  29199=>"101110101",
  29200=>"110111011",
  29201=>"110101000",
  29202=>"010010000",
  29203=>"111010110",
  29204=>"010110010",
  29205=>"001001011",
  29206=>"110101011",
  29207=>"110100010",
  29208=>"000001000",
  29209=>"111101010",
  29210=>"111100110",
  29211=>"011001111",
  29212=>"100110100",
  29213=>"001001110",
  29214=>"011011111",
  29215=>"011001111",
  29216=>"100111011",
  29217=>"011000100",
  29218=>"011100101",
  29219=>"010010001",
  29220=>"111010111",
  29221=>"010000000",
  29222=>"111011110",
  29223=>"000110011",
  29224=>"111100111",
  29225=>"011110000",
  29226=>"100000111",
  29227=>"101011001",
  29228=>"001011000",
  29229=>"000100000",
  29230=>"000010101",
  29231=>"101111000",
  29232=>"111000000",
  29233=>"101011010",
  29234=>"001001111",
  29235=>"111000101",
  29236=>"100011110",
  29237=>"101000010",
  29238=>"000001000",
  29239=>"110110110",
  29240=>"011100101",
  29241=>"110000000",
  29242=>"010100001",
  29243=>"001010000",
  29244=>"000000111",
  29245=>"100011010",
  29246=>"111101000",
  29247=>"010101010",
  29248=>"011110111",
  29249=>"100001111",
  29250=>"100000111",
  29251=>"100110111",
  29252=>"100000100",
  29253=>"100011101",
  29254=>"111001111",
  29255=>"110011001",
  29256=>"110100111",
  29257=>"001101000",
  29258=>"001110001",
  29259=>"100010011",
  29260=>"100110111",
  29261=>"000100000",
  29262=>"110101010",
  29263=>"101010101",
  29264=>"000001000",
  29265=>"000011110",
  29266=>"011011011",
  29267=>"010110001",
  29268=>"101110001",
  29269=>"000010101",
  29270=>"101000110",
  29271=>"111111001",
  29272=>"001000011",
  29273=>"110101011",
  29274=>"100000111",
  29275=>"011001100",
  29276=>"101100111",
  29277=>"000001000",
  29278=>"101011110",
  29279=>"110010000",
  29280=>"100001101",
  29281=>"110001110",
  29282=>"110100011",
  29283=>"010101011",
  29284=>"110111110",
  29285=>"011100001",
  29286=>"011100011",
  29287=>"011101100",
  29288=>"000001000",
  29289=>"101100000",
  29290=>"000000001",
  29291=>"100010001",
  29292=>"011111100",
  29293=>"100001110",
  29294=>"110111010",
  29295=>"001110001",
  29296=>"011110011",
  29297=>"010000100",
  29298=>"010111000",
  29299=>"101101100",
  29300=>"100111011",
  29301=>"000110110",
  29302=>"100100110",
  29303=>"001001000",
  29304=>"011100110",
  29305=>"010110110",
  29306=>"100001011",
  29307=>"001000000",
  29308=>"010100111",
  29309=>"000101111",
  29310=>"011011100",
  29311=>"110100010",
  29312=>"011001111",
  29313=>"010000100",
  29314=>"111100000",
  29315=>"000001010",
  29316=>"000001101",
  29317=>"100011100",
  29318=>"100011010",
  29319=>"000101100",
  29320=>"011010001",
  29321=>"111111001",
  29322=>"101011101",
  29323=>"110010011",
  29324=>"000000011",
  29325=>"010110000",
  29326=>"001010000",
  29327=>"000000000",
  29328=>"011001011",
  29329=>"101010111",
  29330=>"101010010",
  29331=>"000001110",
  29332=>"100010000",
  29333=>"010010011",
  29334=>"010101101",
  29335=>"101001011",
  29336=>"101011001",
  29337=>"101111001",
  29338=>"100100000",
  29339=>"010100111",
  29340=>"011010101",
  29341=>"110111001",
  29342=>"110001011",
  29343=>"010010001",
  29344=>"000011100",
  29345=>"011001001",
  29346=>"110111011",
  29347=>"100000110",
  29348=>"001110111",
  29349=>"010111000",
  29350=>"010000011",
  29351=>"100110000",
  29352=>"101001010",
  29353=>"101000111",
  29354=>"010111000",
  29355=>"101111110",
  29356=>"100000101",
  29357=>"010101010",
  29358=>"100000111",
  29359=>"111101110",
  29360=>"010100000",
  29361=>"000101101",
  29362=>"100100001",
  29363=>"001000100",
  29364=>"100001111",
  29365=>"010100001",
  29366=>"101011100",
  29367=>"000000111",
  29368=>"000100011",
  29369=>"101010000",
  29370=>"101111011",
  29371=>"100010010",
  29372=>"010011110",
  29373=>"011111011",
  29374=>"010011100",
  29375=>"100111100",
  29376=>"001111000",
  29377=>"110100011",
  29378=>"001010100",
  29379=>"001000001",
  29380=>"010101000",
  29381=>"000100110",
  29382=>"001111000",
  29383=>"101001001",
  29384=>"111111110",
  29385=>"010001001",
  29386=>"010100011",
  29387=>"101001111",
  29388=>"110011000",
  29389=>"110011000",
  29390=>"111010110",
  29391=>"111111111",
  29392=>"111111111",
  29393=>"100000001",
  29394=>"000100010",
  29395=>"100111100",
  29396=>"000101001",
  29397=>"000000100",
  29398=>"100000110",
  29399=>"011110000",
  29400=>"000001100",
  29401=>"000011101",
  29402=>"110000101",
  29403=>"100011010",
  29404=>"001101110",
  29405=>"011101011",
  29406=>"101000110",
  29407=>"101000111",
  29408=>"001100101",
  29409=>"010011010",
  29410=>"110110111",
  29411=>"101111111",
  29412=>"111101000",
  29413=>"000010000",
  29414=>"100111010",
  29415=>"000100110",
  29416=>"001000110",
  29417=>"101001011",
  29418=>"101101010",
  29419=>"100110100",
  29420=>"110010101",
  29421=>"101001000",
  29422=>"000000000",
  29423=>"010110100",
  29424=>"010111000",
  29425=>"000000001",
  29426=>"110100011",
  29427=>"011011001",
  29428=>"001011110",
  29429=>"101000001",
  29430=>"000010001",
  29431=>"010111100",
  29432=>"110101101",
  29433=>"101100000",
  29434=>"010010010",
  29435=>"000101110",
  29436=>"010100100",
  29437=>"000000100",
  29438=>"011000110",
  29439=>"000001000",
  29440=>"000000110",
  29441=>"011011011",
  29442=>"011101010",
  29443=>"110111000",
  29444=>"001000100",
  29445=>"000011000",
  29446=>"101001101",
  29447=>"001000000",
  29448=>"101010001",
  29449=>"010010010",
  29450=>"001110110",
  29451=>"101011111",
  29452=>"000011100",
  29453=>"110110110",
  29454=>"101001111",
  29455=>"001001001",
  29456=>"001010010",
  29457=>"001000000",
  29458=>"011100000",
  29459=>"011111001",
  29460=>"110011111",
  29461=>"010011010",
  29462=>"011100111",
  29463=>"101001100",
  29464=>"001100110",
  29465=>"110000100",
  29466=>"110100111",
  29467=>"010010111",
  29468=>"111110111",
  29469=>"001000001",
  29470=>"111010011",
  29471=>"111000101",
  29472=>"000001100",
  29473=>"000001011",
  29474=>"101110011",
  29475=>"001011110",
  29476=>"010100000",
  29477=>"110101011",
  29478=>"010000100",
  29479=>"100100010",
  29480=>"100001110",
  29481=>"110001100",
  29482=>"001110010",
  29483=>"000110100",
  29484=>"100010010",
  29485=>"000011011",
  29486=>"011011111",
  29487=>"011011111",
  29488=>"010101000",
  29489=>"101110000",
  29490=>"110010101",
  29491=>"110100001",
  29492=>"111010001",
  29493=>"101010000",
  29494=>"000010010",
  29495=>"111011110",
  29496=>"010110110",
  29497=>"010000100",
  29498=>"111101110",
  29499=>"010011010",
  29500=>"101101100",
  29501=>"100010011",
  29502=>"101000010",
  29503=>"100011001",
  29504=>"110110000",
  29505=>"101101000",
  29506=>"101001011",
  29507=>"111101001",
  29508=>"001010000",
  29509=>"010001011",
  29510=>"010111000",
  29511=>"010101111",
  29512=>"100111001",
  29513=>"101110001",
  29514=>"010000110",
  29515=>"010001000",
  29516=>"110111000",
  29517=>"011011101",
  29518=>"111000101",
  29519=>"000101110",
  29520=>"001100010",
  29521=>"111110110",
  29522=>"100001001",
  29523=>"001111100",
  29524=>"010010101",
  29525=>"110001110",
  29526=>"001011010",
  29527=>"100010001",
  29528=>"110111001",
  29529=>"110111001",
  29530=>"100001101",
  29531=>"101101110",
  29532=>"111110100",
  29533=>"100001101",
  29534=>"011010100",
  29535=>"100000100",
  29536=>"000011110",
  29537=>"000010111",
  29538=>"010100100",
  29539=>"101101010",
  29540=>"001110111",
  29541=>"011101111",
  29542=>"000001100",
  29543=>"011010100",
  29544=>"001101100",
  29545=>"000001101",
  29546=>"101101110",
  29547=>"101101100",
  29548=>"001011100",
  29549=>"101111010",
  29550=>"101010010",
  29551=>"101010101",
  29552=>"100100101",
  29553=>"011001000",
  29554=>"000111111",
  29555=>"111110101",
  29556=>"111100111",
  29557=>"110110001",
  29558=>"101110011",
  29559=>"000000010",
  29560=>"011000000",
  29561=>"001001011",
  29562=>"101111110",
  29563=>"111000001",
  29564=>"111010100",
  29565=>"101111000",
  29566=>"000000010",
  29567=>"111010010",
  29568=>"000001000",
  29569=>"111010100",
  29570=>"101000011",
  29571=>"010011000",
  29572=>"100000110",
  29573=>"100001010",
  29574=>"101111110",
  29575=>"000001101",
  29576=>"001000111",
  29577=>"110000111",
  29578=>"101110011",
  29579=>"100101011",
  29580=>"010111111",
  29581=>"010111001",
  29582=>"110100010",
  29583=>"100111000",
  29584=>"111101001",
  29585=>"010111111",
  29586=>"100011001",
  29587=>"010111011",
  29588=>"010111101",
  29589=>"001101011",
  29590=>"010101100",
  29591=>"001001001",
  29592=>"010100010",
  29593=>"001101000",
  29594=>"010101000",
  29595=>"000110001",
  29596=>"111011010",
  29597=>"110000000",
  29598=>"110000000",
  29599=>"101010000",
  29600=>"000000110",
  29601=>"011111011",
  29602=>"101011111",
  29603=>"011110101",
  29604=>"001110100",
  29605=>"011111001",
  29606=>"001011011",
  29607=>"010110111",
  29608=>"011010110",
  29609=>"000000111",
  29610=>"111111110",
  29611=>"101010110",
  29612=>"111100010",
  29613=>"010001100",
  29614=>"110101100",
  29615=>"100000001",
  29616=>"001110110",
  29617=>"110001010",
  29618=>"001001110",
  29619=>"110000011",
  29620=>"111100011",
  29621=>"110101100",
  29622=>"101111111",
  29623=>"111111000",
  29624=>"111101101",
  29625=>"110110000",
  29626=>"011111110",
  29627=>"000000110",
  29628=>"101001000",
  29629=>"111010110",
  29630=>"011010100",
  29631=>"011000001",
  29632=>"101011011",
  29633=>"101010001",
  29634=>"000000010",
  29635=>"110110111",
  29636=>"000000100",
  29637=>"101101010",
  29638=>"000100101",
  29639=>"111100000",
  29640=>"100101000",
  29641=>"001100011",
  29642=>"011001101",
  29643=>"100001011",
  29644=>"010010011",
  29645=>"010011100",
  29646=>"110011111",
  29647=>"101100100",
  29648=>"001111011",
  29649=>"110000010",
  29650=>"011101010",
  29651=>"010011001",
  29652=>"000010110",
  29653=>"000001000",
  29654=>"000001001",
  29655=>"011010111",
  29656=>"011101010",
  29657=>"010000101",
  29658=>"011000101",
  29659=>"101101101",
  29660=>"101110010",
  29661=>"101011011",
  29662=>"010010000",
  29663=>"100111010",
  29664=>"000110110",
  29665=>"010101111",
  29666=>"100011111",
  29667=>"110001010",
  29668=>"101101010",
  29669=>"101001101",
  29670=>"000000101",
  29671=>"000010010",
  29672=>"000110101",
  29673=>"100111011",
  29674=>"111110111",
  29675=>"001010010",
  29676=>"111101101",
  29677=>"111000101",
  29678=>"111101100",
  29679=>"011010011",
  29680=>"110111000",
  29681=>"000000110",
  29682=>"111010110",
  29683=>"101110111",
  29684=>"010100100",
  29685=>"100111000",
  29686=>"000110010",
  29687=>"101111101",
  29688=>"110000001",
  29689=>"000010110",
  29690=>"001000001",
  29691=>"111110111",
  29692=>"101001011",
  29693=>"101101100",
  29694=>"101000011",
  29695=>"110000111",
  29696=>"110000001",
  29697=>"110010101",
  29698=>"000111010",
  29699=>"111001000",
  29700=>"100100100",
  29701=>"000110001",
  29702=>"000000011",
  29703=>"111011100",
  29704=>"001000010",
  29705=>"101000011",
  29706=>"011011010",
  29707=>"011011110",
  29708=>"100010011",
  29709=>"000110111",
  29710=>"111000111",
  29711=>"000111000",
  29712=>"000110101",
  29713=>"100110100",
  29714=>"011011101",
  29715=>"000010000",
  29716=>"000101001",
  29717=>"111011100",
  29718=>"110111110",
  29719=>"011000101",
  29720=>"101000000",
  29721=>"000001110",
  29722=>"110110011",
  29723=>"111011100",
  29724=>"011011100",
  29725=>"001000100",
  29726=>"111000001",
  29727=>"101010100",
  29728=>"111000001",
  29729=>"110111100",
  29730=>"111001001",
  29731=>"110000010",
  29732=>"111010000",
  29733=>"110001111",
  29734=>"001011110",
  29735=>"101011010",
  29736=>"111111011",
  29737=>"110000000",
  29738=>"010010111",
  29739=>"100000011",
  29740=>"101111110",
  29741=>"100001011",
  29742=>"000000001",
  29743=>"111001110",
  29744=>"110110111",
  29745=>"111000100",
  29746=>"011100000",
  29747=>"011100101",
  29748=>"101101010",
  29749=>"100100100",
  29750=>"110001100",
  29751=>"010010101",
  29752=>"000000101",
  29753=>"011110000",
  29754=>"000001101",
  29755=>"011101110",
  29756=>"011001100",
  29757=>"000001111",
  29758=>"001111101",
  29759=>"101100011",
  29760=>"100011101",
  29761=>"000010010",
  29762=>"000011110",
  29763=>"111010111",
  29764=>"101001110",
  29765=>"010011111",
  29766=>"111111010",
  29767=>"000000011",
  29768=>"111001001",
  29769=>"110100010",
  29770=>"000000011",
  29771=>"010010010",
  29772=>"111010011",
  29773=>"101001000",
  29774=>"100110111",
  29775=>"010110100",
  29776=>"001000000",
  29777=>"111101111",
  29778=>"111011011",
  29779=>"111100100",
  29780=>"011100011",
  29781=>"000110001",
  29782=>"011000011",
  29783=>"001000100",
  29784=>"001101001",
  29785=>"011011101",
  29786=>"101010011",
  29787=>"111000101",
  29788=>"101110110",
  29789=>"000001100",
  29790=>"010011011",
  29791=>"010111101",
  29792=>"001000101",
  29793=>"000000100",
  29794=>"000000001",
  29795=>"000110001",
  29796=>"111100010",
  29797=>"001100011",
  29798=>"000001100",
  29799=>"000101110",
  29800=>"111001110",
  29801=>"111101110",
  29802=>"000001011",
  29803=>"001101001",
  29804=>"111110000",
  29805=>"000000110",
  29806=>"011100010",
  29807=>"011010100",
  29808=>"010011001",
  29809=>"010000111",
  29810=>"111111001",
  29811=>"101010110",
  29812=>"001011101",
  29813=>"011110000",
  29814=>"110111110",
  29815=>"001101010",
  29816=>"001001110",
  29817=>"101110000",
  29818=>"101101010",
  29819=>"111010011",
  29820=>"101001101",
  29821=>"010000010",
  29822=>"110101100",
  29823=>"010110011",
  29824=>"001100110",
  29825=>"010111110",
  29826=>"001101100",
  29827=>"001100000",
  29828=>"100111001",
  29829=>"010000101",
  29830=>"000010001",
  29831=>"000110011",
  29832=>"101000101",
  29833=>"000011000",
  29834=>"100110100",
  29835=>"110100010",
  29836=>"101100010",
  29837=>"110011000",
  29838=>"111110101",
  29839=>"111111000",
  29840=>"011000100",
  29841=>"100110110",
  29842=>"000100001",
  29843=>"110101001",
  29844=>"000001101",
  29845=>"111110010",
  29846=>"101110010",
  29847=>"101100000",
  29848=>"000010010",
  29849=>"011011111",
  29850=>"000000101",
  29851=>"000000101",
  29852=>"100110110",
  29853=>"000001000",
  29854=>"000011001",
  29855=>"011110000",
  29856=>"011001001",
  29857=>"010001110",
  29858=>"111110001",
  29859=>"001000101",
  29860=>"010001111",
  29861=>"110100000",
  29862=>"010101011",
  29863=>"000111111",
  29864=>"100010010",
  29865=>"111010111",
  29866=>"100001110",
  29867=>"011011100",
  29868=>"100101011",
  29869=>"111101111",
  29870=>"001111010",
  29871=>"011100000",
  29872=>"001110100",
  29873=>"000000000",
  29874=>"110001110",
  29875=>"111111111",
  29876=>"110010101",
  29877=>"000001111",
  29878=>"001101010",
  29879=>"011101101",
  29880=>"010111111",
  29881=>"100101010",
  29882=>"101000100",
  29883=>"101101011",
  29884=>"011001110",
  29885=>"100101110",
  29886=>"010010101",
  29887=>"101000111",
  29888=>"111011100",
  29889=>"011010100",
  29890=>"001010100",
  29891=>"100110001",
  29892=>"111110000",
  29893=>"110011101",
  29894=>"111111111",
  29895=>"111000000",
  29896=>"010000100",
  29897=>"101101011",
  29898=>"000101111",
  29899=>"010100011",
  29900=>"100010010",
  29901=>"110000001",
  29902=>"000000000",
  29903=>"110000011",
  29904=>"110010110",
  29905=>"101001110",
  29906=>"010111111",
  29907=>"110110011",
  29908=>"011101001",
  29909=>"000000110",
  29910=>"000101001",
  29911=>"000101001",
  29912=>"110110000",
  29913=>"000000001",
  29914=>"001100001",
  29915=>"100110010",
  29916=>"000101110",
  29917=>"100010000",
  29918=>"011001000",
  29919=>"001011010",
  29920=>"110000000",
  29921=>"111111111",
  29922=>"000111011",
  29923=>"000111110",
  29924=>"110000110",
  29925=>"000010011",
  29926=>"010011100",
  29927=>"000000100",
  29928=>"010010001",
  29929=>"011011001",
  29930=>"010101010",
  29931=>"011111010",
  29932=>"101111110",
  29933=>"001001011",
  29934=>"111000000",
  29935=>"000110001",
  29936=>"111011101",
  29937=>"001000101",
  29938=>"000011000",
  29939=>"001100001",
  29940=>"001101001",
  29941=>"001100101",
  29942=>"110010011",
  29943=>"001001100",
  29944=>"001011010",
  29945=>"000000110",
  29946=>"111001110",
  29947=>"000001111",
  29948=>"000001100",
  29949=>"011010011",
  29950=>"000010111",
  29951=>"100010101",
  29952=>"011001000",
  29953=>"011010110",
  29954=>"100000100",
  29955=>"100000010",
  29956=>"011000101",
  29957=>"001100100",
  29958=>"101010001",
  29959=>"011011100",
  29960=>"000001001",
  29961=>"010010110",
  29962=>"001101010",
  29963=>"010000101",
  29964=>"001001111",
  29965=>"100011000",
  29966=>"010110001",
  29967=>"110101110",
  29968=>"001000111",
  29969=>"000001011",
  29970=>"001001110",
  29971=>"001110000",
  29972=>"011100010",
  29973=>"110001001",
  29974=>"110100111",
  29975=>"111011111",
  29976=>"001101101",
  29977=>"011010111",
  29978=>"100100100",
  29979=>"110100010",
  29980=>"111000110",
  29981=>"011110000",
  29982=>"000010000",
  29983=>"110101000",
  29984=>"101100111",
  29985=>"011101111",
  29986=>"011001111",
  29987=>"100100010",
  29988=>"110000010",
  29989=>"111100111",
  29990=>"001110100",
  29991=>"010111011",
  29992=>"001111001",
  29993=>"011101100",
  29994=>"100100011",
  29995=>"101111111",
  29996=>"100000101",
  29997=>"010000100",
  29998=>"100000010",
  29999=>"110011110",
  30000=>"100010001",
  30001=>"100011100",
  30002=>"110001010",
  30003=>"000001010",
  30004=>"001000011",
  30005=>"010001000",
  30006=>"100001011",
  30007=>"000111110",
  30008=>"010000111",
  30009=>"100110001",
  30010=>"011010110",
  30011=>"010100111",
  30012=>"000100000",
  30013=>"000011101",
  30014=>"110100001",
  30015=>"111111100",
  30016=>"100111001",
  30017=>"001101000",
  30018=>"110001010",
  30019=>"011010010",
  30020=>"100001111",
  30021=>"110101001",
  30022=>"010000010",
  30023=>"000010111",
  30024=>"011001001",
  30025=>"101001111",
  30026=>"010100111",
  30027=>"000111110",
  30028=>"000111100",
  30029=>"010100111",
  30030=>"100101100",
  30031=>"110110100",
  30032=>"100100110",
  30033=>"111010001",
  30034=>"000010000",
  30035=>"111001011",
  30036=>"011111011",
  30037=>"010110010",
  30038=>"111010110",
  30039=>"100111010",
  30040=>"000100101",
  30041=>"010110010",
  30042=>"110100111",
  30043=>"001111010",
  30044=>"101110000",
  30045=>"110101000",
  30046=>"000000000",
  30047=>"101000010",
  30048=>"111111111",
  30049=>"111101000",
  30050=>"000000010",
  30051=>"010000001",
  30052=>"010111001",
  30053=>"011100010",
  30054=>"110101010",
  30055=>"000110101",
  30056=>"110000010",
  30057=>"000110111",
  30058=>"111011010",
  30059=>"101101101",
  30060=>"011001001",
  30061=>"001001001",
  30062=>"010111110",
  30063=>"011111100",
  30064=>"111000000",
  30065=>"101011100",
  30066=>"111110011",
  30067=>"111101011",
  30068=>"110110101",
  30069=>"011101110",
  30070=>"100111001",
  30071=>"010100001",
  30072=>"111001011",
  30073=>"101000011",
  30074=>"010111011",
  30075=>"010001011",
  30076=>"101110110",
  30077=>"111110111",
  30078=>"111100111",
  30079=>"100100010",
  30080=>"111101111",
  30081=>"110000100",
  30082=>"001111011",
  30083=>"101110100",
  30084=>"010101111",
  30085=>"111010100",
  30086=>"011011111",
  30087=>"111010101",
  30088=>"010111110",
  30089=>"111100110",
  30090=>"100001100",
  30091=>"010100111",
  30092=>"111101001",
  30093=>"001111100",
  30094=>"000110100",
  30095=>"011100101",
  30096=>"001110111",
  30097=>"000010101",
  30098=>"101011100",
  30099=>"010111110",
  30100=>"100110000",
  30101=>"001100111",
  30102=>"000010000",
  30103=>"101001001",
  30104=>"101000101",
  30105=>"110001110",
  30106=>"000001111",
  30107=>"111100111",
  30108=>"011010101",
  30109=>"000000000",
  30110=>"000010011",
  30111=>"010000001",
  30112=>"010010000",
  30113=>"010101010",
  30114=>"001001111",
  30115=>"011000000",
  30116=>"000100100",
  30117=>"000010001",
  30118=>"101011010",
  30119=>"011111100",
  30120=>"100001011",
  30121=>"101111100",
  30122=>"000000000",
  30123=>"100000101",
  30124=>"000011011",
  30125=>"101010001",
  30126=>"110111011",
  30127=>"100110101",
  30128=>"001101101",
  30129=>"111100111",
  30130=>"000011000",
  30131=>"110111011",
  30132=>"001100111",
  30133=>"011011111",
  30134=>"110000101",
  30135=>"001101100",
  30136=>"011101000",
  30137=>"100000111",
  30138=>"001101010",
  30139=>"010011001",
  30140=>"111100010",
  30141=>"111001110",
  30142=>"100101111",
  30143=>"111110101",
  30144=>"001010110",
  30145=>"110011000",
  30146=>"000101010",
  30147=>"111111011",
  30148=>"010110010",
  30149=>"100111100",
  30150=>"111010101",
  30151=>"111000010",
  30152=>"111110011",
  30153=>"001001011",
  30154=>"110001001",
  30155=>"111111100",
  30156=>"111100011",
  30157=>"011001011",
  30158=>"001100101",
  30159=>"010010000",
  30160=>"101110001",
  30161=>"101001100",
  30162=>"010110001",
  30163=>"001010000",
  30164=>"110011110",
  30165=>"110111011",
  30166=>"011000111",
  30167=>"111001100",
  30168=>"000001101",
  30169=>"111111111",
  30170=>"110111011",
  30171=>"110011011",
  30172=>"001101000",
  30173=>"101010110",
  30174=>"010001111",
  30175=>"110110001",
  30176=>"000110110",
  30177=>"000110001",
  30178=>"110101000",
  30179=>"000011100",
  30180=>"100101000",
  30181=>"101100111",
  30182=>"101101110",
  30183=>"101110011",
  30184=>"100101011",
  30185=>"010111000",
  30186=>"101001011",
  30187=>"111110101",
  30188=>"000100100",
  30189=>"000001101",
  30190=>"111100101",
  30191=>"110111111",
  30192=>"001010110",
  30193=>"101100010",
  30194=>"101101110",
  30195=>"000010010",
  30196=>"000001000",
  30197=>"010110100",
  30198=>"000111111",
  30199=>"010001110",
  30200=>"111001000",
  30201=>"110000001",
  30202=>"101011111",
  30203=>"110010011",
  30204=>"111001101",
  30205=>"000101010",
  30206=>"110111001",
  30207=>"101111101",
  30208=>"001000101",
  30209=>"001101110",
  30210=>"110000100",
  30211=>"010110111",
  30212=>"111100111",
  30213=>"000110101",
  30214=>"001101111",
  30215=>"001000110",
  30216=>"001000110",
  30217=>"111111011",
  30218=>"111100100",
  30219=>"000001110",
  30220=>"111001110",
  30221=>"000000100",
  30222=>"111001010",
  30223=>"101111111",
  30224=>"100111011",
  30225=>"000000010",
  30226=>"111101001",
  30227=>"011000001",
  30228=>"001010000",
  30229=>"001100101",
  30230=>"111001101",
  30231=>"010101000",
  30232=>"111101000",
  30233=>"010000111",
  30234=>"001101101",
  30235=>"011110011",
  30236=>"001011010",
  30237=>"001111101",
  30238=>"011001110",
  30239=>"100101101",
  30240=>"011010111",
  30241=>"101010110",
  30242=>"010110000",
  30243=>"000110100",
  30244=>"101010111",
  30245=>"111000001",
  30246=>"001010000",
  30247=>"010011110",
  30248=>"000100000",
  30249=>"110101111",
  30250=>"010001100",
  30251=>"001101100",
  30252=>"011011001",
  30253=>"100100111",
  30254=>"100110111",
  30255=>"000000011",
  30256=>"100100010",
  30257=>"101110110",
  30258=>"001011110",
  30259=>"101110000",
  30260=>"000101110",
  30261=>"011010000",
  30262=>"010100000",
  30263=>"101101101",
  30264=>"001000000",
  30265=>"001011001",
  30266=>"101010001",
  30267=>"001000110",
  30268=>"001111100",
  30269=>"111001000",
  30270=>"011011010",
  30271=>"110101100",
  30272=>"000111110",
  30273=>"001101110",
  30274=>"100110000",
  30275=>"110111110",
  30276=>"010110000",
  30277=>"111010111",
  30278=>"110000100",
  30279=>"110011000",
  30280=>"110110110",
  30281=>"001001000",
  30282=>"001101100",
  30283=>"101000111",
  30284=>"001110110",
  30285=>"011101111",
  30286=>"110010011",
  30287=>"101111010",
  30288=>"000011010",
  30289=>"101101111",
  30290=>"010111101",
  30291=>"000011101",
  30292=>"000100100",
  30293=>"010110010",
  30294=>"100101110",
  30295=>"001010001",
  30296=>"111000010",
  30297=>"111111100",
  30298=>"011001000",
  30299=>"110001000",
  30300=>"000110111",
  30301=>"111111110",
  30302=>"101010001",
  30303=>"000110110",
  30304=>"100001001",
  30305=>"010001000",
  30306=>"111111101",
  30307=>"100011001",
  30308=>"101011101",
  30309=>"010000100",
  30310=>"111011010",
  30311=>"010110101",
  30312=>"110011100",
  30313=>"010100000",
  30314=>"110010111",
  30315=>"111000000",
  30316=>"100010011",
  30317=>"010100111",
  30318=>"101101011",
  30319=>"110111010",
  30320=>"001011000",
  30321=>"001001111",
  30322=>"011010110",
  30323=>"011000101",
  30324=>"110010110",
  30325=>"111101001",
  30326=>"100101100",
  30327=>"000101110",
  30328=>"011011011",
  30329=>"010110110",
  30330=>"111101000",
  30331=>"001001011",
  30332=>"111111110",
  30333=>"101000101",
  30334=>"111010111",
  30335=>"011010000",
  30336=>"101010000",
  30337=>"110101110",
  30338=>"011001011",
  30339=>"101101101",
  30340=>"100001001",
  30341=>"111111001",
  30342=>"000110110",
  30343=>"100101111",
  30344=>"011000011",
  30345=>"011000001",
  30346=>"111010101",
  30347=>"101111001",
  30348=>"000000111",
  30349=>"111111111",
  30350=>"110000001",
  30351=>"011001000",
  30352=>"010111100",
  30353=>"010001000",
  30354=>"001010110",
  30355=>"101001101",
  30356=>"010000111",
  30357=>"000111010",
  30358=>"100000101",
  30359=>"000011100",
  30360=>"110100111",
  30361=>"000111111",
  30362=>"000110100",
  30363=>"110011001",
  30364=>"101001111",
  30365=>"110110111",
  30366=>"000001000",
  30367=>"011011100",
  30368=>"000010000",
  30369=>"001000000",
  30370=>"011101000",
  30371=>"000000010",
  30372=>"101011111",
  30373=>"100010100",
  30374=>"011111000",
  30375=>"000000111",
  30376=>"011011100",
  30377=>"101110110",
  30378=>"000111101",
  30379=>"110001111",
  30380=>"101011010",
  30381=>"101100011",
  30382=>"001101110",
  30383=>"111101101",
  30384=>"000110111",
  30385=>"100100100",
  30386=>"101000110",
  30387=>"110111111",
  30388=>"000000100",
  30389=>"101011111",
  30390=>"110111001",
  30391=>"111000100",
  30392=>"011111011",
  30393=>"110001100",
  30394=>"011011101",
  30395=>"111101011",
  30396=>"111010111",
  30397=>"111000101",
  30398=>"000111101",
  30399=>"100100111",
  30400=>"101000001",
  30401=>"101111101",
  30402=>"111100100",
  30403=>"001000011",
  30404=>"111001110",
  30405=>"101011001",
  30406=>"100011110",
  30407=>"001010011",
  30408=>"011110101",
  30409=>"110101000",
  30410=>"000011100",
  30411=>"000100111",
  30412=>"000001101",
  30413=>"000000101",
  30414=>"001100101",
  30415=>"010001011",
  30416=>"111110100",
  30417=>"101010000",
  30418=>"111010011",
  30419=>"010100100",
  30420=>"001110011",
  30421=>"000111000",
  30422=>"001001000",
  30423=>"001001011",
  30424=>"000011000",
  30425=>"011010011",
  30426=>"111100010",
  30427=>"010101000",
  30428=>"011111000",
  30429=>"010110101",
  30430=>"100110000",
  30431=>"100000011",
  30432=>"001010000",
  30433=>"010010101",
  30434=>"101000110",
  30435=>"100101101",
  30436=>"010001101",
  30437=>"111110101",
  30438=>"110010000",
  30439=>"100101111",
  30440=>"011011111",
  30441=>"001111010",
  30442=>"101000010",
  30443=>"101111110",
  30444=>"011010101",
  30445=>"011101111",
  30446=>"100001011",
  30447=>"100011011",
  30448=>"000011100",
  30449=>"100110000",
  30450=>"100000110",
  30451=>"111010011",
  30452=>"010000010",
  30453=>"100101101",
  30454=>"000010011",
  30455=>"010011001",
  30456=>"101111011",
  30457=>"100010101",
  30458=>"000000110",
  30459=>"000011011",
  30460=>"100111000",
  30461=>"010011110",
  30462=>"001001111",
  30463=>"011111111",
  30464=>"100110000",
  30465=>"011010100",
  30466=>"101110110",
  30467=>"111110100",
  30468=>"110110010",
  30469=>"110111001",
  30470=>"000010110",
  30471=>"001010011",
  30472=>"100100111",
  30473=>"111111110",
  30474=>"110010100",
  30475=>"111110100",
  30476=>"010011010",
  30477=>"001011011",
  30478=>"111100111",
  30479=>"011001100",
  30480=>"010010101",
  30481=>"011100001",
  30482=>"101101011",
  30483=>"011101010",
  30484=>"001010100",
  30485=>"010111110",
  30486=>"000110100",
  30487=>"111111010",
  30488=>"011011010",
  30489=>"010101101",
  30490=>"111011101",
  30491=>"101000100",
  30492=>"111101111",
  30493=>"111111010",
  30494=>"101101101",
  30495=>"101101101",
  30496=>"010101111",
  30497=>"010011011",
  30498=>"111101101",
  30499=>"010011010",
  30500=>"001101011",
  30501=>"111101101",
  30502=>"000111110",
  30503=>"101111110",
  30504=>"010010111",
  30505=>"000000000",
  30506=>"101010011",
  30507=>"000110111",
  30508=>"001011110",
  30509=>"000000011",
  30510=>"010001110",
  30511=>"110100110",
  30512=>"000000000",
  30513=>"110110010",
  30514=>"100000010",
  30515=>"111110110",
  30516=>"110100100",
  30517=>"000001101",
  30518=>"110000010",
  30519=>"011101110",
  30520=>"110011000",
  30521=>"101100011",
  30522=>"111010110",
  30523=>"110000110",
  30524=>"101001100",
  30525=>"011000100",
  30526=>"101000011",
  30527=>"100110110",
  30528=>"011001001",
  30529=>"010111011",
  30530=>"010000000",
  30531=>"110001010",
  30532=>"110110101",
  30533=>"101001101",
  30534=>"011111111",
  30535=>"110110010",
  30536=>"010001001",
  30537=>"101001011",
  30538=>"010100000",
  30539=>"010000100",
  30540=>"000001001",
  30541=>"111011110",
  30542=>"101111001",
  30543=>"110101001",
  30544=>"110000111",
  30545=>"000100011",
  30546=>"101011111",
  30547=>"010011001",
  30548=>"010011111",
  30549=>"000000111",
  30550=>"101010111",
  30551=>"000000010",
  30552=>"101101000",
  30553=>"001010110",
  30554=>"101000111",
  30555=>"000000111",
  30556=>"111111101",
  30557=>"010001011",
  30558=>"000101110",
  30559=>"111001111",
  30560=>"101100111",
  30561=>"110111100",
  30562=>"111011110",
  30563=>"111011101",
  30564=>"010111000",
  30565=>"000010001",
  30566=>"111111010",
  30567=>"110101000",
  30568=>"000101001",
  30569=>"011011100",
  30570=>"010010000",
  30571=>"010110101",
  30572=>"010011011",
  30573=>"111000000",
  30574=>"111111010",
  30575=>"111000000",
  30576=>"110001111",
  30577=>"000001101",
  30578=>"101110100",
  30579=>"010101000",
  30580=>"000010010",
  30581=>"000001100",
  30582=>"011010111",
  30583=>"111011010",
  30584=>"100000000",
  30585=>"001111010",
  30586=>"110111011",
  30587=>"000111011",
  30588=>"000000101",
  30589=>"100000011",
  30590=>"000110010",
  30591=>"001010100",
  30592=>"101111010",
  30593=>"000000110",
  30594=>"001110100",
  30595=>"100000100",
  30596=>"100000010",
  30597=>"110100000",
  30598=>"110101110",
  30599=>"000001100",
  30600=>"010101010",
  30601=>"110111110",
  30602=>"110111111",
  30603=>"000100010",
  30604=>"000111110",
  30605=>"101001000",
  30606=>"111000100",
  30607=>"110001010",
  30608=>"111010011",
  30609=>"111000010",
  30610=>"011101001",
  30611=>"101001000",
  30612=>"011110100",
  30613=>"100011110",
  30614=>"101101001",
  30615=>"100010111",
  30616=>"111000101",
  30617=>"001001001",
  30618=>"010010110",
  30619=>"101000000",
  30620=>"011001111",
  30621=>"111000000",
  30622=>"111010000",
  30623=>"000111011",
  30624=>"010111000",
  30625=>"100110111",
  30626=>"111000000",
  30627=>"111011100",
  30628=>"111110111",
  30629=>"001001010",
  30630=>"111110001",
  30631=>"010111001",
  30632=>"101100111",
  30633=>"000011100",
  30634=>"111111100",
  30635=>"110001010",
  30636=>"001010101",
  30637=>"100001011",
  30638=>"111111111",
  30639=>"011010111",
  30640=>"000100000",
  30641=>"101000101",
  30642=>"010011101",
  30643=>"001000000",
  30644=>"001000100",
  30645=>"110001101",
  30646=>"001100110",
  30647=>"010001101",
  30648=>"111011010",
  30649=>"010010011",
  30650=>"110111111",
  30651=>"110110011",
  30652=>"001000000",
  30653=>"111100110",
  30654=>"111100111",
  30655=>"001001000",
  30656=>"001101000",
  30657=>"101111101",
  30658=>"001101001",
  30659=>"000001010",
  30660=>"101001100",
  30661=>"010010111",
  30662=>"010011001",
  30663=>"000100011",
  30664=>"100010001",
  30665=>"111100101",
  30666=>"011000111",
  30667=>"011010010",
  30668=>"010101010",
  30669=>"100100111",
  30670=>"111011101",
  30671=>"001010000",
  30672=>"011000100",
  30673=>"110001111",
  30674=>"111010011",
  30675=>"100100100",
  30676=>"111011111",
  30677=>"010011000",
  30678=>"000000011",
  30679=>"010001111",
  30680=>"001100111",
  30681=>"000101001",
  30682=>"010100111",
  30683=>"010000110",
  30684=>"110000010",
  30685=>"011001110",
  30686=>"001010010",
  30687=>"000111101",
  30688=>"001110011",
  30689=>"101100101",
  30690=>"011100000",
  30691=>"001101111",
  30692=>"101011111",
  30693=>"000110010",
  30694=>"011111110",
  30695=>"011111011",
  30696=>"000000010",
  30697=>"111101011",
  30698=>"001000001",
  30699=>"011011110",
  30700=>"100110111",
  30701=>"001011110",
  30702=>"101111010",
  30703=>"011011011",
  30704=>"000010011",
  30705=>"111011001",
  30706=>"110111110",
  30707=>"111011100",
  30708=>"100001111",
  30709=>"110111101",
  30710=>"110110011",
  30711=>"111001011",
  30712=>"000010010",
  30713=>"100100101",
  30714=>"000100111",
  30715=>"110101011",
  30716=>"000011111",
  30717=>"001110001",
  30718=>"000000011",
  30719=>"011110101",
  30720=>"001000010",
  30721=>"000110010",
  30722=>"101000000",
  30723=>"011001101",
  30724=>"011011111",
  30725=>"100010111",
  30726=>"011101110",
  30727=>"011010110",
  30728=>"110010010",
  30729=>"110110001",
  30730=>"011010101",
  30731=>"101011000",
  30732=>"110111100",
  30733=>"001001000",
  30734=>"100001011",
  30735=>"111101000",
  30736=>"100001010",
  30737=>"101011000",
  30738=>"101110011",
  30739=>"110110011",
  30740=>"111011101",
  30741=>"111100000",
  30742=>"111001010",
  30743=>"111111010",
  30744=>"100101001",
  30745=>"100110110",
  30746=>"000010101",
  30747=>"001100110",
  30748=>"100110000",
  30749=>"000100010",
  30750=>"011111001",
  30751=>"100110010",
  30752=>"110011011",
  30753=>"111010011",
  30754=>"100110101",
  30755=>"110101011",
  30756=>"001101101",
  30757=>"111111100",
  30758=>"110110111",
  30759=>"101101011",
  30760=>"001101010",
  30761=>"100010101",
  30762=>"000100010",
  30763=>"100001011",
  30764=>"100111010",
  30765=>"111111011",
  30766=>"001111111",
  30767=>"111100111",
  30768=>"001000000",
  30769=>"100111001",
  30770=>"101100000",
  30771=>"100100010",
  30772=>"011111001",
  30773=>"101101000",
  30774=>"010101100",
  30775=>"111101001",
  30776=>"011100011",
  30777=>"001110101",
  30778=>"000101111",
  30779=>"110010111",
  30780=>"011000011",
  30781=>"111001110",
  30782=>"111000000",
  30783=>"101100101",
  30784=>"110001110",
  30785=>"000011101",
  30786=>"110110111",
  30787=>"110000110",
  30788=>"010100001",
  30789=>"010110011",
  30790=>"111101111",
  30791=>"001010010",
  30792=>"001001000",
  30793=>"100111011",
  30794=>"000000000",
  30795=>"100000000",
  30796=>"110010000",
  30797=>"101000111",
  30798=>"111010000",
  30799=>"001110110",
  30800=>"000101011",
  30801=>"111101111",
  30802=>"110100110",
  30803=>"011000010",
  30804=>"000000111",
  30805=>"100111110",
  30806=>"000000010",
  30807=>"000100000",
  30808=>"010001010",
  30809=>"111110101",
  30810=>"000010111",
  30811=>"011100000",
  30812=>"111100110",
  30813=>"111011111",
  30814=>"111110010",
  30815=>"001111111",
  30816=>"000101000",
  30817=>"101100110",
  30818=>"001110111",
  30819=>"100001111",
  30820=>"110011101",
  30821=>"101101111",
  30822=>"100100011",
  30823=>"011010110",
  30824=>"010101101",
  30825=>"001111111",
  30826=>"001100111",
  30827=>"001011100",
  30828=>"011101101",
  30829=>"000001111",
  30830=>"110110111",
  30831=>"100000100",
  30832=>"011001001",
  30833=>"101110111",
  30834=>"111100001",
  30835=>"010010110",
  30836=>"001001011",
  30837=>"110011010",
  30838=>"111010001",
  30839=>"100111011",
  30840=>"011100110",
  30841=>"110101001",
  30842=>"000010100",
  30843=>"010011111",
  30844=>"010000111",
  30845=>"100010011",
  30846=>"111110000",
  30847=>"011100010",
  30848=>"110000010",
  30849=>"110001100",
  30850=>"111011111",
  30851=>"010100100",
  30852=>"011101110",
  30853=>"010110111",
  30854=>"111011111",
  30855=>"101110101",
  30856=>"111100101",
  30857=>"011000110",
  30858=>"001010110",
  30859=>"000100011",
  30860=>"101111110",
  30861=>"100011010",
  30862=>"011000000",
  30863=>"100011000",
  30864=>"000010101",
  30865=>"000010101",
  30866=>"100010000",
  30867=>"001001000",
  30868=>"011001000",
  30869=>"110010000",
  30870=>"110111010",
  30871=>"000111011",
  30872=>"100010010",
  30873=>"011110111",
  30874=>"001001010",
  30875=>"011010001",
  30876=>"010000110",
  30877=>"101111001",
  30878=>"000010101",
  30879=>"011101101",
  30880=>"000110010",
  30881=>"001110010",
  30882=>"110110010",
  30883=>"101011101",
  30884=>"011011001",
  30885=>"001010100",
  30886=>"000100000",
  30887=>"011100011",
  30888=>"111101011",
  30889=>"001111101",
  30890=>"001001100",
  30891=>"101111101",
  30892=>"000110110",
  30893=>"000110011",
  30894=>"111111011",
  30895=>"100111100",
  30896=>"010011101",
  30897=>"111000000",
  30898=>"111010101",
  30899=>"001110000",
  30900=>"111110011",
  30901=>"001011011",
  30902=>"000101001",
  30903=>"100100011",
  30904=>"110100100",
  30905=>"001001010",
  30906=>"111001110",
  30907=>"111001111",
  30908=>"101010110",
  30909=>"101011110",
  30910=>"001010001",
  30911=>"100011100",
  30912=>"001111111",
  30913=>"000010100",
  30914=>"101011111",
  30915=>"011001111",
  30916=>"100101011",
  30917=>"000111101",
  30918=>"010010100",
  30919=>"010010101",
  30920=>"100011111",
  30921=>"111011111",
  30922=>"111001011",
  30923=>"101010110",
  30924=>"110111001",
  30925=>"011110001",
  30926=>"100000010",
  30927=>"110101111",
  30928=>"010010111",
  30929=>"110011111",
  30930=>"110111101",
  30931=>"100010011",
  30932=>"110101011",
  30933=>"100110011",
  30934=>"111110001",
  30935=>"001010000",
  30936=>"111011001",
  30937=>"100000001",
  30938=>"001011100",
  30939=>"110101111",
  30940=>"100011100",
  30941=>"110111010",
  30942=>"001100101",
  30943=>"110101011",
  30944=>"111100111",
  30945=>"001110100",
  30946=>"110110000",
  30947=>"011100100",
  30948=>"000000111",
  30949=>"100010010",
  30950=>"100100101",
  30951=>"000100100",
  30952=>"000100100",
  30953=>"010000101",
  30954=>"001100000",
  30955=>"001110010",
  30956=>"101000010",
  30957=>"001101100",
  30958=>"001111111",
  30959=>"001101000",
  30960=>"001011000",
  30961=>"101001110",
  30962=>"101110000",
  30963=>"001101010",
  30964=>"111110010",
  30965=>"000101010",
  30966=>"100001110",
  30967=>"110001001",
  30968=>"011101110",
  30969=>"001101111",
  30970=>"101100001",
  30971=>"100010100",
  30972=>"100110101",
  30973=>"001100111",
  30974=>"011010000",
  30975=>"101000010",
  30976=>"110011011",
  30977=>"101111101",
  30978=>"010110110",
  30979=>"110111001",
  30980=>"100111011",
  30981=>"011111100",
  30982=>"000011010",
  30983=>"011011111",
  30984=>"010000100",
  30985=>"100100010",
  30986=>"001111011",
  30987=>"001010110",
  30988=>"111100011",
  30989=>"101011001",
  30990=>"000110010",
  30991=>"101111111",
  30992=>"001100101",
  30993=>"010011010",
  30994=>"111000000",
  30995=>"111110100",
  30996=>"110100001",
  30997=>"111110111",
  30998=>"101110100",
  30999=>"101101101",
  31000=>"100111111",
  31001=>"001101000",
  31002=>"011010010",
  31003=>"100110001",
  31004=>"110101011",
  31005=>"011111011",
  31006=>"111101100",
  31007=>"100100010",
  31008=>"000101111",
  31009=>"101111101",
  31010=>"110010110",
  31011=>"100001011",
  31012=>"010100010",
  31013=>"111100100",
  31014=>"010010010",
  31015=>"100011100",
  31016=>"010011011",
  31017=>"000010001",
  31018=>"001100111",
  31019=>"111110100",
  31020=>"001000001",
  31021=>"100110001",
  31022=>"111000111",
  31023=>"100101101",
  31024=>"010010001",
  31025=>"111101011",
  31026=>"001000000",
  31027=>"111111110",
  31028=>"111111101",
  31029=>"000001001",
  31030=>"000110101",
  31031=>"011111110",
  31032=>"001111000",
  31033=>"101111101",
  31034=>"111100111",
  31035=>"110011100",
  31036=>"110100001",
  31037=>"001010011",
  31038=>"001000011",
  31039=>"110001010",
  31040=>"101001011",
  31041=>"110101100",
  31042=>"100101010",
  31043=>"011110010",
  31044=>"110111110",
  31045=>"100011010",
  31046=>"001000011",
  31047=>"101100011",
  31048=>"010010010",
  31049=>"101110111",
  31050=>"110011101",
  31051=>"000000001",
  31052=>"101100101",
  31053=>"110010001",
  31054=>"111101111",
  31055=>"101111111",
  31056=>"011101111",
  31057=>"111000110",
  31058=>"011000111",
  31059=>"110001100",
  31060=>"001111000",
  31061=>"011100101",
  31062=>"101010101",
  31063=>"001000000",
  31064=>"100100110",
  31065=>"011101110",
  31066=>"100101110",
  31067=>"000010111",
  31068=>"101000001",
  31069=>"110000111",
  31070=>"101101111",
  31071=>"000000101",
  31072=>"011111100",
  31073=>"011101010",
  31074=>"111100100",
  31075=>"101011001",
  31076=>"100000101",
  31077=>"000100101",
  31078=>"110111010",
  31079=>"011100011",
  31080=>"000110011",
  31081=>"000000000",
  31082=>"000001011",
  31083=>"000110000",
  31084=>"101111001",
  31085=>"111011010",
  31086=>"000110100",
  31087=>"001010101",
  31088=>"001100101",
  31089=>"111110110",
  31090=>"010111011",
  31091=>"110001001",
  31092=>"110111101",
  31093=>"100001001",
  31094=>"111100110",
  31095=>"011001110",
  31096=>"111001100",
  31097=>"111000100",
  31098=>"001110101",
  31099=>"110010100",
  31100=>"111011101",
  31101=>"001000011",
  31102=>"001111011",
  31103=>"011000100",
  31104=>"000000011",
  31105=>"111001011",
  31106=>"000110010",
  31107=>"111101011",
  31108=>"100110100",
  31109=>"000100010",
  31110=>"000110011",
  31111=>"110000000",
  31112=>"010001011",
  31113=>"111101111",
  31114=>"100010011",
  31115=>"110100000",
  31116=>"000000010",
  31117=>"000110000",
  31118=>"001000110",
  31119=>"100011101",
  31120=>"101011001",
  31121=>"001100010",
  31122=>"110100011",
  31123=>"101110010",
  31124=>"111110101",
  31125=>"010101110",
  31126=>"100001010",
  31127=>"000000011",
  31128=>"100000111",
  31129=>"111110101",
  31130=>"101101000",
  31131=>"111011001",
  31132=>"010010111",
  31133=>"000110110",
  31134=>"001101010",
  31135=>"111000100",
  31136=>"101110111",
  31137=>"101011000",
  31138=>"111010000",
  31139=>"001000001",
  31140=>"000001001",
  31141=>"110000101",
  31142=>"011101001",
  31143=>"000011100",
  31144=>"101000000",
  31145=>"101100111",
  31146=>"110101011",
  31147=>"110001110",
  31148=>"111100011",
  31149=>"000100011",
  31150=>"111110011",
  31151=>"000101110",
  31152=>"100000100",
  31153=>"110110010",
  31154=>"000100010",
  31155=>"011111110",
  31156=>"111001100",
  31157=>"100110111",
  31158=>"111001110",
  31159=>"101010100",
  31160=>"011101101",
  31161=>"001111101",
  31162=>"010010010",
  31163=>"010011010",
  31164=>"100111110",
  31165=>"100110110",
  31166=>"011000110",
  31167=>"111110001",
  31168=>"011111000",
  31169=>"000100110",
  31170=>"010010001",
  31171=>"110111001",
  31172=>"111110011",
  31173=>"000000011",
  31174=>"000010000",
  31175=>"110001001",
  31176=>"000101110",
  31177=>"101101011",
  31178=>"011011111",
  31179=>"100010111",
  31180=>"100111110",
  31181=>"010100101",
  31182=>"001011000",
  31183=>"100110000",
  31184=>"101111111",
  31185=>"100110110",
  31186=>"000110111",
  31187=>"011010110",
  31188=>"101101101",
  31189=>"110001000",
  31190=>"101001001",
  31191=>"000010001",
  31192=>"110011111",
  31193=>"001111000",
  31194=>"000110000",
  31195=>"000000110",
  31196=>"000000010",
  31197=>"000000000",
  31198=>"100110001",
  31199=>"110001000",
  31200=>"111110010",
  31201=>"101110110",
  31202=>"000010000",
  31203=>"001001001",
  31204=>"000010110",
  31205=>"000010000",
  31206=>"010011101",
  31207=>"100001100",
  31208=>"001000000",
  31209=>"110001011",
  31210=>"010010010",
  31211=>"110010001",
  31212=>"010011010",
  31213=>"001000001",
  31214=>"001000110",
  31215=>"001011010",
  31216=>"100001110",
  31217=>"011100101",
  31218=>"111000101",
  31219=>"011111000",
  31220=>"001001101",
  31221=>"010010010",
  31222=>"011000101",
  31223=>"110110101",
  31224=>"010000110",
  31225=>"110101000",
  31226=>"001010101",
  31227=>"101011100",
  31228=>"111001001",
  31229=>"000110001",
  31230=>"010001100",
  31231=>"100110110",
  31232=>"101111101",
  31233=>"001101000",
  31234=>"101011011",
  31235=>"110101011",
  31236=>"111010010",
  31237=>"111010110",
  31238=>"001110001",
  31239=>"111011011",
  31240=>"100000101",
  31241=>"111101100",
  31242=>"000001010",
  31243=>"000000010",
  31244=>"011011110",
  31245=>"000011000",
  31246=>"101001001",
  31247=>"100011010",
  31248=>"101100001",
  31249=>"011010010",
  31250=>"100111110",
  31251=>"011111111",
  31252=>"010001011",
  31253=>"010111100",
  31254=>"010000011",
  31255=>"100110100",
  31256=>"101010101",
  31257=>"011000111",
  31258=>"100100011",
  31259=>"010110001",
  31260=>"111001010",
  31261=>"101100010",
  31262=>"110101111",
  31263=>"101111101",
  31264=>"100101111",
  31265=>"101110110",
  31266=>"101001011",
  31267=>"111100011",
  31268=>"101111110",
  31269=>"000001011",
  31270=>"111000000",
  31271=>"100001010",
  31272=>"010010100",
  31273=>"000000111",
  31274=>"000111011",
  31275=>"000100110",
  31276=>"000110110",
  31277=>"111111111",
  31278=>"000101011",
  31279=>"000001000",
  31280=>"010110101",
  31281=>"101000110",
  31282=>"100001110",
  31283=>"110010100",
  31284=>"111101110",
  31285=>"000110010",
  31286=>"110000001",
  31287=>"101111110",
  31288=>"111101100",
  31289=>"100001001",
  31290=>"010101100",
  31291=>"011011000",
  31292=>"101110100",
  31293=>"110111011",
  31294=>"000000101",
  31295=>"100000100",
  31296=>"101111001",
  31297=>"100010110",
  31298=>"111000011",
  31299=>"111111111",
  31300=>"001110001",
  31301=>"101011100",
  31302=>"000000101",
  31303=>"010100000",
  31304=>"001011001",
  31305=>"011111110",
  31306=>"000010011",
  31307=>"000000110",
  31308=>"100000111",
  31309=>"010011110",
  31310=>"010011011",
  31311=>"110011100",
  31312=>"010000010",
  31313=>"011101100",
  31314=>"010110011",
  31315=>"111111100",
  31316=>"000111111",
  31317=>"000101010",
  31318=>"001111111",
  31319=>"011010100",
  31320=>"011101011",
  31321=>"111000011",
  31322=>"111011101",
  31323=>"111110011",
  31324=>"111111111",
  31325=>"100111011",
  31326=>"011010001",
  31327=>"011101100",
  31328=>"000100011",
  31329=>"001001111",
  31330=>"001000100",
  31331=>"010101101",
  31332=>"111110100",
  31333=>"011100100",
  31334=>"100100110",
  31335=>"000001101",
  31336=>"110010000",
  31337=>"011010110",
  31338=>"100101101",
  31339=>"000101000",
  31340=>"011111101",
  31341=>"100010011",
  31342=>"110111101",
  31343=>"110011100",
  31344=>"100010110",
  31345=>"000001000",
  31346=>"100110111",
  31347=>"010000110",
  31348=>"100011011",
  31349=>"111010101",
  31350=>"111111100",
  31351=>"111110011",
  31352=>"100101000",
  31353=>"111000110",
  31354=>"000010001",
  31355=>"111001001",
  31356=>"110001001",
  31357=>"110111100",
  31358=>"111100001",
  31359=>"101000011",
  31360=>"010000100",
  31361=>"001001001",
  31362=>"111001011",
  31363=>"110111001",
  31364=>"101000011",
  31365=>"101111101",
  31366=>"010110000",
  31367=>"101111110",
  31368=>"110111000",
  31369=>"111000010",
  31370=>"100111010",
  31371=>"000100011",
  31372=>"110001111",
  31373=>"001111111",
  31374=>"111000110",
  31375=>"100111000",
  31376=>"101100111",
  31377=>"111100111",
  31378=>"101101001",
  31379=>"001001100",
  31380=>"000010111",
  31381=>"100111011",
  31382=>"101100100",
  31383=>"100100100",
  31384=>"011110000",
  31385=>"111111001",
  31386=>"010100000",
  31387=>"010110011",
  31388=>"110111100",
  31389=>"010000111",
  31390=>"111101011",
  31391=>"100010110",
  31392=>"000000110",
  31393=>"110100101",
  31394=>"000100010",
  31395=>"101111001",
  31396=>"011110100",
  31397=>"000011110",
  31398=>"011001010",
  31399=>"010000010",
  31400=>"000110000",
  31401=>"011010110",
  31402=>"100000100",
  31403=>"000001000",
  31404=>"110100001",
  31405=>"111111110",
  31406=>"000111011",
  31407=>"111011100",
  31408=>"101010001",
  31409=>"101010001",
  31410=>"001100011",
  31411=>"111000010",
  31412=>"111011100",
  31413=>"111110011",
  31414=>"101100011",
  31415=>"101100110",
  31416=>"110101100",
  31417=>"010000100",
  31418=>"000110000",
  31419=>"111100101",
  31420=>"001100101",
  31421=>"011010111",
  31422=>"100110100",
  31423=>"101110111",
  31424=>"010011111",
  31425=>"010111111",
  31426=>"101000010",
  31427=>"001110000",
  31428=>"000101100",
  31429=>"001100100",
  31430=>"011010001",
  31431=>"111010101",
  31432=>"110011010",
  31433=>"011010011",
  31434=>"001010100",
  31435=>"101110010",
  31436=>"100001000",
  31437=>"000000010",
  31438=>"110100100",
  31439=>"100010101",
  31440=>"101110011",
  31441=>"101110011",
  31442=>"000100100",
  31443=>"100000101",
  31444=>"101011011",
  31445=>"110000011",
  31446=>"101100101",
  31447=>"010011101",
  31448=>"100101101",
  31449=>"011110110",
  31450=>"000000001",
  31451=>"101000010",
  31452=>"111001111",
  31453=>"010010010",
  31454=>"101110010",
  31455=>"100010010",
  31456=>"010111010",
  31457=>"100000110",
  31458=>"010101110",
  31459=>"001000010",
  31460=>"010111110",
  31461=>"010010001",
  31462=>"100001111",
  31463=>"001100110",
  31464=>"110101111",
  31465=>"101000101",
  31466=>"011100010",
  31467=>"110100110",
  31468=>"001001001",
  31469=>"100010000",
  31470=>"000001111",
  31471=>"110001110",
  31472=>"111000110",
  31473=>"100001010",
  31474=>"101001001",
  31475=>"101011000",
  31476=>"010110010",
  31477=>"011010000",
  31478=>"111101001",
  31479=>"111101110",
  31480=>"010000001",
  31481=>"110101111",
  31482=>"100011111",
  31483=>"111011001",
  31484=>"101100100",
  31485=>"100010110",
  31486=>"010001011",
  31487=>"001011110",
  31488=>"011111101",
  31489=>"100010000",
  31490=>"110010010",
  31491=>"110000110",
  31492=>"101100101",
  31493=>"000010000",
  31494=>"100000000",
  31495=>"101010010",
  31496=>"000000000",
  31497=>"111000111",
  31498=>"110010011",
  31499=>"001101000",
  31500=>"011000000",
  31501=>"000101111",
  31502=>"011011000",
  31503=>"111000111",
  31504=>"111001010",
  31505=>"111111010",
  31506=>"001001000",
  31507=>"000010110",
  31508=>"100010101",
  31509=>"111000110",
  31510=>"011000000",
  31511=>"001111111",
  31512=>"111101110",
  31513=>"001111111",
  31514=>"100110100",
  31515=>"101001001",
  31516=>"100001010",
  31517=>"110100101",
  31518=>"010000011",
  31519=>"111111011",
  31520=>"111010001",
  31521=>"000000001",
  31522=>"000101101",
  31523=>"010100001",
  31524=>"100010010",
  31525=>"010000001",
  31526=>"111000010",
  31527=>"110001010",
  31528=>"000110110",
  31529=>"110000110",
  31530=>"000001100",
  31531=>"111000000",
  31532=>"010100011",
  31533=>"111110100",
  31534=>"011101111",
  31535=>"111100100",
  31536=>"111111100",
  31537=>"110000101",
  31538=>"011111110",
  31539=>"111100100",
  31540=>"010100000",
  31541=>"011100110",
  31542=>"110101000",
  31543=>"110111011",
  31544=>"010101001",
  31545=>"001111010",
  31546=>"100000000",
  31547=>"101110100",
  31548=>"001001011",
  31549=>"011110111",
  31550=>"011010101",
  31551=>"000011101",
  31552=>"100110001",
  31553=>"000000000",
  31554=>"001011101",
  31555=>"111010100",
  31556=>"111111010",
  31557=>"000111001",
  31558=>"101011001",
  31559=>"001101111",
  31560=>"000000100",
  31561=>"001010001",
  31562=>"000100110",
  31563=>"000000010",
  31564=>"100000110",
  31565=>"100100011",
  31566=>"011101000",
  31567=>"111110110",
  31568=>"010100111",
  31569=>"000110010",
  31570=>"101010111",
  31571=>"010001000",
  31572=>"101010100",
  31573=>"110011100",
  31574=>"100001111",
  31575=>"100001000",
  31576=>"100100010",
  31577=>"101001010",
  31578=>"011010010",
  31579=>"001110010",
  31580=>"010100000",
  31581=>"000010011",
  31582=>"111111001",
  31583=>"011110111",
  31584=>"000111001",
  31585=>"011111111",
  31586=>"001010110",
  31587=>"111111111",
  31588=>"111110000",
  31589=>"100110010",
  31590=>"010100000",
  31591=>"101011100",
  31592=>"110000000",
  31593=>"001000001",
  31594=>"110100000",
  31595=>"001100101",
  31596=>"010100011",
  31597=>"100111010",
  31598=>"100110001",
  31599=>"101000000",
  31600=>"110110100",
  31601=>"110111011",
  31602=>"110000011",
  31603=>"000101010",
  31604=>"110011010",
  31605=>"000011100",
  31606=>"000010010",
  31607=>"100010001",
  31608=>"101001010",
  31609=>"110110110",
  31610=>"000000101",
  31611=>"011110001",
  31612=>"010101111",
  31613=>"001011011",
  31614=>"100000001",
  31615=>"110110111",
  31616=>"100000010",
  31617=>"001000000",
  31618=>"101101111",
  31619=>"100000001",
  31620=>"111110110",
  31621=>"010110100",
  31622=>"011110000",
  31623=>"001000000",
  31624=>"001101111",
  31625=>"001011010",
  31626=>"000001010",
  31627=>"110110111",
  31628=>"111011111",
  31629=>"110101010",
  31630=>"100010000",
  31631=>"101010111",
  31632=>"111000001",
  31633=>"001001101",
  31634=>"111101111",
  31635=>"111110101",
  31636=>"010111000",
  31637=>"110011010",
  31638=>"001101011",
  31639=>"010101000",
  31640=>"011001011",
  31641=>"010011000",
  31642=>"011100011",
  31643=>"100001000",
  31644=>"111001110",
  31645=>"111111011",
  31646=>"100011101",
  31647=>"101100100",
  31648=>"100010010",
  31649=>"100010101",
  31650=>"100000100",
  31651=>"010101111",
  31652=>"010000000",
  31653=>"111011001",
  31654=>"100101110",
  31655=>"000000010",
  31656=>"101110000",
  31657=>"111101101",
  31658=>"110001111",
  31659=>"100001110",
  31660=>"001010100",
  31661=>"111111111",
  31662=>"111100100",
  31663=>"101101011",
  31664=>"010100010",
  31665=>"001000010",
  31666=>"011001011",
  31667=>"001000100",
  31668=>"010001010",
  31669=>"100011100",
  31670=>"111110001",
  31671=>"010111111",
  31672=>"010001000",
  31673=>"000011000",
  31674=>"101010100",
  31675=>"011101010",
  31676=>"101000011",
  31677=>"001010001",
  31678=>"000011010",
  31679=>"111111111",
  31680=>"100100111",
  31681=>"111111111",
  31682=>"110101100",
  31683=>"110110000",
  31684=>"011111101",
  31685=>"010000000",
  31686=>"011001100",
  31687=>"100100111",
  31688=>"000101101",
  31689=>"110011100",
  31690=>"011001100",
  31691=>"111111010",
  31692=>"100100011",
  31693=>"110111010",
  31694=>"110101101",
  31695=>"001001100",
  31696=>"100110110",
  31697=>"000001101",
  31698=>"111010100",
  31699=>"111011001",
  31700=>"101111110",
  31701=>"110001000",
  31702=>"111110110",
  31703=>"010000101",
  31704=>"000100010",
  31705=>"100111010",
  31706=>"101111010",
  31707=>"001011110",
  31708=>"010010000",
  31709=>"111010101",
  31710=>"000010010",
  31711=>"111001000",
  31712=>"101111110",
  31713=>"110100100",
  31714=>"011000001",
  31715=>"010101100",
  31716=>"110111001",
  31717=>"010010100",
  31718=>"100110100",
  31719=>"110110111",
  31720=>"111100010",
  31721=>"001001110",
  31722=>"100001000",
  31723=>"100011000",
  31724=>"100000010",
  31725=>"110111110",
  31726=>"101011010",
  31727=>"001011000",
  31728=>"101000011",
  31729=>"000101000",
  31730=>"010000110",
  31731=>"100110101",
  31732=>"001001101",
  31733=>"000010111",
  31734=>"001000000",
  31735=>"000110111",
  31736=>"011010111",
  31737=>"111101101",
  31738=>"110111100",
  31739=>"010001001",
  31740=>"010010101",
  31741=>"010111100",
  31742=>"001101110",
  31743=>"010100101",
  31744=>"010101111",
  31745=>"110110100",
  31746=>"011011101",
  31747=>"001001011",
  31748=>"111010100",
  31749=>"110000111",
  31750=>"010010010",
  31751=>"011000100",
  31752=>"000010110",
  31753=>"110101100",
  31754=>"010111011",
  31755=>"010000100",
  31756=>"100000000",
  31757=>"101000100",
  31758=>"000010100",
  31759=>"011111100",
  31760=>"100000111",
  31761=>"011100001",
  31762=>"101101011",
  31763=>"001001111",
  31764=>"011100101",
  31765=>"100110011",
  31766=>"000100111",
  31767=>"010011111",
  31768=>"011100000",
  31769=>"001011110",
  31770=>"000011011",
  31771=>"111100001",
  31772=>"001010010",
  31773=>"111100000",
  31774=>"100100110",
  31775=>"110000000",
  31776=>"111100000",
  31777=>"001101111",
  31778=>"101110101",
  31779=>"001000011",
  31780=>"010111101",
  31781=>"101001110",
  31782=>"011001001",
  31783=>"011101001",
  31784=>"010010100",
  31785=>"110100111",
  31786=>"011010010",
  31787=>"111100100",
  31788=>"110000000",
  31789=>"111000100",
  31790=>"010100010",
  31791=>"000001110",
  31792=>"100010100",
  31793=>"011100111",
  31794=>"101111100",
  31795=>"110101000",
  31796=>"101100101",
  31797=>"111001110",
  31798=>"110100000",
  31799=>"010111110",
  31800=>"100111000",
  31801=>"101010111",
  31802=>"101010101",
  31803=>"110110001",
  31804=>"000001000",
  31805=>"110110111",
  31806=>"011110000",
  31807=>"011010011",
  31808=>"011101100",
  31809=>"010000011",
  31810=>"011110100",
  31811=>"000110011",
  31812=>"001111101",
  31813=>"001101001",
  31814=>"101001011",
  31815=>"101010001",
  31816=>"100100001",
  31817=>"001101111",
  31818=>"110001100",
  31819=>"011001011",
  31820=>"101000001",
  31821=>"010001100",
  31822=>"100111110",
  31823=>"000011100",
  31824=>"000100011",
  31825=>"111111000",
  31826=>"011100101",
  31827=>"011000101",
  31828=>"100010011",
  31829=>"001101111",
  31830=>"111011001",
  31831=>"111110101",
  31832=>"001011100",
  31833=>"100011001",
  31834=>"111111110",
  31835=>"000011111",
  31836=>"010110010",
  31837=>"101010010",
  31838=>"110110000",
  31839=>"111000001",
  31840=>"000101111",
  31841=>"110011011",
  31842=>"111101110",
  31843=>"100111001",
  31844=>"110001101",
  31845=>"110001110",
  31846=>"100100101",
  31847=>"100101011",
  31848=>"101110010",
  31849=>"010101101",
  31850=>"100100000",
  31851=>"111101101",
  31852=>"100001111",
  31853=>"001000000",
  31854=>"101010110",
  31855=>"101000001",
  31856=>"100000111",
  31857=>"001001011",
  31858=>"110000110",
  31859=>"011111100",
  31860=>"111111011",
  31861=>"100001100",
  31862=>"111011110",
  31863=>"001101011",
  31864=>"010011001",
  31865=>"010000111",
  31866=>"101111100",
  31867=>"011001100",
  31868=>"111010111",
  31869=>"110101000",
  31870=>"011011100",
  31871=>"011111010",
  31872=>"010011110",
  31873=>"010101001",
  31874=>"011001110",
  31875=>"111011010",
  31876=>"000011000",
  31877=>"000110100",
  31878=>"000011010",
  31879=>"000111110",
  31880=>"100010111",
  31881=>"100010011",
  31882=>"001101001",
  31883=>"001101000",
  31884=>"010000011",
  31885=>"111000111",
  31886=>"100000001",
  31887=>"001111100",
  31888=>"011000111",
  31889=>"000100111",
  31890=>"011110100",
  31891=>"010110111",
  31892=>"011100111",
  31893=>"111100011",
  31894=>"100010001",
  31895=>"011101001",
  31896=>"011101010",
  31897=>"000011010",
  31898=>"111011001",
  31899=>"010100011",
  31900=>"110100100",
  31901=>"010100000",
  31902=>"110110110",
  31903=>"101000011",
  31904=>"100101000",
  31905=>"111111001",
  31906=>"000010010",
  31907=>"001011010",
  31908=>"011000110",
  31909=>"101001001",
  31910=>"000101001",
  31911=>"000000000",
  31912=>"100100000",
  31913=>"001111100",
  31914=>"000101011",
  31915=>"010011111",
  31916=>"111000001",
  31917=>"101010111",
  31918=>"010000111",
  31919=>"100001000",
  31920=>"000011101",
  31921=>"100010000",
  31922=>"110010010",
  31923=>"000011101",
  31924=>"011010101",
  31925=>"111001110",
  31926=>"110100010",
  31927=>"010100111",
  31928=>"100010101",
  31929=>"010000111",
  31930=>"100110000",
  31931=>"011011011",
  31932=>"001111011",
  31933=>"000111010",
  31934=>"011000010",
  31935=>"101001000",
  31936=>"100110100",
  31937=>"001001110",
  31938=>"010010101",
  31939=>"101100001",
  31940=>"010101110",
  31941=>"001111100",
  31942=>"000101100",
  31943=>"100001110",
  31944=>"001001001",
  31945=>"111111110",
  31946=>"100110101",
  31947=>"110101100",
  31948=>"000100010",
  31949=>"011001100",
  31950=>"011110011",
  31951=>"001100001",
  31952=>"011000011",
  31953=>"101001110",
  31954=>"100110111",
  31955=>"011001011",
  31956=>"110010010",
  31957=>"100011110",
  31958=>"101001001",
  31959=>"110000001",
  31960=>"101001011",
  31961=>"000111001",
  31962=>"110111110",
  31963=>"000101000",
  31964=>"010111000",
  31965=>"011010001",
  31966=>"001100100",
  31967=>"101111011",
  31968=>"110111011",
  31969=>"101000010",
  31970=>"010101110",
  31971=>"111000001",
  31972=>"010101111",
  31973=>"111000111",
  31974=>"111000100",
  31975=>"011111111",
  31976=>"111111001",
  31977=>"111110011",
  31978=>"000111011",
  31979=>"011011111",
  31980=>"110010001",
  31981=>"110000101",
  31982=>"000000111",
  31983=>"000010100",
  31984=>"001001101",
  31985=>"110101000",
  31986=>"010000011",
  31987=>"100010101",
  31988=>"010010000",
  31989=>"010000000",
  31990=>"000001011",
  31991=>"100000111",
  31992=>"000101011",
  31993=>"101000010",
  31994=>"011100111",
  31995=>"100010001",
  31996=>"001101100",
  31997=>"101011010",
  31998=>"111010011",
  31999=>"100001001",
  32000=>"011010001",
  32001=>"100110111",
  32002=>"101001110",
  32003=>"111110001",
  32004=>"100110110",
  32005=>"111101011",
  32006=>"011010101",
  32007=>"111111101",
  32008=>"001110010",
  32009=>"011011101",
  32010=>"110000001",
  32011=>"010000110",
  32012=>"011101111",
  32013=>"010010111",
  32014=>"111101001",
  32015=>"011000111",
  32016=>"101001110",
  32017=>"100100000",
  32018=>"000100010",
  32019=>"100100101",
  32020=>"100101011",
  32021=>"001101010",
  32022=>"000111011",
  32023=>"001110010",
  32024=>"101011100",
  32025=>"101010111",
  32026=>"110001011",
  32027=>"000111010",
  32028=>"110010010",
  32029=>"001001011",
  32030=>"001111000",
  32031=>"100101011",
  32032=>"100010011",
  32033=>"101101011",
  32034=>"110111110",
  32035=>"100010000",
  32036=>"001111010",
  32037=>"001011101",
  32038=>"000011001",
  32039=>"010110010",
  32040=>"000010001",
  32041=>"110100010",
  32042=>"110000111",
  32043=>"001110101",
  32044=>"000000010",
  32045=>"111110000",
  32046=>"100100100",
  32047=>"100111111",
  32048=>"111111011",
  32049=>"010011010",
  32050=>"100010000",
  32051=>"100110011",
  32052=>"111111111",
  32053=>"111111000",
  32054=>"100100100",
  32055=>"011101100",
  32056=>"111101111",
  32057=>"110000101",
  32058=>"010111111",
  32059=>"100001000",
  32060=>"001010000",
  32061=>"111100111",
  32062=>"010101110",
  32063=>"111000000",
  32064=>"111011101",
  32065=>"111101011",
  32066=>"010000111",
  32067=>"000101000",
  32068=>"010111100",
  32069=>"000011110",
  32070=>"000111000",
  32071=>"110110111",
  32072=>"100101000",
  32073=>"110101100",
  32074=>"100110010",
  32075=>"111011001",
  32076=>"000100110",
  32077=>"010011101",
  32078=>"000010100",
  32079=>"110001011",
  32080=>"011101000",
  32081=>"001100000",
  32082=>"100011001",
  32083=>"101100101",
  32084=>"110100110",
  32085=>"001010111",
  32086=>"000110111",
  32087=>"011100101",
  32088=>"010100000",
  32089=>"100010110",
  32090=>"000111101",
  32091=>"100001000",
  32092=>"110101100",
  32093=>"001010111",
  32094=>"100111110",
  32095=>"110100101",
  32096=>"101000001",
  32097=>"010011111",
  32098=>"110011000",
  32099=>"100010111",
  32100=>"101100111",
  32101=>"110010011",
  32102=>"100010010",
  32103=>"010000110",
  32104=>"010001001",
  32105=>"011000011",
  32106=>"011100100",
  32107=>"001100100",
  32108=>"111010011",
  32109=>"010011000",
  32110=>"010000011",
  32111=>"100011111",
  32112=>"010101111",
  32113=>"110100000",
  32114=>"111100010",
  32115=>"100110010",
  32116=>"111101101",
  32117=>"110101100",
  32118=>"101100010",
  32119=>"011100111",
  32120=>"011001101",
  32121=>"011110000",
  32122=>"111101011",
  32123=>"111100111",
  32124=>"100101101",
  32125=>"111001011",
  32126=>"101100110",
  32127=>"101101010",
  32128=>"110011010",
  32129=>"110010100",
  32130=>"110010100",
  32131=>"110111010",
  32132=>"111001010",
  32133=>"100000001",
  32134=>"100011000",
  32135=>"001001110",
  32136=>"111111011",
  32137=>"000000010",
  32138=>"010011001",
  32139=>"110100101",
  32140=>"000011000",
  32141=>"101101011",
  32142=>"101101111",
  32143=>"110011111",
  32144=>"101110111",
  32145=>"111001001",
  32146=>"001010110",
  32147=>"111100101",
  32148=>"101110000",
  32149=>"101100111",
  32150=>"101100101",
  32151=>"011011101",
  32152=>"101000001",
  32153=>"010001100",
  32154=>"000000101",
  32155=>"101100000",
  32156=>"110001100",
  32157=>"101011000",
  32158=>"111001010",
  32159=>"001100100",
  32160=>"100001100",
  32161=>"111000101",
  32162=>"111111001",
  32163=>"001111011",
  32164=>"111101100",
  32165=>"101000100",
  32166=>"100010000",
  32167=>"100101011",
  32168=>"000001011",
  32169=>"011100111",
  32170=>"110111111",
  32171=>"000010110",
  32172=>"110001111",
  32173=>"110100110",
  32174=>"000001110",
  32175=>"100010010",
  32176=>"010110000",
  32177=>"100111110",
  32178=>"011000111",
  32179=>"101100011",
  32180=>"000010110",
  32181=>"000101011",
  32182=>"101011011",
  32183=>"011011011",
  32184=>"111111100",
  32185=>"011000111",
  32186=>"111110110",
  32187=>"001110000",
  32188=>"101100111",
  32189=>"101001010",
  32190=>"111111010",
  32191=>"101111101",
  32192=>"111000100",
  32193=>"010101001",
  32194=>"111011110",
  32195=>"000010110",
  32196=>"011100101",
  32197=>"110100001",
  32198=>"001101011",
  32199=>"011111000",
  32200=>"010101010",
  32201=>"001001110",
  32202=>"111101110",
  32203=>"010000111",
  32204=>"111101100",
  32205=>"001101111",
  32206=>"001011101",
  32207=>"001111111",
  32208=>"000110110",
  32209=>"000000110",
  32210=>"001011111",
  32211=>"000110100",
  32212=>"011001000",
  32213=>"111000100",
  32214=>"001101001",
  32215=>"100100000",
  32216=>"010010011",
  32217=>"110100100",
  32218=>"000010001",
  32219=>"101100000",
  32220=>"000001011",
  32221=>"111101011",
  32222=>"100110001",
  32223=>"101110110",
  32224=>"100011010",
  32225=>"011111110",
  32226=>"010001110",
  32227=>"110000000",
  32228=>"011111111",
  32229=>"010110111",
  32230=>"111110010",
  32231=>"110111101",
  32232=>"110100100",
  32233=>"010101011",
  32234=>"101011011",
  32235=>"010100010",
  32236=>"001000111",
  32237=>"111011110",
  32238=>"101000001",
  32239=>"110000000",
  32240=>"000011010",
  32241=>"101110100",
  32242=>"011100000",
  32243=>"010000000",
  32244=>"110010110",
  32245=>"100010000",
  32246=>"000111110",
  32247=>"000000000",
  32248=>"101000111",
  32249=>"110001000",
  32250=>"000010100",
  32251=>"001001011",
  32252=>"100111100",
  32253=>"000110010",
  32254=>"010111000",
  32255=>"001011001",
  32256=>"000111110",
  32257=>"000001111",
  32258=>"000011110",
  32259=>"100101111",
  32260=>"011000010",
  32261=>"000011111",
  32262=>"110000101",
  32263=>"001100001",
  32264=>"110101111",
  32265=>"100010001",
  32266=>"110001100",
  32267=>"000111011",
  32268=>"010100000",
  32269=>"010000111",
  32270=>"000000111",
  32271=>"001000101",
  32272=>"000110001",
  32273=>"101000000",
  32274=>"110101000",
  32275=>"100101110",
  32276=>"111001110",
  32277=>"000110000",
  32278=>"111011101",
  32279=>"011111100",
  32280=>"010010100",
  32281=>"100000100",
  32282=>"110000001",
  32283=>"111011001",
  32284=>"000111010",
  32285=>"001000101",
  32286=>"111100110",
  32287=>"011100011",
  32288=>"111011110",
  32289=>"001010011",
  32290=>"100101111",
  32291=>"110010011",
  32292=>"010101111",
  32293=>"110001000",
  32294=>"001001001",
  32295=>"000100101",
  32296=>"110101010",
  32297=>"101001011",
  32298=>"100110000",
  32299=>"101000001",
  32300=>"110010011",
  32301=>"010110101",
  32302=>"111001000",
  32303=>"101001000",
  32304=>"001011101",
  32305=>"100111001",
  32306=>"000110000",
  32307=>"110100111",
  32308=>"100000011",
  32309=>"000001010",
  32310=>"001110011",
  32311=>"010101111",
  32312=>"001001011",
  32313=>"111101001",
  32314=>"100000100",
  32315=>"010010111",
  32316=>"001001011",
  32317=>"101101100",
  32318=>"010100100",
  32319=>"000010111",
  32320=>"001011101",
  32321=>"100111000",
  32322=>"000110000",
  32323=>"010100000",
  32324=>"000011010",
  32325=>"001000110",
  32326=>"010111111",
  32327=>"010000100",
  32328=>"111010000",
  32329=>"000100111",
  32330=>"001111101",
  32331=>"000111101",
  32332=>"100010101",
  32333=>"110110001",
  32334=>"111001101",
  32335=>"101010001",
  32336=>"010111000",
  32337=>"010010000",
  32338=>"000001100",
  32339=>"001011010",
  32340=>"111000110",
  32341=>"100001100",
  32342=>"000111011",
  32343=>"000100001",
  32344=>"100100011",
  32345=>"101100011",
  32346=>"000101011",
  32347=>"000100001",
  32348=>"100000000",
  32349=>"101001100",
  32350=>"000000001",
  32351=>"110010101",
  32352=>"101000101",
  32353=>"000000111",
  32354=>"000110101",
  32355=>"010011111",
  32356=>"110010010",
  32357=>"011110111",
  32358=>"010100001",
  32359=>"011010101",
  32360=>"100110110",
  32361=>"101111001",
  32362=>"001101111",
  32363=>"111111111",
  32364=>"000000001",
  32365=>"111110010",
  32366=>"001011001",
  32367=>"000000111",
  32368=>"111010000",
  32369=>"011011000",
  32370=>"101001110",
  32371=>"101011000",
  32372=>"111110000",
  32373=>"000110101",
  32374=>"101111101",
  32375=>"001111000",
  32376=>"011001001",
  32377=>"010110110",
  32378=>"000101111",
  32379=>"110001101",
  32380=>"011011110",
  32381=>"101111001",
  32382=>"111110110",
  32383=>"011001010",
  32384=>"100100001",
  32385=>"000110001",
  32386=>"111001101",
  32387=>"111110000",
  32388=>"110011110",
  32389=>"101101101",
  32390=>"000111111",
  32391=>"000001111",
  32392=>"001001001",
  32393=>"110110110",
  32394=>"111100101",
  32395=>"111110101",
  32396=>"100001111",
  32397=>"011000011",
  32398=>"000101001",
  32399=>"111001000",
  32400=>"000001010",
  32401=>"010001011",
  32402=>"101110001",
  32403=>"111011000",
  32404=>"001010010",
  32405=>"100101011",
  32406=>"011111110",
  32407=>"010001100",
  32408=>"000101010",
  32409=>"000110111",
  32410=>"001101011",
  32411=>"110111111",
  32412=>"000100010",
  32413=>"101111000",
  32414=>"101000110",
  32415=>"001101010",
  32416=>"001000010",
  32417=>"010001011",
  32418=>"101100000",
  32419=>"000011011",
  32420=>"110111000",
  32421=>"111101010",
  32422=>"000111100",
  32423=>"110101010",
  32424=>"000111001",
  32425=>"000011111",
  32426=>"100001011",
  32427=>"001011000",
  32428=>"010001101",
  32429=>"110111011",
  32430=>"110110110",
  32431=>"001101101",
  32432=>"101010000",
  32433=>"111110110",
  32434=>"010100011",
  32435=>"011000010",
  32436=>"111100110",
  32437=>"011110101",
  32438=>"000010111",
  32439=>"110111110",
  32440=>"000111011",
  32441=>"100000110",
  32442=>"100101110",
  32443=>"101010101",
  32444=>"000011011",
  32445=>"011100110",
  32446=>"110000100",
  32447=>"010100000",
  32448=>"100111000",
  32449=>"010001000",
  32450=>"101000000",
  32451=>"100010000",
  32452=>"010010100",
  32453=>"001110010",
  32454=>"000101100",
  32455=>"001111100",
  32456=>"011100011",
  32457=>"010101001",
  32458=>"110011010",
  32459=>"111010000",
  32460=>"111001100",
  32461=>"101000000",
  32462=>"011110110",
  32463=>"001010001",
  32464=>"011000110",
  32465=>"111011000",
  32466=>"111101001",
  32467=>"101101110",
  32468=>"100001111",
  32469=>"011000101",
  32470=>"111011000",
  32471=>"001010111",
  32472=>"110011100",
  32473=>"000111100",
  32474=>"111111101",
  32475=>"000110011",
  32476=>"111101001",
  32477=>"001010000",
  32478=>"110000100",
  32479=>"101111111",
  32480=>"101001001",
  32481=>"111010010",
  32482=>"110111110",
  32483=>"100110000",
  32484=>"011000000",
  32485=>"011101000",
  32486=>"100110010",
  32487=>"000101010",
  32488=>"101111110",
  32489=>"111001000",
  32490=>"000000101",
  32491=>"101001001",
  32492=>"100010111",
  32493=>"001110001",
  32494=>"011000110",
  32495=>"011101011",
  32496=>"000111100",
  32497=>"110110111",
  32498=>"100111100",
  32499=>"010110011",
  32500=>"110011001",
  32501=>"111001101",
  32502=>"110001111",
  32503=>"101110101",
  32504=>"100001111",
  32505=>"101000011",
  32506=>"010101011",
  32507=>"111100101",
  32508=>"000011110",
  32509=>"001101001",
  32510=>"110001000",
  32511=>"111101001",
  32512=>"010000001",
  32513=>"101101011",
  32514=>"011001101",
  32515=>"001001000",
  32516=>"000001110",
  32517=>"101001001",
  32518=>"111100111",
  32519=>"001000110",
  32520=>"110110101",
  32521=>"001101111",
  32522=>"100011100",
  32523=>"011000110",
  32524=>"000100111",
  32525=>"001010001",
  32526=>"000001010",
  32527=>"001001111",
  32528=>"001010110",
  32529=>"101100110",
  32530=>"110100101",
  32531=>"110101000",
  32532=>"111110000",
  32533=>"101001000",
  32534=>"010110000",
  32535=>"011000000",
  32536=>"101111110",
  32537=>"010000001",
  32538=>"110101010",
  32539=>"110000100",
  32540=>"100010001",
  32541=>"110101111",
  32542=>"110100111",
  32543=>"110011110",
  32544=>"101100110",
  32545=>"110111100",
  32546=>"011011000",
  32547=>"111010000",
  32548=>"010001100",
  32549=>"101101000",
  32550=>"001010101",
  32551=>"010010111",
  32552=>"001101110",
  32553=>"001111111",
  32554=>"110111111",
  32555=>"000101101",
  32556=>"011101111",
  32557=>"111001111",
  32558=>"110000110",
  32559=>"110011111",
  32560=>"101000011",
  32561=>"011111011",
  32562=>"111101001",
  32563=>"100101101",
  32564=>"010000010",
  32565=>"100011111",
  32566=>"110011010",
  32567=>"101111001",
  32568=>"000100100",
  32569=>"100111111",
  32570=>"000001000",
  32571=>"100011111",
  32572=>"111011010",
  32573=>"100111100",
  32574=>"000101001",
  32575=>"000000100",
  32576=>"000000100",
  32577=>"111110000",
  32578=>"010001100",
  32579=>"010010101",
  32580=>"101110010",
  32581=>"000100110",
  32582=>"000010100",
  32583=>"110000100",
  32584=>"000011100",
  32585=>"010001111",
  32586=>"111001010",
  32587=>"010101110",
  32588=>"011010111",
  32589=>"110111010",
  32590=>"000100011",
  32591=>"100010001",
  32592=>"101000101",
  32593=>"111001100",
  32594=>"101110000",
  32595=>"000110111",
  32596=>"001010101",
  32597=>"111110000",
  32598=>"100100100",
  32599=>"001101101",
  32600=>"011100100",
  32601=>"011000011",
  32602=>"100010101",
  32603=>"011111101",
  32604=>"000001001",
  32605=>"001100001",
  32606=>"010100000",
  32607=>"110111110",
  32608=>"110001010",
  32609=>"010100100",
  32610=>"111001111",
  32611=>"101011101",
  32612=>"000000101",
  32613=>"101000000",
  32614=>"000110000",
  32615=>"011101010",
  32616=>"100000001",
  32617=>"010100000",
  32618=>"110110101",
  32619=>"000000111",
  32620=>"010001110",
  32621=>"000111011",
  32622=>"001110111",
  32623=>"010000010",
  32624=>"110010010",
  32625=>"011100010",
  32626=>"110000001",
  32627=>"100101001",
  32628=>"000110111",
  32629=>"110000100",
  32630=>"000100100",
  32631=>"101111011",
  32632=>"100001100",
  32633=>"101001110",
  32634=>"011111001",
  32635=>"010100110",
  32636=>"000101110",
  32637=>"000100001",
  32638=>"110110100",
  32639=>"000001011",
  32640=>"001011000",
  32641=>"100001011",
  32642=>"110011101",
  32643=>"101000100",
  32644=>"001110001",
  32645=>"011110001",
  32646=>"010100100",
  32647=>"000010111",
  32648=>"011111010",
  32649=>"000000000",
  32650=>"111010001",
  32651=>"001000111",
  32652=>"010100001",
  32653=>"111000100",
  32654=>"010011111",
  32655=>"110001001",
  32656=>"111100000",
  32657=>"001101010",
  32658=>"000011111",
  32659=>"010011001",
  32660=>"101010010",
  32661=>"101110001",
  32662=>"111011010",
  32663=>"000110100",
  32664=>"101001011",
  32665=>"011110110",
  32666=>"100000011",
  32667=>"111111111",
  32668=>"100001000",
  32669=>"110010110",
  32670=>"001110011",
  32671=>"010001111",
  32672=>"101101100",
  32673=>"000000000",
  32674=>"110101000",
  32675=>"110010001",
  32676=>"111011111",
  32677=>"010010110",
  32678=>"010110101",
  32679=>"001100100",
  32680=>"011100111",
  32681=>"101001101",
  32682=>"000101111",
  32683=>"110010010",
  32684=>"111101001",
  32685=>"000000001",
  32686=>"111110100",
  32687=>"001010101",
  32688=>"111000111",
  32689=>"101001111",
  32690=>"001010010",
  32691=>"111100011",
  32692=>"001010100",
  32693=>"110101010",
  32694=>"011010111",
  32695=>"001011011",
  32696=>"011101111",
  32697=>"010001001",
  32698=>"000010011",
  32699=>"111100010",
  32700=>"000100110",
  32701=>"111001101",
  32702=>"100100010",
  32703=>"001110100",
  32704=>"101011100",
  32705=>"110010100",
  32706=>"000000000",
  32707=>"000001101",
  32708=>"001001011",
  32709=>"111111000",
  32710=>"110101111",
  32711=>"001110110",
  32712=>"100011011",
  32713=>"110101111",
  32714=>"010101100",
  32715=>"110111110",
  32716=>"011010101",
  32717=>"101001101",
  32718=>"010100101",
  32719=>"111011110",
  32720=>"000110011",
  32721=>"101010101",
  32722=>"011011111",
  32723=>"111111111",
  32724=>"010101000",
  32725=>"111010110",
  32726=>"010011101",
  32727=>"110010111",
  32728=>"111111111",
  32729=>"011100011",
  32730=>"010101001",
  32731=>"010100101",
  32732=>"000100101",
  32733=>"000001011",
  32734=>"000000101",
  32735=>"111001111",
  32736=>"111011110",
  32737=>"110010110",
  32738=>"001010101",
  32739=>"100011100",
  32740=>"101100000",
  32741=>"001110111",
  32742=>"110000110",
  32743=>"111001000",
  32744=>"110110001",
  32745=>"100110011",
  32746=>"001100100",
  32747=>"000100111",
  32748=>"011011100",
  32749=>"001011111",
  32750=>"010001001",
  32751=>"001100100",
  32752=>"000001001",
  32753=>"111100111",
  32754=>"101101100",
  32755=>"010000110",
  32756=>"011011100",
  32757=>"100100011",
  32758=>"001011001",
  32759=>"111000101",
  32760=>"010110010",
  32761=>"110001010",
  32762=>"110101110",
  32763=>"000100110",
  32764=>"011101111",
  32765=>"111000001",
  32766=>"011001000",
  32767=>"111001000",
  32768=>"111110011",
  32769=>"101001011",
  32770=>"001001100",
  32771=>"111100010",
  32772=>"100100001",
  32773=>"010010001",
  32774=>"101100111",
  32775=>"101010110",
  32776=>"001000000",
  32777=>"111000000",
  32778=>"111110000",
  32779=>"011011011",
  32780=>"100101110",
  32781=>"000100110",
  32782=>"100001101",
  32783=>"001010110",
  32784=>"100100001",
  32785=>"101101101",
  32786=>"111101101",
  32787=>"100010000",
  32788=>"000000000",
  32789=>"100010110",
  32790=>"101111001",
  32791=>"000101110",
  32792=>"111101011",
  32793=>"010110000",
  32794=>"111001011",
  32795=>"010001000",
  32796=>"101111100",
  32797=>"101000001",
  32798=>"010100111",
  32799=>"101111100",
  32800=>"001001000",
  32801=>"011011101",
  32802=>"001111101",
  32803=>"110010100",
  32804=>"100110011",
  32805=>"110111010",
  32806=>"100010000",
  32807=>"110111000",
  32808=>"010010001",
  32809=>"101101001",
  32810=>"101111100",
  32811=>"100011011",
  32812=>"000000100",
  32813=>"110100111",
  32814=>"111100101",
  32815=>"111100011",
  32816=>"001101111",
  32817=>"110010010",
  32818=>"111111001",
  32819=>"110010000",
  32820=>"110101111",
  32821=>"000110011",
  32822=>"010101110",
  32823=>"000000111",
  32824=>"000011101",
  32825=>"111110111",
  32826=>"001101100",
  32827=>"011100010",
  32828=>"101110100",
  32829=>"001000111",
  32830=>"111111011",
  32831=>"000100010",
  32832=>"010110000",
  32833=>"011111111",
  32834=>"110111000",
  32835=>"010111101",
  32836=>"111011010",
  32837=>"001001100",
  32838=>"010111101",
  32839=>"110001001",
  32840=>"110001101",
  32841=>"110101010",
  32842=>"000101010",
  32843=>"010111001",
  32844=>"100111101",
  32845=>"101110101",
  32846=>"010110010",
  32847=>"110010001",
  32848=>"110001010",
  32849=>"000100001",
  32850=>"000001100",
  32851=>"000011000",
  32852=>"101101000",
  32853=>"111010000",
  32854=>"001000000",
  32855=>"010001000",
  32856=>"010101001",
  32857=>"010000000",
  32858=>"110111000",
  32859=>"100001101",
  32860=>"000110110",
  32861=>"101010000",
  32862=>"000001110",
  32863=>"101101101",
  32864=>"110010010",
  32865=>"100111010",
  32866=>"011001000",
  32867=>"100100001",
  32868=>"111110101",
  32869=>"111110101",
  32870=>"000000101",
  32871=>"101111100",
  32872=>"100001011",
  32873=>"111011011",
  32874=>"011010100",
  32875=>"000101011",
  32876=>"111010010",
  32877=>"101001000",
  32878=>"101110000",
  32879=>"111101111",
  32880=>"001101000",
  32881=>"001111000",
  32882=>"011110110",
  32883=>"000101101",
  32884=>"000010111",
  32885=>"111000110",
  32886=>"011100001",
  32887=>"101000110",
  32888=>"101101001",
  32889=>"101110000",
  32890=>"000100000",
  32891=>"101100000",
  32892=>"011001110",
  32893=>"001010100",
  32894=>"111000111",
  32895=>"000111010",
  32896=>"001111110",
  32897=>"010100001",
  32898=>"000101000",
  32899=>"000011000",
  32900=>"110011111",
  32901=>"111011110",
  32902=>"100011000",
  32903=>"101001001",
  32904=>"011100010",
  32905=>"000100100",
  32906=>"000000000",
  32907=>"000110100",
  32908=>"011000110",
  32909=>"110001010",
  32910=>"101001101",
  32911=>"111111001",
  32912=>"111100010",
  32913=>"011110110",
  32914=>"100010010",
  32915=>"100111010",
  32916=>"101111110",
  32917=>"111011001",
  32918=>"100000010",
  32919=>"001011010",
  32920=>"000010111",
  32921=>"111000001",
  32922=>"100101111",
  32923=>"100100011",
  32924=>"010000111",
  32925=>"010111011",
  32926=>"011100000",
  32927=>"010011011",
  32928=>"110010111",
  32929=>"010100111",
  32930=>"100111110",
  32931=>"110100111",
  32932=>"100100100",
  32933=>"000100101",
  32934=>"000110010",
  32935=>"000001110",
  32936=>"111010000",
  32937=>"001011101",
  32938=>"100011110",
  32939=>"101101100",
  32940=>"110000111",
  32941=>"110001100",
  32942=>"000010000",
  32943=>"000100100",
  32944=>"100111001",
  32945=>"110000010",
  32946=>"000101001",
  32947=>"000100010",
  32948=>"110100010",
  32949=>"100001001",
  32950=>"101111010",
  32951=>"011011110",
  32952=>"110010111",
  32953=>"001100100",
  32954=>"101111101",
  32955=>"111110110",
  32956=>"001110111",
  32957=>"111101101",
  32958=>"101011101",
  32959=>"010011001",
  32960=>"000110111",
  32961=>"110000000",
  32962=>"001110011",
  32963=>"110000100",
  32964=>"010100110",
  32965=>"001100111",
  32966=>"110111001",
  32967=>"011011010",
  32968=>"110100110",
  32969=>"001101110",
  32970=>"010100000",
  32971=>"001001101",
  32972=>"011110010",
  32973=>"010000101",
  32974=>"110000011",
  32975=>"110100101",
  32976=>"011011111",
  32977=>"000101001",
  32978=>"100111101",
  32979=>"111110101",
  32980=>"000000000",
  32981=>"011010101",
  32982=>"000111111",
  32983=>"010010011",
  32984=>"000110111",
  32985=>"010011000",
  32986=>"000111000",
  32987=>"000011110",
  32988=>"001010010",
  32989=>"110010011",
  32990=>"010101010",
  32991=>"110110111",
  32992=>"001000110",
  32993=>"001111000",
  32994=>"101000100",
  32995=>"100111000",
  32996=>"011100011",
  32997=>"000001011",
  32998=>"100110100",
  32999=>"010000010",
  33000=>"100010001",
  33001=>"000010011",
  33002=>"000110100",
  33003=>"111000001",
  33004=>"010110010",
  33005=>"000010100",
  33006=>"110001011",
  33007=>"010001001",
  33008=>"101001011",
  33009=>"100000001",
  33010=>"001010010",
  33011=>"000011111",
  33012=>"000111101",
  33013=>"111000100",
  33014=>"000000110",
  33015=>"100110101",
  33016=>"000001110",
  33017=>"101111110",
  33018=>"111001011",
  33019=>"000101101",
  33020=>"000011000",
  33021=>"000101001",
  33022=>"111000100",
  33023=>"010111101",
  33024=>"110101101",
  33025=>"010000011",
  33026=>"011010110",
  33027=>"001001100",
  33028=>"010000101",
  33029=>"100001011",
  33030=>"000000010",
  33031=>"000110001",
  33032=>"011011100",
  33033=>"111100101",
  33034=>"010001110",
  33035=>"111001111",
  33036=>"101010101",
  33037=>"101001111",
  33038=>"011111011",
  33039=>"011100110",
  33040=>"010101111",
  33041=>"001001100",
  33042=>"100110111",
  33043=>"101100101",
  33044=>"110110011",
  33045=>"111010000",
  33046=>"111011101",
  33047=>"100111101",
  33048=>"010100100",
  33049=>"010000010",
  33050=>"010110000",
  33051=>"111000111",
  33052=>"010000110",
  33053=>"111010011",
  33054=>"111011111",
  33055=>"011111011",
  33056=>"001100000",
  33057=>"010001000",
  33058=>"100110111",
  33059=>"111110010",
  33060=>"111101100",
  33061=>"101010110",
  33062=>"111111000",
  33063=>"100011011",
  33064=>"111101001",
  33065=>"101001000",
  33066=>"110001001",
  33067=>"000011011",
  33068=>"000001011",
  33069=>"101000010",
  33070=>"101000110",
  33071=>"011000000",
  33072=>"101100101",
  33073=>"011100100",
  33074=>"110110111",
  33075=>"001000011",
  33076=>"011110100",
  33077=>"111000100",
  33078=>"011000010",
  33079=>"100011101",
  33080=>"000100001",
  33081=>"101111100",
  33082=>"101000011",
  33083=>"011111011",
  33084=>"000111110",
  33085=>"000101100",
  33086=>"011010111",
  33087=>"011011011",
  33088=>"000011001",
  33089=>"110110101",
  33090=>"111000000",
  33091=>"110011010",
  33092=>"001000001",
  33093=>"011011000",
  33094=>"101000110",
  33095=>"011011001",
  33096=>"110011000",
  33097=>"011100000",
  33098=>"101001001",
  33099=>"001110000",
  33100=>"110000011",
  33101=>"010111010",
  33102=>"000001001",
  33103=>"000001110",
  33104=>"011110000",
  33105=>"011000100",
  33106=>"001010010",
  33107=>"111001000",
  33108=>"001111101",
  33109=>"110001010",
  33110=>"000111010",
  33111=>"001110000",
  33112=>"000001011",
  33113=>"010100111",
  33114=>"101010101",
  33115=>"000001001",
  33116=>"010110010",
  33117=>"001000011",
  33118=>"111011111",
  33119=>"010001101",
  33120=>"100111100",
  33121=>"011101010",
  33122=>"001001001",
  33123=>"000110010",
  33124=>"011000001",
  33125=>"010000100",
  33126=>"110000100",
  33127=>"101010111",
  33128=>"000010011",
  33129=>"000010000",
  33130=>"110111000",
  33131=>"110100001",
  33132=>"011100011",
  33133=>"110100001",
  33134=>"111001010",
  33135=>"101000001",
  33136=>"010010011",
  33137=>"111010011",
  33138=>"000011100",
  33139=>"011111011",
  33140=>"010000001",
  33141=>"000011111",
  33142=>"010100101",
  33143=>"100110111",
  33144=>"000011110",
  33145=>"110000010",
  33146=>"110101010",
  33147=>"110110101",
  33148=>"011011001",
  33149=>"110101100",
  33150=>"010011101",
  33151=>"111111110",
  33152=>"011000101",
  33153=>"011100111",
  33154=>"000000001",
  33155=>"010100001",
  33156=>"011011110",
  33157=>"001010001",
  33158=>"101001111",
  33159=>"100111001",
  33160=>"100101100",
  33161=>"110101001",
  33162=>"011101010",
  33163=>"111011101",
  33164=>"001010100",
  33165=>"000010011",
  33166=>"001110001",
  33167=>"100110000",
  33168=>"111100100",
  33169=>"110010000",
  33170=>"001001000",
  33171=>"011100000",
  33172=>"111011100",
  33173=>"000011000",
  33174=>"000010010",
  33175=>"111111101",
  33176=>"010011101",
  33177=>"101000111",
  33178=>"111001110",
  33179=>"110110100",
  33180=>"111011111",
  33181=>"101101011",
  33182=>"101000000",
  33183=>"100110001",
  33184=>"101100001",
  33185=>"101101000",
  33186=>"111010001",
  33187=>"100000010",
  33188=>"101000110",
  33189=>"001101101",
  33190=>"011100110",
  33191=>"011100100",
  33192=>"111011101",
  33193=>"100011100",
  33194=>"101000001",
  33195=>"010000011",
  33196=>"000001001",
  33197=>"010010101",
  33198=>"000001000",
  33199=>"000111101",
  33200=>"000010011",
  33201=>"011000000",
  33202=>"001010000",
  33203=>"110001101",
  33204=>"111101111",
  33205=>"100011000",
  33206=>"000000110",
  33207=>"111111001",
  33208=>"100101101",
  33209=>"011111001",
  33210=>"001101011",
  33211=>"000010011",
  33212=>"010101010",
  33213=>"001001110",
  33214=>"011001111",
  33215=>"001100101",
  33216=>"000111111",
  33217=>"010010001",
  33218=>"011111011",
  33219=>"101010111",
  33220=>"101000111",
  33221=>"000100010",
  33222=>"101111011",
  33223=>"001010000",
  33224=>"001101001",
  33225=>"001100101",
  33226=>"011000001",
  33227=>"110010111",
  33228=>"010000000",
  33229=>"011010000",
  33230=>"111000000",
  33231=>"101001110",
  33232=>"010000100",
  33233=>"111000110",
  33234=>"001010000",
  33235=>"000100110",
  33236=>"101100001",
  33237=>"000010000",
  33238=>"010101101",
  33239=>"001011010",
  33240=>"011010011",
  33241=>"111011111",
  33242=>"000010100",
  33243=>"101111110",
  33244=>"101011011",
  33245=>"100111100",
  33246=>"100111111",
  33247=>"011101001",
  33248=>"010111101",
  33249=>"000100001",
  33250=>"111100000",
  33251=>"011111000",
  33252=>"001110000",
  33253=>"011010101",
  33254=>"001010000",
  33255=>"100011011",
  33256=>"000011110",
  33257=>"010001111",
  33258=>"011000111",
  33259=>"100101111",
  33260=>"111110011",
  33261=>"011110100",
  33262=>"100000010",
  33263=>"001110000",
  33264=>"110110001",
  33265=>"010100110",
  33266=>"001100100",
  33267=>"011110100",
  33268=>"001110000",
  33269=>"011101000",
  33270=>"110011000",
  33271=>"101100000",
  33272=>"010010100",
  33273=>"111110000",
  33274=>"011100111",
  33275=>"100101001",
  33276=>"000110010",
  33277=>"010101111",
  33278=>"101011100",
  33279=>"111101111",
  33280=>"000110110",
  33281=>"010010001",
  33282=>"010010100",
  33283=>"100000110",
  33284=>"011001100",
  33285=>"111010101",
  33286=>"010000111",
  33287=>"001000110",
  33288=>"101110001",
  33289=>"010000011",
  33290=>"100000111",
  33291=>"100011010",
  33292=>"110110110",
  33293=>"101010110",
  33294=>"010000100",
  33295=>"001111000",
  33296=>"000101110",
  33297=>"100000110",
  33298=>"001111000",
  33299=>"011000110",
  33300=>"111110010",
  33301=>"101100010",
  33302=>"001101111",
  33303=>"110010111",
  33304=>"100011010",
  33305=>"000000001",
  33306=>"011100111",
  33307=>"001100001",
  33308=>"100110101",
  33309=>"001011111",
  33310=>"010101000",
  33311=>"101100000",
  33312=>"111001001",
  33313=>"110110000",
  33314=>"111001010",
  33315=>"000010100",
  33316=>"111111110",
  33317=>"111001111",
  33318=>"111101101",
  33319=>"101011110",
  33320=>"111010111",
  33321=>"010000000",
  33322=>"011110101",
  33323=>"011010111",
  33324=>"011110001",
  33325=>"001001011",
  33326=>"011000110",
  33327=>"000011100",
  33328=>"011100110",
  33329=>"010101011",
  33330=>"100001011",
  33331=>"100001001",
  33332=>"010000111",
  33333=>"100001000",
  33334=>"001010001",
  33335=>"001101001",
  33336=>"111010010",
  33337=>"110000100",
  33338=>"000100100",
  33339=>"011001110",
  33340=>"101011011",
  33341=>"111010000",
  33342=>"101000101",
  33343=>"111101100",
  33344=>"010110111",
  33345=>"000001100",
  33346=>"001110010",
  33347=>"001111101",
  33348=>"111100000",
  33349=>"101101001",
  33350=>"010111101",
  33351=>"011111001",
  33352=>"100110100",
  33353=>"011000111",
  33354=>"000111110",
  33355=>"001000001",
  33356=>"011111101",
  33357=>"111011011",
  33358=>"000101010",
  33359=>"100111011",
  33360=>"101110111",
  33361=>"101011001",
  33362=>"001000011",
  33363=>"100010000",
  33364=>"010010100",
  33365=>"101101001",
  33366=>"001001110",
  33367=>"011001010",
  33368=>"110111101",
  33369=>"111001001",
  33370=>"101100001",
  33371=>"111000000",
  33372=>"111000000",
  33373=>"111011100",
  33374=>"001000101",
  33375=>"001000100",
  33376=>"101000011",
  33377=>"111001100",
  33378=>"100111011",
  33379=>"111110111",
  33380=>"110111011",
  33381=>"110010101",
  33382=>"001100101",
  33383=>"011111100",
  33384=>"000011101",
  33385=>"111110100",
  33386=>"000001111",
  33387=>"011100110",
  33388=>"101000100",
  33389=>"111101100",
  33390=>"101001000",
  33391=>"101101101",
  33392=>"111001101",
  33393=>"100100000",
  33394=>"000001010",
  33395=>"101100100",
  33396=>"101010010",
  33397=>"101101011",
  33398=>"011010001",
  33399=>"100011000",
  33400=>"011010111",
  33401=>"110110001",
  33402=>"111101111",
  33403=>"010101000",
  33404=>"101011000",
  33405=>"111101011",
  33406=>"101111101",
  33407=>"110000000",
  33408=>"010101101",
  33409=>"000011110",
  33410=>"110111101",
  33411=>"001001000",
  33412=>"001001100",
  33413=>"011000010",
  33414=>"000100101",
  33415=>"000101001",
  33416=>"101111110",
  33417=>"001001110",
  33418=>"111101100",
  33419=>"001110010",
  33420=>"111110010",
  33421=>"010000110",
  33422=>"100000100",
  33423=>"111001011",
  33424=>"011111100",
  33425=>"101011101",
  33426=>"110111000",
  33427=>"001111101",
  33428=>"001000011",
  33429=>"101101001",
  33430=>"100111110",
  33431=>"101011001",
  33432=>"011001100",
  33433=>"100101100",
  33434=>"000101111",
  33435=>"110001000",
  33436=>"101011010",
  33437=>"100010111",
  33438=>"000001111",
  33439=>"011111011",
  33440=>"011110000",
  33441=>"110111001",
  33442=>"111110001",
  33443=>"011101010",
  33444=>"110101110",
  33445=>"011011100",
  33446=>"001000100",
  33447=>"010111000",
  33448=>"001111010",
  33449=>"011010110",
  33450=>"011011111",
  33451=>"101111101",
  33452=>"010111001",
  33453=>"001100110",
  33454=>"101000010",
  33455=>"001000111",
  33456=>"100100011",
  33457=>"000000000",
  33458=>"010110000",
  33459=>"001011001",
  33460=>"001011101",
  33461=>"000011100",
  33462=>"101001111",
  33463=>"111010010",
  33464=>"110010101",
  33465=>"011110001",
  33466=>"000110001",
  33467=>"111111100",
  33468=>"011001000",
  33469=>"010101000",
  33470=>"011010101",
  33471=>"001111110",
  33472=>"010101000",
  33473=>"101010111",
  33474=>"110101110",
  33475=>"000110100",
  33476=>"111011011",
  33477=>"001000000",
  33478=>"100111100",
  33479=>"001100011",
  33480=>"011111111",
  33481=>"110100100",
  33482=>"000001011",
  33483=>"100001110",
  33484=>"000010111",
  33485=>"010000111",
  33486=>"011011000",
  33487=>"111110101",
  33488=>"111010010",
  33489=>"111111100",
  33490=>"101100010",
  33491=>"110001110",
  33492=>"000011011",
  33493=>"111110000",
  33494=>"000011101",
  33495=>"010010000",
  33496=>"001100101",
  33497=>"111010101",
  33498=>"011111011",
  33499=>"101000101",
  33500=>"000111100",
  33501=>"010011100",
  33502=>"010010111",
  33503=>"010110000",
  33504=>"111001000",
  33505=>"001111110",
  33506=>"010011010",
  33507=>"111111011",
  33508=>"111000001",
  33509=>"101111010",
  33510=>"001100011",
  33511=>"111101001",
  33512=>"110000010",
  33513=>"101011001",
  33514=>"010110111",
  33515=>"010101010",
  33516=>"110101001",
  33517=>"010011111",
  33518=>"010111010",
  33519=>"101000111",
  33520=>"001100100",
  33521=>"100101110",
  33522=>"101000100",
  33523=>"010100011",
  33524=>"110010010",
  33525=>"100100100",
  33526=>"100011111",
  33527=>"100100101",
  33528=>"000101100",
  33529=>"110011001",
  33530=>"001000010",
  33531=>"100001110",
  33532=>"010010110",
  33533=>"100001000",
  33534=>"010001111",
  33535=>"111111111",
  33536=>"100100000",
  33537=>"110010000",
  33538=>"101110010",
  33539=>"011110110",
  33540=>"011110010",
  33541=>"001101000",
  33542=>"011001110",
  33543=>"011011110",
  33544=>"010000100",
  33545=>"111000000",
  33546=>"100010010",
  33547=>"111111000",
  33548=>"100111010",
  33549=>"101000101",
  33550=>"111100001",
  33551=>"101011101",
  33552=>"010101010",
  33553=>"111000100",
  33554=>"111101010",
  33555=>"111000111",
  33556=>"101100011",
  33557=>"001100011",
  33558=>"011100001",
  33559=>"100000110",
  33560=>"111010011",
  33561=>"010011000",
  33562=>"100111001",
  33563=>"111110000",
  33564=>"101011010",
  33565=>"000001100",
  33566=>"011000000",
  33567=>"010101101",
  33568=>"011011101",
  33569=>"100001110",
  33570=>"011101110",
  33571=>"010001001",
  33572=>"000110011",
  33573=>"001001011",
  33574=>"011000100",
  33575=>"000001101",
  33576=>"000001110",
  33577=>"000111000",
  33578=>"011101111",
  33579=>"001111010",
  33580=>"101000011",
  33581=>"101101001",
  33582=>"101010010",
  33583=>"011010010",
  33584=>"101000010",
  33585=>"000011100",
  33586=>"001010010",
  33587=>"001010001",
  33588=>"010010000",
  33589=>"011001010",
  33590=>"000110100",
  33591=>"011111011",
  33592=>"101001111",
  33593=>"110110111",
  33594=>"010111001",
  33595=>"100101011",
  33596=>"111111001",
  33597=>"010011000",
  33598=>"100111000",
  33599=>"010101101",
  33600=>"011111110",
  33601=>"010011110",
  33602=>"110111110",
  33603=>"110011000",
  33604=>"111110001",
  33605=>"110100000",
  33606=>"111000010",
  33607=>"000111111",
  33608=>"111111110",
  33609=>"110111111",
  33610=>"000111111",
  33611=>"000000010",
  33612=>"100100001",
  33613=>"011101110",
  33614=>"111010110",
  33615=>"010110110",
  33616=>"111001111",
  33617=>"111001010",
  33618=>"000110100",
  33619=>"011101001",
  33620=>"011110111",
  33621=>"010100000",
  33622=>"010000001",
  33623=>"011011110",
  33624=>"110010110",
  33625=>"110010000",
  33626=>"100010010",
  33627=>"100001011",
  33628=>"000101101",
  33629=>"010101010",
  33630=>"110011010",
  33631=>"111001000",
  33632=>"000010000",
  33633=>"010110111",
  33634=>"110000010",
  33635=>"001010111",
  33636=>"101010100",
  33637=>"000011111",
  33638=>"000110011",
  33639=>"111111110",
  33640=>"001011011",
  33641=>"011111100",
  33642=>"000011110",
  33643=>"011011011",
  33644=>"110110001",
  33645=>"001010011",
  33646=>"000011010",
  33647=>"011111010",
  33648=>"000001100",
  33649=>"100001111",
  33650=>"111111101",
  33651=>"011111111",
  33652=>"010110100",
  33653=>"010010100",
  33654=>"111110110",
  33655=>"101111111",
  33656=>"110010010",
  33657=>"011110011",
  33658=>"110110111",
  33659=>"001110011",
  33660=>"001000101",
  33661=>"101111010",
  33662=>"011001110",
  33663=>"010000101",
  33664=>"011010011",
  33665=>"110010100",
  33666=>"110011001",
  33667=>"010001001",
  33668=>"000101001",
  33669=>"101111100",
  33670=>"110000110",
  33671=>"111000000",
  33672=>"100010000",
  33673=>"101111111",
  33674=>"111111001",
  33675=>"111110111",
  33676=>"010100001",
  33677=>"010110100",
  33678=>"111110001",
  33679=>"001001000",
  33680=>"111111110",
  33681=>"010101011",
  33682=>"111001100",
  33683=>"101111111",
  33684=>"100111000",
  33685=>"000101101",
  33686=>"100011111",
  33687=>"111000001",
  33688=>"010111111",
  33689=>"110000100",
  33690=>"101010111",
  33691=>"000011001",
  33692=>"100111101",
  33693=>"001111010",
  33694=>"110111110",
  33695=>"000111000",
  33696=>"101010101",
  33697=>"100100010",
  33698=>"100010110",
  33699=>"111010011",
  33700=>"110010101",
  33701=>"000001000",
  33702=>"111000011",
  33703=>"101010111",
  33704=>"110111101",
  33705=>"100101011",
  33706=>"001100011",
  33707=>"101111101",
  33708=>"001011111",
  33709=>"010110011",
  33710=>"110111110",
  33711=>"001100001",
  33712=>"100101001",
  33713=>"110011110",
  33714=>"010000001",
  33715=>"111001101",
  33716=>"010100000",
  33717=>"011111101",
  33718=>"111101000",
  33719=>"110101100",
  33720=>"000100010",
  33721=>"000110110",
  33722=>"011111110",
  33723=>"110001110",
  33724=>"101100000",
  33725=>"011101010",
  33726=>"010010010",
  33727=>"011011000",
  33728=>"000011100",
  33729=>"111010000",
  33730=>"111011000",
  33731=>"001101101",
  33732=>"100111111",
  33733=>"001011001",
  33734=>"101011011",
  33735=>"100010010",
  33736=>"000101110",
  33737=>"111011110",
  33738=>"100111101",
  33739=>"000010111",
  33740=>"101001100",
  33741=>"100011000",
  33742=>"000101100",
  33743=>"001000101",
  33744=>"001100000",
  33745=>"111111001",
  33746=>"000100100",
  33747=>"001111111",
  33748=>"111010001",
  33749=>"100110100",
  33750=>"001100100",
  33751=>"111001011",
  33752=>"000010001",
  33753=>"110010001",
  33754=>"011011001",
  33755=>"001111110",
  33756=>"001110111",
  33757=>"011101011",
  33758=>"101001000",
  33759=>"100000100",
  33760=>"000100100",
  33761=>"111011000",
  33762=>"000100101",
  33763=>"000100111",
  33764=>"110100111",
  33765=>"111000010",
  33766=>"000110011",
  33767=>"011100111",
  33768=>"111110010",
  33769=>"101100101",
  33770=>"101000100",
  33771=>"100000011",
  33772=>"011101111",
  33773=>"001000111",
  33774=>"000100010",
  33775=>"111001100",
  33776=>"010010011",
  33777=>"010101111",
  33778=>"011001000",
  33779=>"000000010",
  33780=>"101101101",
  33781=>"111001011",
  33782=>"111100011",
  33783=>"011011001",
  33784=>"110100010",
  33785=>"010110110",
  33786=>"101010111",
  33787=>"010111010",
  33788=>"001101000",
  33789=>"011000111",
  33790=>"001001001",
  33791=>"010111010",
  33792=>"010010100",
  33793=>"100101000",
  33794=>"011100010",
  33795=>"001100100",
  33796=>"110010011",
  33797=>"100000100",
  33798=>"111111001",
  33799=>"000011001",
  33800=>"011111010",
  33801=>"000000010",
  33802=>"010111111",
  33803=>"101111000",
  33804=>"111111001",
  33805=>"101100000",
  33806=>"111110001",
  33807=>"000001100",
  33808=>"110101000",
  33809=>"100000111",
  33810=>"010011111",
  33811=>"010100010",
  33812=>"100101011",
  33813=>"011010001",
  33814=>"110111010",
  33815=>"010101010",
  33816=>"111110001",
  33817=>"001100000",
  33818=>"111010011",
  33819=>"110010110",
  33820=>"110001001",
  33821=>"100101011",
  33822=>"111111010",
  33823=>"001001010",
  33824=>"011000000",
  33825=>"111110000",
  33826=>"100001001",
  33827=>"010011011",
  33828=>"110011101",
  33829=>"101011011",
  33830=>"110110001",
  33831=>"100011110",
  33832=>"001101000",
  33833=>"110100100",
  33834=>"110100111",
  33835=>"111010110",
  33836=>"111010000",
  33837=>"001101000",
  33838=>"001000110",
  33839=>"111001100",
  33840=>"010100110",
  33841=>"001000000",
  33842=>"101000001",
  33843=>"000101101",
  33844=>"011001010",
  33845=>"001101001",
  33846=>"101100100",
  33847=>"111111101",
  33848=>"000100100",
  33849=>"001100101",
  33850=>"001100000",
  33851=>"111100111",
  33852=>"001110010",
  33853=>"111011010",
  33854=>"101001000",
  33855=>"101010101",
  33856=>"101000001",
  33857=>"000100000",
  33858=>"011010111",
  33859=>"010000111",
  33860=>"001100110",
  33861=>"001010010",
  33862=>"110001000",
  33863=>"000100101",
  33864=>"110000101",
  33865=>"111001011",
  33866=>"101000000",
  33867=>"101001001",
  33868=>"010000011",
  33869=>"011010001",
  33870=>"011000000",
  33871=>"110000001",
  33872=>"111110010",
  33873=>"111010000",
  33874=>"001011100",
  33875=>"100101110",
  33876=>"110110010",
  33877=>"111101111",
  33878=>"001000000",
  33879=>"010101101",
  33880=>"011000101",
  33881=>"010101110",
  33882=>"000110100",
  33883=>"111110100",
  33884=>"010110011",
  33885=>"100011011",
  33886=>"000100011",
  33887=>"000010111",
  33888=>"000101000",
  33889=>"000111000",
  33890=>"110011101",
  33891=>"110010010",
  33892=>"111001101",
  33893=>"100001000",
  33894=>"101001100",
  33895=>"101001101",
  33896=>"110000011",
  33897=>"000100011",
  33898=>"001100000",
  33899=>"000010001",
  33900=>"111010000",
  33901=>"110100010",
  33902=>"000111011",
  33903=>"100111111",
  33904=>"100011001",
  33905=>"111101011",
  33906=>"100110111",
  33907=>"001001001",
  33908=>"111101111",
  33909=>"010111101",
  33910=>"011001100",
  33911=>"000000010",
  33912=>"101001111",
  33913=>"011011101",
  33914=>"011010011",
  33915=>"000011001",
  33916=>"101110010",
  33917=>"101100010",
  33918=>"111000111",
  33919=>"110011000",
  33920=>"111110101",
  33921=>"011011011",
  33922=>"011001110",
  33923=>"010000001",
  33924=>"010010000",
  33925=>"001001111",
  33926=>"001111011",
  33927=>"111001100",
  33928=>"111101000",
  33929=>"101001100",
  33930=>"001111101",
  33931=>"001111001",
  33932=>"110000111",
  33933=>"110100110",
  33934=>"111101011",
  33935=>"000100000",
  33936=>"110011001",
  33937=>"111011001",
  33938=>"110111011",
  33939=>"011001111",
  33940=>"011111000",
  33941=>"101111011",
  33942=>"111110101",
  33943=>"010100111",
  33944=>"011111101",
  33945=>"111000110",
  33946=>"000010010",
  33947=>"111011010",
  33948=>"001010100",
  33949=>"010000000",
  33950=>"011100000",
  33951=>"110011110",
  33952=>"011110111",
  33953=>"001010001",
  33954=>"110100101",
  33955=>"101110100",
  33956=>"101001011",
  33957=>"101010111",
  33958=>"110101100",
  33959=>"011001110",
  33960=>"101101111",
  33961=>"011010110",
  33962=>"110011100",
  33963=>"000000011",
  33964=>"001100101",
  33965=>"100110011",
  33966=>"001010000",
  33967=>"101011110",
  33968=>"101111000",
  33969=>"011010000",
  33970=>"010001111",
  33971=>"100110011",
  33972=>"001010010",
  33973=>"100111111",
  33974=>"010101100",
  33975=>"010110001",
  33976=>"001011000",
  33977=>"011110111",
  33978=>"110110100",
  33979=>"011101111",
  33980=>"001100100",
  33981=>"000001000",
  33982=>"111111011",
  33983=>"110000111",
  33984=>"001001000",
  33985=>"010001001",
  33986=>"111000100",
  33987=>"001100010",
  33988=>"111010001",
  33989=>"000100010",
  33990=>"101100111",
  33991=>"100001100",
  33992=>"000001001",
  33993=>"110001000",
  33994=>"000101101",
  33995=>"101110011",
  33996=>"000111010",
  33997=>"001100110",
  33998=>"011001100",
  33999=>"010110010",
  34000=>"100110100",
  34001=>"100101000",
  34002=>"011110011",
  34003=>"011111100",
  34004=>"100011010",
  34005=>"001110001",
  34006=>"100110001",
  34007=>"101000001",
  34008=>"111001110",
  34009=>"101011101",
  34010=>"100100000",
  34011=>"011010010",
  34012=>"110000111",
  34013=>"100000101",
  34014=>"110001011",
  34015=>"110111111",
  34016=>"000101110",
  34017=>"000000001",
  34018=>"000011110",
  34019=>"010111011",
  34020=>"100111111",
  34021=>"000001011",
  34022=>"010110011",
  34023=>"110100100",
  34024=>"110101111",
  34025=>"111000100",
  34026=>"101000111",
  34027=>"010100111",
  34028=>"000010000",
  34029=>"111111000",
  34030=>"111100011",
  34031=>"100010000",
  34032=>"100010110",
  34033=>"101101111",
  34034=>"010010100",
  34035=>"000011000",
  34036=>"100110010",
  34037=>"001101110",
  34038=>"111111111",
  34039=>"000110001",
  34040=>"000111010",
  34041=>"011111010",
  34042=>"000100111",
  34043=>"000101011",
  34044=>"010001011",
  34045=>"100001101",
  34046=>"001101101",
  34047=>"111010010",
  34048=>"000100111",
  34049=>"011110010",
  34050=>"111100111",
  34051=>"011100010",
  34052=>"101001000",
  34053=>"001100111",
  34054=>"010010110",
  34055=>"101010011",
  34056=>"001000110",
  34057=>"111000101",
  34058=>"100010101",
  34059=>"011111010",
  34060=>"010111000",
  34061=>"110010110",
  34062=>"110111100",
  34063=>"110100011",
  34064=>"100000001",
  34065=>"111101000",
  34066=>"001110011",
  34067=>"010011011",
  34068=>"000011110",
  34069=>"001111010",
  34070=>"111101000",
  34071=>"111110101",
  34072=>"000101001",
  34073=>"100100100",
  34074=>"000110100",
  34075=>"110101111",
  34076=>"010111010",
  34077=>"000101010",
  34078=>"111111010",
  34079=>"111001100",
  34080=>"001010101",
  34081=>"000000111",
  34082=>"110110101",
  34083=>"111000010",
  34084=>"001110000",
  34085=>"000010111",
  34086=>"001101100",
  34087=>"001110111",
  34088=>"010100111",
  34089=>"100011001",
  34090=>"000011100",
  34091=>"000110111",
  34092=>"001100011",
  34093=>"110000001",
  34094=>"111110000",
  34095=>"101101000",
  34096=>"010110010",
  34097=>"000001010",
  34098=>"001010011",
  34099=>"011010010",
  34100=>"111000110",
  34101=>"010100010",
  34102=>"011110000",
  34103=>"111101100",
  34104=>"110010000",
  34105=>"010111101",
  34106=>"011000010",
  34107=>"101001111",
  34108=>"111011110",
  34109=>"001000101",
  34110=>"000101001",
  34111=>"000001000",
  34112=>"001111011",
  34113=>"110111110",
  34114=>"100001101",
  34115=>"110010011",
  34116=>"101110000",
  34117=>"101100010",
  34118=>"001100111",
  34119=>"011111010",
  34120=>"011101000",
  34121=>"001110011",
  34122=>"110010111",
  34123=>"000111110",
  34124=>"011000011",
  34125=>"000010011",
  34126=>"101001100",
  34127=>"110010100",
  34128=>"000111010",
  34129=>"001000101",
  34130=>"101010010",
  34131=>"101010110",
  34132=>"010111000",
  34133=>"111011001",
  34134=>"000100001",
  34135=>"111110110",
  34136=>"010110110",
  34137=>"000001101",
  34138=>"110101001",
  34139=>"110100011",
  34140=>"011101110",
  34141=>"101101111",
  34142=>"111001001",
  34143=>"001010101",
  34144=>"110000000",
  34145=>"111101100",
  34146=>"011000101",
  34147=>"001101101",
  34148=>"010110000",
  34149=>"000100000",
  34150=>"001011011",
  34151=>"110101000",
  34152=>"001101000",
  34153=>"001110000",
  34154=>"101101101",
  34155=>"100000101",
  34156=>"111110100",
  34157=>"100011111",
  34158=>"101001100",
  34159=>"001110010",
  34160=>"000000101",
  34161=>"000010100",
  34162=>"101001010",
  34163=>"001010101",
  34164=>"101000000",
  34165=>"100001111",
  34166=>"001110001",
  34167=>"110010000",
  34168=>"011010100",
  34169=>"011000011",
  34170=>"001101110",
  34171=>"111011000",
  34172=>"010000011",
  34173=>"011001110",
  34174=>"111011101",
  34175=>"001111010",
  34176=>"111101001",
  34177=>"101011110",
  34178=>"011101101",
  34179=>"010011000",
  34180=>"100101101",
  34181=>"010100111",
  34182=>"001110101",
  34183=>"100100000",
  34184=>"110110110",
  34185=>"011110111",
  34186=>"100110101",
  34187=>"110111101",
  34188=>"010101110",
  34189=>"101101101",
  34190=>"000000000",
  34191=>"111011111",
  34192=>"001100111",
  34193=>"101001110",
  34194=>"111110000",
  34195=>"110100100",
  34196=>"110001010",
  34197=>"011011101",
  34198=>"001001001",
  34199=>"110000010",
  34200=>"011010001",
  34201=>"010110001",
  34202=>"011000011",
  34203=>"001101001",
  34204=>"111111000",
  34205=>"111100101",
  34206=>"110111111",
  34207=>"000110001",
  34208=>"111010100",
  34209=>"110111101",
  34210=>"111010110",
  34211=>"110111111",
  34212=>"101000100",
  34213=>"101111111",
  34214=>"000110000",
  34215=>"000101000",
  34216=>"110110101",
  34217=>"010001111",
  34218=>"100000100",
  34219=>"000000010",
  34220=>"110010110",
  34221=>"011000010",
  34222=>"101001100",
  34223=>"010000001",
  34224=>"011100111",
  34225=>"110010011",
  34226=>"100000010",
  34227=>"011001000",
  34228=>"101101100",
  34229=>"110000101",
  34230=>"110000011",
  34231=>"110100110",
  34232=>"011110111",
  34233=>"000010100",
  34234=>"001100011",
  34235=>"110110110",
  34236=>"101111011",
  34237=>"000000100",
  34238=>"000011111",
  34239=>"100000100",
  34240=>"101100100",
  34241=>"011000100",
  34242=>"011000001",
  34243=>"101000011",
  34244=>"011110001",
  34245=>"011000001",
  34246=>"110111111",
  34247=>"111001110",
  34248=>"011101011",
  34249=>"010001010",
  34250=>"100000010",
  34251=>"111011111",
  34252=>"010100101",
  34253=>"101001010",
  34254=>"010000010",
  34255=>"101100000",
  34256=>"100011010",
  34257=>"101101010",
  34258=>"111111101",
  34259=>"011000100",
  34260=>"100100101",
  34261=>"000001110",
  34262=>"111000011",
  34263=>"011010000",
  34264=>"010111100",
  34265=>"100101010",
  34266=>"111010010",
  34267=>"000100000",
  34268=>"100110011",
  34269=>"000011001",
  34270=>"101101010",
  34271=>"001001011",
  34272=>"110111100",
  34273=>"000011111",
  34274=>"011110000",
  34275=>"010010000",
  34276=>"000100100",
  34277=>"100101101",
  34278=>"101111000",
  34279=>"011001000",
  34280=>"101001010",
  34281=>"010101101",
  34282=>"101010010",
  34283=>"001010001",
  34284=>"010010111",
  34285=>"011100111",
  34286=>"110010010",
  34287=>"010010100",
  34288=>"110001010",
  34289=>"101011001",
  34290=>"100111011",
  34291=>"001101111",
  34292=>"111101101",
  34293=>"111010111",
  34294=>"010000101",
  34295=>"110001111",
  34296=>"100111110",
  34297=>"100111110",
  34298=>"111100110",
  34299=>"001000100",
  34300=>"111010100",
  34301=>"111101011",
  34302=>"000111100",
  34303=>"100110110",
  34304=>"000011010",
  34305=>"100000010",
  34306=>"110101100",
  34307=>"010011101",
  34308=>"000000011",
  34309=>"101110010",
  34310=>"101010000",
  34311=>"101011011",
  34312=>"101011011",
  34313=>"010011001",
  34314=>"101100010",
  34315=>"000010100",
  34316=>"000011001",
  34317=>"001000111",
  34318=>"000000110",
  34319=>"101010000",
  34320=>"010101101",
  34321=>"001110001",
  34322=>"110011111",
  34323=>"010010110",
  34324=>"101110011",
  34325=>"010001010",
  34326=>"110111011",
  34327=>"010101110",
  34328=>"100110111",
  34329=>"100101000",
  34330=>"110011011",
  34331=>"001111110",
  34332=>"100010110",
  34333=>"011010010",
  34334=>"100101001",
  34335=>"110011011",
  34336=>"001001010",
  34337=>"010011100",
  34338=>"100001100",
  34339=>"010011101",
  34340=>"011010101",
  34341=>"010110101",
  34342=>"110001001",
  34343=>"110111001",
  34344=>"101011000",
  34345=>"110100010",
  34346=>"010110011",
  34347=>"010100011",
  34348=>"000010111",
  34349=>"110010010",
  34350=>"011000111",
  34351=>"000011001",
  34352=>"010110011",
  34353=>"000010011",
  34354=>"100001110",
  34355=>"001101000",
  34356=>"110111101",
  34357=>"100011000",
  34358=>"001111010",
  34359=>"111010111",
  34360=>"101100111",
  34361=>"011111000",
  34362=>"011101111",
  34363=>"111101110",
  34364=>"001011001",
  34365=>"010001100",
  34366=>"100001111",
  34367=>"100111101",
  34368=>"001001010",
  34369=>"000001010",
  34370=>"001101001",
  34371=>"111000000",
  34372=>"010111100",
  34373=>"101110111",
  34374=>"101001000",
  34375=>"000110001",
  34376=>"100110011",
  34377=>"011100101",
  34378=>"111110000",
  34379=>"000101001",
  34380=>"110011111",
  34381=>"110001011",
  34382=>"100101010",
  34383=>"110001111",
  34384=>"110111111",
  34385=>"101001000",
  34386=>"000000111",
  34387=>"100011000",
  34388=>"001010000",
  34389=>"101110001",
  34390=>"010001001",
  34391=>"010000000",
  34392=>"101101101",
  34393=>"000110110",
  34394=>"101011001",
  34395=>"110110011",
  34396=>"011001111",
  34397=>"010101101",
  34398=>"011001111",
  34399=>"101100011",
  34400=>"010111011",
  34401=>"000110101",
  34402=>"000100011",
  34403=>"101000000",
  34404=>"001111010",
  34405=>"000110011",
  34406=>"101101000",
  34407=>"010001100",
  34408=>"110001101",
  34409=>"110001001",
  34410=>"111111000",
  34411=>"001111100",
  34412=>"100000111",
  34413=>"011101100",
  34414=>"011011010",
  34415=>"111010110",
  34416=>"101001000",
  34417=>"110000100",
  34418=>"011110110",
  34419=>"110010001",
  34420=>"100101011",
  34421=>"111000000",
  34422=>"011111110",
  34423=>"011001000",
  34424=>"010010110",
  34425=>"100100111",
  34426=>"110111000",
  34427=>"000100001",
  34428=>"011011000",
  34429=>"110011011",
  34430=>"101001000",
  34431=>"000000100",
  34432=>"111110010",
  34433=>"111001010",
  34434=>"100001111",
  34435=>"100010111",
  34436=>"110011101",
  34437=>"101000101",
  34438=>"010011010",
  34439=>"110010111",
  34440=>"010001110",
  34441=>"000010000",
  34442=>"010101111",
  34443=>"110101101",
  34444=>"010101111",
  34445=>"100011000",
  34446=>"011101110",
  34447=>"100010110",
  34448=>"111100101",
  34449=>"110111101",
  34450=>"001011100",
  34451=>"000011101",
  34452=>"000001101",
  34453=>"011101011",
  34454=>"010010101",
  34455=>"010001001",
  34456=>"111011000",
  34457=>"111100100",
  34458=>"000000001",
  34459=>"001010010",
  34460=>"111111100",
  34461=>"001100010",
  34462=>"001011111",
  34463=>"010010011",
  34464=>"000111110",
  34465=>"110010111",
  34466=>"001010001",
  34467=>"000011011",
  34468=>"011100111",
  34469=>"100111011",
  34470=>"100100010",
  34471=>"011110001",
  34472=>"110010100",
  34473=>"110000011",
  34474=>"100100110",
  34475=>"001111000",
  34476=>"001111101",
  34477=>"001101000",
  34478=>"001100000",
  34479=>"100010001",
  34480=>"000000001",
  34481=>"010000011",
  34482=>"001000100",
  34483=>"110101110",
  34484=>"010010010",
  34485=>"110001011",
  34486=>"000000100",
  34487=>"111100010",
  34488=>"011001001",
  34489=>"100010001",
  34490=>"001111110",
  34491=>"011001010",
  34492=>"101101001",
  34493=>"111100110",
  34494=>"101101001",
  34495=>"001101101",
  34496=>"010110110",
  34497=>"111101100",
  34498=>"010010010",
  34499=>"101010100",
  34500=>"111011011",
  34501=>"101010100",
  34502=>"100111010",
  34503=>"111000110",
  34504=>"000001110",
  34505=>"000100110",
  34506=>"001010100",
  34507=>"010011110",
  34508=>"111100011",
  34509=>"110101100",
  34510=>"100000011",
  34511=>"111000111",
  34512=>"000101001",
  34513=>"100111000",
  34514=>"110011110",
  34515=>"000010101",
  34516=>"110110011",
  34517=>"100011000",
  34518=>"011010001",
  34519=>"000011011",
  34520=>"010011011",
  34521=>"101011100",
  34522=>"011000001",
  34523=>"111110011",
  34524=>"100110101",
  34525=>"110001000",
  34526=>"100100110",
  34527=>"011110000",
  34528=>"110110110",
  34529=>"100110001",
  34530=>"101000000",
  34531=>"011100110",
  34532=>"100110110",
  34533=>"011000011",
  34534=>"001111101",
  34535=>"001011011",
  34536=>"010100111",
  34537=>"110000000",
  34538=>"111111001",
  34539=>"000010010",
  34540=>"001010101",
  34541=>"101001100",
  34542=>"011001100",
  34543=>"101000001",
  34544=>"110001101",
  34545=>"100001110",
  34546=>"100111111",
  34547=>"010100011",
  34548=>"110100101",
  34549=>"100111011",
  34550=>"111111111",
  34551=>"111100100",
  34552=>"001110011",
  34553=>"100011110",
  34554=>"010101100",
  34555=>"110000010",
  34556=>"001101001",
  34557=>"011101110",
  34558=>"010001110",
  34559=>"011000110",
  34560=>"100000001",
  34561=>"111100001",
  34562=>"111100101",
  34563=>"011000010",
  34564=>"011010110",
  34565=>"001010010",
  34566=>"110111001",
  34567=>"001111010",
  34568=>"111001100",
  34569=>"000011101",
  34570=>"011000110",
  34571=>"000110101",
  34572=>"011100100",
  34573=>"111000010",
  34574=>"100010000",
  34575=>"000110001",
  34576=>"101110001",
  34577=>"111000010",
  34578=>"101001101",
  34579=>"111000000",
  34580=>"100010010",
  34581=>"001011010",
  34582=>"000100010",
  34583=>"110101000",
  34584=>"101101101",
  34585=>"000101001",
  34586=>"000001101",
  34587=>"110000011",
  34588=>"000110001",
  34589=>"111110111",
  34590=>"011000001",
  34591=>"101101000",
  34592=>"001001100",
  34593=>"010110100",
  34594=>"011011110",
  34595=>"001110000",
  34596=>"011101000",
  34597=>"010101001",
  34598=>"000111011",
  34599=>"011101101",
  34600=>"000001110",
  34601=>"110000110",
  34602=>"010100101",
  34603=>"111010000",
  34604=>"000011100",
  34605=>"011011110",
  34606=>"000111101",
  34607=>"010010001",
  34608=>"110101000",
  34609=>"011010011",
  34610=>"000001011",
  34611=>"000011001",
  34612=>"110101110",
  34613=>"101011011",
  34614=>"011110101",
  34615=>"110101100",
  34616=>"111101110",
  34617=>"000001001",
  34618=>"011010000",
  34619=>"010000100",
  34620=>"101011010",
  34621=>"100010010",
  34622=>"001100000",
  34623=>"001011010",
  34624=>"000110100",
  34625=>"101110100",
  34626=>"111010001",
  34627=>"001011111",
  34628=>"011000001",
  34629=>"000101010",
  34630=>"010011000",
  34631=>"000011110",
  34632=>"011001111",
  34633=>"000100010",
  34634=>"100001100",
  34635=>"001101111",
  34636=>"001001100",
  34637=>"000000111",
  34638=>"100110011",
  34639=>"011001100",
  34640=>"111011100",
  34641=>"001110000",
  34642=>"110111011",
  34643=>"010111011",
  34644=>"001010011",
  34645=>"010101110",
  34646=>"111010101",
  34647=>"110011010",
  34648=>"110010001",
  34649=>"010101011",
  34650=>"000001111",
  34651=>"111111110",
  34652=>"110011000",
  34653=>"101100110",
  34654=>"111011010",
  34655=>"101100100",
  34656=>"100001110",
  34657=>"010101001",
  34658=>"000001111",
  34659=>"010010111",
  34660=>"010111011",
  34661=>"000101001",
  34662=>"001101110",
  34663=>"000101110",
  34664=>"100110100",
  34665=>"111111010",
  34666=>"111011001",
  34667=>"101001010",
  34668=>"001100000",
  34669=>"011010000",
  34670=>"111101011",
  34671=>"011101010",
  34672=>"101010100",
  34673=>"000000101",
  34674=>"111110000",
  34675=>"010011110",
  34676=>"001010001",
  34677=>"010010011",
  34678=>"100000011",
  34679=>"011100101",
  34680=>"011111011",
  34681=>"000010111",
  34682=>"101110110",
  34683=>"101110110",
  34684=>"011001111",
  34685=>"100101101",
  34686=>"011110000",
  34687=>"101010111",
  34688=>"100000001",
  34689=>"011001011",
  34690=>"000100000",
  34691=>"110111101",
  34692=>"000100010",
  34693=>"001010010",
  34694=>"100110001",
  34695=>"110010001",
  34696=>"001001000",
  34697=>"011000101",
  34698=>"000100100",
  34699=>"001100000",
  34700=>"011100111",
  34701=>"111110101",
  34702=>"000001001",
  34703=>"000100101",
  34704=>"001110100",
  34705=>"011111011",
  34706=>"000100101",
  34707=>"110110010",
  34708=>"101110001",
  34709=>"011111111",
  34710=>"101101110",
  34711=>"001000100",
  34712=>"111000111",
  34713=>"011011101",
  34714=>"000101101",
  34715=>"010111111",
  34716=>"111100101",
  34717=>"000100010",
  34718=>"101111110",
  34719=>"100000010",
  34720=>"110000010",
  34721=>"100011100",
  34722=>"001111011",
  34723=>"011001011",
  34724=>"001001111",
  34725=>"101010010",
  34726=>"110100001",
  34727=>"111101010",
  34728=>"000011001",
  34729=>"111101001",
  34730=>"110001010",
  34731=>"001101010",
  34732=>"001010100",
  34733=>"111000001",
  34734=>"011001110",
  34735=>"111011111",
  34736=>"010000000",
  34737=>"110100100",
  34738=>"000001001",
  34739=>"000111000",
  34740=>"011010100",
  34741=>"011100110",
  34742=>"011100011",
  34743=>"001000110",
  34744=>"011010001",
  34745=>"101001001",
  34746=>"001111110",
  34747=>"010101011",
  34748=>"111101111",
  34749=>"010011110",
  34750=>"000100110",
  34751=>"101000111",
  34752=>"001011010",
  34753=>"111000111",
  34754=>"000001011",
  34755=>"111100100",
  34756=>"110111111",
  34757=>"101011101",
  34758=>"011110110",
  34759=>"101110101",
  34760=>"101001100",
  34761=>"100000001",
  34762=>"011101101",
  34763=>"010000100",
  34764=>"001111000",
  34765=>"010000010",
  34766=>"110010010",
  34767=>"100011111",
  34768=>"111101011",
  34769=>"000001101",
  34770=>"010101100",
  34771=>"001011010",
  34772=>"101000000",
  34773=>"000001010",
  34774=>"100010010",
  34775=>"000010011",
  34776=>"000110110",
  34777=>"110111100",
  34778=>"001110111",
  34779=>"010100100",
  34780=>"001111101",
  34781=>"001011000",
  34782=>"000000010",
  34783=>"010000110",
  34784=>"100011101",
  34785=>"101011011",
  34786=>"001001111",
  34787=>"010001000",
  34788=>"111001001",
  34789=>"011001010",
  34790=>"101110001",
  34791=>"001101110",
  34792=>"001001011",
  34793=>"010011101",
  34794=>"011100100",
  34795=>"001101100",
  34796=>"011010001",
  34797=>"000101001",
  34798=>"011101101",
  34799=>"011111010",
  34800=>"101000101",
  34801=>"111101110",
  34802=>"010101101",
  34803=>"001000011",
  34804=>"001100011",
  34805=>"001000011",
  34806=>"001000000",
  34807=>"000001011",
  34808=>"000000010",
  34809=>"101110001",
  34810=>"010100001",
  34811=>"101110111",
  34812=>"010011110",
  34813=>"110101110",
  34814=>"010011101",
  34815=>"001110011",
  34816=>"101000001",
  34817=>"111111110",
  34818=>"001000100",
  34819=>"101000000",
  34820=>"110001010",
  34821=>"100010010",
  34822=>"000100110",
  34823=>"100110000",
  34824=>"001010001",
  34825=>"001010101",
  34826=>"111101000",
  34827=>"001101011",
  34828=>"001001011",
  34829=>"101100000",
  34830=>"001011100",
  34831=>"110000111",
  34832=>"101111001",
  34833=>"101000110",
  34834=>"111111010",
  34835=>"111011001",
  34836=>"111100101",
  34837=>"011001000",
  34838=>"101011100",
  34839=>"101100010",
  34840=>"110010111",
  34841=>"101100100",
  34842=>"000111001",
  34843=>"011000110",
  34844=>"111000010",
  34845=>"000010100",
  34846=>"111010011",
  34847=>"000001000",
  34848=>"111100011",
  34849=>"000111000",
  34850=>"001010000",
  34851=>"011110111",
  34852=>"110111110",
  34853=>"010101101",
  34854=>"110000101",
  34855=>"110110001",
  34856=>"101010100",
  34857=>"011001111",
  34858=>"100111010",
  34859=>"010000111",
  34860=>"101011111",
  34861=>"010001010",
  34862=>"001001000",
  34863=>"111111110",
  34864=>"010001101",
  34865=>"011010100",
  34866=>"001101010",
  34867=>"010011011",
  34868=>"000000000",
  34869=>"010111000",
  34870=>"111010000",
  34871=>"001010010",
  34872=>"101110010",
  34873=>"010010001",
  34874=>"110110101",
  34875=>"111000100",
  34876=>"100110010",
  34877=>"011010100",
  34878=>"110100000",
  34879=>"110110111",
  34880=>"110000011",
  34881=>"001000001",
  34882=>"011011000",
  34883=>"000000110",
  34884=>"010111110",
  34885=>"010110100",
  34886=>"101001011",
  34887=>"010111101",
  34888=>"000001100",
  34889=>"001001101",
  34890=>"010110011",
  34891=>"100111100",
  34892=>"111000100",
  34893=>"010011111",
  34894=>"100001110",
  34895=>"011001001",
  34896=>"001000100",
  34897=>"010001011",
  34898=>"100001111",
  34899=>"010110011",
  34900=>"001111011",
  34901=>"110010011",
  34902=>"100100101",
  34903=>"101010001",
  34904=>"111000100",
  34905=>"111000001",
  34906=>"111011111",
  34907=>"110101000",
  34908=>"100000000",
  34909=>"001010110",
  34910=>"110110101",
  34911=>"011111010",
  34912=>"111000001",
  34913=>"101101100",
  34914=>"001111111",
  34915=>"110100111",
  34916=>"110101001",
  34917=>"100000001",
  34918=>"100000111",
  34919=>"010000101",
  34920=>"101000000",
  34921=>"100100010",
  34922=>"011001010",
  34923=>"100001011",
  34924=>"011110011",
  34925=>"010001000",
  34926=>"111100010",
  34927=>"010010010",
  34928=>"111011011",
  34929=>"000000100",
  34930=>"001010100",
  34931=>"001011010",
  34932=>"000011011",
  34933=>"011111100",
  34934=>"010111101",
  34935=>"011010111",
  34936=>"010100010",
  34937=>"010110001",
  34938=>"000101010",
  34939=>"010010110",
  34940=>"000011111",
  34941=>"110110111",
  34942=>"100000010",
  34943=>"001100011",
  34944=>"100101111",
  34945=>"010010111",
  34946=>"111101110",
  34947=>"111010100",
  34948=>"110011011",
  34949=>"100101010",
  34950=>"001001110",
  34951=>"101000000",
  34952=>"011110100",
  34953=>"110111011",
  34954=>"110011011",
  34955=>"000101111",
  34956=>"100101110",
  34957=>"010011000",
  34958=>"000011001",
  34959=>"011110100",
  34960=>"101101011",
  34961=>"101000101",
  34962=>"010110111",
  34963=>"110100101",
  34964=>"000100101",
  34965=>"100101101",
  34966=>"010110001",
  34967=>"111010000",
  34968=>"001000000",
  34969=>"001000101",
  34970=>"001010111",
  34971=>"000110000",
  34972=>"010111101",
  34973=>"001001100",
  34974=>"011100011",
  34975=>"110001100",
  34976=>"111000010",
  34977=>"100100100",
  34978=>"101101110",
  34979=>"111000111",
  34980=>"100111011",
  34981=>"010001001",
  34982=>"111100000",
  34983=>"101011011",
  34984=>"110101100",
  34985=>"100000100",
  34986=>"111000011",
  34987=>"111111111",
  34988=>"110101111",
  34989=>"111001001",
  34990=>"000000110",
  34991=>"111001011",
  34992=>"110101110",
  34993=>"010001100",
  34994=>"001100111",
  34995=>"001000011",
  34996=>"000011111",
  34997=>"010100111",
  34998=>"001111011",
  34999=>"111011011",
  35000=>"011000010",
  35001=>"000011111",
  35002=>"110011010",
  35003=>"000101011",
  35004=>"111001001",
  35005=>"000110001",
  35006=>"011111110",
  35007=>"101111011",
  35008=>"101110101",
  35009=>"011010101",
  35010=>"101101111",
  35011=>"001111110",
  35012=>"100110011",
  35013=>"000001101",
  35014=>"111001001",
  35015=>"110011010",
  35016=>"010101001",
  35017=>"101011001",
  35018=>"001101101",
  35019=>"000111011",
  35020=>"110100110",
  35021=>"000000010",
  35022=>"001111010",
  35023=>"111110111",
  35024=>"110100100",
  35025=>"010111101",
  35026=>"000000010",
  35027=>"001010101",
  35028=>"000111100",
  35029=>"111010101",
  35030=>"111111011",
  35031=>"110110101",
  35032=>"000011001",
  35033=>"100011100",
  35034=>"110011001",
  35035=>"011010101",
  35036=>"000011000",
  35037=>"101011110",
  35038=>"010100110",
  35039=>"100101101",
  35040=>"111111110",
  35041=>"110111000",
  35042=>"100110001",
  35043=>"000010011",
  35044=>"000011110",
  35045=>"100110110",
  35046=>"000101100",
  35047=>"110111000",
  35048=>"010100101",
  35049=>"001001100",
  35050=>"001100111",
  35051=>"000101110",
  35052=>"011010101",
  35053=>"001011000",
  35054=>"001011110",
  35055=>"011111110",
  35056=>"101110000",
  35057=>"000011001",
  35058=>"010001001",
  35059=>"010111000",
  35060=>"111101001",
  35061=>"110111100",
  35062=>"100000101",
  35063=>"010000010",
  35064=>"001100110",
  35065=>"111101110",
  35066=>"101110001",
  35067=>"010011001",
  35068=>"100111010",
  35069=>"000101100",
  35070=>"101000001",
  35071=>"000111011",
  35072=>"000111001",
  35073=>"110010011",
  35074=>"001000101",
  35075=>"001100101",
  35076=>"010011000",
  35077=>"111010000",
  35078=>"010010111",
  35079=>"000111011",
  35080=>"010000000",
  35081=>"010001110",
  35082=>"000100101",
  35083=>"100110110",
  35084=>"001011001",
  35085=>"010101110",
  35086=>"011100111",
  35087=>"001101111",
  35088=>"001000110",
  35089=>"010111011",
  35090=>"001110011",
  35091=>"111101101",
  35092=>"111001010",
  35093=>"110111011",
  35094=>"011010010",
  35095=>"000000001",
  35096=>"110010000",
  35097=>"101010010",
  35098=>"010111011",
  35099=>"010101010",
  35100=>"001011011",
  35101=>"110011001",
  35102=>"100110011",
  35103=>"110000110",
  35104=>"110101100",
  35105=>"111100100",
  35106=>"001001110",
  35107=>"000110101",
  35108=>"001100011",
  35109=>"111110000",
  35110=>"011111101",
  35111=>"110001011",
  35112=>"100010011",
  35113=>"000010100",
  35114=>"110110100",
  35115=>"010100000",
  35116=>"010010010",
  35117=>"110011101",
  35118=>"000101111",
  35119=>"010101100",
  35120=>"110110010",
  35121=>"010111111",
  35122=>"000010100",
  35123=>"011110111",
  35124=>"011000110",
  35125=>"011000110",
  35126=>"101010110",
  35127=>"111101001",
  35128=>"101001000",
  35129=>"111110010",
  35130=>"101101110",
  35131=>"100100001",
  35132=>"111011110",
  35133=>"010011111",
  35134=>"001000010",
  35135=>"111010010",
  35136=>"111011000",
  35137=>"010101111",
  35138=>"100010100",
  35139=>"101001011",
  35140=>"101001000",
  35141=>"111000100",
  35142=>"100100100",
  35143=>"000000110",
  35144=>"100110000",
  35145=>"100110011",
  35146=>"001110010",
  35147=>"001101011",
  35148=>"100010001",
  35149=>"101011101",
  35150=>"000011011",
  35151=>"001011110",
  35152=>"111101000",
  35153=>"101000110",
  35154=>"111101101",
  35155=>"100001010",
  35156=>"001001100",
  35157=>"111011000",
  35158=>"110111111",
  35159=>"100111101",
  35160=>"011101110",
  35161=>"011111100",
  35162=>"111100101",
  35163=>"110001100",
  35164=>"111111000",
  35165=>"100110101",
  35166=>"011011010",
  35167=>"111001010",
  35168=>"100000111",
  35169=>"110001001",
  35170=>"000100011",
  35171=>"100100100",
  35172=>"010010011",
  35173=>"011111001",
  35174=>"001101111",
  35175=>"011001000",
  35176=>"110111010",
  35177=>"110001011",
  35178=>"110010100",
  35179=>"001110010",
  35180=>"111000101",
  35181=>"010010101",
  35182=>"100011100",
  35183=>"011001100",
  35184=>"010001100",
  35185=>"110111111",
  35186=>"110011000",
  35187=>"100100011",
  35188=>"001111001",
  35189=>"001110010",
  35190=>"100010111",
  35191=>"001101101",
  35192=>"010110000",
  35193=>"100100000",
  35194=>"101100011",
  35195=>"001100101",
  35196=>"010001000",
  35197=>"111111101",
  35198=>"110111010",
  35199=>"101110011",
  35200=>"100010101",
  35201=>"010011100",
  35202=>"000100010",
  35203=>"010010011",
  35204=>"110010011",
  35205=>"111000000",
  35206=>"100010011",
  35207=>"001011010",
  35208=>"010011000",
  35209=>"000101000",
  35210=>"011110001",
  35211=>"111011011",
  35212=>"110001100",
  35213=>"011010000",
  35214=>"111010011",
  35215=>"100010100",
  35216=>"111000101",
  35217=>"010000100",
  35218=>"010000110",
  35219=>"101000100",
  35220=>"011000011",
  35221=>"100101010",
  35222=>"001010000",
  35223=>"000100000",
  35224=>"111110011",
  35225=>"000001111",
  35226=>"011001100",
  35227=>"011010001",
  35228=>"000010010",
  35229=>"011111101",
  35230=>"011000100",
  35231=>"110101000",
  35232=>"010011011",
  35233=>"101001011",
  35234=>"010011000",
  35235=>"000000010",
  35236=>"011110011",
  35237=>"100000111",
  35238=>"000001110",
  35239=>"001001010",
  35240=>"000101111",
  35241=>"100010001",
  35242=>"000000110",
  35243=>"110110110",
  35244=>"000001110",
  35245=>"001100001",
  35246=>"101010010",
  35247=>"110010101",
  35248=>"010101101",
  35249=>"010101000",
  35250=>"110011011",
  35251=>"110111010",
  35252=>"100001100",
  35253=>"000101110",
  35254=>"110011001",
  35255=>"000110001",
  35256=>"101010111",
  35257=>"000101010",
  35258=>"100001101",
  35259=>"000000111",
  35260=>"110001001",
  35261=>"001101011",
  35262=>"010101001",
  35263=>"000000110",
  35264=>"101001000",
  35265=>"000111111",
  35266=>"011000100",
  35267=>"100110000",
  35268=>"001000011",
  35269=>"011110110",
  35270=>"111001011",
  35271=>"101001000",
  35272=>"101110110",
  35273=>"001111101",
  35274=>"011001101",
  35275=>"100111100",
  35276=>"101001101",
  35277=>"110001100",
  35278=>"001011000",
  35279=>"010011110",
  35280=>"110001001",
  35281=>"000010101",
  35282=>"010110001",
  35283=>"101011001",
  35284=>"010010000",
  35285=>"001010110",
  35286=>"110110010",
  35287=>"001100000",
  35288=>"111101111",
  35289=>"100100001",
  35290=>"111110011",
  35291=>"110000100",
  35292=>"010000001",
  35293=>"001000010",
  35294=>"001000001",
  35295=>"011100101",
  35296=>"000110001",
  35297=>"100011111",
  35298=>"000001111",
  35299=>"010111001",
  35300=>"000000100",
  35301=>"100110111",
  35302=>"000001001",
  35303=>"000010010",
  35304=>"110000011",
  35305=>"000100111",
  35306=>"100011011",
  35307=>"000100100",
  35308=>"001001000",
  35309=>"110000110",
  35310=>"001100011",
  35311=>"011001001",
  35312=>"100000011",
  35313=>"101111100",
  35314=>"010111001",
  35315=>"001100000",
  35316=>"011010101",
  35317=>"001100111",
  35318=>"001001010",
  35319=>"010100111",
  35320=>"101001010",
  35321=>"011100100",
  35322=>"100110000",
  35323=>"101111000",
  35324=>"100111111",
  35325=>"000001111",
  35326=>"000100011",
  35327=>"010110010",
  35328=>"111111101",
  35329=>"111000010",
  35330=>"001011011",
  35331=>"100001100",
  35332=>"001011111",
  35333=>"011000011",
  35334=>"111010111",
  35335=>"101111010",
  35336=>"110100001",
  35337=>"000000111",
  35338=>"111100000",
  35339=>"011111100",
  35340=>"010111111",
  35341=>"111100111",
  35342=>"001000001",
  35343=>"000001010",
  35344=>"110111111",
  35345=>"111000000",
  35346=>"011011111",
  35347=>"001000010",
  35348=>"000100100",
  35349=>"101011000",
  35350=>"111010000",
  35351=>"111111110",
  35352=>"000100010",
  35353=>"110101110",
  35354=>"111000001",
  35355=>"101110101",
  35356=>"010000001",
  35357=>"101000100",
  35358=>"001011100",
  35359=>"101001110",
  35360=>"110110001",
  35361=>"101001101",
  35362=>"000110001",
  35363=>"000000011",
  35364=>"111011010",
  35365=>"011111111",
  35366=>"011010010",
  35367=>"001001011",
  35368=>"100100001",
  35369=>"001110111",
  35370=>"111100000",
  35371=>"000100001",
  35372=>"011111110",
  35373=>"001111110",
  35374=>"101001000",
  35375=>"100011001",
  35376=>"000100100",
  35377=>"011011110",
  35378=>"100100110",
  35379=>"111011101",
  35380=>"000001011",
  35381=>"100100111",
  35382=>"010100000",
  35383=>"110111110",
  35384=>"111010111",
  35385=>"010101010",
  35386=>"010110111",
  35387=>"111101110",
  35388=>"010111111",
  35389=>"110000100",
  35390=>"101000011",
  35391=>"100000010",
  35392=>"011111011",
  35393=>"100101011",
  35394=>"111111110",
  35395=>"100101100",
  35396=>"000010111",
  35397=>"000010101",
  35398=>"101010010",
  35399=>"111010000",
  35400=>"110001011",
  35401=>"110010110",
  35402=>"000111011",
  35403=>"001011100",
  35404=>"111001110",
  35405=>"100000010",
  35406=>"000100110",
  35407=>"100111100",
  35408=>"011001110",
  35409=>"010000111",
  35410=>"110101001",
  35411=>"011001111",
  35412=>"100100010",
  35413=>"100000100",
  35414=>"001010110",
  35415=>"010000111",
  35416=>"000111010",
  35417=>"001111011",
  35418=>"110111001",
  35419=>"011101001",
  35420=>"000010101",
  35421=>"110001000",
  35422=>"001111011",
  35423=>"111100101",
  35424=>"100011111",
  35425=>"001110000",
  35426=>"001011011",
  35427=>"000010000",
  35428=>"111100110",
  35429=>"100000110",
  35430=>"111011111",
  35431=>"110110110",
  35432=>"000010011",
  35433=>"110101111",
  35434=>"001001000",
  35435=>"011011000",
  35436=>"110101010",
  35437=>"000110111",
  35438=>"011001001",
  35439=>"011111111",
  35440=>"111000001",
  35441=>"000110100",
  35442=>"011111101",
  35443=>"100100110",
  35444=>"100001110",
  35445=>"111010101",
  35446=>"110010111",
  35447=>"100110000",
  35448=>"100011000",
  35449=>"001111011",
  35450=>"000101010",
  35451=>"001111001",
  35452=>"101001000",
  35453=>"000111011",
  35454=>"111001011",
  35455=>"111110101",
  35456=>"101010000",
  35457=>"001001001",
  35458=>"010100101",
  35459=>"011100111",
  35460=>"101110100",
  35461=>"000001000",
  35462=>"000100111",
  35463=>"110111010",
  35464=>"010000111",
  35465=>"110110011",
  35466=>"010111000",
  35467=>"100110111",
  35468=>"010011111",
  35469=>"111010110",
  35470=>"010101000",
  35471=>"100001011",
  35472=>"100011001",
  35473=>"110110011",
  35474=>"111101110",
  35475=>"101110000",
  35476=>"100011101",
  35477=>"010100101",
  35478=>"100110111",
  35479=>"110110000",
  35480=>"000100000",
  35481=>"010100110",
  35482=>"011001000",
  35483=>"000000101",
  35484=>"111011011",
  35485=>"001000000",
  35486=>"111010101",
  35487=>"001110110",
  35488=>"001010110",
  35489=>"101000100",
  35490=>"111000000",
  35491=>"010001000",
  35492=>"010100110",
  35493=>"001001111",
  35494=>"011101011",
  35495=>"100000011",
  35496=>"111111100",
  35497=>"011101000",
  35498=>"001001000",
  35499=>"110111000",
  35500=>"010010000",
  35501=>"001000011",
  35502=>"101011011",
  35503=>"110111001",
  35504=>"010011001",
  35505=>"001100100",
  35506=>"101110110",
  35507=>"010001101",
  35508=>"001001101",
  35509=>"101011101",
  35510=>"010011011",
  35511=>"000100101",
  35512=>"100000000",
  35513=>"011111000",
  35514=>"101110010",
  35515=>"001010000",
  35516=>"101111111",
  35517=>"011110010",
  35518=>"011100100",
  35519=>"101010111",
  35520=>"111011100",
  35521=>"010001111",
  35522=>"000000000",
  35523=>"000001101",
  35524=>"000101101",
  35525=>"000010010",
  35526=>"101001101",
  35527=>"001001011",
  35528=>"010010100",
  35529=>"100000000",
  35530=>"111001100",
  35531=>"011010000",
  35532=>"010011010",
  35533=>"001111001",
  35534=>"110101111",
  35535=>"011011110",
  35536=>"100100010",
  35537=>"111110101",
  35538=>"001000100",
  35539=>"100110010",
  35540=>"100000111",
  35541=>"000010010",
  35542=>"111100001",
  35543=>"011101111",
  35544=>"011101111",
  35545=>"010111000",
  35546=>"011010101",
  35547=>"111010010",
  35548=>"000100111",
  35549=>"100001100",
  35550=>"001110101",
  35551=>"000000111",
  35552=>"111101111",
  35553=>"100000101",
  35554=>"001100100",
  35555=>"011110001",
  35556=>"001100001",
  35557=>"101001011",
  35558=>"010011011",
  35559=>"100100001",
  35560=>"001111101",
  35561=>"011011001",
  35562=>"001101110",
  35563=>"010000000",
  35564=>"110101101",
  35565=>"100001101",
  35566=>"111110001",
  35567=>"100101001",
  35568=>"101010111",
  35569=>"111000100",
  35570=>"010011111",
  35571=>"000100110",
  35572=>"010101000",
  35573=>"111101110",
  35574=>"111100101",
  35575=>"010010111",
  35576=>"101111110",
  35577=>"111101111",
  35578=>"111101001",
  35579=>"000011111",
  35580=>"110010110",
  35581=>"110101110",
  35582=>"111001100",
  35583=>"100001001",
  35584=>"101110010",
  35585=>"000010100",
  35586=>"011110010",
  35587=>"100000010",
  35588=>"001101101",
  35589=>"011001000",
  35590=>"000101111",
  35591=>"011101111",
  35592=>"100000010",
  35593=>"101010001",
  35594=>"110000000",
  35595=>"101100111",
  35596=>"101001101",
  35597=>"011111101",
  35598=>"000001001",
  35599=>"010010100",
  35600=>"101001010",
  35601=>"111111100",
  35602=>"010000100",
  35603=>"100011001",
  35604=>"101000110",
  35605=>"111000010",
  35606=>"111011111",
  35607=>"000101101",
  35608=>"000100000",
  35609=>"100001110",
  35610=>"000011111",
  35611=>"000101111",
  35612=>"101100000",
  35613=>"001110111",
  35614=>"100101000",
  35615=>"110100000",
  35616=>"001001110",
  35617=>"010111001",
  35618=>"000011011",
  35619=>"011111100",
  35620=>"010101100",
  35621=>"011011011",
  35622=>"111011001",
  35623=>"001001000",
  35624=>"010101000",
  35625=>"111001010",
  35626=>"011001000",
  35627=>"110000010",
  35628=>"111000011",
  35629=>"010010010",
  35630=>"111111011",
  35631=>"000000000",
  35632=>"010011000",
  35633=>"100000101",
  35634=>"001000110",
  35635=>"101011110",
  35636=>"000111011",
  35637=>"111100011",
  35638=>"001101110",
  35639=>"001011111",
  35640=>"000110101",
  35641=>"011100101",
  35642=>"010111101",
  35643=>"011110011",
  35644=>"110111010",
  35645=>"000111001",
  35646=>"011011111",
  35647=>"100100110",
  35648=>"100010000",
  35649=>"011010010",
  35650=>"110011101",
  35651=>"100001000",
  35652=>"001011011",
  35653=>"111001010",
  35654=>"100001101",
  35655=>"111011000",
  35656=>"100101000",
  35657=>"101100000",
  35658=>"001111101",
  35659=>"001101111",
  35660=>"100011111",
  35661=>"010001001",
  35662=>"111111011",
  35663=>"101001101",
  35664=>"000001011",
  35665=>"111110010",
  35666=>"011010111",
  35667=>"001010010",
  35668=>"101101111",
  35669=>"010010010",
  35670=>"010101100",
  35671=>"111101100",
  35672=>"111111001",
  35673=>"101100101",
  35674=>"111100011",
  35675=>"001001001",
  35676=>"001111000",
  35677=>"000010011",
  35678=>"100001011",
  35679=>"001100001",
  35680=>"010011001",
  35681=>"011010001",
  35682=>"101101100",
  35683=>"110100111",
  35684=>"110100101",
  35685=>"101100111",
  35686=>"100100110",
  35687=>"110111011",
  35688=>"011000110",
  35689=>"010001010",
  35690=>"010110101",
  35691=>"000010011",
  35692=>"010111000",
  35693=>"110011100",
  35694=>"111100000",
  35695=>"111010110",
  35696=>"110101110",
  35697=>"111011000",
  35698=>"011000010",
  35699=>"101101000",
  35700=>"010111010",
  35701=>"000001010",
  35702=>"010111101",
  35703=>"111111001",
  35704=>"111101111",
  35705=>"011001000",
  35706=>"100100101",
  35707=>"000101111",
  35708=>"100010000",
  35709=>"000000110",
  35710=>"111101100",
  35711=>"100100010",
  35712=>"000001101",
  35713=>"001011111",
  35714=>"001100110",
  35715=>"010110001",
  35716=>"100100110",
  35717=>"011110001",
  35718=>"000110110",
  35719=>"011011000",
  35720=>"110000011",
  35721=>"000011000",
  35722=>"011100010",
  35723=>"010110110",
  35724=>"110100101",
  35725=>"000100110",
  35726=>"011011111",
  35727=>"101000111",
  35728=>"110100110",
  35729=>"101001001",
  35730=>"000100001",
  35731=>"111010011",
  35732=>"010110111",
  35733=>"101001001",
  35734=>"101111011",
  35735=>"101010101",
  35736=>"011001100",
  35737=>"010101110",
  35738=>"000010101",
  35739=>"010101100",
  35740=>"000111011",
  35741=>"101010101",
  35742=>"110100110",
  35743=>"111100000",
  35744=>"101101101",
  35745=>"111111111",
  35746=>"001100100",
  35747=>"000001101",
  35748=>"110000101",
  35749=>"111001110",
  35750=>"110011000",
  35751=>"010111110",
  35752=>"110100000",
  35753=>"010011011",
  35754=>"001011010",
  35755=>"000001101",
  35756=>"100010001",
  35757=>"001100101",
  35758=>"010010101",
  35759=>"000001000",
  35760=>"010101100",
  35761=>"011101011",
  35762=>"100110110",
  35763=>"011000101",
  35764=>"111100110",
  35765=>"000111100",
  35766=>"111011110",
  35767=>"110000000",
  35768=>"110110011",
  35769=>"011110110",
  35770=>"100101110",
  35771=>"110000000",
  35772=>"001110100",
  35773=>"001011100",
  35774=>"101001001",
  35775=>"000010000",
  35776=>"001111100",
  35777=>"111110110",
  35778=>"000111110",
  35779=>"000011110",
  35780=>"101000010",
  35781=>"001000101",
  35782=>"010001000",
  35783=>"100011100",
  35784=>"001110101",
  35785=>"111001111",
  35786=>"010011101",
  35787=>"011000010",
  35788=>"110100011",
  35789=>"000110011",
  35790=>"101011000",
  35791=>"010111000",
  35792=>"000010111",
  35793=>"111010011",
  35794=>"001011000",
  35795=>"100101000",
  35796=>"100111001",
  35797=>"000001110",
  35798=>"111011111",
  35799=>"000110101",
  35800=>"001000101",
  35801=>"010010110",
  35802=>"100001000",
  35803=>"101111010",
  35804=>"000010011",
  35805=>"111111110",
  35806=>"001111001",
  35807=>"000111111",
  35808=>"111110100",
  35809=>"011100111",
  35810=>"001111000",
  35811=>"001001110",
  35812=>"010001001",
  35813=>"111000000",
  35814=>"001010010",
  35815=>"010001010",
  35816=>"100101110",
  35817=>"010011100",
  35818=>"010000101",
  35819=>"100100101",
  35820=>"110010111",
  35821=>"101010010",
  35822=>"110011001",
  35823=>"101101100",
  35824=>"110111010",
  35825=>"100010101",
  35826=>"110100111",
  35827=>"011110100",
  35828=>"010110000",
  35829=>"000111110",
  35830=>"000111101",
  35831=>"000000010",
  35832=>"100100000",
  35833=>"001010001",
  35834=>"000000010",
  35835=>"101011110",
  35836=>"000101111",
  35837=>"100111100",
  35838=>"111110110",
  35839=>"001000101",
  35840=>"101100100",
  35841=>"010101000",
  35842=>"111110101",
  35843=>"001100111",
  35844=>"101111010",
  35845=>"010010010",
  35846=>"001101001",
  35847=>"100000111",
  35848=>"110110011",
  35849=>"100101001",
  35850=>"111100000",
  35851=>"111000110",
  35852=>"100110001",
  35853=>"111010001",
  35854=>"110001001",
  35855=>"001000011",
  35856=>"010010101",
  35857=>"010100000",
  35858=>"100000000",
  35859=>"010110011",
  35860=>"011000001",
  35861=>"100010000",
  35862=>"100001001",
  35863=>"101011011",
  35864=>"111101101",
  35865=>"111110000",
  35866=>"000101110",
  35867=>"001111111",
  35868=>"100010010",
  35869=>"000001101",
  35870=>"100001100",
  35871=>"110000110",
  35872=>"110111011",
  35873=>"100110011",
  35874=>"100010101",
  35875=>"101110111",
  35876=>"000000100",
  35877=>"011101010",
  35878=>"000110011",
  35879=>"010101011",
  35880=>"101100101",
  35881=>"000001010",
  35882=>"000010011",
  35883=>"110100101",
  35884=>"011001100",
  35885=>"010000101",
  35886=>"101001000",
  35887=>"100000110",
  35888=>"101011011",
  35889=>"000001111",
  35890=>"010011110",
  35891=>"011101111",
  35892=>"011011010",
  35893=>"101111101",
  35894=>"100101010",
  35895=>"001111010",
  35896=>"001011010",
  35897=>"011101101",
  35898=>"111000011",
  35899=>"101111111",
  35900=>"010001011",
  35901=>"111000000",
  35902=>"010001001",
  35903=>"010101010",
  35904=>"011001111",
  35905=>"100011110",
  35906=>"010111111",
  35907=>"000100101",
  35908=>"111011110",
  35909=>"001101011",
  35910=>"001111010",
  35911=>"000000100",
  35912=>"011100000",
  35913=>"100110011",
  35914=>"100000101",
  35915=>"111101110",
  35916=>"110011000",
  35917=>"101100010",
  35918=>"101110111",
  35919=>"011110111",
  35920=>"010000001",
  35921=>"100110000",
  35922=>"100101000",
  35923=>"010001110",
  35924=>"010111000",
  35925=>"011111100",
  35926=>"110000010",
  35927=>"001101001",
  35928=>"111011110",
  35929=>"001101101",
  35930=>"100010111",
  35931=>"111010100",
  35932=>"111000100",
  35933=>"000100100",
  35934=>"000110101",
  35935=>"100011110",
  35936=>"011011001",
  35937=>"101101001",
  35938=>"010110111",
  35939=>"111010111",
  35940=>"000101100",
  35941=>"000000001",
  35942=>"101010000",
  35943=>"010101111",
  35944=>"101110001",
  35945=>"011001011",
  35946=>"111101111",
  35947=>"001110000",
  35948=>"111110001",
  35949=>"000110101",
  35950=>"100011011",
  35951=>"110111001",
  35952=>"111110011",
  35953=>"000111100",
  35954=>"001011011",
  35955=>"010001001",
  35956=>"001100101",
  35957=>"001100100",
  35958=>"111000101",
  35959=>"000100111",
  35960=>"110100101",
  35961=>"100110000",
  35962=>"100110111",
  35963=>"001011001",
  35964=>"110000101",
  35965=>"111100101",
  35966=>"011110001",
  35967=>"111011101",
  35968=>"111010011",
  35969=>"101011001",
  35970=>"001010011",
  35971=>"000111101",
  35972=>"110101110",
  35973=>"000110100",
  35974=>"101110101",
  35975=>"000101101",
  35976=>"000011000",
  35977=>"101111100",
  35978=>"111110101",
  35979=>"011000000",
  35980=>"011101000",
  35981=>"101010111",
  35982=>"011111110",
  35983=>"100101110",
  35984=>"000001100",
  35985=>"000001100",
  35986=>"100110011",
  35987=>"101011101",
  35988=>"110101000",
  35989=>"101000000",
  35990=>"101100100",
  35991=>"000000000",
  35992=>"010101111",
  35993=>"111110110",
  35994=>"001001100",
  35995=>"001100110",
  35996=>"011101100",
  35997=>"101101111",
  35998=>"001111001",
  35999=>"100000101",
  36000=>"111001000",
  36001=>"010001011",
  36002=>"000010111",
  36003=>"110100111",
  36004=>"010110101",
  36005=>"101111111",
  36006=>"001010000",
  36007=>"101011000",
  36008=>"100011110",
  36009=>"011110100",
  36010=>"110000111",
  36011=>"101111000",
  36012=>"111001101",
  36013=>"011110011",
  36014=>"110101011",
  36015=>"101001101",
  36016=>"011011100",
  36017=>"111000001",
  36018=>"111101100",
  36019=>"101000110",
  36020=>"111100101",
  36021=>"010011101",
  36022=>"101111011",
  36023=>"110100010",
  36024=>"011011111",
  36025=>"001000101",
  36026=>"111000101",
  36027=>"011000010",
  36028=>"101010011",
  36029=>"000101010",
  36030=>"111010010",
  36031=>"011000011",
  36032=>"010001111",
  36033=>"001101001",
  36034=>"110011000",
  36035=>"000110110",
  36036=>"110111011",
  36037=>"000111101",
  36038=>"101001010",
  36039=>"111100011",
  36040=>"111011111",
  36041=>"111011110",
  36042=>"100011111",
  36043=>"100110000",
  36044=>"001111010",
  36045=>"011110100",
  36046=>"011010111",
  36047=>"111110110",
  36048=>"000010001",
  36049=>"011001001",
  36050=>"010000010",
  36051=>"001010111",
  36052=>"101001011",
  36053=>"110111101",
  36054=>"010110001",
  36055=>"001101101",
  36056=>"110010000",
  36057=>"000001110",
  36058=>"100110010",
  36059=>"101010111",
  36060=>"111111000",
  36061=>"100001100",
  36062=>"111100111",
  36063=>"010000100",
  36064=>"111100010",
  36065=>"010110011",
  36066=>"000011110",
  36067=>"011101000",
  36068=>"110100011",
  36069=>"101011101",
  36070=>"101001001",
  36071=>"001100100",
  36072=>"110111001",
  36073=>"011001100",
  36074=>"110001010",
  36075=>"100010111",
  36076=>"011101100",
  36077=>"111010100",
  36078=>"110100001",
  36079=>"111100101",
  36080=>"011011001",
  36081=>"111101011",
  36082=>"000111100",
  36083=>"010000010",
  36084=>"100111111",
  36085=>"000100000",
  36086=>"001001001",
  36087=>"011011000",
  36088=>"011100001",
  36089=>"100000001",
  36090=>"100101000",
  36091=>"001111001",
  36092=>"101000111",
  36093=>"101000010",
  36094=>"101001100",
  36095=>"000110100",
  36096=>"110001101",
  36097=>"011111110",
  36098=>"100101110",
  36099=>"000101111",
  36100=>"000011001",
  36101=>"010001110",
  36102=>"011111011",
  36103=>"110101000",
  36104=>"111110000",
  36105=>"100111001",
  36106=>"001000110",
  36107=>"010010101",
  36108=>"000010001",
  36109=>"001001101",
  36110=>"011101000",
  36111=>"011011011",
  36112=>"101101011",
  36113=>"110010000",
  36114=>"011111000",
  36115=>"110010101",
  36116=>"111010111",
  36117=>"110010110",
  36118=>"100111000",
  36119=>"000001001",
  36120=>"010011101",
  36121=>"001001001",
  36122=>"101011001",
  36123=>"011110000",
  36124=>"100110111",
  36125=>"110010110",
  36126=>"110111011",
  36127=>"111110000",
  36128=>"111001100",
  36129=>"101001010",
  36130=>"100011011",
  36131=>"110110111",
  36132=>"011000011",
  36133=>"111011010",
  36134=>"011101100",
  36135=>"111001010",
  36136=>"111001100",
  36137=>"001111000",
  36138=>"100110100",
  36139=>"110101101",
  36140=>"010011100",
  36141=>"101101001",
  36142=>"001110100",
  36143=>"110010101",
  36144=>"000110111",
  36145=>"011101000",
  36146=>"101111100",
  36147=>"111101111",
  36148=>"010110010",
  36149=>"010000010",
  36150=>"110111101",
  36151=>"010111011",
  36152=>"000110001",
  36153=>"100111011",
  36154=>"001100000",
  36155=>"000000101",
  36156=>"100100101",
  36157=>"001101001",
  36158=>"100111010",
  36159=>"100111111",
  36160=>"111101000",
  36161=>"011101111",
  36162=>"001011101",
  36163=>"110011010",
  36164=>"001011100",
  36165=>"010010111",
  36166=>"000100111",
  36167=>"100101000",
  36168=>"100000011",
  36169=>"101100101",
  36170=>"111111101",
  36171=>"110110011",
  36172=>"000001010",
  36173=>"000000111",
  36174=>"011001111",
  36175=>"101111010",
  36176=>"101100010",
  36177=>"001100100",
  36178=>"110000101",
  36179=>"101101000",
  36180=>"101100110",
  36181=>"011001000",
  36182=>"100011001",
  36183=>"110000010",
  36184=>"011110111",
  36185=>"001001110",
  36186=>"111011010",
  36187=>"110011110",
  36188=>"101100000",
  36189=>"001100111",
  36190=>"001110000",
  36191=>"100111101",
  36192=>"000001000",
  36193=>"110101001",
  36194=>"001101011",
  36195=>"000011101",
  36196=>"010001101",
  36197=>"000100010",
  36198=>"000000100",
  36199=>"011110101",
  36200=>"111110100",
  36201=>"010000100",
  36202=>"010010111",
  36203=>"111111110",
  36204=>"111011001",
  36205=>"101100000",
  36206=>"001001011",
  36207=>"001000100",
  36208=>"010001101",
  36209=>"100111111",
  36210=>"000011011",
  36211=>"111101000",
  36212=>"000011101",
  36213=>"011001100",
  36214=>"000000101",
  36215=>"111110010",
  36216=>"100011111",
  36217=>"111000000",
  36218=>"100011100",
  36219=>"000000110",
  36220=>"010111000",
  36221=>"010000000",
  36222=>"001010011",
  36223=>"100111001",
  36224=>"010001010",
  36225=>"101101110",
  36226=>"100110110",
  36227=>"011001001",
  36228=>"011001100",
  36229=>"111011111",
  36230=>"110100010",
  36231=>"101010000",
  36232=>"101010111",
  36233=>"101001000",
  36234=>"110111010",
  36235=>"000110010",
  36236=>"110101101",
  36237=>"000010001",
  36238=>"100000110",
  36239=>"110010010",
  36240=>"101110110",
  36241=>"100101100",
  36242=>"011000110",
  36243=>"010111110",
  36244=>"110101111",
  36245=>"000111101",
  36246=>"000000010",
  36247=>"001000001",
  36248=>"110001100",
  36249=>"001011100",
  36250=>"111111110",
  36251=>"001110101",
  36252=>"111000101",
  36253=>"111100000",
  36254=>"101001111",
  36255=>"111110111",
  36256=>"001101101",
  36257=>"111101101",
  36258=>"111011001",
  36259=>"101100011",
  36260=>"111100101",
  36261=>"000010101",
  36262=>"011000110",
  36263=>"110101010",
  36264=>"111001001",
  36265=>"000001011",
  36266=>"000101101",
  36267=>"110101101",
  36268=>"001011010",
  36269=>"111111100",
  36270=>"001110100",
  36271=>"111011001",
  36272=>"000001011",
  36273=>"010010101",
  36274=>"001010010",
  36275=>"011101100",
  36276=>"110101110",
  36277=>"001100101",
  36278=>"000000110",
  36279=>"110111000",
  36280=>"101111001",
  36281=>"010000110",
  36282=>"001101100",
  36283=>"100000111",
  36284=>"110100110",
  36285=>"001100101",
  36286=>"011001100",
  36287=>"001011000",
  36288=>"111110011",
  36289=>"100111111",
  36290=>"011101010",
  36291=>"000111001",
  36292=>"000001100",
  36293=>"010101100",
  36294=>"010111000",
  36295=>"111110000",
  36296=>"011101110",
  36297=>"100100001",
  36298=>"000011110",
  36299=>"110000010",
  36300=>"000100001",
  36301=>"000111001",
  36302=>"110010110",
  36303=>"110000111",
  36304=>"110111011",
  36305=>"000100101",
  36306=>"111011001",
  36307=>"111110111",
  36308=>"010110001",
  36309=>"111001001",
  36310=>"111000001",
  36311=>"110000111",
  36312=>"001111101",
  36313=>"000111100",
  36314=>"101110111",
  36315=>"100111000",
  36316=>"100110011",
  36317=>"000010100",
  36318=>"000000101",
  36319=>"000011101",
  36320=>"110101110",
  36321=>"011000011",
  36322=>"111110111",
  36323=>"000001111",
  36324=>"010110000",
  36325=>"101110001",
  36326=>"111110000",
  36327=>"100001100",
  36328=>"011111111",
  36329=>"111110010",
  36330=>"110011001",
  36331=>"011111101",
  36332=>"000000000",
  36333=>"101110000",
  36334=>"100110110",
  36335=>"111101010",
  36336=>"101110100",
  36337=>"000001000",
  36338=>"110101010",
  36339=>"000011011",
  36340=>"000011111",
  36341=>"011101011",
  36342=>"101001001",
  36343=>"001010001",
  36344=>"011100110",
  36345=>"100110001",
  36346=>"000111010",
  36347=>"001100101",
  36348=>"000111011",
  36349=>"010111000",
  36350=>"010111111",
  36351=>"001011111",
  36352=>"010100001",
  36353=>"010011011",
  36354=>"111101001",
  36355=>"010000011",
  36356=>"101001011",
  36357=>"100010100",
  36358=>"100010110",
  36359=>"101010010",
  36360=>"010110000",
  36361=>"010101101",
  36362=>"100101110",
  36363=>"001101111",
  36364=>"110101011",
  36365=>"101001001",
  36366=>"111110000",
  36367=>"110010111",
  36368=>"001000101",
  36369=>"011011011",
  36370=>"101011101",
  36371=>"000100111",
  36372=>"111001100",
  36373=>"111010100",
  36374=>"111001110",
  36375=>"110010010",
  36376=>"111001000",
  36377=>"001100001",
  36378=>"101010001",
  36379=>"101000110",
  36380=>"111001110",
  36381=>"111111001",
  36382=>"000101100",
  36383=>"001011111",
  36384=>"101101011",
  36385=>"011110010",
  36386=>"001011000",
  36387=>"101111110",
  36388=>"001100010",
  36389=>"001000110",
  36390=>"010110010",
  36391=>"000000010",
  36392=>"010000001",
  36393=>"110100000",
  36394=>"110010001",
  36395=>"000100010",
  36396=>"101011111",
  36397=>"100101001",
  36398=>"000111000",
  36399=>"011100101",
  36400=>"010001001",
  36401=>"110011010",
  36402=>"000001011",
  36403=>"000001000",
  36404=>"100101101",
  36405=>"111011001",
  36406=>"001111010",
  36407=>"010111000",
  36408=>"000111011",
  36409=>"101000101",
  36410=>"100110011",
  36411=>"000011000",
  36412=>"000110101",
  36413=>"010011101",
  36414=>"000100011",
  36415=>"111110001",
  36416=>"111001100",
  36417=>"100001101",
  36418=>"011111110",
  36419=>"011100101",
  36420=>"100110000",
  36421=>"111001111",
  36422=>"111010111",
  36423=>"110001001",
  36424=>"001101011",
  36425=>"111010110",
  36426=>"010011010",
  36427=>"100101001",
  36428=>"011100011",
  36429=>"010101101",
  36430=>"111100101",
  36431=>"110110110",
  36432=>"000011011",
  36433=>"101010101",
  36434=>"101110110",
  36435=>"110001000",
  36436=>"001100111",
  36437=>"000000010",
  36438=>"110111111",
  36439=>"100101001",
  36440=>"110100100",
  36441=>"010010100",
  36442=>"101111111",
  36443=>"001101111",
  36444=>"000010111",
  36445=>"110000111",
  36446=>"101101000",
  36447=>"110100100",
  36448=>"000011011",
  36449=>"100100011",
  36450=>"001010111",
  36451=>"010010011",
  36452=>"001110000",
  36453=>"000000110",
  36454=>"101100101",
  36455=>"011011110",
  36456=>"111111001",
  36457=>"001001111",
  36458=>"010111011",
  36459=>"100000101",
  36460=>"101110010",
  36461=>"110111111",
  36462=>"100001000",
  36463=>"111011000",
  36464=>"000101111",
  36465=>"101001100",
  36466=>"100101000",
  36467=>"111011111",
  36468=>"001010010",
  36469=>"011001000",
  36470=>"111111010",
  36471=>"001011111",
  36472=>"111010101",
  36473=>"101100110",
  36474=>"101011111",
  36475=>"100000100",
  36476=>"100011011",
  36477=>"000001001",
  36478=>"000101001",
  36479=>"010110100",
  36480=>"100001000",
  36481=>"001011110",
  36482=>"010001100",
  36483=>"010010111",
  36484=>"101110100",
  36485=>"100011110",
  36486=>"000010011",
  36487=>"000000001",
  36488=>"110000011",
  36489=>"000010110",
  36490=>"001110111",
  36491=>"001110100",
  36492=>"001100111",
  36493=>"001011000",
  36494=>"100100010",
  36495=>"010111001",
  36496=>"010011001",
  36497=>"101011001",
  36498=>"101110010",
  36499=>"101110000",
  36500=>"000001001",
  36501=>"101010101",
  36502=>"010001100",
  36503=>"001101011",
  36504=>"001110001",
  36505=>"010111001",
  36506=>"000110001",
  36507=>"100101110",
  36508=>"111000000",
  36509=>"100100101",
  36510=>"001100010",
  36511=>"110001000",
  36512=>"010101100",
  36513=>"001011001",
  36514=>"011000111",
  36515=>"111101000",
  36516=>"101000100",
  36517=>"000010011",
  36518=>"000110111",
  36519=>"000110111",
  36520=>"001010100",
  36521=>"010100000",
  36522=>"001001001",
  36523=>"110110110",
  36524=>"011111000",
  36525=>"110000111",
  36526=>"111000101",
  36527=>"111010100",
  36528=>"111110111",
  36529=>"011101010",
  36530=>"111000001",
  36531=>"100101000",
  36532=>"100101100",
  36533=>"100011100",
  36534=>"101111010",
  36535=>"001110110",
  36536=>"110101010",
  36537=>"101001101",
  36538=>"100101111",
  36539=>"100001110",
  36540=>"000111001",
  36541=>"011011110",
  36542=>"111010010",
  36543=>"000010001",
  36544=>"111101000",
  36545=>"111110011",
  36546=>"111010100",
  36547=>"011100000",
  36548=>"111101010",
  36549=>"001011001",
  36550=>"111110010",
  36551=>"100000110",
  36552=>"111111101",
  36553=>"001111001",
  36554=>"010101001",
  36555=>"101110111",
  36556=>"000110100",
  36557=>"011100100",
  36558=>"010001010",
  36559=>"001000001",
  36560=>"110101011",
  36561=>"001100100",
  36562=>"111111010",
  36563=>"010000000",
  36564=>"100111101",
  36565=>"101010101",
  36566=>"011010010",
  36567=>"000101110",
  36568=>"111000101",
  36569=>"011000100",
  36570=>"110000100",
  36571=>"010000100",
  36572=>"101111011",
  36573=>"101101110",
  36574=>"100110001",
  36575=>"100101010",
  36576=>"100010011",
  36577=>"010001100",
  36578=>"010100010",
  36579=>"100000000",
  36580=>"001111010",
  36581=>"111010110",
  36582=>"110011001",
  36583=>"100100001",
  36584=>"011011100",
  36585=>"101011010",
  36586=>"111110110",
  36587=>"001000111",
  36588=>"000010110",
  36589=>"000001111",
  36590=>"100000010",
  36591=>"111011010",
  36592=>"111101111",
  36593=>"011101101",
  36594=>"110001001",
  36595=>"101010001",
  36596=>"101100110",
  36597=>"001111011",
  36598=>"011111001",
  36599=>"101001001",
  36600=>"011100110",
  36601=>"000101010",
  36602=>"011111111",
  36603=>"010000100",
  36604=>"011110100",
  36605=>"000111000",
  36606=>"010000101",
  36607=>"100100011",
  36608=>"100011000",
  36609=>"111010101",
  36610=>"111000100",
  36611=>"000010011",
  36612=>"010011000",
  36613=>"111111010",
  36614=>"000101111",
  36615=>"010110000",
  36616=>"100001110",
  36617=>"101110101",
  36618=>"000100001",
  36619=>"100101110",
  36620=>"001110001",
  36621=>"100011110",
  36622=>"111000000",
  36623=>"011000010",
  36624=>"000000110",
  36625=>"101011100",
  36626=>"011111001",
  36627=>"000011101",
  36628=>"100101100",
  36629=>"001100011",
  36630=>"101110001",
  36631=>"100110011",
  36632=>"101011111",
  36633=>"010100001",
  36634=>"001000111",
  36635=>"001110111",
  36636=>"110100111",
  36637=>"001111111",
  36638=>"101111011",
  36639=>"001100010",
  36640=>"010110000",
  36641=>"010001000",
  36642=>"100110011",
  36643=>"100010000",
  36644=>"111010111",
  36645=>"111010001",
  36646=>"100101101",
  36647=>"001001100",
  36648=>"000100101",
  36649=>"111001111",
  36650=>"101010110",
  36651=>"110111010",
  36652=>"000011001",
  36653=>"111011110",
  36654=>"101101010",
  36655=>"100010010",
  36656=>"010101001",
  36657=>"101010000",
  36658=>"100100111",
  36659=>"110110010",
  36660=>"111101011",
  36661=>"001101110",
  36662=>"100111111",
  36663=>"100001111",
  36664=>"000000101",
  36665=>"010000000",
  36666=>"001110110",
  36667=>"111000011",
  36668=>"111111111",
  36669=>"111011011",
  36670=>"011001011",
  36671=>"000010000",
  36672=>"001000000",
  36673=>"000101110",
  36674=>"110000000",
  36675=>"000111001",
  36676=>"001011110",
  36677=>"001111101",
  36678=>"010011100",
  36679=>"000101110",
  36680=>"001110000",
  36681=>"000001000",
  36682=>"011111110",
  36683=>"001100001",
  36684=>"111110100",
  36685=>"010010010",
  36686=>"111111010",
  36687=>"011000011",
  36688=>"001010000",
  36689=>"100110100",
  36690=>"110001010",
  36691=>"110010000",
  36692=>"011111110",
  36693=>"100010010",
  36694=>"000001111",
  36695=>"011111101",
  36696=>"010010100",
  36697=>"110011001",
  36698=>"010100100",
  36699=>"010010111",
  36700=>"000001011",
  36701=>"000110010",
  36702=>"001000111",
  36703=>"100100101",
  36704=>"110001011",
  36705=>"101000001",
  36706=>"000101111",
  36707=>"011001010",
  36708=>"101101010",
  36709=>"101001111",
  36710=>"111101101",
  36711=>"111111100",
  36712=>"111101110",
  36713=>"100110011",
  36714=>"111110000",
  36715=>"100011010",
  36716=>"101111001",
  36717=>"001000111",
  36718=>"010010110",
  36719=>"101111011",
  36720=>"011110100",
  36721=>"101111110",
  36722=>"110101101",
  36723=>"000110001",
  36724=>"100111010",
  36725=>"101011110",
  36726=>"110000011",
  36727=>"000010100",
  36728=>"011011011",
  36729=>"110100000",
  36730=>"001010101",
  36731=>"011100001",
  36732=>"111011000",
  36733=>"100111101",
  36734=>"111011001",
  36735=>"001110001",
  36736=>"000011010",
  36737=>"000001011",
  36738=>"101110010",
  36739=>"111110110",
  36740=>"001100100",
  36741=>"110011001",
  36742=>"001001100",
  36743=>"000010000",
  36744=>"001101110",
  36745=>"000000111",
  36746=>"110110110",
  36747=>"011001011",
  36748=>"011101001",
  36749=>"001110010",
  36750=>"011111101",
  36751=>"101100001",
  36752=>"101110101",
  36753=>"100100100",
  36754=>"111000000",
  36755=>"111111000",
  36756=>"011011001",
  36757=>"101011101",
  36758=>"001101111",
  36759=>"101111010",
  36760=>"111011110",
  36761=>"111010000",
  36762=>"000110000",
  36763=>"100010111",
  36764=>"001100010",
  36765=>"011111100",
  36766=>"111010011",
  36767=>"111111001",
  36768=>"111100011",
  36769=>"010000001",
  36770=>"010001001",
  36771=>"110110111",
  36772=>"000001111",
  36773=>"011011010",
  36774=>"001101010",
  36775=>"010111111",
  36776=>"000000001",
  36777=>"101010100",
  36778=>"001111000",
  36779=>"010000101",
  36780=>"011001110",
  36781=>"011010001",
  36782=>"100100110",
  36783=>"001100101",
  36784=>"000000100",
  36785=>"110101101",
  36786=>"100011001",
  36787=>"000000011",
  36788=>"110101000",
  36789=>"010011100",
  36790=>"000101011",
  36791=>"010001000",
  36792=>"000000100",
  36793=>"010110011",
  36794=>"111000101",
  36795=>"111000000",
  36796=>"001101111",
  36797=>"011010101",
  36798=>"000101111",
  36799=>"100001101",
  36800=>"111100100",
  36801=>"010101110",
  36802=>"100001100",
  36803=>"110011100",
  36804=>"100100000",
  36805=>"110011001",
  36806=>"100101011",
  36807=>"001001000",
  36808=>"111100011",
  36809=>"110110001",
  36810=>"100001010",
  36811=>"101010001",
  36812=>"110001010",
  36813=>"100001010",
  36814=>"110110111",
  36815=>"000101100",
  36816=>"000010011",
  36817=>"111011111",
  36818=>"100011000",
  36819=>"110100010",
  36820=>"000001001",
  36821=>"100011011",
  36822=>"011001100",
  36823=>"011110100",
  36824=>"000011101",
  36825=>"100001100",
  36826=>"111101111",
  36827=>"111101001",
  36828=>"100000001",
  36829=>"000110000",
  36830=>"010000010",
  36831=>"100010100",
  36832=>"011011111",
  36833=>"100000011",
  36834=>"111011000",
  36835=>"111000101",
  36836=>"011101001",
  36837=>"011100001",
  36838=>"110000100",
  36839=>"100101101",
  36840=>"000001100",
  36841=>"110110010",
  36842=>"001011000",
  36843=>"000010001",
  36844=>"010111110",
  36845=>"011011011",
  36846=>"000011001",
  36847=>"111101110",
  36848=>"000111011",
  36849=>"001101100",
  36850=>"000010101",
  36851=>"110110101",
  36852=>"111010100",
  36853=>"001011110",
  36854=>"010101111",
  36855=>"010101100",
  36856=>"101010111",
  36857=>"001101101",
  36858=>"111110111",
  36859=>"110100111",
  36860=>"101111000",
  36861=>"111111001",
  36862=>"010001100",
  36863=>"011101011",
  36864=>"001101110",
  36865=>"010000111",
  36866=>"101101001",
  36867=>"011111011",
  36868=>"101100111",
  36869=>"101011011",
  36870=>"111100010",
  36871=>"011011100",
  36872=>"001011101",
  36873=>"000110000",
  36874=>"110110101",
  36875=>"011001001",
  36876=>"110000100",
  36877=>"011010001",
  36878=>"011001111",
  36879=>"110110101",
  36880=>"001001110",
  36881=>"100100111",
  36882=>"111111100",
  36883=>"101001010",
  36884=>"111001100",
  36885=>"011100111",
  36886=>"011111000",
  36887=>"000001101",
  36888=>"101101000",
  36889=>"000011111",
  36890=>"111011000",
  36891=>"110000001",
  36892=>"001010110",
  36893=>"111111011",
  36894=>"111111000",
  36895=>"000010000",
  36896=>"110101100",
  36897=>"110000011",
  36898=>"111000000",
  36899=>"000100110",
  36900=>"110000010",
  36901=>"011010111",
  36902=>"000101001",
  36903=>"111111110",
  36904=>"101001010",
  36905=>"000010110",
  36906=>"010100001",
  36907=>"110100101",
  36908=>"011100100",
  36909=>"111101011",
  36910=>"000101101",
  36911=>"010001111",
  36912=>"110110100",
  36913=>"001010000",
  36914=>"101100011",
  36915=>"000100111",
  36916=>"010011011",
  36917=>"001101000",
  36918=>"101010100",
  36919=>"000001111",
  36920=>"000001101",
  36921=>"110111110",
  36922=>"111001100",
  36923=>"101010111",
  36924=>"110101100",
  36925=>"010000110",
  36926=>"001100001",
  36927=>"001110000",
  36928=>"100010010",
  36929=>"000000110",
  36930=>"101100000",
  36931=>"101000001",
  36932=>"111010011",
  36933=>"101001010",
  36934=>"000001000",
  36935=>"000101111",
  36936=>"110111110",
  36937=>"110101011",
  36938=>"111101001",
  36939=>"011010100",
  36940=>"001101000",
  36941=>"001101100",
  36942=>"110010101",
  36943=>"000110011",
  36944=>"010011011",
  36945=>"000010001",
  36946=>"100110101",
  36947=>"100111101",
  36948=>"110011010",
  36949=>"000011000",
  36950=>"010111101",
  36951=>"101100111",
  36952=>"001101001",
  36953=>"100010001",
  36954=>"010101011",
  36955=>"100011000",
  36956=>"000000001",
  36957=>"111010101",
  36958=>"111101000",
  36959=>"101000000",
  36960=>"010001111",
  36961=>"110011101",
  36962=>"100001110",
  36963=>"000100101",
  36964=>"101110101",
  36965=>"101010110",
  36966=>"011100001",
  36967=>"111010101",
  36968=>"010100101",
  36969=>"111101101",
  36970=>"110001010",
  36971=>"011010111",
  36972=>"101101101",
  36973=>"000011000",
  36974=>"010110000",
  36975=>"111000001",
  36976=>"101011101",
  36977=>"000011111",
  36978=>"100101110",
  36979=>"010101101",
  36980=>"011110100",
  36981=>"011011010",
  36982=>"111000000",
  36983=>"111000001",
  36984=>"111101001",
  36985=>"000000011",
  36986=>"111111101",
  36987=>"101111000",
  36988=>"111000111",
  36989=>"010001010",
  36990=>"100001111",
  36991=>"100110010",
  36992=>"010101110",
  36993=>"110001001",
  36994=>"000101110",
  36995=>"101010000",
  36996=>"010001000",
  36997=>"111011110",
  36998=>"001100011",
  36999=>"010101101",
  37000=>"010111001",
  37001=>"010011001",
  37002=>"001111101",
  37003=>"010001101",
  37004=>"101011100",
  37005=>"011011111",
  37006=>"001101110",
  37007=>"101100000",
  37008=>"010001111",
  37009=>"101000001",
  37010=>"000111011",
  37011=>"110101110",
  37012=>"101101110",
  37013=>"100011110",
  37014=>"011101100",
  37015=>"101100101",
  37016=>"000101000",
  37017=>"111111110",
  37018=>"100100111",
  37019=>"000110000",
  37020=>"000000000",
  37021=>"101110110",
  37022=>"100111101",
  37023=>"010111001",
  37024=>"100110111",
  37025=>"101000000",
  37026=>"000100111",
  37027=>"111001101",
  37028=>"101100000",
  37029=>"111111010",
  37030=>"011001010",
  37031=>"000110000",
  37032=>"011110110",
  37033=>"000011011",
  37034=>"010011110",
  37035=>"001101100",
  37036=>"001100100",
  37037=>"100000111",
  37038=>"011111000",
  37039=>"111001010",
  37040=>"010101100",
  37041=>"000100110",
  37042=>"000110010",
  37043=>"010110100",
  37044=>"101111111",
  37045=>"101111000",
  37046=>"010100000",
  37047=>"010101000",
  37048=>"111001010",
  37049=>"111000101",
  37050=>"000101001",
  37051=>"011001010",
  37052=>"101111000",
  37053=>"110100100",
  37054=>"111010011",
  37055=>"111111111",
  37056=>"010001100",
  37057=>"100011011",
  37058=>"001011100",
  37059=>"101111101",
  37060=>"000000001",
  37061=>"010101101",
  37062=>"110010100",
  37063=>"100001111",
  37064=>"101101011",
  37065=>"101011101",
  37066=>"100010101",
  37067=>"110100111",
  37068=>"001010100",
  37069=>"110010011",
  37070=>"111011100",
  37071=>"111011011",
  37072=>"001100000",
  37073=>"100011000",
  37074=>"000000111",
  37075=>"111110111",
  37076=>"010000010",
  37077=>"000100100",
  37078=>"001101111",
  37079=>"101101010",
  37080=>"111101000",
  37081=>"110011011",
  37082=>"110011001",
  37083=>"001011111",
  37084=>"110000000",
  37085=>"011100010",
  37086=>"100101001",
  37087=>"001100101",
  37088=>"011010111",
  37089=>"000001101",
  37090=>"010010100",
  37091=>"110100000",
  37092=>"110010101",
  37093=>"011000010",
  37094=>"000100010",
  37095=>"011101101",
  37096=>"101111011",
  37097=>"110000110",
  37098=>"110001001",
  37099=>"000000011",
  37100=>"110110110",
  37101=>"101101111",
  37102=>"110000010",
  37103=>"001101000",
  37104=>"000010010",
  37105=>"111010001",
  37106=>"000101101",
  37107=>"010110000",
  37108=>"101010110",
  37109=>"000100111",
  37110=>"001010100",
  37111=>"000000100",
  37112=>"101101010",
  37113=>"010101100",
  37114=>"010010101",
  37115=>"011010110",
  37116=>"110010000",
  37117=>"000010100",
  37118=>"110010110",
  37119=>"110000111",
  37120=>"111101001",
  37121=>"101010000",
  37122=>"000001100",
  37123=>"101011101",
  37124=>"110000000",
  37125=>"110100000",
  37126=>"011001010",
  37127=>"011000011",
  37128=>"000000100",
  37129=>"000101010",
  37130=>"101001100",
  37131=>"000010101",
  37132=>"101100110",
  37133=>"011010010",
  37134=>"111100010",
  37135=>"001110011",
  37136=>"100010011",
  37137=>"001010110",
  37138=>"011001110",
  37139=>"101011110",
  37140=>"110100001",
  37141=>"001101011",
  37142=>"011111001",
  37143=>"011011001",
  37144=>"100000001",
  37145=>"101110010",
  37146=>"000000101",
  37147=>"011000001",
  37148=>"111110000",
  37149=>"110010110",
  37150=>"011001001",
  37151=>"110000101",
  37152=>"001001101",
  37153=>"111010000",
  37154=>"101111011",
  37155=>"001110111",
  37156=>"000001111",
  37157=>"001110111",
  37158=>"010011111",
  37159=>"000111010",
  37160=>"101011001",
  37161=>"011100001",
  37162=>"110100001",
  37163=>"101111000",
  37164=>"001010100",
  37165=>"111100101",
  37166=>"100010110",
  37167=>"100011011",
  37168=>"101000111",
  37169=>"011011001",
  37170=>"000101111",
  37171=>"111000110",
  37172=>"001010100",
  37173=>"001011000",
  37174=>"101111100",
  37175=>"101100101",
  37176=>"100010100",
  37177=>"111011101",
  37178=>"101010010",
  37179=>"001001000",
  37180=>"111100001",
  37181=>"000010000",
  37182=>"011110000",
  37183=>"001100011",
  37184=>"100010100",
  37185=>"010000011",
  37186=>"000111111",
  37187=>"001100110",
  37188=>"011010100",
  37189=>"110101110",
  37190=>"011000100",
  37191=>"111000000",
  37192=>"110001110",
  37193=>"010001000",
  37194=>"011011011",
  37195=>"001101101",
  37196=>"111001001",
  37197=>"101011101",
  37198=>"000111000",
  37199=>"101101001",
  37200=>"100011111",
  37201=>"100011101",
  37202=>"111010100",
  37203=>"000011101",
  37204=>"001110001",
  37205=>"010110111",
  37206=>"100000101",
  37207=>"010100110",
  37208=>"100100111",
  37209=>"101000000",
  37210=>"011011010",
  37211=>"011000110",
  37212=>"110101011",
  37213=>"101001100",
  37214=>"100111100",
  37215=>"101000011",
  37216=>"101011010",
  37217=>"011110100",
  37218=>"100111101",
  37219=>"001001101",
  37220=>"100011110",
  37221=>"001001010",
  37222=>"111110010",
  37223=>"011011111",
  37224=>"000111011",
  37225=>"111010001",
  37226=>"001000011",
  37227=>"001101101",
  37228=>"100000111",
  37229=>"000001100",
  37230=>"001000101",
  37231=>"011101000",
  37232=>"001001100",
  37233=>"000000001",
  37234=>"001101011",
  37235=>"000011110",
  37236=>"101101011",
  37237=>"110100111",
  37238=>"000000100",
  37239=>"000011110",
  37240=>"001011011",
  37241=>"101010110",
  37242=>"011010100",
  37243=>"011000100",
  37244=>"001001000",
  37245=>"000001110",
  37246=>"000000000",
  37247=>"000001000",
  37248=>"001101100",
  37249=>"001100000",
  37250=>"011001110",
  37251=>"110010110",
  37252=>"100110010",
  37253=>"110001101",
  37254=>"000111011",
  37255=>"010001101",
  37256=>"100000000",
  37257=>"001101001",
  37258=>"001100111",
  37259=>"111000011",
  37260=>"100100000",
  37261=>"011101000",
  37262=>"001110110",
  37263=>"111100111",
  37264=>"101000101",
  37265=>"111101101",
  37266=>"011010000",
  37267=>"010101110",
  37268=>"001100110",
  37269=>"111010001",
  37270=>"000110111",
  37271=>"110110010",
  37272=>"100110011",
  37273=>"010101011",
  37274=>"111000100",
  37275=>"111010010",
  37276=>"101101101",
  37277=>"011101001",
  37278=>"010001111",
  37279=>"100110001",
  37280=>"111100010",
  37281=>"011000011",
  37282=>"000000001",
  37283=>"110010100",
  37284=>"001001100",
  37285=>"001110000",
  37286=>"100101101",
  37287=>"100110010",
  37288=>"011000000",
  37289=>"100011001",
  37290=>"100011110",
  37291=>"100010110",
  37292=>"100101111",
  37293=>"011010101",
  37294=>"000101001",
  37295=>"000110111",
  37296=>"111000011",
  37297=>"001111011",
  37298=>"000110000",
  37299=>"100111010",
  37300=>"011110010",
  37301=>"101110111",
  37302=>"011001011",
  37303=>"010001000",
  37304=>"010011100",
  37305=>"101000010",
  37306=>"111100111",
  37307=>"101001110",
  37308=>"000110101",
  37309=>"100000110",
  37310=>"001101111",
  37311=>"100010010",
  37312=>"100110011",
  37313=>"011100100",
  37314=>"011110110",
  37315=>"111011000",
  37316=>"001111111",
  37317=>"001101100",
  37318=>"111101011",
  37319=>"001100101",
  37320=>"000101110",
  37321=>"010101001",
  37322=>"000100011",
  37323=>"111111011",
  37324=>"111000111",
  37325=>"000110100",
  37326=>"001011011",
  37327=>"111010110",
  37328=>"000110111",
  37329=>"010010001",
  37330=>"001100011",
  37331=>"111110010",
  37332=>"001100110",
  37333=>"000101001",
  37334=>"000011010",
  37335=>"111100000",
  37336=>"000001101",
  37337=>"100011100",
  37338=>"010100001",
  37339=>"001111010",
  37340=>"110101111",
  37341=>"010111010",
  37342=>"010001101",
  37343=>"100001001",
  37344=>"111100101",
  37345=>"100110011",
  37346=>"110111101",
  37347=>"011011000",
  37348=>"000011100",
  37349=>"000001010",
  37350=>"110101101",
  37351=>"010110001",
  37352=>"110010000",
  37353=>"000101111",
  37354=>"110100100",
  37355=>"000101101",
  37356=>"011100000",
  37357=>"110111001",
  37358=>"101100100",
  37359=>"101101011",
  37360=>"111111110",
  37361=>"001011110",
  37362=>"100010111",
  37363=>"000011011",
  37364=>"110001100",
  37365=>"100001001",
  37366=>"100111000",
  37367=>"101000100",
  37368=>"001010000",
  37369=>"100111011",
  37370=>"101100110",
  37371=>"011111101",
  37372=>"100110010",
  37373=>"010001111",
  37374=>"100011000",
  37375=>"110010100",
  37376=>"111000101",
  37377=>"001110011",
  37378=>"100000011",
  37379=>"110010010",
  37380=>"100010100",
  37381=>"110101101",
  37382=>"111110111",
  37383=>"100111001",
  37384=>"110111000",
  37385=>"101101010",
  37386=>"100000110",
  37387=>"100010111",
  37388=>"011111111",
  37389=>"001011000",
  37390=>"100100010",
  37391=>"001011110",
  37392=>"110000101",
  37393=>"110111101",
  37394=>"010010101",
  37395=>"111000000",
  37396=>"000001000",
  37397=>"111010000",
  37398=>"100111010",
  37399=>"000001110",
  37400=>"100100111",
  37401=>"010011000",
  37402=>"100110101",
  37403=>"110100001",
  37404=>"010010001",
  37405=>"111100101",
  37406=>"001101001",
  37407=>"100001101",
  37408=>"100101011",
  37409=>"010000111",
  37410=>"001010000",
  37411=>"011110110",
  37412=>"110000100",
  37413=>"000110111",
  37414=>"011101010",
  37415=>"111011010",
  37416=>"111111110",
  37417=>"111111101",
  37418=>"011001000",
  37419=>"010001111",
  37420=>"010111000",
  37421=>"001100111",
  37422=>"100101010",
  37423=>"001101100",
  37424=>"001111010",
  37425=>"100011011",
  37426=>"010011000",
  37427=>"100001000",
  37428=>"111000110",
  37429=>"001011110",
  37430=>"001101101",
  37431=>"001100111",
  37432=>"101011110",
  37433=>"011101110",
  37434=>"100001110",
  37435=>"011110011",
  37436=>"011110000",
  37437=>"001110111",
  37438=>"010110111",
  37439=>"001010111",
  37440=>"000000010",
  37441=>"100011111",
  37442=>"100101010",
  37443=>"010010101",
  37444=>"010001001",
  37445=>"100001110",
  37446=>"000010001",
  37447=>"010111011",
  37448=>"100010100",
  37449=>"000101101",
  37450=>"101110000",
  37451=>"100000110",
  37452=>"101010100",
  37453=>"001010011",
  37454=>"010111000",
  37455=>"011110010",
  37456=>"010101100",
  37457=>"100010110",
  37458=>"110100111",
  37459=>"101010111",
  37460=>"000000110",
  37461=>"110000100",
  37462=>"000100101",
  37463=>"000001011",
  37464=>"110011101",
  37465=>"101101000",
  37466=>"011100000",
  37467=>"100010001",
  37468=>"010000000",
  37469=>"000100100",
  37470=>"100001101",
  37471=>"011010000",
  37472=>"000011111",
  37473=>"100001110",
  37474=>"100000000",
  37475=>"100010010",
  37476=>"011010010",
  37477=>"010000101",
  37478=>"110011110",
  37479=>"100101111",
  37480=>"110001001",
  37481=>"101110101",
  37482=>"010101000",
  37483=>"001001101",
  37484=>"110010100",
  37485=>"001010111",
  37486=>"011111000",
  37487=>"010001110",
  37488=>"100001010",
  37489=>"101000101",
  37490=>"111011001",
  37491=>"010000110",
  37492=>"001111010",
  37493=>"010010110",
  37494=>"000001011",
  37495=>"100110001",
  37496=>"011011100",
  37497=>"111100101",
  37498=>"110000101",
  37499=>"111110100",
  37500=>"011001011",
  37501=>"110011000",
  37502=>"010010011",
  37503=>"101100011",
  37504=>"101011010",
  37505=>"011001100",
  37506=>"101111010",
  37507=>"111001000",
  37508=>"110010101",
  37509=>"001000100",
  37510=>"111101110",
  37511=>"110111011",
  37512=>"000100111",
  37513=>"011100001",
  37514=>"110100001",
  37515=>"101010111",
  37516=>"010110100",
  37517=>"100000101",
  37518=>"101100001",
  37519=>"001000100",
  37520=>"111110101",
  37521=>"111001111",
  37522=>"101111010",
  37523=>"100000100",
  37524=>"100001101",
  37525=>"101101111",
  37526=>"101100000",
  37527=>"010011010",
  37528=>"011101010",
  37529=>"110000100",
  37530=>"000110111",
  37531=>"100100000",
  37532=>"000001000",
  37533=>"101011111",
  37534=>"111111001",
  37535=>"011010001",
  37536=>"010010111",
  37537=>"011011110",
  37538=>"111110100",
  37539=>"011101110",
  37540=>"010001001",
  37541=>"100011101",
  37542=>"010100111",
  37543=>"010010000",
  37544=>"000000010",
  37545=>"000011010",
  37546=>"100001001",
  37547=>"110101001",
  37548=>"010111101",
  37549=>"110000111",
  37550=>"000110110",
  37551=>"001000000",
  37552=>"111000110",
  37553=>"010100110",
  37554=>"101011011",
  37555=>"010011100",
  37556=>"000101110",
  37557=>"010001010",
  37558=>"111101111",
  37559=>"100110100",
  37560=>"001101011",
  37561=>"111110111",
  37562=>"100001100",
  37563=>"111100100",
  37564=>"000000111",
  37565=>"010110000",
  37566=>"010100101",
  37567=>"101010000",
  37568=>"010001111",
  37569=>"100000011",
  37570=>"101000101",
  37571=>"001011000",
  37572=>"010110010",
  37573=>"100001111",
  37574=>"011110101",
  37575=>"101111110",
  37576=>"001011100",
  37577=>"001100110",
  37578=>"111100101",
  37579=>"001001001",
  37580=>"101001101",
  37581=>"011111000",
  37582=>"110000001",
  37583=>"010000111",
  37584=>"100111111",
  37585=>"001111000",
  37586=>"110011000",
  37587=>"101110110",
  37588=>"001010001",
  37589=>"010001001",
  37590=>"111111111",
  37591=>"010001001",
  37592=>"000001011",
  37593=>"110100101",
  37594=>"010001101",
  37595=>"010010001",
  37596=>"001100000",
  37597=>"000110010",
  37598=>"000110001",
  37599=>"100111010",
  37600=>"011001000",
  37601=>"110111011",
  37602=>"001010001",
  37603=>"101100010",
  37604=>"000111011",
  37605=>"000100100",
  37606=>"000001000",
  37607=>"111001011",
  37608=>"101100001",
  37609=>"111000001",
  37610=>"001001101",
  37611=>"101100010",
  37612=>"100010010",
  37613=>"111010111",
  37614=>"101100111",
  37615=>"110101000",
  37616=>"111001100",
  37617=>"001100110",
  37618=>"100111001",
  37619=>"111010111",
  37620=>"010001010",
  37621=>"010110001",
  37622=>"100110011",
  37623=>"111100101",
  37624=>"011110111",
  37625=>"011101001",
  37626=>"000100010",
  37627=>"101000100",
  37628=>"111010011",
  37629=>"011100101",
  37630=>"110011000",
  37631=>"001110011",
  37632=>"011110111",
  37633=>"101010000",
  37634=>"100000110",
  37635=>"011000010",
  37636=>"111011101",
  37637=>"001100101",
  37638=>"010000011",
  37639=>"011000001",
  37640=>"011010000",
  37641=>"000110000",
  37642=>"100110010",
  37643=>"001000000",
  37644=>"011010111",
  37645=>"110011000",
  37646=>"010100000",
  37647=>"001110000",
  37648=>"110010110",
  37649=>"001001010",
  37650=>"101010110",
  37651=>"010010100",
  37652=>"011001110",
  37653=>"110100000",
  37654=>"001111100",
  37655=>"000000011",
  37656=>"010100010",
  37657=>"000100000",
  37658=>"111001110",
  37659=>"101010000",
  37660=>"000000001",
  37661=>"011101111",
  37662=>"000011110",
  37663=>"110001000",
  37664=>"000000110",
  37665=>"001010011",
  37666=>"110010111",
  37667=>"101101000",
  37668=>"101011111",
  37669=>"110110000",
  37670=>"110111101",
  37671=>"001110111",
  37672=>"110011110",
  37673=>"010000101",
  37674=>"100111101",
  37675=>"100110010",
  37676=>"101101110",
  37677=>"111001100",
  37678=>"101000111",
  37679=>"110000011",
  37680=>"110010101",
  37681=>"011100110",
  37682=>"101001001",
  37683=>"101101000",
  37684=>"100010001",
  37685=>"010010011",
  37686=>"001100100",
  37687=>"111101010",
  37688=>"010000010",
  37689=>"000000101",
  37690=>"001000001",
  37691=>"010100000",
  37692=>"000010010",
  37693=>"111001010",
  37694=>"111010010",
  37695=>"101101111",
  37696=>"000110000",
  37697=>"010001111",
  37698=>"001011010",
  37699=>"100010101",
  37700=>"010101000",
  37701=>"101100011",
  37702=>"010011100",
  37703=>"101101100",
  37704=>"101110101",
  37705=>"100111110",
  37706=>"111101011",
  37707=>"111111011",
  37708=>"110001100",
  37709=>"010001111",
  37710=>"001001010",
  37711=>"011000000",
  37712=>"100100000",
  37713=>"100011001",
  37714=>"010010111",
  37715=>"000011111",
  37716=>"010111001",
  37717=>"010011101",
  37718=>"100100000",
  37719=>"010011111",
  37720=>"001001011",
  37721=>"001101000",
  37722=>"101110110",
  37723=>"101000011",
  37724=>"110011011",
  37725=>"011001100",
  37726=>"000000100",
  37727=>"011101111",
  37728=>"010000001",
  37729=>"000101101",
  37730=>"100001101",
  37731=>"011001001",
  37732=>"111010010",
  37733=>"101000101",
  37734=>"001000110",
  37735=>"001010011",
  37736=>"001110000",
  37737=>"111001101",
  37738=>"000101100",
  37739=>"010010100",
  37740=>"101011000",
  37741=>"010100001",
  37742=>"000001100",
  37743=>"001000011",
  37744=>"010001110",
  37745=>"100000111",
  37746=>"110010100",
  37747=>"111111101",
  37748=>"111010001",
  37749=>"100000101",
  37750=>"000001011",
  37751=>"111111011",
  37752=>"100100110",
  37753=>"111110100",
  37754=>"010011000",
  37755=>"010000101",
  37756=>"000001011",
  37757=>"010101101",
  37758=>"111010001",
  37759=>"101000001",
  37760=>"001000010",
  37761=>"001110110",
  37762=>"001111100",
  37763=>"010101010",
  37764=>"111100101",
  37765=>"111001101",
  37766=>"110111010",
  37767=>"001011011",
  37768=>"001111101",
  37769=>"011100100",
  37770=>"110000111",
  37771=>"010010110",
  37772=>"000000111",
  37773=>"000110100",
  37774=>"101101100",
  37775=>"000111011",
  37776=>"100111100",
  37777=>"110011001",
  37778=>"000010011",
  37779=>"110111000",
  37780=>"111010001",
  37781=>"100110111",
  37782=>"010010110",
  37783=>"110110010",
  37784=>"100100111",
  37785=>"110101000",
  37786=>"100011110",
  37787=>"001010000",
  37788=>"010010100",
  37789=>"001101011",
  37790=>"010010010",
  37791=>"010100111",
  37792=>"100011010",
  37793=>"111010100",
  37794=>"000110010",
  37795=>"011001010",
  37796=>"011011000",
  37797=>"100011011",
  37798=>"011100001",
  37799=>"011101110",
  37800=>"011110100",
  37801=>"101111001",
  37802=>"111010001",
  37803=>"110010000",
  37804=>"100101100",
  37805=>"011100111",
  37806=>"000101001",
  37807=>"011100100",
  37808=>"010100111",
  37809=>"000001000",
  37810=>"001110110",
  37811=>"100010000",
  37812=>"000101000",
  37813=>"111111011",
  37814=>"101100001",
  37815=>"110000001",
  37816=>"000111001",
  37817=>"100101001",
  37818=>"000001000",
  37819=>"110001010",
  37820=>"011101001",
  37821=>"101110110",
  37822=>"101101010",
  37823=>"111011110",
  37824=>"011110111",
  37825=>"101010100",
  37826=>"101100100",
  37827=>"001111101",
  37828=>"110000001",
  37829=>"000001111",
  37830=>"100011100",
  37831=>"111110111",
  37832=>"000110000",
  37833=>"111110010",
  37834=>"110010100",
  37835=>"010111111",
  37836=>"001010010",
  37837=>"111001001",
  37838=>"110001111",
  37839=>"101111001",
  37840=>"110010110",
  37841=>"010000010",
  37842=>"001111101",
  37843=>"000000100",
  37844=>"100111110",
  37845=>"111110111",
  37846=>"000011111",
  37847=>"001100110",
  37848=>"111101110",
  37849=>"110101101",
  37850=>"010001010",
  37851=>"000001011",
  37852=>"111000100",
  37853=>"111000111",
  37854=>"010111101",
  37855=>"101000011",
  37856=>"101111000",
  37857=>"111110101",
  37858=>"111011110",
  37859=>"011100000",
  37860=>"000000101",
  37861=>"111101010",
  37862=>"010110001",
  37863=>"111000100",
  37864=>"001000011",
  37865=>"011000011",
  37866=>"110011000",
  37867=>"010001101",
  37868=>"111111101",
  37869=>"000000010",
  37870=>"010001100",
  37871=>"111011010",
  37872=>"100111010",
  37873=>"011101110",
  37874=>"100110100",
  37875=>"010000100",
  37876=>"101111111",
  37877=>"000001111",
  37878=>"010011000",
  37879=>"110000101",
  37880=>"001000010",
  37881=>"010011000",
  37882=>"010000111",
  37883=>"110100001",
  37884=>"011101100",
  37885=>"111010101",
  37886=>"000100110",
  37887=>"011101001",
  37888=>"110110111",
  37889=>"001000101",
  37890=>"101000111",
  37891=>"101101100",
  37892=>"100111110",
  37893=>"000100000",
  37894=>"101111000",
  37895=>"000111010",
  37896=>"110010000",
  37897=>"001101001",
  37898=>"111101101",
  37899=>"101001000",
  37900=>"101110111",
  37901=>"011000100",
  37902=>"100101001",
  37903=>"111000101",
  37904=>"010000100",
  37905=>"001100110",
  37906=>"111011110",
  37907=>"000011101",
  37908=>"000110101",
  37909=>"110001101",
  37910=>"000100100",
  37911=>"001010010",
  37912=>"001000110",
  37913=>"100011100",
  37914=>"011101011",
  37915=>"100101110",
  37916=>"101101000",
  37917=>"010000011",
  37918=>"110001101",
  37919=>"010001001",
  37920=>"110000000",
  37921=>"110000110",
  37922=>"000010000",
  37923=>"011001101",
  37924=>"010111101",
  37925=>"110101001",
  37926=>"011000001",
  37927=>"100101111",
  37928=>"101111101",
  37929=>"010101111",
  37930=>"010100111",
  37931=>"111111000",
  37932=>"010100111",
  37933=>"000011110",
  37934=>"011111001",
  37935=>"100100000",
  37936=>"100011001",
  37937=>"010011010",
  37938=>"000101000",
  37939=>"011111100",
  37940=>"010111101",
  37941=>"101100000",
  37942=>"000101101",
  37943=>"111101110",
  37944=>"110110101",
  37945=>"001110010",
  37946=>"100010010",
  37947=>"000100101",
  37948=>"011110100",
  37949=>"001110110",
  37950=>"111000011",
  37951=>"001110111",
  37952=>"001001100",
  37953=>"000000011",
  37954=>"101000001",
  37955=>"100101000",
  37956=>"000100011",
  37957=>"001011101",
  37958=>"110100010",
  37959=>"100001000",
  37960=>"000110000",
  37961=>"010010010",
  37962=>"110110011",
  37963=>"010001100",
  37964=>"011011111",
  37965=>"110000101",
  37966=>"111101111",
  37967=>"111111101",
  37968=>"010110000",
  37969=>"011111011",
  37970=>"111100001",
  37971=>"111111011",
  37972=>"010001111",
  37973=>"110011000",
  37974=>"010011011",
  37975=>"100100110",
  37976=>"110001000",
  37977=>"111011111",
  37978=>"010111010",
  37979=>"001000000",
  37980=>"011110010",
  37981=>"001011111",
  37982=>"000011110",
  37983=>"000000011",
  37984=>"111100101",
  37985=>"111111001",
  37986=>"100110101",
  37987=>"100000100",
  37988=>"110110100",
  37989=>"100000101",
  37990=>"111001101",
  37991=>"000110010",
  37992=>"010001101",
  37993=>"011100100",
  37994=>"010100000",
  37995=>"000011101",
  37996=>"010101001",
  37997=>"011100101",
  37998=>"010111000",
  37999=>"010010001",
  38000=>"111000111",
  38001=>"111101100",
  38002=>"000101001",
  38003=>"111001100",
  38004=>"010101100",
  38005=>"010100111",
  38006=>"101010010",
  38007=>"111010111",
  38008=>"101111101",
  38009=>"001111101",
  38010=>"110100011",
  38011=>"101110111",
  38012=>"000010001",
  38013=>"100010101",
  38014=>"100110110",
  38015=>"101111010",
  38016=>"000010001",
  38017=>"101001100",
  38018=>"110011000",
  38019=>"110100000",
  38020=>"001101000",
  38021=>"000011101",
  38022=>"100110000",
  38023=>"100011110",
  38024=>"101101110",
  38025=>"100001100",
  38026=>"001010010",
  38027=>"011000010",
  38028=>"110010000",
  38029=>"100000000",
  38030=>"110100010",
  38031=>"100000111",
  38032=>"110011101",
  38033=>"010100111",
  38034=>"101011111",
  38035=>"111110110",
  38036=>"000111001",
  38037=>"011111001",
  38038=>"111100001",
  38039=>"011000110",
  38040=>"101101010",
  38041=>"001101111",
  38042=>"110111101",
  38043=>"111011110",
  38044=>"000100000",
  38045=>"111000000",
  38046=>"010001000",
  38047=>"000110100",
  38048=>"001000100",
  38049=>"100110001",
  38050=>"010101100",
  38051=>"101000101",
  38052=>"110110000",
  38053=>"010100011",
  38054=>"100000101",
  38055=>"111110100",
  38056=>"011001101",
  38057=>"001000000",
  38058=>"101100010",
  38059=>"111101101",
  38060=>"101000010",
  38061=>"000111001",
  38062=>"101111111",
  38063=>"110000111",
  38064=>"010001110",
  38065=>"010011110",
  38066=>"010011000",
  38067=>"001001011",
  38068=>"100110001",
  38069=>"000001010",
  38070=>"111100100",
  38071=>"011000000",
  38072=>"110001100",
  38073=>"011001001",
  38074=>"011100011",
  38075=>"110111000",
  38076=>"111100111",
  38077=>"111011000",
  38078=>"110100100",
  38079=>"100001110",
  38080=>"011100010",
  38081=>"000000111",
  38082=>"011010010",
  38083=>"011010111",
  38084=>"111111111",
  38085=>"001101110",
  38086=>"010011101",
  38087=>"000100001",
  38088=>"001011100",
  38089=>"001100110",
  38090=>"100110111",
  38091=>"101111111",
  38092=>"011101111",
  38093=>"100000010",
  38094=>"011100011",
  38095=>"111100010",
  38096=>"000001100",
  38097=>"010010010",
  38098=>"100111101",
  38099=>"101011010",
  38100=>"000011001",
  38101=>"000111100",
  38102=>"011011010",
  38103=>"001000001",
  38104=>"010110010",
  38105=>"110000110",
  38106=>"011010010",
  38107=>"101110111",
  38108=>"110011110",
  38109=>"111011010",
  38110=>"010111010",
  38111=>"011110110",
  38112=>"110101000",
  38113=>"100000000",
  38114=>"001010100",
  38115=>"001111101",
  38116=>"110000011",
  38117=>"111110001",
  38118=>"100111100",
  38119=>"001110110",
  38120=>"001000000",
  38121=>"010000101",
  38122=>"000100000",
  38123=>"001010010",
  38124=>"000000010",
  38125=>"111111110",
  38126=>"100101100",
  38127=>"100011100",
  38128=>"110011101",
  38129=>"110100101",
  38130=>"011010100",
  38131=>"010101110",
  38132=>"010000100",
  38133=>"101010010",
  38134=>"111100110",
  38135=>"110001110",
  38136=>"111011000",
  38137=>"111001111",
  38138=>"011000001",
  38139=>"000100111",
  38140=>"110010100",
  38141=>"110001000",
  38142=>"101111111",
  38143=>"011011110",
  38144=>"100010101",
  38145=>"100111011",
  38146=>"101110011",
  38147=>"100110000",
  38148=>"010000100",
  38149=>"001001110",
  38150=>"011101001",
  38151=>"011101100",
  38152=>"010101001",
  38153=>"111101111",
  38154=>"110100010",
  38155=>"010100010",
  38156=>"110000100",
  38157=>"010010101",
  38158=>"000010000",
  38159=>"110111000",
  38160=>"110000101",
  38161=>"110111001",
  38162=>"111110100",
  38163=>"011010101",
  38164=>"010010001",
  38165=>"001110000",
  38166=>"101010100",
  38167=>"101100101",
  38168=>"001000011",
  38169=>"010010111",
  38170=>"011101010",
  38171=>"010101101",
  38172=>"000110111",
  38173=>"011101101",
  38174=>"101101100",
  38175=>"100001100",
  38176=>"000100011",
  38177=>"001001110",
  38178=>"101111000",
  38179=>"110110010",
  38180=>"000101101",
  38181=>"001100000",
  38182=>"001000110",
  38183=>"001100101",
  38184=>"110101010",
  38185=>"101111101",
  38186=>"110110101",
  38187=>"011000001",
  38188=>"101111111",
  38189=>"101111111",
  38190=>"100000001",
  38191=>"111000111",
  38192=>"101001101",
  38193=>"011010100",
  38194=>"101101101",
  38195=>"000001000",
  38196=>"000011110",
  38197=>"010111001",
  38198=>"100010000",
  38199=>"011100101",
  38200=>"011010000",
  38201=>"101101001",
  38202=>"110011110",
  38203=>"001001001",
  38204=>"101110110",
  38205=>"011100110",
  38206=>"110011101",
  38207=>"000110010",
  38208=>"000110100",
  38209=>"100001011",
  38210=>"101101101",
  38211=>"010100101",
  38212=>"111111000",
  38213=>"001001011",
  38214=>"110010011",
  38215=>"101101001",
  38216=>"110011110",
  38217=>"000001101",
  38218=>"000110110",
  38219=>"111111110",
  38220=>"111010000",
  38221=>"100101111",
  38222=>"110001000",
  38223=>"000001100",
  38224=>"101001010",
  38225=>"011101011",
  38226=>"111010010",
  38227=>"000100011",
  38228=>"000011000",
  38229=>"101001001",
  38230=>"010111010",
  38231=>"011111000",
  38232=>"100111111",
  38233=>"000010011",
  38234=>"010000101",
  38235=>"100100011",
  38236=>"110000011",
  38237=>"111000101",
  38238=>"110100110",
  38239=>"100001100",
  38240=>"011101000",
  38241=>"101110100",
  38242=>"000100111",
  38243=>"011110111",
  38244=>"100110110",
  38245=>"101001000",
  38246=>"111100100",
  38247=>"001011001",
  38248=>"111010111",
  38249=>"101101110",
  38250=>"001001010",
  38251=>"011011110",
  38252=>"110110100",
  38253=>"000000011",
  38254=>"101101110",
  38255=>"000101100",
  38256=>"111011000",
  38257=>"100100101",
  38258=>"110001110",
  38259=>"000100000",
  38260=>"011001110",
  38261=>"110010100",
  38262=>"011001111",
  38263=>"100101001",
  38264=>"010100111",
  38265=>"100101011",
  38266=>"011011011",
  38267=>"000100110",
  38268=>"110110001",
  38269=>"111101100",
  38270=>"011001110",
  38271=>"110011000",
  38272=>"111111000",
  38273=>"111100101",
  38274=>"111100011",
  38275=>"100010000",
  38276=>"000000111",
  38277=>"001111010",
  38278=>"011011101",
  38279=>"000001100",
  38280=>"101010001",
  38281=>"111001111",
  38282=>"101100111",
  38283=>"100000101",
  38284=>"110110110",
  38285=>"101001000",
  38286=>"011111011",
  38287=>"010010111",
  38288=>"111100111",
  38289=>"000101000",
  38290=>"000010111",
  38291=>"011000100",
  38292=>"111011101",
  38293=>"011100011",
  38294=>"111110100",
  38295=>"010110001",
  38296=>"100010000",
  38297=>"000000001",
  38298=>"000111001",
  38299=>"110000001",
  38300=>"110011000",
  38301=>"101001100",
  38302=>"111111111",
  38303=>"100001111",
  38304=>"001101011",
  38305=>"010100011",
  38306=>"000010000",
  38307=>"100011100",
  38308=>"010111001",
  38309=>"011011101",
  38310=>"111011010",
  38311=>"001100100",
  38312=>"111000110",
  38313=>"100101110",
  38314=>"000110010",
  38315=>"001111110",
  38316=>"010110100",
  38317=>"011011101",
  38318=>"000111010",
  38319=>"000011100",
  38320=>"000110010",
  38321=>"110111101",
  38322=>"011010101",
  38323=>"111111011",
  38324=>"101010100",
  38325=>"110100110",
  38326=>"100011010",
  38327=>"010111111",
  38328=>"010111111",
  38329=>"110010000",
  38330=>"101011010",
  38331=>"110111111",
  38332=>"111010111",
  38333=>"011010110",
  38334=>"101111110",
  38335=>"110011000",
  38336=>"010010001",
  38337=>"100011111",
  38338=>"000110101",
  38339=>"001001011",
  38340=>"100011110",
  38341=>"011011011",
  38342=>"000011000",
  38343=>"010110000",
  38344=>"010001100",
  38345=>"111000100",
  38346=>"100001001",
  38347=>"101101111",
  38348=>"110000010",
  38349=>"111101000",
  38350=>"111101100",
  38351=>"001010101",
  38352=>"101000011",
  38353=>"011111010",
  38354=>"100100100",
  38355=>"101000000",
  38356=>"110000011",
  38357=>"111110010",
  38358=>"111000100",
  38359=>"011101101",
  38360=>"100100001",
  38361=>"000001000",
  38362=>"000101000",
  38363=>"110011100",
  38364=>"110111011",
  38365=>"010010011",
  38366=>"101011100",
  38367=>"001110100",
  38368=>"001000000",
  38369=>"001001101",
  38370=>"110100011",
  38371=>"000010001",
  38372=>"010110001",
  38373=>"001011010",
  38374=>"011111101",
  38375=>"001000000",
  38376=>"100110011",
  38377=>"111101011",
  38378=>"101010010",
  38379=>"000011000",
  38380=>"100100011",
  38381=>"000000011",
  38382=>"010101000",
  38383=>"011101100",
  38384=>"000110001",
  38385=>"001011101",
  38386=>"010001010",
  38387=>"111011010",
  38388=>"101100111",
  38389=>"001100010",
  38390=>"010010110",
  38391=>"101011111",
  38392=>"000011111",
  38393=>"000100111",
  38394=>"111111111",
  38395=>"110011010",
  38396=>"110010101",
  38397=>"010010110",
  38398=>"111001100",
  38399=>"111100011",
  38400=>"011001001",
  38401=>"001110110",
  38402=>"001110001",
  38403=>"101000011",
  38404=>"101110111",
  38405=>"111001110",
  38406=>"001000110",
  38407=>"000010001",
  38408=>"010111001",
  38409=>"101010110",
  38410=>"100010010",
  38411=>"110010110",
  38412=>"000010011",
  38413=>"100001000",
  38414=>"110111001",
  38415=>"111111111",
  38416=>"100111011",
  38417=>"110010010",
  38418=>"010100011",
  38419=>"000000100",
  38420=>"001111101",
  38421=>"000001000",
  38422=>"001010111",
  38423=>"111001111",
  38424=>"101010011",
  38425=>"001011001",
  38426=>"101000001",
  38427=>"101110001",
  38428=>"111110010",
  38429=>"010111010",
  38430=>"110111101",
  38431=>"010011110",
  38432=>"011010001",
  38433=>"110000100",
  38434=>"000001100",
  38435=>"000110010",
  38436=>"011011111",
  38437=>"010100110",
  38438=>"111001111",
  38439=>"110000100",
  38440=>"000001001",
  38441=>"001111101",
  38442=>"010010110",
  38443=>"001011011",
  38444=>"000000000",
  38445=>"101100110",
  38446=>"011100100",
  38447=>"111100101",
  38448=>"101001011",
  38449=>"110110110",
  38450=>"110000010",
  38451=>"000000010",
  38452=>"011010001",
  38453=>"111011010",
  38454=>"010111111",
  38455=>"010000001",
  38456=>"100110100",
  38457=>"001111011",
  38458=>"000010100",
  38459=>"110011101",
  38460=>"110101100",
  38461=>"001000101",
  38462=>"100011101",
  38463=>"011001000",
  38464=>"110000100",
  38465=>"111110111",
  38466=>"100011000",
  38467=>"011000010",
  38468=>"111001100",
  38469=>"101110000",
  38470=>"010011000",
  38471=>"011110111",
  38472=>"001000001",
  38473=>"111000110",
  38474=>"100110001",
  38475=>"100011001",
  38476=>"010001010",
  38477=>"011100110",
  38478=>"110000001",
  38479=>"000111010",
  38480=>"100111101",
  38481=>"100001000",
  38482=>"101100101",
  38483=>"100100100",
  38484=>"100100010",
  38485=>"100000111",
  38486=>"110000101",
  38487=>"010000110",
  38488=>"001110100",
  38489=>"101100110",
  38490=>"000010000",
  38491=>"010110100",
  38492=>"110010011",
  38493=>"101110110",
  38494=>"000000101",
  38495=>"000100000",
  38496=>"001110011",
  38497=>"000000101",
  38498=>"111100010",
  38499=>"000001001",
  38500=>"100011000",
  38501=>"110000001",
  38502=>"001011100",
  38503=>"111101011",
  38504=>"100001001",
  38505=>"101010110",
  38506=>"110100101",
  38507=>"001001001",
  38508=>"010100110",
  38509=>"010001100",
  38510=>"110101001",
  38511=>"100101101",
  38512=>"010110011",
  38513=>"011010100",
  38514=>"100101101",
  38515=>"111001110",
  38516=>"100111000",
  38517=>"000111100",
  38518=>"010000000",
  38519=>"110010010",
  38520=>"011000110",
  38521=>"010100100",
  38522=>"111011010",
  38523=>"100100100",
  38524=>"100011100",
  38525=>"101001111",
  38526=>"011101001",
  38527=>"001111100",
  38528=>"111110111",
  38529=>"110100000",
  38530=>"001011000",
  38531=>"010110000",
  38532=>"111011101",
  38533=>"110011110",
  38534=>"101001100",
  38535=>"011001011",
  38536=>"101111010",
  38537=>"010010011",
  38538=>"011011011",
  38539=>"111111111",
  38540=>"001001100",
  38541=>"010011000",
  38542=>"100000110",
  38543=>"001000110",
  38544=>"111110110",
  38545=>"000010001",
  38546=>"111111000",
  38547=>"011000101",
  38548=>"111110000",
  38549=>"110110001",
  38550=>"011010010",
  38551=>"011110110",
  38552=>"011100000",
  38553=>"101000111",
  38554=>"101011010",
  38555=>"111110111",
  38556=>"111010011",
  38557=>"001000111",
  38558=>"011000011",
  38559=>"111111111",
  38560=>"110101000",
  38561=>"000000110",
  38562=>"111111010",
  38563=>"000010000",
  38564=>"010000111",
  38565=>"000100111",
  38566=>"111001001",
  38567=>"010010000",
  38568=>"000100010",
  38569=>"110011011",
  38570=>"000001011",
  38571=>"001011010",
  38572=>"010100111",
  38573=>"001001100",
  38574=>"111000000",
  38575=>"001111101",
  38576=>"101111010",
  38577=>"110101111",
  38578=>"000101010",
  38579=>"110110110",
  38580=>"110101000",
  38581=>"100111000",
  38582=>"011111010",
  38583=>"101100111",
  38584=>"010011001",
  38585=>"110100111",
  38586=>"111010110",
  38587=>"001001111",
  38588=>"100011111",
  38589=>"111101000",
  38590=>"001001010",
  38591=>"000100110",
  38592=>"101001111",
  38593=>"110110001",
  38594=>"110001011",
  38595=>"110101111",
  38596=>"001011011",
  38597=>"010111011",
  38598=>"100110101",
  38599=>"110011100",
  38600=>"101111000",
  38601=>"010011100",
  38602=>"011110100",
  38603=>"100000010",
  38604=>"001111010",
  38605=>"111111000",
  38606=>"010011101",
  38607=>"100011110",
  38608=>"101010000",
  38609=>"010100001",
  38610=>"101000000",
  38611=>"100010110",
  38612=>"100101000",
  38613=>"001111101",
  38614=>"101000101",
  38615=>"001111111",
  38616=>"111011111",
  38617=>"011011001",
  38618=>"110001001",
  38619=>"000100001",
  38620=>"011000010",
  38621=>"000010000",
  38622=>"000001001",
  38623=>"010011110",
  38624=>"110100101",
  38625=>"101000001",
  38626=>"001110011",
  38627=>"111001111",
  38628=>"111111100",
  38629=>"101000001",
  38630=>"101110110",
  38631=>"101111110",
  38632=>"000101011",
  38633=>"110010101",
  38634=>"100101101",
  38635=>"010000100",
  38636=>"010000011",
  38637=>"001010111",
  38638=>"001111110",
  38639=>"010100000",
  38640=>"111011011",
  38641=>"010101111",
  38642=>"000110110",
  38643=>"100000101",
  38644=>"101111111",
  38645=>"101110101",
  38646=>"000001101",
  38647=>"000010000",
  38648=>"011100011",
  38649=>"111010100",
  38650=>"000000010",
  38651=>"100000001",
  38652=>"011101111",
  38653=>"101111000",
  38654=>"000101011",
  38655=>"000010110",
  38656=>"000010110",
  38657=>"110011110",
  38658=>"001000010",
  38659=>"111001001",
  38660=>"000001100",
  38661=>"000000010",
  38662=>"001100000",
  38663=>"101011101",
  38664=>"100011000",
  38665=>"010001000",
  38666=>"000100110",
  38667=>"001101001",
  38668=>"110011100",
  38669=>"000000100",
  38670=>"000011101",
  38671=>"101101111",
  38672=>"110100110",
  38673=>"011110011",
  38674=>"010111111",
  38675=>"000000111",
  38676=>"010001001",
  38677=>"001001000",
  38678=>"110101011",
  38679=>"000110010",
  38680=>"000001001",
  38681=>"001101100",
  38682=>"011110111",
  38683=>"001011010",
  38684=>"100101100",
  38685=>"111110001",
  38686=>"101000011",
  38687=>"001001100",
  38688=>"011110000",
  38689=>"011000101",
  38690=>"111111000",
  38691=>"101110111",
  38692=>"000011010",
  38693=>"000101010",
  38694=>"000101111",
  38695=>"000111110",
  38696=>"111000111",
  38697=>"011111101",
  38698=>"101100100",
  38699=>"000110010",
  38700=>"000101010",
  38701=>"111101111",
  38702=>"001011001",
  38703=>"101011000",
  38704=>"111000101",
  38705=>"111000010",
  38706=>"110110010",
  38707=>"011010001",
  38708=>"101010101",
  38709=>"000000011",
  38710=>"001001111",
  38711=>"011101101",
  38712=>"111110110",
  38713=>"100000110",
  38714=>"011000000",
  38715=>"010101000",
  38716=>"111011010",
  38717=>"111111111",
  38718=>"111110101",
  38719=>"000000110",
  38720=>"010101001",
  38721=>"101000111",
  38722=>"100010001",
  38723=>"010000001",
  38724=>"011100111",
  38725=>"001011000",
  38726=>"100000111",
  38727=>"100001001",
  38728=>"110101000",
  38729=>"011101010",
  38730=>"101001010",
  38731=>"000010000",
  38732=>"100001000",
  38733=>"001011001",
  38734=>"010111110",
  38735=>"101100101",
  38736=>"111101000",
  38737=>"011100010",
  38738=>"110101001",
  38739=>"100010110",
  38740=>"101000001",
  38741=>"011010001",
  38742=>"101111111",
  38743=>"001001100",
  38744=>"101100010",
  38745=>"100010010",
  38746=>"111110010",
  38747=>"011101101",
  38748=>"110001010",
  38749=>"110111101",
  38750=>"111100011",
  38751=>"100001100",
  38752=>"001000001",
  38753=>"000100110",
  38754=>"110000100",
  38755=>"100010110",
  38756=>"010001010",
  38757=>"010010001",
  38758=>"001011110",
  38759=>"110011011",
  38760=>"101110111",
  38761=>"101001011",
  38762=>"011001010",
  38763=>"001010011",
  38764=>"101011000",
  38765=>"011110111",
  38766=>"000000000",
  38767=>"101001111",
  38768=>"010010001",
  38769=>"001011101",
  38770=>"011001000",
  38771=>"000100111",
  38772=>"010000110",
  38773=>"100111001",
  38774=>"100110001",
  38775=>"101011110",
  38776=>"001100011",
  38777=>"000110011",
  38778=>"111100011",
  38779=>"000011011",
  38780=>"101101101",
  38781=>"101010100",
  38782=>"101010011",
  38783=>"101111000",
  38784=>"010111000",
  38785=>"011110011",
  38786=>"011000111",
  38787=>"100000110",
  38788=>"100010101",
  38789=>"011000101",
  38790=>"011101010",
  38791=>"000010100",
  38792=>"010001100",
  38793=>"001101101",
  38794=>"001000000",
  38795=>"000000000",
  38796=>"000000111",
  38797=>"101111001",
  38798=>"001101110",
  38799=>"011011001",
  38800=>"011100000",
  38801=>"000011011",
  38802=>"010011100",
  38803=>"111001010",
  38804=>"000011101",
  38805=>"000011101",
  38806=>"101011001",
  38807=>"001011111",
  38808=>"000011000",
  38809=>"101011110",
  38810=>"000101110",
  38811=>"001001101",
  38812=>"110000111",
  38813=>"101111000",
  38814=>"000001100",
  38815=>"100111101",
  38816=>"000100100",
  38817=>"111101001",
  38818=>"101101111",
  38819=>"001111010",
  38820=>"001011111",
  38821=>"010110010",
  38822=>"101000001",
  38823=>"111101000",
  38824=>"001000010",
  38825=>"011010000",
  38826=>"111010101",
  38827=>"010101001",
  38828=>"100010010",
  38829=>"010101101",
  38830=>"000001100",
  38831=>"010111011",
  38832=>"010100110",
  38833=>"111111110",
  38834=>"010111010",
  38835=>"110001011",
  38836=>"010000001",
  38837=>"011100000",
  38838=>"101001011",
  38839=>"111000100",
  38840=>"111010011",
  38841=>"111001111",
  38842=>"111110011",
  38843=>"001110000",
  38844=>"011110001",
  38845=>"101000100",
  38846=>"011100011",
  38847=>"100100000",
  38848=>"101001011",
  38849=>"010111111",
  38850=>"111111110",
  38851=>"101011000",
  38852=>"010111010",
  38853=>"101101001",
  38854=>"010000100",
  38855=>"111110100",
  38856=>"011100101",
  38857=>"111010110",
  38858=>"111110001",
  38859=>"101110111",
  38860=>"000101110",
  38861=>"011111011",
  38862=>"101111010",
  38863=>"100000000",
  38864=>"011001001",
  38865=>"010100000",
  38866=>"010100111",
  38867=>"001101111",
  38868=>"001010001",
  38869=>"101001101",
  38870=>"110000011",
  38871=>"100111010",
  38872=>"100100101",
  38873=>"011111011",
  38874=>"100010101",
  38875=>"011111101",
  38876=>"001101001",
  38877=>"000101010",
  38878=>"001001110",
  38879=>"001011000",
  38880=>"111001100",
  38881=>"001001011",
  38882=>"111000101",
  38883=>"100001111",
  38884=>"001101010",
  38885=>"111101100",
  38886=>"000011101",
  38887=>"010101101",
  38888=>"000111011",
  38889=>"000010000",
  38890=>"010100001",
  38891=>"111100101",
  38892=>"001001111",
  38893=>"111001011",
  38894=>"101011110",
  38895=>"100111111",
  38896=>"010110110",
  38897=>"100010010",
  38898=>"011111111",
  38899=>"000011110",
  38900=>"101010001",
  38901=>"111001110",
  38902=>"101011110",
  38903=>"001100000",
  38904=>"001001001",
  38905=>"101101100",
  38906=>"011100110",
  38907=>"000011000",
  38908=>"100110011",
  38909=>"000010010",
  38910=>"000111010",
  38911=>"111111011",
  38912=>"100000011",
  38913=>"101110001",
  38914=>"100001110",
  38915=>"110010100",
  38916=>"111111111",
  38917=>"111001111",
  38918=>"001010011",
  38919=>"111111111",
  38920=>"100011010",
  38921=>"111011011",
  38922=>"001011000",
  38923=>"000110100",
  38924=>"100101101",
  38925=>"100000011",
  38926=>"111101001",
  38927=>"001111010",
  38928=>"000000011",
  38929=>"000000000",
  38930=>"101111000",
  38931=>"010001101",
  38932=>"110011101",
  38933=>"110011000",
  38934=>"100001010",
  38935=>"100001111",
  38936=>"010011100",
  38937=>"100010001",
  38938=>"000001111",
  38939=>"001110100",
  38940=>"110110110",
  38941=>"000101011",
  38942=>"000101101",
  38943=>"001011000",
  38944=>"100000001",
  38945=>"111111110",
  38946=>"100000000",
  38947=>"010110001",
  38948=>"100111111",
  38949=>"110010101",
  38950=>"100110000",
  38951=>"111001001",
  38952=>"001100100",
  38953=>"000111101",
  38954=>"010001111",
  38955=>"011110110",
  38956=>"001000101",
  38957=>"010001001",
  38958=>"111010010",
  38959=>"001011100",
  38960=>"110110110",
  38961=>"010000010",
  38962=>"111100100",
  38963=>"110110001",
  38964=>"111110111",
  38965=>"110101100",
  38966=>"000010100",
  38967=>"011101101",
  38968=>"000011000",
  38969=>"001000111",
  38970=>"000000101",
  38971=>"101001000",
  38972=>"000000011",
  38973=>"110011101",
  38974=>"101101011",
  38975=>"110111000",
  38976=>"100111011",
  38977=>"001001010",
  38978=>"111111100",
  38979=>"011101101",
  38980=>"100010001",
  38981=>"111011100",
  38982=>"001110101",
  38983=>"110110010",
  38984=>"010110001",
  38985=>"110000101",
  38986=>"101101110",
  38987=>"010001101",
  38988=>"111011010",
  38989=>"101000000",
  38990=>"111101101",
  38991=>"111100110",
  38992=>"011100110",
  38993=>"111110111",
  38994=>"111001001",
  38995=>"101111010",
  38996=>"001111110",
  38997=>"010101110",
  38998=>"010011111",
  38999=>"001111001",
  39000=>"001110100",
  39001=>"101011111",
  39002=>"011100001",
  39003=>"000110010",
  39004=>"001101111",
  39005=>"000001101",
  39006=>"010110010",
  39007=>"010000011",
  39008=>"000000101",
  39009=>"100101001",
  39010=>"011010100",
  39011=>"000100011",
  39012=>"100001010",
  39013=>"111000100",
  39014=>"100001000",
  39015=>"101101010",
  39016=>"101110001",
  39017=>"111101000",
  39018=>"110011101",
  39019=>"101110010",
  39020=>"010101101",
  39021=>"000001100",
  39022=>"101011011",
  39023=>"011010011",
  39024=>"101110101",
  39025=>"101010111",
  39026=>"110100110",
  39027=>"011110101",
  39028=>"011101000",
  39029=>"100110010",
  39030=>"111110111",
  39031=>"111011010",
  39032=>"001001111",
  39033=>"110000111",
  39034=>"101100110",
  39035=>"111111000",
  39036=>"001110011",
  39037=>"010010100",
  39038=>"011001111",
  39039=>"100100111",
  39040=>"001110000",
  39041=>"111111111",
  39042=>"111001001",
  39043=>"010010010",
  39044=>"100111111",
  39045=>"001100001",
  39046=>"010011001",
  39047=>"100111110",
  39048=>"100111111",
  39049=>"001000000",
  39050=>"010100000",
  39051=>"100001000",
  39052=>"110011011",
  39053=>"101100001",
  39054=>"110100111",
  39055=>"111110101",
  39056=>"001111110",
  39057=>"010101110",
  39058=>"010101000",
  39059=>"111101111",
  39060=>"110111011",
  39061=>"011111111",
  39062=>"000101001",
  39063=>"001100000",
  39064=>"111111111",
  39065=>"001111010",
  39066=>"100110110",
  39067=>"010100100",
  39068=>"101100000",
  39069=>"100011000",
  39070=>"101100101",
  39071=>"100001010",
  39072=>"100101000",
  39073=>"011101010",
  39074=>"110100010",
  39075=>"100110001",
  39076=>"111010111",
  39077=>"010011110",
  39078=>"111111111",
  39079=>"011110110",
  39080=>"001111001",
  39081=>"010001101",
  39082=>"100011010",
  39083=>"110111111",
  39084=>"101100011",
  39085=>"011100101",
  39086=>"110011011",
  39087=>"001111010",
  39088=>"011010000",
  39089=>"001000110",
  39090=>"101000010",
  39091=>"011011110",
  39092=>"011000011",
  39093=>"001000000",
  39094=>"000100010",
  39095=>"010010001",
  39096=>"100011101",
  39097=>"010000001",
  39098=>"010111000",
  39099=>"111001000",
  39100=>"000001000",
  39101=>"011110010",
  39102=>"110001000",
  39103=>"100110000",
  39104=>"001111001",
  39105=>"000000010",
  39106=>"010111101",
  39107=>"011000010",
  39108=>"001001110",
  39109=>"100111001",
  39110=>"010000110",
  39111=>"100101011",
  39112=>"001001011",
  39113=>"101111011",
  39114=>"010001110",
  39115=>"010010100",
  39116=>"110111010",
  39117=>"010001100",
  39118=>"000010100",
  39119=>"001000110",
  39120=>"000100100",
  39121=>"001000110",
  39122=>"000011101",
  39123=>"011001111",
  39124=>"101101001",
  39125=>"100101001",
  39126=>"011001111",
  39127=>"010000100",
  39128=>"101010100",
  39129=>"110010010",
  39130=>"111010001",
  39131=>"011100000",
  39132=>"011010100",
  39133=>"001010110",
  39134=>"101001001",
  39135=>"011011110",
  39136=>"001001011",
  39137=>"001111101",
  39138=>"100100110",
  39139=>"101001110",
  39140=>"111000111",
  39141=>"111010010",
  39142=>"101000110",
  39143=>"100000100",
  39144=>"100111101",
  39145=>"101001110",
  39146=>"001100011",
  39147=>"001001110",
  39148=>"010111010",
  39149=>"111010010",
  39150=>"111111100",
  39151=>"010011000",
  39152=>"100001101",
  39153=>"010100111",
  39154=>"110111101",
  39155=>"010111110",
  39156=>"111110011",
  39157=>"000110101",
  39158=>"110001000",
  39159=>"101010100",
  39160=>"011111011",
  39161=>"011011110",
  39162=>"000000000",
  39163=>"101001101",
  39164=>"100110001",
  39165=>"011110101",
  39166=>"011111010",
  39167=>"010101010",
  39168=>"101000011",
  39169=>"110011011",
  39170=>"100000001",
  39171=>"000110001",
  39172=>"001110011",
  39173=>"111011100",
  39174=>"000010100",
  39175=>"100100000",
  39176=>"000100010",
  39177=>"000001111",
  39178=>"101011010",
  39179=>"111100010",
  39180=>"001000011",
  39181=>"001101000",
  39182=>"000100010",
  39183=>"000100100",
  39184=>"111000110",
  39185=>"100001001",
  39186=>"010101111",
  39187=>"110010000",
  39188=>"001011110",
  39189=>"000110100",
  39190=>"010111011",
  39191=>"011101001",
  39192=>"011101011",
  39193=>"001001101",
  39194=>"000000000",
  39195=>"111001101",
  39196=>"110011000",
  39197=>"110101010",
  39198=>"101010101",
  39199=>"000011001",
  39200=>"100111000",
  39201=>"100000101",
  39202=>"000011000",
  39203=>"001101101",
  39204=>"101001001",
  39205=>"010000000",
  39206=>"110011011",
  39207=>"110010011",
  39208=>"101001110",
  39209=>"001100000",
  39210=>"010011001",
  39211=>"100000101",
  39212=>"100101000",
  39213=>"101110100",
  39214=>"001000100",
  39215=>"101011110",
  39216=>"111000000",
  39217=>"010111011",
  39218=>"001000000",
  39219=>"001001100",
  39220=>"010010001",
  39221=>"011100110",
  39222=>"101000010",
  39223=>"101010011",
  39224=>"100001001",
  39225=>"011110000",
  39226=>"100100000",
  39227=>"001000010",
  39228=>"011101101",
  39229=>"101011010",
  39230=>"111001101",
  39231=>"100000101",
  39232=>"001110100",
  39233=>"011000001",
  39234=>"101100011",
  39235=>"100110010",
  39236=>"110101111",
  39237=>"010110101",
  39238=>"101000011",
  39239=>"101111011",
  39240=>"111110011",
  39241=>"001001010",
  39242=>"000010110",
  39243=>"000011011",
  39244=>"110001010",
  39245=>"101011001",
  39246=>"110001000",
  39247=>"110010111",
  39248=>"001110001",
  39249=>"110101010",
  39250=>"100011110",
  39251=>"011100110",
  39252=>"010111000",
  39253=>"110000001",
  39254=>"101000010",
  39255=>"011011110",
  39256=>"111010011",
  39257=>"100100001",
  39258=>"101111101",
  39259=>"001011101",
  39260=>"000101111",
  39261=>"000111100",
  39262=>"101001111",
  39263=>"001100001",
  39264=>"111100101",
  39265=>"001011111",
  39266=>"000111110",
  39267=>"000101110",
  39268=>"001011111",
  39269=>"011100010",
  39270=>"011010011",
  39271=>"111111001",
  39272=>"110010010",
  39273=>"000001101",
  39274=>"011110111",
  39275=>"110011101",
  39276=>"100101011",
  39277=>"100110000",
  39278=>"001001000",
  39279=>"000101000",
  39280=>"001000010",
  39281=>"010011001",
  39282=>"100100000",
  39283=>"111111111",
  39284=>"001000010",
  39285=>"110011110",
  39286=>"100000011",
  39287=>"111101010",
  39288=>"100010101",
  39289=>"000011100",
  39290=>"110111100",
  39291=>"001111001",
  39292=>"100010100",
  39293=>"111010001",
  39294=>"011000000",
  39295=>"010000010",
  39296=>"100000101",
  39297=>"011110101",
  39298=>"101101000",
  39299=>"011110010",
  39300=>"010010111",
  39301=>"110100101",
  39302=>"001011010",
  39303=>"001000110",
  39304=>"011100001",
  39305=>"011110110",
  39306=>"000110101",
  39307=>"010111010",
  39308=>"010000001",
  39309=>"101111101",
  39310=>"000110101",
  39311=>"010110011",
  39312=>"011001110",
  39313=>"111111111",
  39314=>"111000111",
  39315=>"011110111",
  39316=>"110011101",
  39317=>"100010110",
  39318=>"001101100",
  39319=>"110000101",
  39320=>"000000101",
  39321=>"101010000",
  39322=>"001000111",
  39323=>"011000000",
  39324=>"100011011",
  39325=>"000101001",
  39326=>"101110000",
  39327=>"110110010",
  39328=>"111001111",
  39329=>"000000011",
  39330=>"000101111",
  39331=>"100011101",
  39332=>"111110101",
  39333=>"001010100",
  39334=>"110010100",
  39335=>"111000000",
  39336=>"110011111",
  39337=>"011001011",
  39338=>"001111000",
  39339=>"110100011",
  39340=>"101000011",
  39341=>"001111000",
  39342=>"010001000",
  39343=>"101000011",
  39344=>"000000100",
  39345=>"011010111",
  39346=>"111100000",
  39347=>"011001000",
  39348=>"000001111",
  39349=>"101101110",
  39350=>"100111110",
  39351=>"101101101",
  39352=>"101010000",
  39353=>"010001110",
  39354=>"101111011",
  39355=>"110111000",
  39356=>"010111110",
  39357=>"111100010",
  39358=>"011110110",
  39359=>"001001110",
  39360=>"111100010",
  39361=>"101000101",
  39362=>"101001010",
  39363=>"110001000",
  39364=>"000010011",
  39365=>"111000000",
  39366=>"010010001",
  39367=>"001101110",
  39368=>"011000111",
  39369=>"000000001",
  39370=>"110010001",
  39371=>"101101110",
  39372=>"100110100",
  39373=>"001010000",
  39374=>"000011010",
  39375=>"000101100",
  39376=>"100001000",
  39377=>"001111001",
  39378=>"001110111",
  39379=>"001001100",
  39380=>"111101111",
  39381=>"000011100",
  39382=>"100011001",
  39383=>"100001000",
  39384=>"001010011",
  39385=>"110001011",
  39386=>"110111111",
  39387=>"101111110",
  39388=>"000110011",
  39389=>"100011000",
  39390=>"100110011",
  39391=>"100011011",
  39392=>"100101101",
  39393=>"111011101",
  39394=>"111110110",
  39395=>"111011100",
  39396=>"101000101",
  39397=>"101110011",
  39398=>"110100001",
  39399=>"001010010",
  39400=>"111011111",
  39401=>"011110000",
  39402=>"000110100",
  39403=>"111010110",
  39404=>"000010010",
  39405=>"001000000",
  39406=>"111010110",
  39407=>"011001111",
  39408=>"010010011",
  39409=>"111001110",
  39410=>"011000000",
  39411=>"000101001",
  39412=>"000111010",
  39413=>"000010010",
  39414=>"101001000",
  39415=>"010110110",
  39416=>"000101111",
  39417=>"001011110",
  39418=>"101101011",
  39419=>"110001001",
  39420=>"001001101",
  39421=>"111101001",
  39422=>"101110011",
  39423=>"101111010",
  39424=>"100010101",
  39425=>"011100100",
  39426=>"100110000",
  39427=>"101001100",
  39428=>"000101101",
  39429=>"111110001",
  39430=>"011000010",
  39431=>"011110110",
  39432=>"001000000",
  39433=>"111011101",
  39434=>"001111000",
  39435=>"001100100",
  39436=>"010100000",
  39437=>"100100000",
  39438=>"000001001",
  39439=>"011111000",
  39440=>"111111001",
  39441=>"110011100",
  39442=>"100110111",
  39443=>"111101001",
  39444=>"100100100",
  39445=>"110101001",
  39446=>"000100100",
  39447=>"101100011",
  39448=>"001101000",
  39449=>"101101000",
  39450=>"010110011",
  39451=>"111000010",
  39452=>"111011101",
  39453=>"111111111",
  39454=>"000100010",
  39455=>"011100010",
  39456=>"000000011",
  39457=>"111111010",
  39458=>"001000001",
  39459=>"011000010",
  39460=>"010010110",
  39461=>"011000001",
  39462=>"110001010",
  39463=>"100101000",
  39464=>"000100110",
  39465=>"111111100",
  39466=>"100100000",
  39467=>"101011100",
  39468=>"101011011",
  39469=>"001001000",
  39470=>"000101111",
  39471=>"001101011",
  39472=>"001101010",
  39473=>"110100100",
  39474=>"111000111",
  39475=>"110100011",
  39476=>"010011010",
  39477=>"001110100",
  39478=>"010111110",
  39479=>"001111110",
  39480=>"010101001",
  39481=>"011001000",
  39482=>"000001100",
  39483=>"110100010",
  39484=>"101110010",
  39485=>"010101111",
  39486=>"001111101",
  39487=>"110001100",
  39488=>"110110000",
  39489=>"111100110",
  39490=>"011100011",
  39491=>"011000001",
  39492=>"001101000",
  39493=>"101101100",
  39494=>"110111010",
  39495=>"000011101",
  39496=>"110100101",
  39497=>"001000001",
  39498=>"001011111",
  39499=>"011011001",
  39500=>"111000010",
  39501=>"100001010",
  39502=>"111010000",
  39503=>"100110100",
  39504=>"111101101",
  39505=>"110011001",
  39506=>"101100100",
  39507=>"110101110",
  39508=>"111000101",
  39509=>"011010101",
  39510=>"011011101",
  39511=>"001100111",
  39512=>"010000001",
  39513=>"100001101",
  39514=>"000110101",
  39515=>"011111000",
  39516=>"101111110",
  39517=>"011001100",
  39518=>"001110110",
  39519=>"100111000",
  39520=>"000000010",
  39521=>"110111001",
  39522=>"010011100",
  39523=>"001111010",
  39524=>"011010000",
  39525=>"111011100",
  39526=>"010101011",
  39527=>"110010000",
  39528=>"011110110",
  39529=>"110100110",
  39530=>"011100010",
  39531=>"111000101",
  39532=>"101010011",
  39533=>"100111011",
  39534=>"010110011",
  39535=>"100110011",
  39536=>"110001110",
  39537=>"011001000",
  39538=>"000101100",
  39539=>"111110000",
  39540=>"111001100",
  39541=>"101000000",
  39542=>"011010000",
  39543=>"111010011",
  39544=>"110000101",
  39545=>"011001101",
  39546=>"001100100",
  39547=>"001101011",
  39548=>"110110100",
  39549=>"001000100",
  39550=>"111111110",
  39551=>"000001111",
  39552=>"101110110",
  39553=>"010110100",
  39554=>"110010110",
  39555=>"000000001",
  39556=>"001110110",
  39557=>"011011011",
  39558=>"101110101",
  39559=>"011010100",
  39560=>"011100011",
  39561=>"111001001",
  39562=>"011110011",
  39563=>"011011111",
  39564=>"100100011",
  39565=>"110111100",
  39566=>"111010001",
  39567=>"110111111",
  39568=>"111110101",
  39569=>"010011001",
  39570=>"100110001",
  39571=>"001100111",
  39572=>"000010101",
  39573=>"110100111",
  39574=>"000001001",
  39575=>"110101110",
  39576=>"010000010",
  39577=>"111111111",
  39578=>"110001110",
  39579=>"011111111",
  39580=>"100011111",
  39581=>"000010010",
  39582=>"111110100",
  39583=>"000110001",
  39584=>"111100101",
  39585=>"101001000",
  39586=>"011101011",
  39587=>"110010000",
  39588=>"100101001",
  39589=>"111000111",
  39590=>"110100101",
  39591=>"010100000",
  39592=>"000100001",
  39593=>"101011111",
  39594=>"101101100",
  39595=>"100010111",
  39596=>"001001110",
  39597=>"001010111",
  39598=>"001010000",
  39599=>"111010000",
  39600=>"011100110",
  39601=>"101001001",
  39602=>"011010010",
  39603=>"000101101",
  39604=>"100100000",
  39605=>"010100001",
  39606=>"111110101",
  39607=>"101000100",
  39608=>"011110111",
  39609=>"000100111",
  39610=>"111111100",
  39611=>"000101111",
  39612=>"110110110",
  39613=>"110011000",
  39614=>"000010001",
  39615=>"101000010",
  39616=>"100101000",
  39617=>"100011111",
  39618=>"011111001",
  39619=>"001001001",
  39620=>"000011100",
  39621=>"011101111",
  39622=>"100111010",
  39623=>"000100000",
  39624=>"100100000",
  39625=>"011000111",
  39626=>"111111111",
  39627=>"110110011",
  39628=>"011111101",
  39629=>"101001011",
  39630=>"110110111",
  39631=>"010100110",
  39632=>"000011101",
  39633=>"001100111",
  39634=>"010100000",
  39635=>"010100000",
  39636=>"111110001",
  39637=>"101000111",
  39638=>"110000011",
  39639=>"110111110",
  39640=>"000100000",
  39641=>"101001011",
  39642=>"111001100",
  39643=>"011101101",
  39644=>"100000101",
  39645=>"000001010",
  39646=>"000110010",
  39647=>"100011011",
  39648=>"101010000",
  39649=>"010011100",
  39650=>"001011000",
  39651=>"011101010",
  39652=>"101100111",
  39653=>"011011011",
  39654=>"001000001",
  39655=>"100010110",
  39656=>"010101111",
  39657=>"110011000",
  39658=>"000000010",
  39659=>"110011111",
  39660=>"000110000",
  39661=>"100000101",
  39662=>"010111011",
  39663=>"100110100",
  39664=>"100001001",
  39665=>"110101010",
  39666=>"011110110",
  39667=>"101111010",
  39668=>"111111110",
  39669=>"110100111",
  39670=>"100001100",
  39671=>"100001101",
  39672=>"101011101",
  39673=>"100011101",
  39674=>"000111001",
  39675=>"100110011",
  39676=>"101010101",
  39677=>"010010010",
  39678=>"110110101",
  39679=>"000001010",
  39680=>"110000000",
  39681=>"000000011",
  39682=>"110101010",
  39683=>"100011111",
  39684=>"100111101",
  39685=>"111111100",
  39686=>"001000011",
  39687=>"001111111",
  39688=>"000010001",
  39689=>"010001001",
  39690=>"011111010",
  39691=>"000000010",
  39692=>"000000000",
  39693=>"011110011",
  39694=>"110111011",
  39695=>"011001110",
  39696=>"101011110",
  39697=>"100000100",
  39698=>"101111001",
  39699=>"011010011",
  39700=>"100001110",
  39701=>"010101000",
  39702=>"111100110",
  39703=>"010111011",
  39704=>"010010010",
  39705=>"100010010",
  39706=>"111111010",
  39707=>"010011011",
  39708=>"100101100",
  39709=>"110011010",
  39710=>"011000101",
  39711=>"111101111",
  39712=>"010000110",
  39713=>"111100100",
  39714=>"001010100",
  39715=>"110100110",
  39716=>"110100000",
  39717=>"111011111",
  39718=>"110011001",
  39719=>"111000000",
  39720=>"010000000",
  39721=>"000111100",
  39722=>"110100010",
  39723=>"111101111",
  39724=>"010010010",
  39725=>"000100110",
  39726=>"000001011",
  39727=>"110110111",
  39728=>"100101011",
  39729=>"010110101",
  39730=>"100100001",
  39731=>"000111111",
  39732=>"000111000",
  39733=>"100001111",
  39734=>"100011111",
  39735=>"001111010",
  39736=>"111000110",
  39737=>"100100011",
  39738=>"010111000",
  39739=>"011001010",
  39740=>"000001010",
  39741=>"101101000",
  39742=>"001101011",
  39743=>"111000010",
  39744=>"010011011",
  39745=>"011000001",
  39746=>"111111011",
  39747=>"010100001",
  39748=>"100101100",
  39749=>"100101000",
  39750=>"001111101",
  39751=>"110100000",
  39752=>"011010001",
  39753=>"010110111",
  39754=>"010101000",
  39755=>"100100101",
  39756=>"010100100",
  39757=>"111000011",
  39758=>"001010110",
  39759=>"001101000",
  39760=>"110101111",
  39761=>"101000011",
  39762=>"000111100",
  39763=>"111110101",
  39764=>"010010011",
  39765=>"000011010",
  39766=>"010101000",
  39767=>"000000111",
  39768=>"111100000",
  39769=>"011110110",
  39770=>"111000110",
  39771=>"100001001",
  39772=>"111111000",
  39773=>"111000000",
  39774=>"101100111",
  39775=>"100111100",
  39776=>"000100011",
  39777=>"000011001",
  39778=>"011111100",
  39779=>"000001100",
  39780=>"110100100",
  39781=>"111100011",
  39782=>"101001010",
  39783=>"001110101",
  39784=>"010010000",
  39785=>"100000000",
  39786=>"011101011",
  39787=>"110010000",
  39788=>"111110101",
  39789=>"100001010",
  39790=>"111100111",
  39791=>"011100110",
  39792=>"110000111",
  39793=>"111110011",
  39794=>"000011001",
  39795=>"011110001",
  39796=>"010010000",
  39797=>"101011100",
  39798=>"100010111",
  39799=>"111001100",
  39800=>"010011111",
  39801=>"110001001",
  39802=>"100010010",
  39803=>"111010111",
  39804=>"011000100",
  39805=>"011010011",
  39806=>"101110111",
  39807=>"101010001",
  39808=>"000110111",
  39809=>"101011011",
  39810=>"000011000",
  39811=>"010010011",
  39812=>"000000111",
  39813=>"110001001",
  39814=>"010101001",
  39815=>"011100001",
  39816=>"000010110",
  39817=>"001101101",
  39818=>"001000000",
  39819=>"111011000",
  39820=>"111111110",
  39821=>"001111010",
  39822=>"101000000",
  39823=>"100000010",
  39824=>"011010101",
  39825=>"111010001",
  39826=>"000101100",
  39827=>"110011101",
  39828=>"011011011",
  39829=>"000010011",
  39830=>"001010010",
  39831=>"110001001",
  39832=>"111011010",
  39833=>"100000101",
  39834=>"001001111",
  39835=>"010001100",
  39836=>"000010000",
  39837=>"001001011",
  39838=>"000010010",
  39839=>"111001001",
  39840=>"000010111",
  39841=>"100100000",
  39842=>"001001000",
  39843=>"110110101",
  39844=>"001011001",
  39845=>"111101000",
  39846=>"000010010",
  39847=>"010010100",
  39848=>"011001101",
  39849=>"110101000",
  39850=>"111100111",
  39851=>"001011001",
  39852=>"000010110",
  39853=>"100110100",
  39854=>"011111101",
  39855=>"001000110",
  39856=>"011000101",
  39857=>"111011111",
  39858=>"010010001",
  39859=>"011010000",
  39860=>"000010010",
  39861=>"011100001",
  39862=>"111011100",
  39863=>"111110010",
  39864=>"111111011",
  39865=>"000001011",
  39866=>"111001100",
  39867=>"010110000",
  39868=>"010110001",
  39869=>"101100111",
  39870=>"101101110",
  39871=>"001000001",
  39872=>"111000100",
  39873=>"011101111",
  39874=>"111111110",
  39875=>"100010001",
  39876=>"010101000",
  39877=>"101100100",
  39878=>"111100101",
  39879=>"011011000",
  39880=>"010010000",
  39881=>"000010000",
  39882=>"111101100",
  39883=>"111100011",
  39884=>"110100010",
  39885=>"001100111",
  39886=>"010001000",
  39887=>"101001111",
  39888=>"001110111",
  39889=>"000100100",
  39890=>"110011101",
  39891=>"001001000",
  39892=>"010110000",
  39893=>"001100000",
  39894=>"101110011",
  39895=>"011100100",
  39896=>"001100111",
  39897=>"001000011",
  39898=>"001011101",
  39899=>"101100100",
  39900=>"110010001",
  39901=>"110010101",
  39902=>"111100001",
  39903=>"101000010",
  39904=>"111000010",
  39905=>"000010000",
  39906=>"010001100",
  39907=>"011111010",
  39908=>"101111100",
  39909=>"100000100",
  39910=>"110101110",
  39911=>"100110111",
  39912=>"001000000",
  39913=>"100010001",
  39914=>"001110111",
  39915=>"110101110",
  39916=>"001111000",
  39917=>"101100011",
  39918=>"011000101",
  39919=>"010001011",
  39920=>"101001011",
  39921=>"011100110",
  39922=>"001110101",
  39923=>"000101001",
  39924=>"100100000",
  39925=>"001100011",
  39926=>"110000011",
  39927=>"001100111",
  39928=>"100010000",
  39929=>"111000001",
  39930=>"010111110",
  39931=>"100100110",
  39932=>"000010001",
  39933=>"110010001",
  39934=>"111011010",
  39935=>"111111011",
  39936=>"011110001",
  39937=>"010010110",
  39938=>"111101110",
  39939=>"111010110",
  39940=>"011010011",
  39941=>"100111111",
  39942=>"000011011",
  39943=>"000100000",
  39944=>"010101001",
  39945=>"110010100",
  39946=>"000011111",
  39947=>"110100001",
  39948=>"001000001",
  39949=>"110110000",
  39950=>"001101000",
  39951=>"010110000",
  39952=>"100100100",
  39953=>"100011110",
  39954=>"010010100",
  39955=>"101111101",
  39956=>"011110110",
  39957=>"010101111",
  39958=>"111101100",
  39959=>"010100110",
  39960=>"010010010",
  39961=>"000010000",
  39962=>"100010000",
  39963=>"100100000",
  39964=>"011110111",
  39965=>"100001000",
  39966=>"011111111",
  39967=>"111111101",
  39968=>"101100100",
  39969=>"001111000",
  39970=>"101010011",
  39971=>"110100000",
  39972=>"011001000",
  39973=>"101110001",
  39974=>"000000110",
  39975=>"000100011",
  39976=>"001110011",
  39977=>"000001111",
  39978=>"001000100",
  39979=>"000000010",
  39980=>"000010000",
  39981=>"100101110",
  39982=>"000110011",
  39983=>"000100101",
  39984=>"110000010",
  39985=>"101011001",
  39986=>"001011010",
  39987=>"100111100",
  39988=>"101111010",
  39989=>"011001101",
  39990=>"010100110",
  39991=>"100101100",
  39992=>"011100101",
  39993=>"111000010",
  39994=>"011010101",
  39995=>"011101101",
  39996=>"011001001",
  39997=>"100011100",
  39998=>"111101000",
  39999=>"100001011",
  40000=>"111000111",
  40001=>"001111000",
  40002=>"010011101",
  40003=>"001011101",
  40004=>"010110111",
  40005=>"100010001",
  40006=>"011100000",
  40007=>"100001001",
  40008=>"101110100",
  40009=>"110010010",
  40010=>"101111001",
  40011=>"011110100",
  40012=>"100111000",
  40013=>"011100001",
  40014=>"101111000",
  40015=>"010111111",
  40016=>"110000011",
  40017=>"001110100",
  40018=>"011101010",
  40019=>"010011010",
  40020=>"010100101",
  40021=>"010001010",
  40022=>"100001101",
  40023=>"001000110",
  40024=>"000000000",
  40025=>"111101011",
  40026=>"100010100",
  40027=>"000101100",
  40028=>"101100011",
  40029=>"000100001",
  40030=>"011000110",
  40031=>"110101010",
  40032=>"011100111",
  40033=>"110100111",
  40034=>"000001101",
  40035=>"000000101",
  40036=>"010110010",
  40037=>"100101000",
  40038=>"010101001",
  40039=>"100101011",
  40040=>"000101001",
  40041=>"011010111",
  40042=>"000010011",
  40043=>"010101001",
  40044=>"101001100",
  40045=>"001001001",
  40046=>"000000000",
  40047=>"000011001",
  40048=>"000011111",
  40049=>"001010010",
  40050=>"011011111",
  40051=>"110100010",
  40052=>"101110011",
  40053=>"001000010",
  40054=>"111011000",
  40055=>"100101111",
  40056=>"101110110",
  40057=>"000010101",
  40058=>"010011011",
  40059=>"110100100",
  40060=>"110010010",
  40061=>"010100010",
  40062=>"110110000",
  40063=>"100000000",
  40064=>"101101100",
  40065=>"001001010",
  40066=>"101100001",
  40067=>"001001001",
  40068=>"010011000",
  40069=>"110011111",
  40070=>"010101001",
  40071=>"010010101",
  40072=>"100011111",
  40073=>"111011011",
  40074=>"101111010",
  40075=>"001011000",
  40076=>"000111001",
  40077=>"001101100",
  40078=>"001100010",
  40079=>"100001011",
  40080=>"001001100",
  40081=>"110111100",
  40082=>"111111010",
  40083=>"101000011",
  40084=>"011000110",
  40085=>"001000001",
  40086=>"100100111",
  40087=>"011100100",
  40088=>"010001010",
  40089=>"010011011",
  40090=>"111110111",
  40091=>"101011010",
  40092=>"011000101",
  40093=>"010001100",
  40094=>"011110111",
  40095=>"001101011",
  40096=>"110001000",
  40097=>"011001010",
  40098=>"001001110",
  40099=>"010001001",
  40100=>"010111101",
  40101=>"011000000",
  40102=>"100100010",
  40103=>"101101011",
  40104=>"000001111",
  40105=>"010010001",
  40106=>"111111101",
  40107=>"011011011",
  40108=>"010011010",
  40109=>"100110011",
  40110=>"000111001",
  40111=>"000111110",
  40112=>"110011100",
  40113=>"000010110",
  40114=>"101011110",
  40115=>"011111100",
  40116=>"010110000",
  40117=>"101010000",
  40118=>"111001010",
  40119=>"000000000",
  40120=>"001001011",
  40121=>"011011011",
  40122=>"111010001",
  40123=>"000101111",
  40124=>"110000000",
  40125=>"101111110",
  40126=>"000110001",
  40127=>"000110000",
  40128=>"010010110",
  40129=>"000000011",
  40130=>"100100010",
  40131=>"101010101",
  40132=>"110101101",
  40133=>"010011001",
  40134=>"111110001",
  40135=>"001001111",
  40136=>"010101000",
  40137=>"101110000",
  40138=>"010011101",
  40139=>"111011000",
  40140=>"010111000",
  40141=>"111110010",
  40142=>"010101110",
  40143=>"110101111",
  40144=>"001111010",
  40145=>"000101001",
  40146=>"010100100",
  40147=>"011000001",
  40148=>"111101001",
  40149=>"100001010",
  40150=>"000000000",
  40151=>"000111010",
  40152=>"110110101",
  40153=>"101110000",
  40154=>"111101001",
  40155=>"000000100",
  40156=>"010101101",
  40157=>"110101000",
  40158=>"011100011",
  40159=>"000110011",
  40160=>"111110011",
  40161=>"001010110",
  40162=>"101010101",
  40163=>"001001001",
  40164=>"101111010",
  40165=>"111101010",
  40166=>"111010110",
  40167=>"001011110",
  40168=>"100101100",
  40169=>"110001100",
  40170=>"100000110",
  40171=>"001011110",
  40172=>"001010000",
  40173=>"011111100",
  40174=>"011110100",
  40175=>"111010110",
  40176=>"100110101",
  40177=>"011011001",
  40178=>"000110110",
  40179=>"000000100",
  40180=>"110110100",
  40181=>"110011010",
  40182=>"000010011",
  40183=>"001101000",
  40184=>"111101010",
  40185=>"110001000",
  40186=>"000111100",
  40187=>"000100100",
  40188=>"101001001",
  40189=>"000011110",
  40190=>"100010111",
  40191=>"101111110",
  40192=>"100011101",
  40193=>"000101001",
  40194=>"010100110",
  40195=>"011100111",
  40196=>"101011101",
  40197=>"100001101",
  40198=>"101010101",
  40199=>"010111101",
  40200=>"100100111",
  40201=>"100000001",
  40202=>"101001100",
  40203=>"111000010",
  40204=>"111101101",
  40205=>"010100111",
  40206=>"001100011",
  40207=>"001111011",
  40208=>"100111110",
  40209=>"111010100",
  40210=>"101010100",
  40211=>"001010000",
  40212=>"000001100",
  40213=>"101011110",
  40214=>"111001100",
  40215=>"000000100",
  40216=>"101001001",
  40217=>"001100000",
  40218=>"110000011",
  40219=>"100101000",
  40220=>"000100010",
  40221=>"011011001",
  40222=>"010011111",
  40223=>"011100110",
  40224=>"100001011",
  40225=>"101000110",
  40226=>"111001011",
  40227=>"001101111",
  40228=>"111001010",
  40229=>"111101111",
  40230=>"001010100",
  40231=>"100110001",
  40232=>"011010111",
  40233=>"101101010",
  40234=>"000100110",
  40235=>"111010000",
  40236=>"000011101",
  40237=>"000000010",
  40238=>"000000000",
  40239=>"001011101",
  40240=>"011011001",
  40241=>"010000111",
  40242=>"011100101",
  40243=>"100011001",
  40244=>"101101001",
  40245=>"010100100",
  40246=>"101100101",
  40247=>"111010000",
  40248=>"111111111",
  40249=>"111010100",
  40250=>"001110111",
  40251=>"110111010",
  40252=>"101011100",
  40253=>"110000110",
  40254=>"110001001",
  40255=>"111111111",
  40256=>"001011101",
  40257=>"110101110",
  40258=>"110111010",
  40259=>"100000010",
  40260=>"111100011",
  40261=>"011011100",
  40262=>"000101010",
  40263=>"110010100",
  40264=>"010011111",
  40265=>"000011101",
  40266=>"101101000",
  40267=>"011001000",
  40268=>"011100011",
  40269=>"001010010",
  40270=>"111101011",
  40271=>"001111111",
  40272=>"100011011",
  40273=>"010100000",
  40274=>"111010000",
  40275=>"100110001",
  40276=>"101111000",
  40277=>"010001011",
  40278=>"000000010",
  40279=>"000100010",
  40280=>"011000111",
  40281=>"001101000",
  40282=>"110110010",
  40283=>"101001101",
  40284=>"010001111",
  40285=>"100101100",
  40286=>"010011100",
  40287=>"001101101",
  40288=>"000000110",
  40289=>"011011011",
  40290=>"011111100",
  40291=>"010101001",
  40292=>"101100000",
  40293=>"010100000",
  40294=>"101011011",
  40295=>"011101101",
  40296=>"010011100",
  40297=>"000000000",
  40298=>"101101001",
  40299=>"000001000",
  40300=>"011010101",
  40301=>"000101101",
  40302=>"001011000",
  40303=>"011010011",
  40304=>"010011110",
  40305=>"000011010",
  40306=>"101001100",
  40307=>"111110100",
  40308=>"111100001",
  40309=>"111001100",
  40310=>"111010110",
  40311=>"111101101",
  40312=>"100010100",
  40313=>"011111100",
  40314=>"011100000",
  40315=>"010011011",
  40316=>"111011111",
  40317=>"001001010",
  40318=>"110110000",
  40319=>"000001101",
  40320=>"100010101",
  40321=>"100110011",
  40322=>"101110111",
  40323=>"100011010",
  40324=>"010100100",
  40325=>"011111110",
  40326=>"011100111",
  40327=>"111101100",
  40328=>"101100001",
  40329=>"111011011",
  40330=>"010000010",
  40331=>"100110101",
  40332=>"001001011",
  40333=>"110110101",
  40334=>"100011110",
  40335=>"111111000",
  40336=>"011110000",
  40337=>"000100100",
  40338=>"100011001",
  40339=>"111011111",
  40340=>"000010110",
  40341=>"011100001",
  40342=>"010001101",
  40343=>"001011011",
  40344=>"100001111",
  40345=>"100111011",
  40346=>"000111100",
  40347=>"011100100",
  40348=>"001000001",
  40349=>"000010001",
  40350=>"110011101",
  40351=>"000011010",
  40352=>"000001100",
  40353=>"000110111",
  40354=>"100111110",
  40355=>"100111011",
  40356=>"110010111",
  40357=>"110100011",
  40358=>"111001100",
  40359=>"001000000",
  40360=>"000011110",
  40361=>"110010000",
  40362=>"011101001",
  40363=>"111101000",
  40364=>"001011111",
  40365=>"110011110",
  40366=>"010011000",
  40367=>"100111101",
  40368=>"110011011",
  40369=>"000010100",
  40370=>"111111100",
  40371=>"000111001",
  40372=>"100111101",
  40373=>"101010011",
  40374=>"101101100",
  40375=>"101100111",
  40376=>"000000010",
  40377=>"101111010",
  40378=>"010110000",
  40379=>"010011001",
  40380=>"101111001",
  40381=>"001101100",
  40382=>"111111010",
  40383=>"101111000",
  40384=>"000001011",
  40385=>"111010111",
  40386=>"001111110",
  40387=>"100011111",
  40388=>"100110111",
  40389=>"001001011",
  40390=>"110100001",
  40391=>"111111011",
  40392=>"100111001",
  40393=>"011100011",
  40394=>"110110011",
  40395=>"000100010",
  40396=>"001101000",
  40397=>"010110101",
  40398=>"100111010",
  40399=>"110010100",
  40400=>"111110110",
  40401=>"100110011",
  40402=>"011010001",
  40403=>"100111111",
  40404=>"111100000",
  40405=>"101000110",
  40406=>"001111011",
  40407=>"100001000",
  40408=>"000000011",
  40409=>"111011111",
  40410=>"110001111",
  40411=>"101011101",
  40412=>"010110111",
  40413=>"110000111",
  40414=>"000110111",
  40415=>"010111010",
  40416=>"111111101",
  40417=>"101001000",
  40418=>"101100100",
  40419=>"111001011",
  40420=>"001111110",
  40421=>"100011111",
  40422=>"010001100",
  40423=>"101110111",
  40424=>"000001101",
  40425=>"100100110",
  40426=>"010101000",
  40427=>"001100110",
  40428=>"111101111",
  40429=>"100011110",
  40430=>"101001101",
  40431=>"101110110",
  40432=>"011101011",
  40433=>"101011000",
  40434=>"111111010",
  40435=>"000010110",
  40436=>"010010001",
  40437=>"100011001",
  40438=>"110011101",
  40439=>"100010001",
  40440=>"101101111",
  40441=>"010011101",
  40442=>"011101011",
  40443=>"000100111",
  40444=>"110011001",
  40445=>"111100000",
  40446=>"001100000",
  40447=>"000010111",
  40448=>"000101110",
  40449=>"000001000",
  40450=>"001111010",
  40451=>"010010110",
  40452=>"000000111",
  40453=>"011000000",
  40454=>"001010100",
  40455=>"101010001",
  40456=>"010010010",
  40457=>"011011001",
  40458=>"111110100",
  40459=>"000000101",
  40460=>"111010110",
  40461=>"100011111",
  40462=>"000010000",
  40463=>"101110001",
  40464=>"101111111",
  40465=>"110011100",
  40466=>"011111011",
  40467=>"110110011",
  40468=>"011100000",
  40469=>"100010001",
  40470=>"010101011",
  40471=>"010111010",
  40472=>"101100110",
  40473=>"010101101",
  40474=>"000001001",
  40475=>"001100110",
  40476=>"010010000",
  40477=>"100110000",
  40478=>"011100100",
  40479=>"110011011",
  40480=>"000001111",
  40481=>"111001110",
  40482=>"010001111",
  40483=>"111100100",
  40484=>"110010010",
  40485=>"110101000",
  40486=>"100110110",
  40487=>"011111000",
  40488=>"000100100",
  40489=>"101000110",
  40490=>"111000100",
  40491=>"100111001",
  40492=>"010001011",
  40493=>"101111000",
  40494=>"010000001",
  40495=>"011010001",
  40496=>"000011111",
  40497=>"110110101",
  40498=>"010001111",
  40499=>"110101101",
  40500=>"001111011",
  40501=>"111111111",
  40502=>"010100111",
  40503=>"100011000",
  40504=>"100011010",
  40505=>"110111010",
  40506=>"101001100",
  40507=>"011111011",
  40508=>"101110111",
  40509=>"101110110",
  40510=>"111110111",
  40511=>"011101001",
  40512=>"000001100",
  40513=>"100011111",
  40514=>"010000111",
  40515=>"000010101",
  40516=>"001100100",
  40517=>"101001111",
  40518=>"000001000",
  40519=>"101001111",
  40520=>"111100101",
  40521=>"001100011",
  40522=>"010111011",
  40523=>"111111100",
  40524=>"100010001",
  40525=>"010110001",
  40526=>"011010001",
  40527=>"100010001",
  40528=>"100001000",
  40529=>"100011011",
  40530=>"010010010",
  40531=>"000010010",
  40532=>"000110000",
  40533=>"000110101",
  40534=>"101011000",
  40535=>"011110100",
  40536=>"000001001",
  40537=>"101000100",
  40538=>"111111111",
  40539=>"110101110",
  40540=>"001110001",
  40541=>"110111000",
  40542=>"000111111",
  40543=>"001001100",
  40544=>"110000100",
  40545=>"011011001",
  40546=>"000010111",
  40547=>"111011110",
  40548=>"111000110",
  40549=>"111010110",
  40550=>"010101111",
  40551=>"000000100",
  40552=>"001000101",
  40553=>"001000001",
  40554=>"011111001",
  40555=>"010010000",
  40556=>"101000101",
  40557=>"010010101",
  40558=>"001011001",
  40559=>"001011110",
  40560=>"011101110",
  40561=>"001111111",
  40562=>"001110011",
  40563=>"011110000",
  40564=>"101001100",
  40565=>"010110010",
  40566=>"001011000",
  40567=>"111010110",
  40568=>"101110100",
  40569=>"100011100",
  40570=>"100010111",
  40571=>"111011101",
  40572=>"010011110",
  40573=>"011111011",
  40574=>"011001010",
  40575=>"011001001",
  40576=>"100011101",
  40577=>"101000111",
  40578=>"100000101",
  40579=>"111001101",
  40580=>"111101110",
  40581=>"100000101",
  40582=>"000011111",
  40583=>"101000000",
  40584=>"111000100",
  40585=>"000001101",
  40586=>"011111101",
  40587=>"101110001",
  40588=>"000001101",
  40589=>"011011111",
  40590=>"101111111",
  40591=>"011100000",
  40592=>"101100110",
  40593=>"001000110",
  40594=>"101001000",
  40595=>"100100011",
  40596=>"100111100",
  40597=>"111110001",
  40598=>"111111111",
  40599=>"000100001",
  40600=>"010010111",
  40601=>"101110001",
  40602=>"111001100",
  40603=>"110110001",
  40604=>"010111100",
  40605=>"100010100",
  40606=>"100101001",
  40607=>"001101000",
  40608=>"111001010",
  40609=>"111101000",
  40610=>"111011110",
  40611=>"010111011",
  40612=>"000111010",
  40613=>"111110101",
  40614=>"111111010",
  40615=>"101101001",
  40616=>"110000100",
  40617=>"010000100",
  40618=>"001111010",
  40619=>"000100010",
  40620=>"010111111",
  40621=>"110000100",
  40622=>"101100001",
  40623=>"101110100",
  40624=>"100011011",
  40625=>"111100001",
  40626=>"111111001",
  40627=>"101111101",
  40628=>"111101000",
  40629=>"110000011",
  40630=>"000110111",
  40631=>"100011000",
  40632=>"110111001",
  40633=>"001010001",
  40634=>"010000000",
  40635=>"011000001",
  40636=>"001110111",
  40637=>"101111000",
  40638=>"111110001",
  40639=>"111100100",
  40640=>"101100011",
  40641=>"001111111",
  40642=>"101110111",
  40643=>"010010101",
  40644=>"011111110",
  40645=>"011111011",
  40646=>"000001010",
  40647=>"111010100",
  40648=>"101101010",
  40649=>"000011010",
  40650=>"101111100",
  40651=>"101111001",
  40652=>"011110011",
  40653=>"101111111",
  40654=>"001111100",
  40655=>"100011011",
  40656=>"011010101",
  40657=>"011101111",
  40658=>"011111011",
  40659=>"100111110",
  40660=>"100110011",
  40661=>"010011101",
  40662=>"111011100",
  40663=>"110111000",
  40664=>"110001001",
  40665=>"010111100",
  40666=>"011101000",
  40667=>"110100110",
  40668=>"111110010",
  40669=>"100001110",
  40670=>"000111110",
  40671=>"010001101",
  40672=>"000000100",
  40673=>"010000110",
  40674=>"111110101",
  40675=>"101111001",
  40676=>"010100110",
  40677=>"100001101",
  40678=>"010111000",
  40679=>"011010000",
  40680=>"001111100",
  40681=>"010010010",
  40682=>"110001000",
  40683=>"111011111",
  40684=>"101111011",
  40685=>"101111111",
  40686=>"101000000",
  40687=>"011010011",
  40688=>"111101010",
  40689=>"100001001",
  40690=>"111011111",
  40691=>"011111011",
  40692=>"010111111",
  40693=>"111011011",
  40694=>"000000001",
  40695=>"011110001",
  40696=>"001001000",
  40697=>"011010101",
  40698=>"101101001",
  40699=>"110110010",
  40700=>"100111110",
  40701=>"000000010",
  40702=>"100000011",
  40703=>"110010010",
  40704=>"001111001",
  40705=>"001110000",
  40706=>"111011101",
  40707=>"010001001",
  40708=>"101110101",
  40709=>"110011100",
  40710=>"110000110",
  40711=>"111101100",
  40712=>"111011111",
  40713=>"010101010",
  40714=>"011110001",
  40715=>"010001111",
  40716=>"100010000",
  40717=>"100111000",
  40718=>"110010000",
  40719=>"010011101",
  40720=>"001101100",
  40721=>"010100011",
  40722=>"011101000",
  40723=>"111001100",
  40724=>"110011100",
  40725=>"111010011",
  40726=>"111111101",
  40727=>"001001101",
  40728=>"111100110",
  40729=>"110000000",
  40730=>"100111101",
  40731=>"001000111",
  40732=>"010101000",
  40733=>"010001101",
  40734=>"100010010",
  40735=>"110101100",
  40736=>"101101111",
  40737=>"010010100",
  40738=>"011101101",
  40739=>"110100010",
  40740=>"000000000",
  40741=>"100001100",
  40742=>"010100100",
  40743=>"100101100",
  40744=>"011011110",
  40745=>"110001010",
  40746=>"111000110",
  40747=>"111100011",
  40748=>"100111110",
  40749=>"100001010",
  40750=>"001010111",
  40751=>"010100000",
  40752=>"001010100",
  40753=>"000100010",
  40754=>"101000101",
  40755=>"010010000",
  40756=>"000100110",
  40757=>"000001010",
  40758=>"000010011",
  40759=>"010000011",
  40760=>"111010000",
  40761=>"100011000",
  40762=>"101100100",
  40763=>"110101011",
  40764=>"111101101",
  40765=>"001000100",
  40766=>"110010101",
  40767=>"110001111",
  40768=>"110001011",
  40769=>"000111001",
  40770=>"011001011",
  40771=>"011011011",
  40772=>"111101111",
  40773=>"111001000",
  40774=>"111111001",
  40775=>"100100010",
  40776=>"110100100",
  40777=>"111110100",
  40778=>"010100001",
  40779=>"110110000",
  40780=>"011100111",
  40781=>"111100001",
  40782=>"100001101",
  40783=>"001010010",
  40784=>"100000100",
  40785=>"000011000",
  40786=>"110001011",
  40787=>"110001000",
  40788=>"110111110",
  40789=>"101101110",
  40790=>"011001100",
  40791=>"111101100",
  40792=>"010100000",
  40793=>"101011000",
  40794=>"111010101",
  40795=>"000100101",
  40796=>"010110011",
  40797=>"111011010",
  40798=>"110010101",
  40799=>"010001010",
  40800=>"011010010",
  40801=>"101011001",
  40802=>"110100101",
  40803=>"101111010",
  40804=>"011011011",
  40805=>"101001111",
  40806=>"011000100",
  40807=>"110110101",
  40808=>"001010010",
  40809=>"100101000",
  40810=>"101110100",
  40811=>"100110000",
  40812=>"001111101",
  40813=>"100101000",
  40814=>"001001011",
  40815=>"101111011",
  40816=>"001111011",
  40817=>"110100111",
  40818=>"010001101",
  40819=>"111011011",
  40820=>"000000110",
  40821=>"111101001",
  40822=>"001110000",
  40823=>"100110000",
  40824=>"011000101",
  40825=>"101111001",
  40826=>"101100111",
  40827=>"110111101",
  40828=>"111010001",
  40829=>"111110110",
  40830=>"100011101",
  40831=>"001001000",
  40832=>"101001001",
  40833=>"110100000",
  40834=>"111100000",
  40835=>"100010000",
  40836=>"111000001",
  40837=>"001000010",
  40838=>"101100001",
  40839=>"010010100",
  40840=>"011110111",
  40841=>"000110101",
  40842=>"010100001",
  40843=>"011110011",
  40844=>"111011111",
  40845=>"111001001",
  40846=>"111001111",
  40847=>"011100110",
  40848=>"110001111",
  40849=>"110010011",
  40850=>"101111010",
  40851=>"000111101",
  40852=>"010101110",
  40853=>"111000011",
  40854=>"001110111",
  40855=>"000011000",
  40856=>"011000000",
  40857=>"010000010",
  40858=>"001011000",
  40859=>"111010100",
  40860=>"100010101",
  40861=>"000101101",
  40862=>"001000100",
  40863=>"000101110",
  40864=>"100000101",
  40865=>"001001010",
  40866=>"110100101",
  40867=>"110110111",
  40868=>"010110011",
  40869=>"011001110",
  40870=>"011100111",
  40871=>"000111101",
  40872=>"000110010",
  40873=>"111111011",
  40874=>"011101000",
  40875=>"011100011",
  40876=>"000110101",
  40877=>"000000000",
  40878=>"101001001",
  40879=>"001110011",
  40880=>"000011100",
  40881=>"001101010",
  40882=>"110010001",
  40883=>"010000010",
  40884=>"010111011",
  40885=>"110101111",
  40886=>"100000110",
  40887=>"101000110",
  40888=>"010101100",
  40889=>"111101110",
  40890=>"101000110",
  40891=>"101100011",
  40892=>"101000100",
  40893=>"101010000",
  40894=>"111111001",
  40895=>"000110111",
  40896=>"110000000",
  40897=>"000110101",
  40898=>"100011010",
  40899=>"001000001",
  40900=>"110110000",
  40901=>"101011101",
  40902=>"110101110",
  40903=>"000110011",
  40904=>"100010100",
  40905=>"010001101",
  40906=>"110111010",
  40907=>"010000010",
  40908=>"100110100",
  40909=>"100110101",
  40910=>"011110110",
  40911=>"000000000",
  40912=>"010111010",
  40913=>"011101011",
  40914=>"110010011",
  40915=>"010101010",
  40916=>"000011011",
  40917=>"000010011",
  40918=>"100111011",
  40919=>"011110110",
  40920=>"111011001",
  40921=>"010101100",
  40922=>"111111011",
  40923=>"110101111",
  40924=>"011111000",
  40925=>"100011100",
  40926=>"110000110",
  40927=>"110100111",
  40928=>"000010000",
  40929=>"111110001",
  40930=>"110110000",
  40931=>"110111011",
  40932=>"111010110",
  40933=>"000110001",
  40934=>"010110000",
  40935=>"100011010",
  40936=>"100110010",
  40937=>"001011100",
  40938=>"110111110",
  40939=>"010111001",
  40940=>"101111110",
  40941=>"001000101",
  40942=>"011000000",
  40943=>"000111010",
  40944=>"100001110",
  40945=>"100110010",
  40946=>"101100011",
  40947=>"101000001",
  40948=>"000011000",
  40949=>"111000111",
  40950=>"010110110",
  40951=>"111011101",
  40952=>"110111111",
  40953=>"111011010",
  40954=>"110011010",
  40955=>"010110000",
  40956=>"101101101",
  40957=>"001000001",
  40958=>"110011111",
  40959=>"110110111",
  40960=>"001010001",
  40961=>"010000011",
  40962=>"011001101",
  40963=>"000111101",
  40964=>"101110110",
  40965=>"001010111",
  40966=>"000100000",
  40967=>"011111000",
  40968=>"100101100",
  40969=>"001010011",
  40970=>"011110000",
  40971=>"011100001",
  40972=>"111100101",
  40973=>"100010011",
  40974=>"100110000",
  40975=>"010110111",
  40976=>"101000110",
  40977=>"101100111",
  40978=>"000110101",
  40979=>"110111101",
  40980=>"000101100",
  40981=>"001100000",
  40982=>"001011110",
  40983=>"000101000",
  40984=>"000000010",
  40985=>"001110010",
  40986=>"101110011",
  40987=>"101011010",
  40988=>"111000001",
  40989=>"011001000",
  40990=>"001101100",
  40991=>"010000110",
  40992=>"110101000",
  40993=>"101010110",
  40994=>"111000100",
  40995=>"010110000",
  40996=>"101100010",
  40997=>"100101000",
  40998=>"100011100",
  40999=>"011101000",
  41000=>"101100110",
  41001=>"100101111",
  41002=>"110000100",
  41003=>"101000100",
  41004=>"001110100",
  41005=>"000011111",
  41006=>"111100000",
  41007=>"001101000",
  41008=>"001000000",
  41009=>"011101001",
  41010=>"000000011",
  41011=>"100011101",
  41012=>"000010001",
  41013=>"101001110",
  41014=>"010010010",
  41015=>"110010111",
  41016=>"011100000",
  41017=>"110010011",
  41018=>"000100101",
  41019=>"011111110",
  41020=>"100101101",
  41021=>"000011001",
  41022=>"101101000",
  41023=>"110100100",
  41024=>"110011110",
  41025=>"001000110",
  41026=>"110000001",
  41027=>"101111001",
  41028=>"101010000",
  41029=>"000011100",
  41030=>"111101101",
  41031=>"010000110",
  41032=>"101001010",
  41033=>"011100001",
  41034=>"010110011",
  41035=>"000101011",
  41036=>"101110001",
  41037=>"101000100",
  41038=>"000101110",
  41039=>"010010111",
  41040=>"000010101",
  41041=>"000001101",
  41042=>"011110111",
  41043=>"010010010",
  41044=>"111001111",
  41045=>"000001010",
  41046=>"110011011",
  41047=>"111101111",
  41048=>"000000010",
  41049=>"110001000",
  41050=>"010111010",
  41051=>"110001000",
  41052=>"000100001",
  41053=>"110011111",
  41054=>"110110010",
  41055=>"000011101",
  41056=>"001010000",
  41057=>"111111100",
  41058=>"010011100",
  41059=>"011100110",
  41060=>"110011000",
  41061=>"001100000",
  41062=>"100000011",
  41063=>"100101100",
  41064=>"011111001",
  41065=>"100000100",
  41066=>"110000101",
  41067=>"011101000",
  41068=>"110111011",
  41069=>"010000000",
  41070=>"101100111",
  41071=>"001001110",
  41072=>"110101011",
  41073=>"011111000",
  41074=>"100110100",
  41075=>"111111100",
  41076=>"000010011",
  41077=>"001010010",
  41078=>"100100101",
  41079=>"011000110",
  41080=>"111011001",
  41081=>"100110000",
  41082=>"001011111",
  41083=>"010000000",
  41084=>"000101111",
  41085=>"011010011",
  41086=>"011000111",
  41087=>"000000111",
  41088=>"010001011",
  41089=>"001101110",
  41090=>"101101110",
  41091=>"001001001",
  41092=>"001001111",
  41093=>"111010110",
  41094=>"101101111",
  41095=>"101110001",
  41096=>"010111011",
  41097=>"000100101",
  41098=>"000111101",
  41099=>"110011001",
  41100=>"000011010",
  41101=>"110000110",
  41102=>"010000011",
  41103=>"010100110",
  41104=>"110101001",
  41105=>"101111011",
  41106=>"000000101",
  41107=>"000111110",
  41108=>"101101111",
  41109=>"000011101",
  41110=>"001101111",
  41111=>"001001101",
  41112=>"111000110",
  41113=>"000100101",
  41114=>"110111001",
  41115=>"011011011",
  41116=>"110111011",
  41117=>"000001110",
  41118=>"101011111",
  41119=>"000011100",
  41120=>"001010000",
  41121=>"100011010",
  41122=>"110010111",
  41123=>"010101101",
  41124=>"100010000",
  41125=>"100110111",
  41126=>"000110001",
  41127=>"010100100",
  41128=>"010000100",
  41129=>"110010011",
  41130=>"100001010",
  41131=>"110100010",
  41132=>"011101011",
  41133=>"101111101",
  41134=>"101101011",
  41135=>"110000110",
  41136=>"100010100",
  41137=>"000010000",
  41138=>"111001111",
  41139=>"000001100",
  41140=>"001000011",
  41141=>"110100010",
  41142=>"110011000",
  41143=>"010001001",
  41144=>"010010000",
  41145=>"110000010",
  41146=>"010010110",
  41147=>"011010110",
  41148=>"100010101",
  41149=>"110110001",
  41150=>"000010011",
  41151=>"111110000",
  41152=>"010111111",
  41153=>"010100011",
  41154=>"001111101",
  41155=>"001001100",
  41156=>"111011001",
  41157=>"010111010",
  41158=>"000011000",
  41159=>"010000011",
  41160=>"010100111",
  41161=>"000101001",
  41162=>"101110001",
  41163=>"011111010",
  41164=>"110011110",
  41165=>"010000100",
  41166=>"111011101",
  41167=>"010100111",
  41168=>"000000010",
  41169=>"011111010",
  41170=>"011100000",
  41171=>"000010111",
  41172=>"100001110",
  41173=>"100100000",
  41174=>"111111100",
  41175=>"111110011",
  41176=>"110111100",
  41177=>"001100010",
  41178=>"100000011",
  41179=>"010110101",
  41180=>"100000110",
  41181=>"100111001",
  41182=>"001100100",
  41183=>"100110011",
  41184=>"111111100",
  41185=>"010011100",
  41186=>"000001100",
  41187=>"110011100",
  41188=>"111111010",
  41189=>"011011101",
  41190=>"011110111",
  41191=>"110000010",
  41192=>"100101010",
  41193=>"111110011",
  41194=>"101101101",
  41195=>"111000010",
  41196=>"000110000",
  41197=>"011000100",
  41198=>"000011111",
  41199=>"111110100",
  41200=>"010001100",
  41201=>"010101101",
  41202=>"011010001",
  41203=>"100100000",
  41204=>"100001001",
  41205=>"010101111",
  41206=>"110111101",
  41207=>"100001000",
  41208=>"000011010",
  41209=>"001111000",
  41210=>"100101000",
  41211=>"000000001",
  41212=>"001000001",
  41213=>"110110000",
  41214=>"110111011",
  41215=>"000011000",
  41216=>"000011010",
  41217=>"111000100",
  41218=>"000010110",
  41219=>"010010010",
  41220=>"001100101",
  41221=>"111011000",
  41222=>"110111111",
  41223=>"011010010",
  41224=>"000100000",
  41225=>"000101011",
  41226=>"011100110",
  41227=>"001010111",
  41228=>"111100101",
  41229=>"100100000",
  41230=>"001100011",
  41231=>"000000011",
  41232=>"111000101",
  41233=>"100011100",
  41234=>"111110100",
  41235=>"001101110",
  41236=>"000101010",
  41237=>"011011001",
  41238=>"001100110",
  41239=>"000011100",
  41240=>"111100100",
  41241=>"000110000",
  41242=>"010111100",
  41243=>"010000000",
  41244=>"010101001",
  41245=>"111001101",
  41246=>"111001011",
  41247=>"010011100",
  41248=>"100000100",
  41249=>"010100100",
  41250=>"000010001",
  41251=>"000011111",
  41252=>"111101001",
  41253=>"010101111",
  41254=>"001101010",
  41255=>"100110111",
  41256=>"010000010",
  41257=>"010110011",
  41258=>"111010011",
  41259=>"100100110",
  41260=>"100001011",
  41261=>"100010000",
  41262=>"000100000",
  41263=>"001010000",
  41264=>"010100110",
  41265=>"100000001",
  41266=>"110100010",
  41267=>"101000111",
  41268=>"110011010",
  41269=>"101011110",
  41270=>"000110011",
  41271=>"000000001",
  41272=>"001001001",
  41273=>"110110100",
  41274=>"101110101",
  41275=>"110000010",
  41276=>"000111101",
  41277=>"000101011",
  41278=>"111100111",
  41279=>"000101001",
  41280=>"101000100",
  41281=>"111000011",
  41282=>"010001111",
  41283=>"110110101",
  41284=>"111000111",
  41285=>"111100111",
  41286=>"100000101",
  41287=>"000000000",
  41288=>"101000001",
  41289=>"111011101",
  41290=>"000000100",
  41291=>"110000000",
  41292=>"000000010",
  41293=>"101111100",
  41294=>"110110001",
  41295=>"110111110",
  41296=>"001000001",
  41297=>"110111001",
  41298=>"101001010",
  41299=>"100010100",
  41300=>"011000011",
  41301=>"011110110",
  41302=>"110011000",
  41303=>"110111101",
  41304=>"000100101",
  41305=>"110110000",
  41306=>"000010000",
  41307=>"110110001",
  41308=>"100010111",
  41309=>"101100000",
  41310=>"011010000",
  41311=>"101111111",
  41312=>"100110110",
  41313=>"111010100",
  41314=>"111101101",
  41315=>"110011000",
  41316=>"000111010",
  41317=>"111010001",
  41318=>"001011000",
  41319=>"001110111",
  41320=>"100000101",
  41321=>"010100000",
  41322=>"011110100",
  41323=>"000101100",
  41324=>"100100000",
  41325=>"111001110",
  41326=>"100100111",
  41327=>"110110101",
  41328=>"010111111",
  41329=>"001001100",
  41330=>"011011000",
  41331=>"111100111",
  41332=>"100101010",
  41333=>"100110001",
  41334=>"001111111",
  41335=>"111010100",
  41336=>"111110100",
  41337=>"100110001",
  41338=>"001000010",
  41339=>"101000001",
  41340=>"000001100",
  41341=>"001010100",
  41342=>"000011101",
  41343=>"000011100",
  41344=>"010100001",
  41345=>"000100100",
  41346=>"001101010",
  41347=>"111110111",
  41348=>"011001001",
  41349=>"100011101",
  41350=>"111101001",
  41351=>"110100011",
  41352=>"111111000",
  41353=>"011000101",
  41354=>"110110001",
  41355=>"000000101",
  41356=>"101011010",
  41357=>"011111111",
  41358=>"011111110",
  41359=>"010110101",
  41360=>"101011010",
  41361=>"100001100",
  41362=>"111010010",
  41363=>"110011010",
  41364=>"110001011",
  41365=>"111011111",
  41366=>"011001110",
  41367=>"011101010",
  41368=>"110111010",
  41369=>"010010100",
  41370=>"001110011",
  41371=>"100001010",
  41372=>"011110111",
  41373=>"110100111",
  41374=>"010111010",
  41375=>"100001110",
  41376=>"000011111",
  41377=>"110110011",
  41378=>"011011111",
  41379=>"000000000",
  41380=>"001000110",
  41381=>"101001011",
  41382=>"101110010",
  41383=>"101011011",
  41384=>"001111100",
  41385=>"111010101",
  41386=>"101010010",
  41387=>"000011101",
  41388=>"100111110",
  41389=>"101000100",
  41390=>"101110010",
  41391=>"011101000",
  41392=>"010001110",
  41393=>"110111100",
  41394=>"011111010",
  41395=>"010110111",
  41396=>"010000101",
  41397=>"111100110",
  41398=>"010010101",
  41399=>"110000000",
  41400=>"111101001",
  41401=>"010100001",
  41402=>"000100010",
  41403=>"010100010",
  41404=>"101000100",
  41405=>"011111010",
  41406=>"000011001",
  41407=>"110011100",
  41408=>"010001001",
  41409=>"101011011",
  41410=>"000111111",
  41411=>"010010001",
  41412=>"000111110",
  41413=>"100000001",
  41414=>"111100100",
  41415=>"010110010",
  41416=>"111010010",
  41417=>"011010001",
  41418=>"011110111",
  41419=>"010010010",
  41420=>"001100110",
  41421=>"010101111",
  41422=>"111011000",
  41423=>"100110011",
  41424=>"111110001",
  41425=>"010100000",
  41426=>"011010101",
  41427=>"111110011",
  41428=>"110001101",
  41429=>"010111110",
  41430=>"101101001",
  41431=>"110111111",
  41432=>"111000001",
  41433=>"011111001",
  41434=>"011100001",
  41435=>"111001111",
  41436=>"011100011",
  41437=>"000101000",
  41438=>"110100111",
  41439=>"010110010",
  41440=>"011011010",
  41441=>"110110010",
  41442=>"000100110",
  41443=>"111011100",
  41444=>"110110001",
  41445=>"111111010",
  41446=>"000100100",
  41447=>"001011000",
  41448=>"011010101",
  41449=>"010001010",
  41450=>"111001100",
  41451=>"100101001",
  41452=>"010001010",
  41453=>"000101001",
  41454=>"100100100",
  41455=>"100110110",
  41456=>"100100110",
  41457=>"111111101",
  41458=>"101011000",
  41459=>"011101100",
  41460=>"001110100",
  41461=>"100001110",
  41462=>"011000001",
  41463=>"101101000",
  41464=>"111110010",
  41465=>"101101100",
  41466=>"000000010",
  41467=>"011101000",
  41468=>"001101000",
  41469=>"010001000",
  41470=>"110011001",
  41471=>"100110111",
  41472=>"011010101",
  41473=>"000101100",
  41474=>"001000011",
  41475=>"101000100",
  41476=>"010101001",
  41477=>"010100001",
  41478=>"011001001",
  41479=>"010100010",
  41480=>"101111011",
  41481=>"100011101",
  41482=>"100010010",
  41483=>"000100010",
  41484=>"001111101",
  41485=>"101010010",
  41486=>"001111110",
  41487=>"100000000",
  41488=>"011111110",
  41489=>"100100100",
  41490=>"110111100",
  41491=>"010100000",
  41492=>"100010011",
  41493=>"111011111",
  41494=>"000011100",
  41495=>"011111010",
  41496=>"101010000",
  41497=>"011100110",
  41498=>"011001111",
  41499=>"001001110",
  41500=>"110110101",
  41501=>"101011011",
  41502=>"111101010",
  41503=>"101000100",
  41504=>"011010111",
  41505=>"000111110",
  41506=>"011010111",
  41507=>"000111111",
  41508=>"111011011",
  41509=>"000011011",
  41510=>"010001000",
  41511=>"010111111",
  41512=>"000001010",
  41513=>"010101110",
  41514=>"010110100",
  41515=>"100010101",
  41516=>"001110101",
  41517=>"000101000",
  41518=>"010101010",
  41519=>"100001001",
  41520=>"110001100",
  41521=>"101010010",
  41522=>"001110001",
  41523=>"010101000",
  41524=>"011000001",
  41525=>"101001011",
  41526=>"011010011",
  41527=>"001001110",
  41528=>"001011110",
  41529=>"101101111",
  41530=>"110010000",
  41531=>"010000000",
  41532=>"101100110",
  41533=>"001011000",
  41534=>"110000000",
  41535=>"111111111",
  41536=>"000010111",
  41537=>"101110011",
  41538=>"000111001",
  41539=>"101100101",
  41540=>"001011101",
  41541=>"010110111",
  41542=>"111010111",
  41543=>"001111000",
  41544=>"000101001",
  41545=>"101111111",
  41546=>"010110111",
  41547=>"000110111",
  41548=>"010000000",
  41549=>"110010011",
  41550=>"101110110",
  41551=>"001001000",
  41552=>"000010100",
  41553=>"011001110",
  41554=>"001010110",
  41555=>"010111000",
  41556=>"001000001",
  41557=>"100001000",
  41558=>"000100000",
  41559=>"101011110",
  41560=>"010010111",
  41561=>"101110001",
  41562=>"001110011",
  41563=>"011000110",
  41564=>"000010111",
  41565=>"000011011",
  41566=>"111101000",
  41567=>"101001010",
  41568=>"111011000",
  41569=>"000111101",
  41570=>"010001110",
  41571=>"001110100",
  41572=>"000100100",
  41573=>"111110101",
  41574=>"100110100",
  41575=>"001001101",
  41576=>"011100100",
  41577=>"001111100",
  41578=>"010110001",
  41579=>"100110101",
  41580=>"010100111",
  41581=>"111010010",
  41582=>"010111000",
  41583=>"101011111",
  41584=>"101110000",
  41585=>"001000100",
  41586=>"001100110",
  41587=>"001010101",
  41588=>"101110101",
  41589=>"011010000",
  41590=>"011111111",
  41591=>"001000011",
  41592=>"001011000",
  41593=>"001110001",
  41594=>"000011111",
  41595=>"011000101",
  41596=>"101010111",
  41597=>"010100000",
  41598=>"100100010",
  41599=>"011000001",
  41600=>"000000001",
  41601=>"100001011",
  41602=>"010101000",
  41603=>"011001011",
  41604=>"101010110",
  41605=>"100101010",
  41606=>"001100010",
  41607=>"111111111",
  41608=>"010000001",
  41609=>"011101111",
  41610=>"110010010",
  41611=>"110011100",
  41612=>"011101111",
  41613=>"010010010",
  41614=>"100101001",
  41615=>"101001101",
  41616=>"110010111",
  41617=>"001010110",
  41618=>"111001011",
  41619=>"111001110",
  41620=>"101100011",
  41621=>"011100011",
  41622=>"111100111",
  41623=>"000011010",
  41624=>"001110001",
  41625=>"001000001",
  41626=>"011101011",
  41627=>"111101110",
  41628=>"010111110",
  41629=>"111101001",
  41630=>"101000011",
  41631=>"000100000",
  41632=>"010000000",
  41633=>"111111110",
  41634=>"111000000",
  41635=>"001100011",
  41636=>"111100111",
  41637=>"111101101",
  41638=>"000011101",
  41639=>"100000001",
  41640=>"110101010",
  41641=>"000000111",
  41642=>"010101010",
  41643=>"111000110",
  41644=>"001010100",
  41645=>"110100111",
  41646=>"100100000",
  41647=>"010000001",
  41648=>"100001011",
  41649=>"011000000",
  41650=>"100010001",
  41651=>"010000001",
  41652=>"000010000",
  41653=>"111100101",
  41654=>"011100101",
  41655=>"111101001",
  41656=>"011101001",
  41657=>"110010010",
  41658=>"111010010",
  41659=>"011110000",
  41660=>"011100010",
  41661=>"011000010",
  41662=>"001001001",
  41663=>"101000100",
  41664=>"001111001",
  41665=>"101010000",
  41666=>"100000000",
  41667=>"000110101",
  41668=>"010110010",
  41669=>"100001110",
  41670=>"001110011",
  41671=>"001111100",
  41672=>"000010101",
  41673=>"111000110",
  41674=>"101011001",
  41675=>"001000111",
  41676=>"101001001",
  41677=>"011110110",
  41678=>"000100001",
  41679=>"100111110",
  41680=>"100010001",
  41681=>"001100001",
  41682=>"011001100",
  41683=>"010010011",
  41684=>"000000011",
  41685=>"011011111",
  41686=>"101001010",
  41687=>"110100001",
  41688=>"101011010",
  41689=>"111000010",
  41690=>"010011101",
  41691=>"000011000",
  41692=>"101110111",
  41693=>"010100111",
  41694=>"100111011",
  41695=>"010011011",
  41696=>"000010011",
  41697=>"010001000",
  41698=>"000110111",
  41699=>"000101001",
  41700=>"100011010",
  41701=>"100100001",
  41702=>"000001101",
  41703=>"111100110",
  41704=>"010000101",
  41705=>"010111101",
  41706=>"110000010",
  41707=>"001001000",
  41708=>"110100111",
  41709=>"000001100",
  41710=>"110111110",
  41711=>"010110010",
  41712=>"001010011",
  41713=>"001101111",
  41714=>"011101111",
  41715=>"000011010",
  41716=>"100011001",
  41717=>"110000000",
  41718=>"000100001",
  41719=>"110100010",
  41720=>"100010001",
  41721=>"101011011",
  41722=>"110000101",
  41723=>"011001000",
  41724=>"111000101",
  41725=>"000000001",
  41726=>"000001011",
  41727=>"001101001",
  41728=>"001110000",
  41729=>"110111111",
  41730=>"101110110",
  41731=>"010010010",
  41732=>"101011000",
  41733=>"010100000",
  41734=>"100001100",
  41735=>"010101011",
  41736=>"011111111",
  41737=>"100010000",
  41738=>"110001111",
  41739=>"100100110",
  41740=>"100101000",
  41741=>"110010000",
  41742=>"101101000",
  41743=>"001010001",
  41744=>"100010111",
  41745=>"100010100",
  41746=>"111001011",
  41747=>"100010100",
  41748=>"110110110",
  41749=>"100001010",
  41750=>"010100010",
  41751=>"000100111",
  41752=>"000101010",
  41753=>"001100100",
  41754=>"100011011",
  41755=>"011100111",
  41756=>"101111001",
  41757=>"110010010",
  41758=>"100111011",
  41759=>"000010110",
  41760=>"111001010",
  41761=>"100000010",
  41762=>"110101011",
  41763=>"100010101",
  41764=>"111011111",
  41765=>"100100010",
  41766=>"100000011",
  41767=>"110001100",
  41768=>"010010100",
  41769=>"010110100",
  41770=>"110100010",
  41771=>"011110001",
  41772=>"011110010",
  41773=>"000100011",
  41774=>"110111111",
  41775=>"101111010",
  41776=>"110110001",
  41777=>"010000110",
  41778=>"000001011",
  41779=>"100111011",
  41780=>"010011001",
  41781=>"111110000",
  41782=>"000100100",
  41783=>"101101011",
  41784=>"101110110",
  41785=>"100101100",
  41786=>"010000011",
  41787=>"111011110",
  41788=>"011001100",
  41789=>"101101100",
  41790=>"100000000",
  41791=>"111010100",
  41792=>"110000001",
  41793=>"010011011",
  41794=>"011001010",
  41795=>"111110001",
  41796=>"101001111",
  41797=>"111100011",
  41798=>"011111010",
  41799=>"100011001",
  41800=>"111011001",
  41801=>"100110001",
  41802=>"111001011",
  41803=>"111100011",
  41804=>"100011010",
  41805=>"101011010",
  41806=>"101100001",
  41807=>"101100111",
  41808=>"100011000",
  41809=>"101101110",
  41810=>"100101100",
  41811=>"011110010",
  41812=>"100010111",
  41813=>"111101101",
  41814=>"001111111",
  41815=>"100110000",
  41816=>"100011110",
  41817=>"111011011",
  41818=>"100011111",
  41819=>"111101010",
  41820=>"010011101",
  41821=>"100001100",
  41822=>"000010011",
  41823=>"100001100",
  41824=>"111001111",
  41825=>"010001101",
  41826=>"101000001",
  41827=>"000101010",
  41828=>"011001101",
  41829=>"011000110",
  41830=>"101100001",
  41831=>"101010011",
  41832=>"101010111",
  41833=>"000100110",
  41834=>"111010011",
  41835=>"101100110",
  41836=>"101010001",
  41837=>"101001101",
  41838=>"101110010",
  41839=>"110110101",
  41840=>"010100010",
  41841=>"000100101",
  41842=>"111000001",
  41843=>"110001111",
  41844=>"001110101",
  41845=>"111000100",
  41846=>"101111111",
  41847=>"111011000",
  41848=>"001010111",
  41849=>"110011110",
  41850=>"100001100",
  41851=>"101011001",
  41852=>"000010011",
  41853=>"110101001",
  41854=>"100101110",
  41855=>"111011100",
  41856=>"001110010",
  41857=>"111101100",
  41858=>"111100111",
  41859=>"000010100",
  41860=>"011000101",
  41861=>"100101000",
  41862=>"101100011",
  41863=>"010111110",
  41864=>"001001110",
  41865=>"001011011",
  41866=>"111011101",
  41867=>"000111010",
  41868=>"110100010",
  41869=>"000010001",
  41870=>"000100010",
  41871=>"000010010",
  41872=>"100110001",
  41873=>"011100000",
  41874=>"000111000",
  41875=>"010101100",
  41876=>"001110111",
  41877=>"010010101",
  41878=>"000110010",
  41879=>"011110011",
  41880=>"111100100",
  41881=>"011101101",
  41882=>"001011100",
  41883=>"100110000",
  41884=>"111101011",
  41885=>"001011110",
  41886=>"110000000",
  41887=>"110000101",
  41888=>"010101110",
  41889=>"110101000",
  41890=>"011110111",
  41891=>"111000011",
  41892=>"001110010",
  41893=>"011110111",
  41894=>"010100000",
  41895=>"111111011",
  41896=>"010110101",
  41897=>"101100010",
  41898=>"001110110",
  41899=>"001011111",
  41900=>"010110000",
  41901=>"010111010",
  41902=>"011000000",
  41903=>"100001011",
  41904=>"001111000",
  41905=>"101011000",
  41906=>"111101101",
  41907=>"100011010",
  41908=>"100001111",
  41909=>"110101001",
  41910=>"000101101",
  41911=>"001001100",
  41912=>"001010011",
  41913=>"000001001",
  41914=>"010100010",
  41915=>"011011110",
  41916=>"000101000",
  41917=>"010010000",
  41918=>"110010110",
  41919=>"010110101",
  41920=>"110110000",
  41921=>"011110110",
  41922=>"110100011",
  41923=>"011001000",
  41924=>"000011011",
  41925=>"100010110",
  41926=>"110000011",
  41927=>"111101011",
  41928=>"000101011",
  41929=>"000110000",
  41930=>"010101010",
  41931=>"010011011",
  41932=>"111101111",
  41933=>"101000000",
  41934=>"000010010",
  41935=>"101110000",
  41936=>"000111110",
  41937=>"110111101",
  41938=>"111101101",
  41939=>"110110000",
  41940=>"111111111",
  41941=>"111000011",
  41942=>"101100110",
  41943=>"111010101",
  41944=>"101000000",
  41945=>"001000110",
  41946=>"010001111",
  41947=>"011000111",
  41948=>"101110101",
  41949=>"100010010",
  41950=>"010100100",
  41951=>"000101100",
  41952=>"111111101",
  41953=>"111100110",
  41954=>"011100000",
  41955=>"110110000",
  41956=>"010111100",
  41957=>"001011100",
  41958=>"100001010",
  41959=>"100100000",
  41960=>"011010011",
  41961=>"111010010",
  41962=>"100000111",
  41963=>"001101001",
  41964=>"001000110",
  41965=>"011010000",
  41966=>"010000010",
  41967=>"001110010",
  41968=>"111111100",
  41969=>"000100100",
  41970=>"000100101",
  41971=>"001000001",
  41972=>"101100010",
  41973=>"111100000",
  41974=>"011000100",
  41975=>"101111111",
  41976=>"001111010",
  41977=>"000111011",
  41978=>"110001101",
  41979=>"100000011",
  41980=>"000011001",
  41981=>"010100011",
  41982=>"100010001",
  41983=>"100000111",
  41984=>"100001000",
  41985=>"101000101",
  41986=>"110000011",
  41987=>"011001001",
  41988=>"001010000",
  41989=>"000011011",
  41990=>"101110010",
  41991=>"110010000",
  41992=>"011011101",
  41993=>"000001110",
  41994=>"001100110",
  41995=>"010001111",
  41996=>"010101101",
  41997=>"000110100",
  41998=>"110001010",
  41999=>"000110010",
  42000=>"101111100",
  42001=>"101010000",
  42002=>"000011101",
  42003=>"101011100",
  42004=>"000101111",
  42005=>"111000101",
  42006=>"101011101",
  42007=>"110010101",
  42008=>"000011101",
  42009=>"010100010",
  42010=>"001011000",
  42011=>"111001011",
  42012=>"101101000",
  42013=>"111001101",
  42014=>"001011001",
  42015=>"000101000",
  42016=>"000001000",
  42017=>"010100100",
  42018=>"111001100",
  42019=>"010101111",
  42020=>"111111111",
  42021=>"110000101",
  42022=>"100110000",
  42023=>"010011001",
  42024=>"101110001",
  42025=>"011111011",
  42026=>"111001000",
  42027=>"000110110",
  42028=>"110110011",
  42029=>"000010110",
  42030=>"010100000",
  42031=>"110101111",
  42032=>"100110111",
  42033=>"011101101",
  42034=>"011100101",
  42035=>"101010001",
  42036=>"001011101",
  42037=>"000011110",
  42038=>"111001001",
  42039=>"010001011",
  42040=>"101111110",
  42041=>"111000100",
  42042=>"111010100",
  42043=>"101000111",
  42044=>"001000001",
  42045=>"000111001",
  42046=>"101110111",
  42047=>"100111100",
  42048=>"000101111",
  42049=>"000010110",
  42050=>"010011100",
  42051=>"101100111",
  42052=>"111001001",
  42053=>"010101110",
  42054=>"101011000",
  42055=>"100101001",
  42056=>"011101001",
  42057=>"010111010",
  42058=>"001100110",
  42059=>"011100110",
  42060=>"100000111",
  42061=>"000111101",
  42062=>"111110011",
  42063=>"110111011",
  42064=>"001000111",
  42065=>"111101111",
  42066=>"000111101",
  42067=>"001011110",
  42068=>"111100000",
  42069=>"010000011",
  42070=>"110001100",
  42071=>"101101001",
  42072=>"110010001",
  42073=>"101101111",
  42074=>"100111110",
  42075=>"000001000",
  42076=>"010110110",
  42077=>"011110010",
  42078=>"101111001",
  42079=>"110010010",
  42080=>"001101000",
  42081=>"101100110",
  42082=>"000011010",
  42083=>"000000001",
  42084=>"001000010",
  42085=>"010000000",
  42086=>"011100000",
  42087=>"000010010",
  42088=>"010000000",
  42089=>"110100101",
  42090=>"100101010",
  42091=>"100000011",
  42092=>"011101101",
  42093=>"111010111",
  42094=>"010100001",
  42095=>"000010000",
  42096=>"100100000",
  42097=>"110000111",
  42098=>"111111001",
  42099=>"000010110",
  42100=>"000110011",
  42101=>"000111101",
  42102=>"111101101",
  42103=>"000101000",
  42104=>"101000100",
  42105=>"000110110",
  42106=>"001001010",
  42107=>"100010000",
  42108=>"010000110",
  42109=>"110011011",
  42110=>"000001000",
  42111=>"001110100",
  42112=>"010001101",
  42113=>"001001111",
  42114=>"110001111",
  42115=>"111001010",
  42116=>"000111000",
  42117=>"101011111",
  42118=>"000000011",
  42119=>"100011011",
  42120=>"001010101",
  42121=>"000000110",
  42122=>"001010000",
  42123=>"111110111",
  42124=>"101111110",
  42125=>"010010000",
  42126=>"110111111",
  42127=>"110101010",
  42128=>"111110011",
  42129=>"010111001",
  42130=>"010101101",
  42131=>"111000111",
  42132=>"000000000",
  42133=>"001100001",
  42134=>"011011111",
  42135=>"010000000",
  42136=>"000011110",
  42137=>"000110111",
  42138=>"000110010",
  42139=>"000110000",
  42140=>"110010111",
  42141=>"000011000",
  42142=>"000110000",
  42143=>"110110111",
  42144=>"001010000",
  42145=>"111010110",
  42146=>"001000101",
  42147=>"001000000",
  42148=>"010111111",
  42149=>"011010100",
  42150=>"010011101",
  42151=>"010001110",
  42152=>"010110000",
  42153=>"010100000",
  42154=>"101100101",
  42155=>"010110010",
  42156=>"000000110",
  42157=>"001011101",
  42158=>"011000110",
  42159=>"101000010",
  42160=>"110110011",
  42161=>"100001011",
  42162=>"111111111",
  42163=>"001110001",
  42164=>"110111100",
  42165=>"110111111",
  42166=>"000100010",
  42167=>"001001100",
  42168=>"111011010",
  42169=>"011101011",
  42170=>"100100011",
  42171=>"011101100",
  42172=>"000010010",
  42173=>"100010111",
  42174=>"000101110",
  42175=>"000100000",
  42176=>"010010001",
  42177=>"111011111",
  42178=>"000011010",
  42179=>"010010011",
  42180=>"111111000",
  42181=>"110000111",
  42182=>"110101010",
  42183=>"000011111",
  42184=>"101110101",
  42185=>"000010111",
  42186=>"011111110",
  42187=>"010101000",
  42188=>"111001000",
  42189=>"111010101",
  42190=>"110000000",
  42191=>"010000110",
  42192=>"100000001",
  42193=>"000000110",
  42194=>"000111011",
  42195=>"010111011",
  42196=>"010000011",
  42197=>"010111110",
  42198=>"111010110",
  42199=>"111111100",
  42200=>"101111011",
  42201=>"110111001",
  42202=>"100110100",
  42203=>"100011011",
  42204=>"100110111",
  42205=>"111011111",
  42206=>"100000001",
  42207=>"100001110",
  42208=>"101110010",
  42209=>"110101010",
  42210=>"011000100",
  42211=>"111110111",
  42212=>"111000000",
  42213=>"101001110",
  42214=>"110000000",
  42215=>"111010011",
  42216=>"111111100",
  42217=>"010111000",
  42218=>"000110101",
  42219=>"100110000",
  42220=>"000001101",
  42221=>"101010011",
  42222=>"100001010",
  42223=>"100111100",
  42224=>"111111010",
  42225=>"000111101",
  42226=>"101000110",
  42227=>"001000111",
  42228=>"000001111",
  42229=>"011001111",
  42230=>"001110010",
  42231=>"001001110",
  42232=>"000111000",
  42233=>"000100011",
  42234=>"111100111",
  42235=>"110100101",
  42236=>"001001000",
  42237=>"011101010",
  42238=>"111001101",
  42239=>"101100111",
  42240=>"111110001",
  42241=>"110101101",
  42242=>"001000001",
  42243=>"011111010",
  42244=>"000110110",
  42245=>"101101100",
  42246=>"001110111",
  42247=>"101101011",
  42248=>"011111000",
  42249=>"001100100",
  42250=>"011011000",
  42251=>"010111000",
  42252=>"010001011",
  42253=>"000010001",
  42254=>"000001001",
  42255=>"010110100",
  42256=>"010111100",
  42257=>"100010010",
  42258=>"001111111",
  42259=>"101010000",
  42260=>"111010111",
  42261=>"001101101",
  42262=>"000111001",
  42263=>"101101010",
  42264=>"000000101",
  42265=>"111011001",
  42266=>"001110110",
  42267=>"100111011",
  42268=>"111111011",
  42269=>"100111100",
  42270=>"000110010",
  42271=>"000000011",
  42272=>"111111111",
  42273=>"011111111",
  42274=>"011001010",
  42275=>"110110000",
  42276=>"101011100",
  42277=>"100101000",
  42278=>"001000111",
  42279=>"101110111",
  42280=>"010110000",
  42281=>"011010101",
  42282=>"010011010",
  42283=>"000101010",
  42284=>"011100000",
  42285=>"000110010",
  42286=>"100010110",
  42287=>"110001111",
  42288=>"101010001",
  42289=>"100000000",
  42290=>"110010110",
  42291=>"000101101",
  42292=>"010011010",
  42293=>"010000101",
  42294=>"100001011",
  42295=>"000111000",
  42296=>"100011110",
  42297=>"111011010",
  42298=>"111101101",
  42299=>"100001011",
  42300=>"001101111",
  42301=>"010010001",
  42302=>"011001001",
  42303=>"111111101",
  42304=>"110000101",
  42305=>"011111010",
  42306=>"101100101",
  42307=>"000111000",
  42308=>"011100111",
  42309=>"011011100",
  42310=>"100111100",
  42311=>"101111011",
  42312=>"001010111",
  42313=>"111010111",
  42314=>"010101100",
  42315=>"110111111",
  42316=>"111001000",
  42317=>"111101100",
  42318=>"110001000",
  42319=>"110101100",
  42320=>"000000010",
  42321=>"011010100",
  42322=>"010010100",
  42323=>"100111100",
  42324=>"001111010",
  42325=>"011010110",
  42326=>"011000111",
  42327=>"111010001",
  42328=>"001110001",
  42329=>"100101111",
  42330=>"110011001",
  42331=>"000011001",
  42332=>"111010011",
  42333=>"101100101",
  42334=>"110000011",
  42335=>"101110100",
  42336=>"111010100",
  42337=>"111101011",
  42338=>"010011001",
  42339=>"000000001",
  42340=>"000000101",
  42341=>"110010101",
  42342=>"010111011",
  42343=>"000110010",
  42344=>"111111010",
  42345=>"001010001",
  42346=>"011000101",
  42347=>"001001110",
  42348=>"111110000",
  42349=>"001000000",
  42350=>"110001010",
  42351=>"001000010",
  42352=>"000111011",
  42353=>"011111101",
  42354=>"111011110",
  42355=>"111100010",
  42356=>"111101110",
  42357=>"000011110",
  42358=>"011000010",
  42359=>"110110100",
  42360=>"001001011",
  42361=>"110100110",
  42362=>"010111010",
  42363=>"101101000",
  42364=>"111011111",
  42365=>"111011001",
  42366=>"010100000",
  42367=>"111011110",
  42368=>"111001001",
  42369=>"100111101",
  42370=>"100100101",
  42371=>"010011011",
  42372=>"010011001",
  42373=>"110111011",
  42374=>"001101010",
  42375=>"111101111",
  42376=>"010011011",
  42377=>"110111010",
  42378=>"111111100",
  42379=>"111001000",
  42380=>"001101001",
  42381=>"100110111",
  42382=>"100111000",
  42383=>"010011011",
  42384=>"011110011",
  42385=>"000000011",
  42386=>"111001110",
  42387=>"000001111",
  42388=>"100010000",
  42389=>"111000011",
  42390=>"111011000",
  42391=>"010110010",
  42392=>"110000011",
  42393=>"010100100",
  42394=>"110100110",
  42395=>"111011111",
  42396=>"010000000",
  42397=>"110101011",
  42398=>"111111111",
  42399=>"010100000",
  42400=>"110101000",
  42401=>"110101000",
  42402=>"001101111",
  42403=>"000101100",
  42404=>"111011001",
  42405=>"010000100",
  42406=>"000011010",
  42407=>"011100110",
  42408=>"010010000",
  42409=>"100100010",
  42410=>"101000000",
  42411=>"100110010",
  42412=>"000110111",
  42413=>"001001000",
  42414=>"000101010",
  42415=>"010110111",
  42416=>"001111111",
  42417=>"111110110",
  42418=>"000110101",
  42419=>"111010101",
  42420=>"000001001",
  42421=>"111110011",
  42422=>"000000001",
  42423=>"011100011",
  42424=>"111101101",
  42425=>"100110111",
  42426=>"011101110",
  42427=>"111110011",
  42428=>"011101111",
  42429=>"111111011",
  42430=>"100000111",
  42431=>"101111010",
  42432=>"010101011",
  42433=>"100001101",
  42434=>"010011101",
  42435=>"101000001",
  42436=>"000100000",
  42437=>"101111000",
  42438=>"110011000",
  42439=>"000000100",
  42440=>"011101100",
  42441=>"001011100",
  42442=>"000000000",
  42443=>"001110011",
  42444=>"000001101",
  42445=>"001010111",
  42446=>"011100011",
  42447=>"100010001",
  42448=>"011110101",
  42449=>"110000011",
  42450=>"000010000",
  42451=>"110011111",
  42452=>"000010000",
  42453=>"011011101",
  42454=>"011001010",
  42455=>"001011001",
  42456=>"000111111",
  42457=>"011110011",
  42458=>"001101110",
  42459=>"111101000",
  42460=>"111110100",
  42461=>"010100011",
  42462=>"001111000",
  42463=>"110100011",
  42464=>"110110110",
  42465=>"001100001",
  42466=>"110011011",
  42467=>"001011010",
  42468=>"100110101",
  42469=>"111011011",
  42470=>"110101100",
  42471=>"010101110",
  42472=>"000101110",
  42473=>"011011110",
  42474=>"000110001",
  42475=>"101111100",
  42476=>"110110111",
  42477=>"101110011",
  42478=>"010110001",
  42479=>"001111011",
  42480=>"110101001",
  42481=>"111011110",
  42482=>"000001110",
  42483=>"111100111",
  42484=>"100001111",
  42485=>"001011110",
  42486=>"010001011",
  42487=>"111001010",
  42488=>"110101010",
  42489=>"110001010",
  42490=>"100111000",
  42491=>"100111000",
  42492=>"101100001",
  42493=>"000000100",
  42494=>"001100001",
  42495=>"001111111",
  42496=>"100001001",
  42497=>"110000001",
  42498=>"010010111",
  42499=>"100100100",
  42500=>"111011110",
  42501=>"110101100",
  42502=>"000011110",
  42503=>"100011000",
  42504=>"001001111",
  42505=>"100010111",
  42506=>"111010111",
  42507=>"110101111",
  42508=>"111110111",
  42509=>"101110000",
  42510=>"010000100",
  42511=>"000010100",
  42512=>"011000111",
  42513=>"101001110",
  42514=>"000111011",
  42515=>"100111111",
  42516=>"111101110",
  42517=>"000110001",
  42518=>"000100010",
  42519=>"010111100",
  42520=>"110101111",
  42521=>"101100001",
  42522=>"111110010",
  42523=>"111010000",
  42524=>"110000001",
  42525=>"110001001",
  42526=>"001100011",
  42527=>"010110001",
  42528=>"110110101",
  42529=>"101000001",
  42530=>"000000101",
  42531=>"000011110",
  42532=>"110110100",
  42533=>"000010110",
  42534=>"100101110",
  42535=>"000010100",
  42536=>"001010001",
  42537=>"010100001",
  42538=>"011101111",
  42539=>"110101010",
  42540=>"000111010",
  42541=>"000010111",
  42542=>"100000010",
  42543=>"000111010",
  42544=>"011111111",
  42545=>"010011111",
  42546=>"111110010",
  42547=>"101001100",
  42548=>"000001000",
  42549=>"101001010",
  42550=>"111110100",
  42551=>"110100001",
  42552=>"100000010",
  42553=>"000010011",
  42554=>"011001101",
  42555=>"000101001",
  42556=>"110001111",
  42557=>"011001111",
  42558=>"100010100",
  42559=>"010010101",
  42560=>"111011111",
  42561=>"011001010",
  42562=>"110110101",
  42563=>"110001101",
  42564=>"010101000",
  42565=>"011100100",
  42566=>"010000000",
  42567=>"010110110",
  42568=>"001000000",
  42569=>"101000100",
  42570=>"010010110",
  42571=>"011110010",
  42572=>"010111001",
  42573=>"101100011",
  42574=>"110111101",
  42575=>"001111101",
  42576=>"000100010",
  42577=>"011100111",
  42578=>"000110111",
  42579=>"100100100",
  42580=>"010011011",
  42581=>"101011001",
  42582=>"101101110",
  42583=>"110011011",
  42584=>"100101111",
  42585=>"111000011",
  42586=>"100001001",
  42587=>"000000111",
  42588=>"000110101",
  42589=>"000101100",
  42590=>"100000101",
  42591=>"000000000",
  42592=>"000000010",
  42593=>"011111001",
  42594=>"001001010",
  42595=>"100101011",
  42596=>"101000110",
  42597=>"100100111",
  42598=>"000010010",
  42599=>"111111011",
  42600=>"101110111",
  42601=>"000110000",
  42602=>"111111010",
  42603=>"111110100",
  42604=>"111111111",
  42605=>"010001001",
  42606=>"100100000",
  42607=>"011010110",
  42608=>"100010110",
  42609=>"110111101",
  42610=>"000011111",
  42611=>"000000111",
  42612=>"111000011",
  42613=>"011001000",
  42614=>"001100111",
  42615=>"110000000",
  42616=>"101001111",
  42617=>"111111110",
  42618=>"110111000",
  42619=>"001101011",
  42620=>"000000000",
  42621=>"010010100",
  42622=>"110110101",
  42623=>"011010011",
  42624=>"000000110",
  42625=>"011000011",
  42626=>"000001001",
  42627=>"011001000",
  42628=>"010011011",
  42629=>"010001100",
  42630=>"000000100",
  42631=>"001001101",
  42632=>"001110011",
  42633=>"000000011",
  42634=>"101010011",
  42635=>"100110111",
  42636=>"010110000",
  42637=>"110111111",
  42638=>"000000011",
  42639=>"100010011",
  42640=>"010011000",
  42641=>"111100110",
  42642=>"101110101",
  42643=>"111100100",
  42644=>"101111101",
  42645=>"110010100",
  42646=>"000100100",
  42647=>"100010101",
  42648=>"111011110",
  42649=>"001110110",
  42650=>"101101000",
  42651=>"101011010",
  42652=>"100011010",
  42653=>"011000110",
  42654=>"000100011",
  42655=>"011000011",
  42656=>"101010100",
  42657=>"100010001",
  42658=>"111111101",
  42659=>"000101011",
  42660=>"101101000",
  42661=>"011011011",
  42662=>"000111100",
  42663=>"000011110",
  42664=>"111111110",
  42665=>"101111101",
  42666=>"000010100",
  42667=>"111111011",
  42668=>"100111111",
  42669=>"011000101",
  42670=>"111100010",
  42671=>"101011101",
  42672=>"010111000",
  42673=>"000011000",
  42674=>"100010101",
  42675=>"001100100",
  42676=>"111100111",
  42677=>"110011110",
  42678=>"001001010",
  42679=>"110001101",
  42680=>"000111000",
  42681=>"000110010",
  42682=>"110100010",
  42683=>"000101011",
  42684=>"111000011",
  42685=>"100101000",
  42686=>"001100101",
  42687=>"000101110",
  42688=>"101110110",
  42689=>"110100111",
  42690=>"101110101",
  42691=>"100100111",
  42692=>"101010011",
  42693=>"111001000",
  42694=>"110001111",
  42695=>"100111101",
  42696=>"101000111",
  42697=>"001011000",
  42698=>"111101101",
  42699=>"000001111",
  42700=>"100000010",
  42701=>"110110000",
  42702=>"100011100",
  42703=>"011000100",
  42704=>"000101001",
  42705=>"011100100",
  42706=>"110001110",
  42707=>"000111001",
  42708=>"000001011",
  42709=>"010010010",
  42710=>"011110111",
  42711=>"010000111",
  42712=>"011101000",
  42713=>"011110100",
  42714=>"100100000",
  42715=>"000100000",
  42716=>"001010000",
  42717=>"000010010",
  42718=>"110110010",
  42719=>"101100111",
  42720=>"010110111",
  42721=>"011000000",
  42722=>"110000111",
  42723=>"111111100",
  42724=>"111111100",
  42725=>"010000000",
  42726=>"000101110",
  42727=>"000100111",
  42728=>"010111000",
  42729=>"011110110",
  42730=>"011100110",
  42731=>"101101110",
  42732=>"111001011",
  42733=>"010011000",
  42734=>"111111011",
  42735=>"100010011",
  42736=>"110001111",
  42737=>"001001011",
  42738=>"100000111",
  42739=>"110000111",
  42740=>"100011101",
  42741=>"111000111",
  42742=>"100010111",
  42743=>"110101100",
  42744=>"000110101",
  42745=>"110101110",
  42746=>"100011001",
  42747=>"000101100",
  42748=>"011010100",
  42749=>"011011001",
  42750=>"010001010",
  42751=>"110000101",
  42752=>"001101111",
  42753=>"110000001",
  42754=>"111110010",
  42755=>"011001011",
  42756=>"100000010",
  42757=>"001110011",
  42758=>"010000000",
  42759=>"100111100",
  42760=>"011010001",
  42761=>"111101111",
  42762=>"111011001",
  42763=>"000000001",
  42764=>"000010110",
  42765=>"001110110",
  42766=>"000000011",
  42767=>"011011111",
  42768=>"010010111",
  42769=>"101010010",
  42770=>"101111110",
  42771=>"111110000",
  42772=>"001001101",
  42773=>"000110011",
  42774=>"101010011",
  42775=>"011000000",
  42776=>"001110110",
  42777=>"000101110",
  42778=>"110100100",
  42779=>"011100011",
  42780=>"111011011",
  42781=>"110010000",
  42782=>"000100111",
  42783=>"000101001",
  42784=>"111100001",
  42785=>"000110111",
  42786=>"111111110",
  42787=>"101000010",
  42788=>"111100100",
  42789=>"100001111",
  42790=>"000110010",
  42791=>"110010101",
  42792=>"101000010",
  42793=>"000110000",
  42794=>"111111111",
  42795=>"100011001",
  42796=>"000000100",
  42797=>"000101110",
  42798=>"111011101",
  42799=>"101101110",
  42800=>"000000011",
  42801=>"000110011",
  42802=>"101101001",
  42803=>"001101100",
  42804=>"110101111",
  42805=>"110111001",
  42806=>"110000110",
  42807=>"111000010",
  42808=>"000000111",
  42809=>"111110000",
  42810=>"001100001",
  42811=>"010111101",
  42812=>"111100000",
  42813=>"000100010",
  42814=>"111100111",
  42815=>"011001100",
  42816=>"000010101",
  42817=>"001001111",
  42818=>"001010011",
  42819=>"111011010",
  42820=>"000001110",
  42821=>"011000101",
  42822=>"110001000",
  42823=>"110001101",
  42824=>"100100000",
  42825=>"110111101",
  42826=>"100011000",
  42827=>"010100010",
  42828=>"101000001",
  42829=>"001111011",
  42830=>"010011100",
  42831=>"010111001",
  42832=>"010010111",
  42833=>"111100111",
  42834=>"000100011",
  42835=>"111101100",
  42836=>"100100010",
  42837=>"011000000",
  42838=>"111001111",
  42839=>"000010111",
  42840=>"000110011",
  42841=>"100111101",
  42842=>"010011001",
  42843=>"110000001",
  42844=>"111001111",
  42845=>"100111010",
  42846=>"110000111",
  42847=>"111100111",
  42848=>"110001010",
  42849=>"110010101",
  42850=>"110000110",
  42851=>"110011000",
  42852=>"111111010",
  42853=>"001001001",
  42854=>"101000100",
  42855=>"011110001",
  42856=>"010000010",
  42857=>"001101001",
  42858=>"010101110",
  42859=>"001101000",
  42860=>"011100000",
  42861=>"011101111",
  42862=>"000001000",
  42863=>"100111100",
  42864=>"100100000",
  42865=>"101100111",
  42866=>"100010110",
  42867=>"000111010",
  42868=>"100101010",
  42869=>"000101111",
  42870=>"010000100",
  42871=>"001001101",
  42872=>"101011100",
  42873=>"101101011",
  42874=>"010100111",
  42875=>"000000010",
  42876=>"001001100",
  42877=>"000011101",
  42878=>"110111110",
  42879=>"001100010",
  42880=>"000110101",
  42881=>"110000101",
  42882=>"010000111",
  42883=>"010011111",
  42884=>"101111110",
  42885=>"000110100",
  42886=>"001001001",
  42887=>"000011110",
  42888=>"111111101",
  42889=>"000110011",
  42890=>"000100000",
  42891=>"000000010",
  42892=>"010100111",
  42893=>"010100101",
  42894=>"000001001",
  42895=>"101100000",
  42896=>"100000110",
  42897=>"110011100",
  42898=>"001100000",
  42899=>"001000010",
  42900=>"100111001",
  42901=>"010111011",
  42902=>"100011000",
  42903=>"010100100",
  42904=>"111110100",
  42905=>"111010110",
  42906=>"010101010",
  42907=>"011110010",
  42908=>"000010001",
  42909=>"111111111",
  42910=>"111000100",
  42911=>"101110001",
  42912=>"110101110",
  42913=>"010011110",
  42914=>"001110011",
  42915=>"100010010",
  42916=>"000110111",
  42917=>"111000101",
  42918=>"111001111",
  42919=>"100000000",
  42920=>"111101110",
  42921=>"100111000",
  42922=>"001111110",
  42923=>"000000001",
  42924=>"010010010",
  42925=>"001001110",
  42926=>"110001110",
  42927=>"100000111",
  42928=>"110100101",
  42929=>"111110000",
  42930=>"011001110",
  42931=>"001010010",
  42932=>"001110001",
  42933=>"000011010",
  42934=>"011001101",
  42935=>"101001110",
  42936=>"101100011",
  42937=>"101000100",
  42938=>"101111111",
  42939=>"011101101",
  42940=>"101101000",
  42941=>"000101100",
  42942=>"000011010",
  42943=>"110101000",
  42944=>"000011001",
  42945=>"100010100",
  42946=>"100111000",
  42947=>"000101111",
  42948=>"101001101",
  42949=>"001111101",
  42950=>"110100011",
  42951=>"011101010",
  42952=>"001111001",
  42953=>"000101000",
  42954=>"010111000",
  42955=>"010101111",
  42956=>"010111011",
  42957=>"101010011",
  42958=>"100100000",
  42959=>"000101100",
  42960=>"001111010",
  42961=>"101111001",
  42962=>"000100100",
  42963=>"011100000",
  42964=>"000001100",
  42965=>"110101110",
  42966=>"010000001",
  42967=>"011010110",
  42968=>"011000000",
  42969=>"000011000",
  42970=>"000101111",
  42971=>"010000110",
  42972=>"111011010",
  42973=>"000000101",
  42974=>"000000010",
  42975=>"111000000",
  42976=>"111010000",
  42977=>"101010011",
  42978=>"000001110",
  42979=>"010000111",
  42980=>"011000100",
  42981=>"000101000",
  42982=>"011001101",
  42983=>"110111001",
  42984=>"101100000",
  42985=>"010010100",
  42986=>"010010010",
  42987=>"011101000",
  42988=>"000111111",
  42989=>"011101001",
  42990=>"010110000",
  42991=>"011000010",
  42992=>"010110111",
  42993=>"111000000",
  42994=>"101000110",
  42995=>"011111111",
  42996=>"100011010",
  42997=>"101101000",
  42998=>"000001011",
  42999=>"111111110",
  43000=>"011100001",
  43001=>"110001001",
  43002=>"111000101",
  43003=>"011101110",
  43004=>"110001000",
  43005=>"011100000",
  43006=>"001000000",
  43007=>"111100100",
  43008=>"101000100",
  43009=>"111001110",
  43010=>"010100101",
  43011=>"001111010",
  43012=>"010010101",
  43013=>"110101100",
  43014=>"000100010",
  43015=>"010000101",
  43016=>"000010100",
  43017=>"101001000",
  43018=>"101001111",
  43019=>"110111100",
  43020=>"101111110",
  43021=>"100100100",
  43022=>"010001001",
  43023=>"010100001",
  43024=>"011101110",
  43025=>"010000111",
  43026=>"001100011",
  43027=>"001001111",
  43028=>"100010000",
  43029=>"101011000",
  43030=>"111010110",
  43031=>"010111100",
  43032=>"000101000",
  43033=>"001010111",
  43034=>"111111011",
  43035=>"111010101",
  43036=>"101010000",
  43037=>"010010001",
  43038=>"011100101",
  43039=>"110011010",
  43040=>"111001100",
  43041=>"000010011",
  43042=>"100111110",
  43043=>"110100111",
  43044=>"011100110",
  43045=>"111001001",
  43046=>"010101100",
  43047=>"001110011",
  43048=>"110110101",
  43049=>"000010110",
  43050=>"000010000",
  43051=>"111111110",
  43052=>"010101100",
  43053=>"110001111",
  43054=>"111100011",
  43055=>"110000011",
  43056=>"001111101",
  43057=>"000100101",
  43058=>"011110111",
  43059=>"110011110",
  43060=>"000010000",
  43061=>"000101000",
  43062=>"111101100",
  43063=>"010101010",
  43064=>"111101011",
  43065=>"000101001",
  43066=>"100000101",
  43067=>"000000001",
  43068=>"000000000",
  43069=>"101000100",
  43070=>"011000011",
  43071=>"101011011",
  43072=>"101010000",
  43073=>"000110101",
  43074=>"111011010",
  43075=>"011110110",
  43076=>"111001001",
  43077=>"111011110",
  43078=>"011101110",
  43079=>"111011000",
  43080=>"110011101",
  43081=>"000110110",
  43082=>"100001000",
  43083=>"010001101",
  43084=>"000100110",
  43085=>"101100000",
  43086=>"111010111",
  43087=>"101110011",
  43088=>"100101101",
  43089=>"101001101",
  43090=>"000111100",
  43091=>"101000100",
  43092=>"010011111",
  43093=>"100000101",
  43094=>"101100111",
  43095=>"001110011",
  43096=>"000111001",
  43097=>"001111111",
  43098=>"000011111",
  43099=>"011010011",
  43100=>"110100101",
  43101=>"000100010",
  43102=>"111011011",
  43103=>"000100101",
  43104=>"001111011",
  43105=>"000101011",
  43106=>"111011111",
  43107=>"101000001",
  43108=>"000010001",
  43109=>"000101101",
  43110=>"110110100",
  43111=>"000111111",
  43112=>"100011101",
  43113=>"110010010",
  43114=>"100101001",
  43115=>"111000111",
  43116=>"000111111",
  43117=>"000010011",
  43118=>"010111010",
  43119=>"101010100",
  43120=>"000100000",
  43121=>"000011011",
  43122=>"010111110",
  43123=>"111001100",
  43124=>"110011000",
  43125=>"000110101",
  43126=>"010110000",
  43127=>"010011001",
  43128=>"001010001",
  43129=>"100000010",
  43130=>"000000101",
  43131=>"101000101",
  43132=>"010110011",
  43133=>"111101001",
  43134=>"000011100",
  43135=>"000001100",
  43136=>"000111001",
  43137=>"001011011",
  43138=>"101001010",
  43139=>"010110100",
  43140=>"011011001",
  43141=>"101111100",
  43142=>"110101100",
  43143=>"111111101",
  43144=>"101100101",
  43145=>"110010000",
  43146=>"101011001",
  43147=>"011110111",
  43148=>"110010001",
  43149=>"110111100",
  43150=>"111000000",
  43151=>"111100011",
  43152=>"000001111",
  43153=>"011101000",
  43154=>"000111100",
  43155=>"110110111",
  43156=>"100111001",
  43157=>"100010110",
  43158=>"101100111",
  43159=>"011101000",
  43160=>"101100000",
  43161=>"111100000",
  43162=>"110110011",
  43163=>"001100000",
  43164=>"101111000",
  43165=>"101010000",
  43166=>"101000010",
  43167=>"101111011",
  43168=>"000001110",
  43169=>"001011000",
  43170=>"000110010",
  43171=>"011110000",
  43172=>"101000011",
  43173=>"010000010",
  43174=>"010000010",
  43175=>"000000000",
  43176=>"111011001",
  43177=>"100110110",
  43178=>"110001111",
  43179=>"101011000",
  43180=>"110101100",
  43181=>"001111111",
  43182=>"010100000",
  43183=>"010011100",
  43184=>"000001000",
  43185=>"000111010",
  43186=>"010111100",
  43187=>"011000111",
  43188=>"101001010",
  43189=>"011100110",
  43190=>"111011001",
  43191=>"010111111",
  43192=>"010110001",
  43193=>"100011001",
  43194=>"100100001",
  43195=>"100001001",
  43196=>"100000111",
  43197=>"111110101",
  43198=>"111001111",
  43199=>"101010001",
  43200=>"100101110",
  43201=>"011101011",
  43202=>"010101110",
  43203=>"101100010",
  43204=>"111010001",
  43205=>"101100101",
  43206=>"010110010",
  43207=>"010011110",
  43208=>"100111100",
  43209=>"000100111",
  43210=>"100111101",
  43211=>"111111111",
  43212=>"001001110",
  43213=>"100101100",
  43214=>"110011100",
  43215=>"011111110",
  43216=>"000001111",
  43217=>"001111110",
  43218=>"101011111",
  43219=>"101000000",
  43220=>"101111101",
  43221=>"101000100",
  43222=>"011011011",
  43223=>"010111110",
  43224=>"000011111",
  43225=>"111011111",
  43226=>"110000110",
  43227=>"101110111",
  43228=>"111011010",
  43229=>"111001000",
  43230=>"100000100",
  43231=>"100111100",
  43232=>"000111111",
  43233=>"101001000",
  43234=>"110100001",
  43235=>"010000000",
  43236=>"101001000",
  43237=>"101110111",
  43238=>"011011010",
  43239=>"101001111",
  43240=>"111000011",
  43241=>"011111010",
  43242=>"110000000",
  43243=>"001111101",
  43244=>"101110001",
  43245=>"110010110",
  43246=>"101000000",
  43247=>"110100000",
  43248=>"000001111",
  43249=>"100000001",
  43250=>"111111100",
  43251=>"000001100",
  43252=>"111111111",
  43253=>"010101110",
  43254=>"000011100",
  43255=>"011000111",
  43256=>"010110110",
  43257=>"101000000",
  43258=>"010000001",
  43259=>"111100000",
  43260=>"011010010",
  43261=>"001101001",
  43262=>"011011100",
  43263=>"111111100",
  43264=>"101110100",
  43265=>"101010011",
  43266=>"010100000",
  43267=>"110000000",
  43268=>"000110001",
  43269=>"001011001",
  43270=>"111100001",
  43271=>"010011110",
  43272=>"100111000",
  43273=>"111101110",
  43274=>"011110010",
  43275=>"101100110",
  43276=>"010011000",
  43277=>"111110110",
  43278=>"101010101",
  43279=>"110110111",
  43280=>"110100101",
  43281=>"011011010",
  43282=>"111101111",
  43283=>"111110100",
  43284=>"101101110",
  43285=>"010011101",
  43286=>"001001110",
  43287=>"111110111",
  43288=>"000111111",
  43289=>"110111011",
  43290=>"010010000",
  43291=>"111010000",
  43292=>"000101010",
  43293=>"100000011",
  43294=>"101110111",
  43295=>"100001101",
  43296=>"000101011",
  43297=>"111001100",
  43298=>"010011011",
  43299=>"000010110",
  43300=>"010000101",
  43301=>"101011010",
  43302=>"100100000",
  43303=>"001111010",
  43304=>"001100101",
  43305=>"000010001",
  43306=>"010010011",
  43307=>"110000100",
  43308=>"110010111",
  43309=>"011111100",
  43310=>"000000100",
  43311=>"110010100",
  43312=>"110010010",
  43313=>"110001001",
  43314=>"111111000",
  43315=>"010000110",
  43316=>"000011111",
  43317=>"000000001",
  43318=>"101101010",
  43319=>"111111100",
  43320=>"101110001",
  43321=>"111110111",
  43322=>"000111011",
  43323=>"001001011",
  43324=>"001000000",
  43325=>"100011100",
  43326=>"001010100",
  43327=>"000010011",
  43328=>"010100101",
  43329=>"011000101",
  43330=>"101010000",
  43331=>"111001011",
  43332=>"110101100",
  43333=>"100100100",
  43334=>"110011101",
  43335=>"111011101",
  43336=>"000100110",
  43337=>"001010110",
  43338=>"000001011",
  43339=>"101111100",
  43340=>"011000001",
  43341=>"111001001",
  43342=>"010110100",
  43343=>"000110001",
  43344=>"101111000",
  43345=>"111100010",
  43346=>"111100111",
  43347=>"101100111",
  43348=>"111111011",
  43349=>"000001001",
  43350=>"111111100",
  43351=>"111001011",
  43352=>"111000001",
  43353=>"011101010",
  43354=>"010010010",
  43355=>"111000001",
  43356=>"100111011",
  43357=>"100100001",
  43358=>"000101000",
  43359=>"010011001",
  43360=>"111100100",
  43361=>"111001010",
  43362=>"011111100",
  43363=>"000010110",
  43364=>"101010111",
  43365=>"100111100",
  43366=>"000101001",
  43367=>"001111011",
  43368=>"001101101",
  43369=>"001011100",
  43370=>"001000011",
  43371=>"100111111",
  43372=>"101000011",
  43373=>"110000010",
  43374=>"010100111",
  43375=>"010100011",
  43376=>"111111001",
  43377=>"100100111",
  43378=>"010100101",
  43379=>"110000001",
  43380=>"000010100",
  43381=>"000110000",
  43382=>"000011100",
  43383=>"110000100",
  43384=>"111010101",
  43385=>"101110011",
  43386=>"001010000",
  43387=>"101110001",
  43388=>"111000001",
  43389=>"000110100",
  43390=>"111010010",
  43391=>"100111110",
  43392=>"101010001",
  43393=>"101001000",
  43394=>"011001010",
  43395=>"000010001",
  43396=>"000000000",
  43397=>"101100111",
  43398=>"010111111",
  43399=>"000010000",
  43400=>"100101001",
  43401=>"010010100",
  43402=>"001000011",
  43403=>"001000110",
  43404=>"100111101",
  43405=>"010010111",
  43406=>"101100110",
  43407=>"110100010",
  43408=>"010111110",
  43409=>"010110101",
  43410=>"010000000",
  43411=>"110111111",
  43412=>"111010011",
  43413=>"100000011",
  43414=>"000110111",
  43415=>"111000001",
  43416=>"000001110",
  43417=>"100000100",
  43418=>"111110000",
  43419=>"111000011",
  43420=>"011101110",
  43421=>"110100011",
  43422=>"100011110",
  43423=>"001000101",
  43424=>"111111110",
  43425=>"000010000",
  43426=>"011000001",
  43427=>"100101111",
  43428=>"010110111",
  43429=>"001001010",
  43430=>"111001101",
  43431=>"000100000",
  43432=>"011110111",
  43433=>"100100011",
  43434=>"000111000",
  43435=>"111000000",
  43436=>"010100011",
  43437=>"100001100",
  43438=>"011000111",
  43439=>"011110010",
  43440=>"110010001",
  43441=>"000011000",
  43442=>"011000100",
  43443=>"001011100",
  43444=>"010001010",
  43445=>"110000011",
  43446=>"001111011",
  43447=>"011101100",
  43448=>"011101111",
  43449=>"010101110",
  43450=>"000001010",
  43451=>"010011000",
  43452=>"101110101",
  43453=>"100100011",
  43454=>"011011100",
  43455=>"000011010",
  43456=>"111001100",
  43457=>"001101101",
  43458=>"111001111",
  43459=>"000111000",
  43460=>"010111111",
  43461=>"000100000",
  43462=>"110100011",
  43463=>"110010001",
  43464=>"111110000",
  43465=>"111011000",
  43466=>"001000001",
  43467=>"011000000",
  43468=>"011100101",
  43469=>"110111100",
  43470=>"100010001",
  43471=>"111101111",
  43472=>"010011001",
  43473=>"111000110",
  43474=>"101110110",
  43475=>"110010111",
  43476=>"011010011",
  43477=>"011011110",
  43478=>"000111000",
  43479=>"011100010",
  43480=>"110101000",
  43481=>"111010011",
  43482=>"010001110",
  43483=>"001100001",
  43484=>"001001001",
  43485=>"111100100",
  43486=>"000011101",
  43487=>"101001111",
  43488=>"101111011",
  43489=>"000100111",
  43490=>"111010101",
  43491=>"001100110",
  43492=>"011001010",
  43493=>"111000000",
  43494=>"011001000",
  43495=>"101101011",
  43496=>"001011101",
  43497=>"110000100",
  43498=>"101111100",
  43499=>"010100010",
  43500=>"110111111",
  43501=>"110101100",
  43502=>"110100000",
  43503=>"001001110",
  43504=>"010011111",
  43505=>"110111011",
  43506=>"001111000",
  43507=>"010011000",
  43508=>"111001000",
  43509=>"011100011",
  43510=>"100001001",
  43511=>"011000011",
  43512=>"110100110",
  43513=>"100101101",
  43514=>"000011011",
  43515=>"110110100",
  43516=>"110010001",
  43517=>"111111110",
  43518=>"100010101",
  43519=>"110010011",
  43520=>"100100010",
  43521=>"110001010",
  43522=>"001101100",
  43523=>"010100001",
  43524=>"011110011",
  43525=>"110010101",
  43526=>"010010111",
  43527=>"111011100",
  43528=>"101011110",
  43529=>"110011111",
  43530=>"100011011",
  43531=>"101110100",
  43532=>"010101111",
  43533=>"111010000",
  43534=>"001100110",
  43535=>"010001010",
  43536=>"011100110",
  43537=>"000001001",
  43538=>"111111001",
  43539=>"111001000",
  43540=>"001001000",
  43541=>"010010101",
  43542=>"000001110",
  43543=>"010010001",
  43544=>"110011000",
  43545=>"011000000",
  43546=>"001000000",
  43547=>"010100100",
  43548=>"110001100",
  43549=>"101011001",
  43550=>"101000101",
  43551=>"110110110",
  43552=>"110010001",
  43553=>"010001101",
  43554=>"101111101",
  43555=>"101111010",
  43556=>"011000110",
  43557=>"001001001",
  43558=>"011100001",
  43559=>"111110000",
  43560=>"111100101",
  43561=>"101001000",
  43562=>"011000110",
  43563=>"000010010",
  43564=>"100001001",
  43565=>"110001000",
  43566=>"101101110",
  43567=>"000000001",
  43568=>"000010010",
  43569=>"011011000",
  43570=>"100100101",
  43571=>"100001110",
  43572=>"110011100",
  43573=>"000001011",
  43574=>"110101111",
  43575=>"000001101",
  43576=>"011010110",
  43577=>"101010100",
  43578=>"001010010",
  43579=>"010000110",
  43580=>"000010100",
  43581=>"001101110",
  43582=>"110101001",
  43583=>"000101101",
  43584=>"001011000",
  43585=>"011111110",
  43586=>"010001000",
  43587=>"010101111",
  43588=>"011101000",
  43589=>"000011110",
  43590=>"000010000",
  43591=>"111101111",
  43592=>"000111110",
  43593=>"100111000",
  43594=>"001000010",
  43595=>"001111000",
  43596=>"110101011",
  43597=>"101100111",
  43598=>"001001110",
  43599=>"101010001",
  43600=>"100101001",
  43601=>"110010111",
  43602=>"111101110",
  43603=>"011110000",
  43604=>"010100011",
  43605=>"101101000",
  43606=>"001101101",
  43607=>"110111010",
  43608=>"010011010",
  43609=>"100110111",
  43610=>"000011001",
  43611=>"100010000",
  43612=>"100010000",
  43613=>"001010010",
  43614=>"011010010",
  43615=>"110010010",
  43616=>"101110110",
  43617=>"001001010",
  43618=>"000010011",
  43619=>"101111111",
  43620=>"001001011",
  43621=>"100000010",
  43622=>"100000000",
  43623=>"011100001",
  43624=>"000001000",
  43625=>"111000011",
  43626=>"111101011",
  43627=>"001010110",
  43628=>"001111010",
  43629=>"101011101",
  43630=>"011101100",
  43631=>"000100111",
  43632=>"001111000",
  43633=>"010100001",
  43634=>"011101110",
  43635=>"100100011",
  43636=>"001100000",
  43637=>"011111111",
  43638=>"001100110",
  43639=>"001100000",
  43640=>"101010010",
  43641=>"100010000",
  43642=>"110111101",
  43643=>"111010101",
  43644=>"001111100",
  43645=>"001110101",
  43646=>"000010111",
  43647=>"110100000",
  43648=>"101000100",
  43649=>"111001101",
  43650=>"101110111",
  43651=>"001001100",
  43652=>"001011101",
  43653=>"011011101",
  43654=>"001000110",
  43655=>"111001101",
  43656=>"001001001",
  43657=>"100100000",
  43658=>"111000111",
  43659=>"100011011",
  43660=>"010010000",
  43661=>"000101001",
  43662=>"101111001",
  43663=>"111000000",
  43664=>"101110100",
  43665=>"101111001",
  43666=>"111101011",
  43667=>"101111100",
  43668=>"100011100",
  43669=>"101010011",
  43670=>"110001110",
  43671=>"100100010",
  43672=>"110000100",
  43673=>"011100111",
  43674=>"110101010",
  43675=>"101101101",
  43676=>"110101000",
  43677=>"101010010",
  43678=>"110100110",
  43679=>"000100111",
  43680=>"101111111",
  43681=>"100100101",
  43682=>"110010110",
  43683=>"111001100",
  43684=>"110000100",
  43685=>"011010000",
  43686=>"011100111",
  43687=>"001101110",
  43688=>"010100000",
  43689=>"100101100",
  43690=>"100000000",
  43691=>"001011101",
  43692=>"110110111",
  43693=>"101100011",
  43694=>"110100101",
  43695=>"100010110",
  43696=>"011111111",
  43697=>"111100011",
  43698=>"011000110",
  43699=>"011010001",
  43700=>"000001111",
  43701=>"011100111",
  43702=>"111100010",
  43703=>"011101000",
  43704=>"011011100",
  43705=>"110011100",
  43706=>"011011010",
  43707=>"000000001",
  43708=>"100010001",
  43709=>"010011000",
  43710=>"000000000",
  43711=>"101000100",
  43712=>"110100101",
  43713=>"010010000",
  43714=>"001110100",
  43715=>"101101011",
  43716=>"011001001",
  43717=>"011110000",
  43718=>"001111111",
  43719=>"001011110",
  43720=>"111100001",
  43721=>"101011100",
  43722=>"101100110",
  43723=>"001011111",
  43724=>"101101011",
  43725=>"100000110",
  43726=>"001010011",
  43727=>"110111001",
  43728=>"000000101",
  43729=>"101000011",
  43730=>"000000111",
  43731=>"000101000",
  43732=>"101001001",
  43733=>"010001110",
  43734=>"101100111",
  43735=>"110110000",
  43736=>"000110010",
  43737=>"001000011",
  43738=>"111011010",
  43739=>"010011110",
  43740=>"100001111",
  43741=>"001010100",
  43742=>"001011000",
  43743=>"010010110",
  43744=>"000011111",
  43745=>"011011000",
  43746=>"111110100",
  43747=>"000001111",
  43748=>"100010101",
  43749=>"100011111",
  43750=>"000110100",
  43751=>"011110000",
  43752=>"010010000",
  43753=>"001110100",
  43754=>"100010001",
  43755=>"111101111",
  43756=>"011100101",
  43757=>"001101100",
  43758=>"101000011",
  43759=>"111100101",
  43760=>"011101111",
  43761=>"001010001",
  43762=>"110100110",
  43763=>"010110010",
  43764=>"000001011",
  43765=>"111011111",
  43766=>"111011000",
  43767=>"000101001",
  43768=>"111000110",
  43769=>"111111111",
  43770=>"111010110",
  43771=>"101100000",
  43772=>"100000011",
  43773=>"111000100",
  43774=>"111010100",
  43775=>"111111100",
  43776=>"101101111",
  43777=>"100001111",
  43778=>"000101011",
  43779=>"111100101",
  43780=>"111111110",
  43781=>"101010001",
  43782=>"010101111",
  43783=>"010111011",
  43784=>"000001000",
  43785=>"010110110",
  43786=>"000000100",
  43787=>"100001011",
  43788=>"110001101",
  43789=>"100101011",
  43790=>"101010010",
  43791=>"100100111",
  43792=>"111011000",
  43793=>"100000010",
  43794=>"001101011",
  43795=>"010100101",
  43796=>"011001110",
  43797=>"101110011",
  43798=>"010011010",
  43799=>"000000011",
  43800=>"110011110",
  43801=>"101000000",
  43802=>"000000011",
  43803=>"011011111",
  43804=>"000010101",
  43805=>"001110110",
  43806=>"001011111",
  43807=>"011111111",
  43808=>"011100111",
  43809=>"011000101",
  43810=>"101000111",
  43811=>"101110101",
  43812=>"001101111",
  43813=>"011100100",
  43814=>"000001101",
  43815=>"011111010",
  43816=>"001100111",
  43817=>"111010111",
  43818=>"011100100",
  43819=>"011110010",
  43820=>"100001000",
  43821=>"010110000",
  43822=>"110100111",
  43823=>"100111011",
  43824=>"101101010",
  43825=>"101111011",
  43826=>"100101000",
  43827=>"100100101",
  43828=>"010100010",
  43829=>"000001101",
  43830=>"000000101",
  43831=>"110001011",
  43832=>"101110111",
  43833=>"101000000",
  43834=>"111010000",
  43835=>"100111110",
  43836=>"111000011",
  43837=>"001001100",
  43838=>"010100101",
  43839=>"111110101",
  43840=>"000011011",
  43841=>"001000001",
  43842=>"100110011",
  43843=>"111001101",
  43844=>"010111100",
  43845=>"011011001",
  43846=>"110001111",
  43847=>"101000010",
  43848=>"100010110",
  43849=>"000101100",
  43850=>"000000010",
  43851=>"111110001",
  43852=>"111100110",
  43853=>"110011011",
  43854=>"111100000",
  43855=>"001011101",
  43856=>"111110010",
  43857=>"101111000",
  43858=>"001111000",
  43859=>"010000100",
  43860=>"010000100",
  43861=>"110010110",
  43862=>"010101010",
  43863=>"101100101",
  43864=>"010011101",
  43865=>"110000111",
  43866=>"101111001",
  43867=>"101101011",
  43868=>"001101011",
  43869=>"001111111",
  43870=>"001000001",
  43871=>"000010110",
  43872=>"111100110",
  43873=>"101111111",
  43874=>"001000100",
  43875=>"000000010",
  43876=>"100110100",
  43877=>"101010011",
  43878=>"101000110",
  43879=>"100001101",
  43880=>"110100100",
  43881=>"100001010",
  43882=>"100010010",
  43883=>"101000111",
  43884=>"010110001",
  43885=>"111110111",
  43886=>"000111001",
  43887=>"110010011",
  43888=>"100111010",
  43889=>"110110111",
  43890=>"101111010",
  43891=>"100110010",
  43892=>"011000000",
  43893=>"100011011",
  43894=>"101011000",
  43895=>"111111100",
  43896=>"011010100",
  43897=>"101001001",
  43898=>"111010110",
  43899=>"001100100",
  43900=>"110000110",
  43901=>"101011110",
  43902=>"010001100",
  43903=>"110111110",
  43904=>"000110110",
  43905=>"010011000",
  43906=>"000011000",
  43907=>"100101000",
  43908=>"010110111",
  43909=>"100000011",
  43910=>"001111010",
  43911=>"110000011",
  43912=>"110101100",
  43913=>"111010000",
  43914=>"001000001",
  43915=>"110011100",
  43916=>"110101111",
  43917=>"110111100",
  43918=>"000000100",
  43919=>"110110110",
  43920=>"000011111",
  43921=>"101000000",
  43922=>"001100000",
  43923=>"011010100",
  43924=>"111100011",
  43925=>"101011000",
  43926=>"100100110",
  43927=>"100110100",
  43928=>"110100100",
  43929=>"111101010",
  43930=>"110101111",
  43931=>"100001110",
  43932=>"011010110",
  43933=>"010101111",
  43934=>"010011001",
  43935=>"111000100",
  43936=>"111000000",
  43937=>"101011111",
  43938=>"001001101",
  43939=>"010010011",
  43940=>"111100111",
  43941=>"101011111",
  43942=>"001011110",
  43943=>"110010011",
  43944=>"010001100",
  43945=>"111010111",
  43946=>"110010010",
  43947=>"001101000",
  43948=>"100111101",
  43949=>"100001101",
  43950=>"100110100",
  43951=>"110110011",
  43952=>"001010000",
  43953=>"010001101",
  43954=>"000110100",
  43955=>"010111111",
  43956=>"111110110",
  43957=>"111011100",
  43958=>"001001101",
  43959=>"000110111",
  43960=>"000101010",
  43961=>"111010101",
  43962=>"110000010",
  43963=>"101001101",
  43964=>"110110111",
  43965=>"100101101",
  43966=>"001011000",
  43967=>"000000000",
  43968=>"001110110",
  43969=>"111111000",
  43970=>"001001110",
  43971=>"111011111",
  43972=>"111110101",
  43973=>"110010100",
  43974=>"110001111",
  43975=>"111000100",
  43976=>"100110110",
  43977=>"010010011",
  43978=>"011000111",
  43979=>"010110011",
  43980=>"111111010",
  43981=>"111110001",
  43982=>"100010100",
  43983=>"101100011",
  43984=>"101000111",
  43985=>"000001000",
  43986=>"101100010",
  43987=>"000000100",
  43988=>"100011111",
  43989=>"001011111",
  43990=>"001011001",
  43991=>"101001110",
  43992=>"001001111",
  43993=>"011111111",
  43994=>"101000010",
  43995=>"011011110",
  43996=>"000101101",
  43997=>"010100101",
  43998=>"111001111",
  43999=>"111111010",
  44000=>"010100101",
  44001=>"011000011",
  44002=>"001001111",
  44003=>"000101000",
  44004=>"010000100",
  44005=>"111001011",
  44006=>"101000111",
  44007=>"111100101",
  44008=>"001111010",
  44009=>"101110100",
  44010=>"100010100",
  44011=>"001010101",
  44012=>"100000010",
  44013=>"111001010",
  44014=>"011100101",
  44015=>"101000100",
  44016=>"000100000",
  44017=>"000010010",
  44018=>"011101110",
  44019=>"001010100",
  44020=>"111011101",
  44021=>"100010011",
  44022=>"100001110",
  44023=>"111011101",
  44024=>"010110010",
  44025=>"001011111",
  44026=>"011111110",
  44027=>"000110100",
  44028=>"111101111",
  44029=>"000010011",
  44030=>"101010001",
  44031=>"100111110",
  44032=>"001000110",
  44033=>"001101000",
  44034=>"101110110",
  44035=>"101110101",
  44036=>"010111010",
  44037=>"001100000",
  44038=>"101110010",
  44039=>"110000000",
  44040=>"110010011",
  44041=>"001010010",
  44042=>"000110001",
  44043=>"111110011",
  44044=>"011111100",
  44045=>"000000000",
  44046=>"110100001",
  44047=>"111111011",
  44048=>"110010001",
  44049=>"100111111",
  44050=>"000100010",
  44051=>"110011101",
  44052=>"011000010",
  44053=>"011000010",
  44054=>"101101111",
  44055=>"001000111",
  44056=>"101101101",
  44057=>"000100101",
  44058=>"100011110",
  44059=>"010110111",
  44060=>"001110001",
  44061=>"001100011",
  44062=>"001100101",
  44063=>"000011001",
  44064=>"110100001",
  44065=>"100011110",
  44066=>"001000111",
  44067=>"000001010",
  44068=>"001111111",
  44069=>"110111100",
  44070=>"010101101",
  44071=>"100000100",
  44072=>"010111011",
  44073=>"101101100",
  44074=>"000101000",
  44075=>"110100101",
  44076=>"100110010",
  44077=>"010100011",
  44078=>"111100101",
  44079=>"101001111",
  44080=>"101100010",
  44081=>"101001101",
  44082=>"001101111",
  44083=>"111101010",
  44084=>"110000101",
  44085=>"001101001",
  44086=>"011100000",
  44087=>"011001111",
  44088=>"101101000",
  44089=>"110111010",
  44090=>"000010001",
  44091=>"000011000",
  44092=>"000100101",
  44093=>"100101001",
  44094=>"100101001",
  44095=>"111100010",
  44096=>"000001010",
  44097=>"000001011",
  44098=>"010111111",
  44099=>"100011101",
  44100=>"010111000",
  44101=>"001001001",
  44102=>"010011100",
  44103=>"001011111",
  44104=>"111101100",
  44105=>"101011011",
  44106=>"001011010",
  44107=>"111011110",
  44108=>"100011110",
  44109=>"110010100",
  44110=>"110001011",
  44111=>"110000010",
  44112=>"110001001",
  44113=>"110110011",
  44114=>"011100100",
  44115=>"010010101",
  44116=>"011001000",
  44117=>"111111000",
  44118=>"011001110",
  44119=>"001011011",
  44120=>"101010011",
  44121=>"100110100",
  44122=>"001011011",
  44123=>"011101110",
  44124=>"001000001",
  44125=>"010100001",
  44126=>"010110011",
  44127=>"101000101",
  44128=>"010001011",
  44129=>"100110001",
  44130=>"010001100",
  44131=>"001111111",
  44132=>"110111000",
  44133=>"000001010",
  44134=>"001101000",
  44135=>"110011100",
  44136=>"001001110",
  44137=>"001110011",
  44138=>"001111100",
  44139=>"110011010",
  44140=>"101011110",
  44141=>"000000000",
  44142=>"100101011",
  44143=>"000001101",
  44144=>"000000011",
  44145=>"101111111",
  44146=>"000001000",
  44147=>"010001010",
  44148=>"101110101",
  44149=>"001111101",
  44150=>"110100001",
  44151=>"110000011",
  44152=>"000111101",
  44153=>"001010001",
  44154=>"101000001",
  44155=>"100001100",
  44156=>"111011100",
  44157=>"110001101",
  44158=>"101110110",
  44159=>"000110000",
  44160=>"100111010",
  44161=>"110111010",
  44162=>"010100011",
  44163=>"000010011",
  44164=>"101100110",
  44165=>"111111110",
  44166=>"100100111",
  44167=>"001011100",
  44168=>"101110110",
  44169=>"111100100",
  44170=>"100100010",
  44171=>"001011011",
  44172=>"111100100",
  44173=>"100000010",
  44174=>"001100011",
  44175=>"001110010",
  44176=>"011000010",
  44177=>"101100100",
  44178=>"110111000",
  44179=>"010001011",
  44180=>"010100101",
  44181=>"100011110",
  44182=>"011101010",
  44183=>"011101001",
  44184=>"010010110",
  44185=>"001110110",
  44186=>"011101111",
  44187=>"110001010",
  44188=>"100111001",
  44189=>"110000010",
  44190=>"110100100",
  44191=>"110001010",
  44192=>"101101011",
  44193=>"111001001",
  44194=>"010101011",
  44195=>"101101110",
  44196=>"011001100",
  44197=>"010001000",
  44198=>"000101001",
  44199=>"010111000",
  44200=>"010000100",
  44201=>"011100110",
  44202=>"000101011",
  44203=>"101101110",
  44204=>"001111001",
  44205=>"101100001",
  44206=>"001101101",
  44207=>"101000000",
  44208=>"101101100",
  44209=>"000111000",
  44210=>"000101111",
  44211=>"100111110",
  44212=>"000001010",
  44213=>"001000000",
  44214=>"011000001",
  44215=>"100111001",
  44216=>"011011111",
  44217=>"100001000",
  44218=>"111111101",
  44219=>"001000010",
  44220=>"011010001",
  44221=>"001100111",
  44222=>"001110111",
  44223=>"011111000",
  44224=>"110100011",
  44225=>"000110011",
  44226=>"001100001",
  44227=>"111101001",
  44228=>"110001110",
  44229=>"001000011",
  44230=>"111000001",
  44231=>"100101001",
  44232=>"111111101",
  44233=>"111110011",
  44234=>"000011001",
  44235=>"100100001",
  44236=>"011011100",
  44237=>"100110101",
  44238=>"000101001",
  44239=>"001101111",
  44240=>"000100111",
  44241=>"100101100",
  44242=>"101110001",
  44243=>"001010000",
  44244=>"110000001",
  44245=>"001110001",
  44246=>"010001100",
  44247=>"111010001",
  44248=>"100010010",
  44249=>"000110010",
  44250=>"011110010",
  44251=>"010001011",
  44252=>"000011110",
  44253=>"010001010",
  44254=>"010000001",
  44255=>"010001111",
  44256=>"000100101",
  44257=>"101101001",
  44258=>"010101101",
  44259=>"111000011",
  44260=>"111101000",
  44261=>"111101101",
  44262=>"011011101",
  44263=>"101100101",
  44264=>"000001010",
  44265=>"100101011",
  44266=>"001001111",
  44267=>"011001001",
  44268=>"111001010",
  44269=>"001100100",
  44270=>"100001011",
  44271=>"111110111",
  44272=>"100001111",
  44273=>"110011010",
  44274=>"001111011",
  44275=>"000101001",
  44276=>"101100101",
  44277=>"001001000",
  44278=>"100011100",
  44279=>"001000010",
  44280=>"000011000",
  44281=>"001111001",
  44282=>"100011111",
  44283=>"100101011",
  44284=>"110000110",
  44285=>"111011010",
  44286=>"110111101",
  44287=>"111100100",
  44288=>"001110101",
  44289=>"101000111",
  44290=>"111110001",
  44291=>"100000110",
  44292=>"110100101",
  44293=>"110001000",
  44294=>"101011000",
  44295=>"101100101",
  44296=>"000001010",
  44297=>"001111101",
  44298=>"111100100",
  44299=>"110000111",
  44300=>"000100000",
  44301=>"010101100",
  44302=>"000000000",
  44303=>"011110000",
  44304=>"011101100",
  44305=>"110011110",
  44306=>"100000001",
  44307=>"010111100",
  44308=>"000101100",
  44309=>"000101010",
  44310=>"010000010",
  44311=>"000011001",
  44312=>"011100101",
  44313=>"101111011",
  44314=>"000001101",
  44315=>"111011000",
  44316=>"100110010",
  44317=>"101111111",
  44318=>"110001001",
  44319=>"011000100",
  44320=>"011011100",
  44321=>"110111010",
  44322=>"000101110",
  44323=>"101011110",
  44324=>"110110101",
  44325=>"111111010",
  44326=>"101001000",
  44327=>"100111011",
  44328=>"010101010",
  44329=>"101010101",
  44330=>"001100100",
  44331=>"101011001",
  44332=>"101001001",
  44333=>"001110100",
  44334=>"110100001",
  44335=>"000101001",
  44336=>"100011010",
  44337=>"010110000",
  44338=>"101100110",
  44339=>"001010000",
  44340=>"000011100",
  44341=>"100000010",
  44342=>"110010110",
  44343=>"101111111",
  44344=>"100100011",
  44345=>"111000110",
  44346=>"000110011",
  44347=>"011100101",
  44348=>"000000111",
  44349=>"010110110",
  44350=>"011010100",
  44351=>"010101100",
  44352=>"011101111",
  44353=>"001011010",
  44354=>"011111001",
  44355=>"000001101",
  44356=>"111111101",
  44357=>"000110001",
  44358=>"010111010",
  44359=>"110100100",
  44360=>"010001010",
  44361=>"000000100",
  44362=>"111111001",
  44363=>"110111101",
  44364=>"011100011",
  44365=>"010001000",
  44366=>"001010001",
  44367=>"100100100",
  44368=>"000011001",
  44369=>"001110010",
  44370=>"110111010",
  44371=>"000011110",
  44372=>"101001001",
  44373=>"100101011",
  44374=>"101001011",
  44375=>"011101100",
  44376=>"110000001",
  44377=>"001101000",
  44378=>"011111011",
  44379=>"001001100",
  44380=>"000101001",
  44381=>"101111101",
  44382=>"011100100",
  44383=>"010111111",
  44384=>"111010011",
  44385=>"110010010",
  44386=>"010100010",
  44387=>"111111011",
  44388=>"110001100",
  44389=>"100111101",
  44390=>"100000001",
  44391=>"010101111",
  44392=>"001010010",
  44393=>"111110110",
  44394=>"011100110",
  44395=>"011101101",
  44396=>"010001000",
  44397=>"001011111",
  44398=>"111110110",
  44399=>"001000100",
  44400=>"000111011",
  44401=>"001100000",
  44402=>"110001101",
  44403=>"010101100",
  44404=>"000110100",
  44405=>"101010011",
  44406=>"111111110",
  44407=>"100101101",
  44408=>"010110101",
  44409=>"100001011",
  44410=>"010010101",
  44411=>"001111001",
  44412=>"011011100",
  44413=>"001101010",
  44414=>"001110111",
  44415=>"110000101",
  44416=>"111101000",
  44417=>"000101000",
  44418=>"011101010",
  44419=>"000111110",
  44420=>"000100101",
  44421=>"000000011",
  44422=>"010011001",
  44423=>"110100001",
  44424=>"001100011",
  44425=>"100111010",
  44426=>"101010001",
  44427=>"111001000",
  44428=>"000000011",
  44429=>"010111010",
  44430=>"000000011",
  44431=>"100011011",
  44432=>"001001110",
  44433=>"000001011",
  44434=>"010010011",
  44435=>"000011111",
  44436=>"111101110",
  44437=>"010111101",
  44438=>"000000000",
  44439=>"000111001",
  44440=>"001110100",
  44441=>"100010110",
  44442=>"000110110",
  44443=>"101100001",
  44444=>"110000111",
  44445=>"001010100",
  44446=>"001100011",
  44447=>"001001010",
  44448=>"101000001",
  44449=>"000011001",
  44450=>"010001100",
  44451=>"101101010",
  44452=>"011000110",
  44453=>"100010010",
  44454=>"111000110",
  44455=>"100110011",
  44456=>"000110001",
  44457=>"001100111",
  44458=>"100011001",
  44459=>"000011101",
  44460=>"101100000",
  44461=>"100000001",
  44462=>"000111010",
  44463=>"100001100",
  44464=>"011110110",
  44465=>"010000001",
  44466=>"101110001",
  44467=>"101000011",
  44468=>"010110110",
  44469=>"111110101",
  44470=>"010110010",
  44471=>"100011101",
  44472=>"101001000",
  44473=>"011000000",
  44474=>"011110110",
  44475=>"110110111",
  44476=>"101101001",
  44477=>"000010011",
  44478=>"001000011",
  44479=>"110001111",
  44480=>"111100110",
  44481=>"001110001",
  44482=>"011101011",
  44483=>"111101110",
  44484=>"011010000",
  44485=>"110111110",
  44486=>"001010010",
  44487=>"100101111",
  44488=>"101001001",
  44489=>"010000100",
  44490=>"001100110",
  44491=>"010110011",
  44492=>"111011101",
  44493=>"110011101",
  44494=>"101011110",
  44495=>"110101111",
  44496=>"110000111",
  44497=>"000001111",
  44498=>"010111110",
  44499=>"100100111",
  44500=>"100111011",
  44501=>"010101111",
  44502=>"100101101",
  44503=>"010011000",
  44504=>"010011100",
  44505=>"000001010",
  44506=>"010111000",
  44507=>"101010010",
  44508=>"011010011",
  44509=>"100001001",
  44510=>"101001000",
  44511=>"000000000",
  44512=>"111010010",
  44513=>"011010000",
  44514=>"100010001",
  44515=>"110011111",
  44516=>"000111100",
  44517=>"100101010",
  44518=>"011010001",
  44519=>"111001110",
  44520=>"001101011",
  44521=>"100010111",
  44522=>"010110001",
  44523=>"010011011",
  44524=>"011001110",
  44525=>"000100001",
  44526=>"110010100",
  44527=>"011010101",
  44528=>"111011011",
  44529=>"111111111",
  44530=>"101111010",
  44531=>"101100000",
  44532=>"010100110",
  44533=>"011000101",
  44534=>"110011100",
  44535=>"110110110",
  44536=>"001010111",
  44537=>"100010001",
  44538=>"100100000",
  44539=>"011101100",
  44540=>"011100000",
  44541=>"100001000",
  44542=>"110000110",
  44543=>"111001011",
  44544=>"101011001",
  44545=>"001010110",
  44546=>"010111000",
  44547=>"011000101",
  44548=>"011110100",
  44549=>"101101100",
  44550=>"110111100",
  44551=>"011100100",
  44552=>"010000001",
  44553=>"000101001",
  44554=>"101101101",
  44555=>"101101010",
  44556=>"100000101",
  44557=>"101001111",
  44558=>"000000010",
  44559=>"000000110",
  44560=>"001011000",
  44561=>"101110000",
  44562=>"000000011",
  44563=>"100111010",
  44564=>"011011011",
  44565=>"010001001",
  44566=>"110001100",
  44567=>"010000010",
  44568=>"100010100",
  44569=>"100000011",
  44570=>"001000111",
  44571=>"110010000",
  44572=>"000101100",
  44573=>"011010101",
  44574=>"010010010",
  44575=>"100101111",
  44576=>"110100000",
  44577=>"101000000",
  44578=>"000101111",
  44579=>"011110000",
  44580=>"111111010",
  44581=>"001100100",
  44582=>"000001000",
  44583=>"011101000",
  44584=>"100100010",
  44585=>"111111001",
  44586=>"011111011",
  44587=>"111010001",
  44588=>"101111111",
  44589=>"000110100",
  44590=>"000010111",
  44591=>"010001100",
  44592=>"011111010",
  44593=>"011010111",
  44594=>"011100001",
  44595=>"111000010",
  44596=>"110001110",
  44597=>"010010110",
  44598=>"101011001",
  44599=>"101111111",
  44600=>"011110010",
  44601=>"111111111",
  44602=>"001011011",
  44603=>"100110000",
  44604=>"110111110",
  44605=>"110000110",
  44606=>"011110101",
  44607=>"110101101",
  44608=>"101111101",
  44609=>"000010111",
  44610=>"001101010",
  44611=>"010001110",
  44612=>"010011001",
  44613=>"101001000",
  44614=>"001111111",
  44615=>"111111110",
  44616=>"011101010",
  44617=>"011010011",
  44618=>"111000111",
  44619=>"010111000",
  44620=>"000111011",
  44621=>"001100001",
  44622=>"110000000",
  44623=>"010101110",
  44624=>"011001000",
  44625=>"110011101",
  44626=>"011001001",
  44627=>"001011111",
  44628=>"011101010",
  44629=>"011010001",
  44630=>"111101001",
  44631=>"110100111",
  44632=>"111100011",
  44633=>"110001000",
  44634=>"100001101",
  44635=>"011111100",
  44636=>"100100100",
  44637=>"100101110",
  44638=>"111000000",
  44639=>"011010110",
  44640=>"100011100",
  44641=>"001011011",
  44642=>"100010011",
  44643=>"010010110",
  44644=>"010111010",
  44645=>"101110101",
  44646=>"001000100",
  44647=>"010001010",
  44648=>"001000011",
  44649=>"001111100",
  44650=>"011010011",
  44651=>"001111111",
  44652=>"010011011",
  44653=>"001011101",
  44654=>"000101000",
  44655=>"111100000",
  44656=>"100111011",
  44657=>"001101000",
  44658=>"011000110",
  44659=>"010011110",
  44660=>"100011010",
  44661=>"001001100",
  44662=>"000000010",
  44663=>"111011010",
  44664=>"010010111",
  44665=>"101001000",
  44666=>"101011010",
  44667=>"001101111",
  44668=>"010111011",
  44669=>"101101100",
  44670=>"101111100",
  44671=>"101000001",
  44672=>"101100000",
  44673=>"101110101",
  44674=>"010101000",
  44675=>"010111111",
  44676=>"111011100",
  44677=>"001110001",
  44678=>"111011001",
  44679=>"111011010",
  44680=>"001000010",
  44681=>"001011010",
  44682=>"100010001",
  44683=>"010011000",
  44684=>"101110000",
  44685=>"100010000",
  44686=>"000000010",
  44687=>"000101101",
  44688=>"001101101",
  44689=>"011000101",
  44690=>"011000110",
  44691=>"010011110",
  44692=>"111110001",
  44693=>"100000100",
  44694=>"010001111",
  44695=>"100100111",
  44696=>"001111010",
  44697=>"011000101",
  44698=>"000001101",
  44699=>"111111001",
  44700=>"010010110",
  44701=>"101110110",
  44702=>"010000001",
  44703=>"110010100",
  44704=>"010011001",
  44705=>"010001110",
  44706=>"111110000",
  44707=>"101000011",
  44708=>"111011010",
  44709=>"000011101",
  44710=>"000000100",
  44711=>"001001000",
  44712=>"010110100",
  44713=>"000000001",
  44714=>"000101110",
  44715=>"000100000",
  44716=>"101110010",
  44717=>"101010000",
  44718=>"000000100",
  44719=>"011001110",
  44720=>"001111110",
  44721=>"001101110",
  44722=>"011110011",
  44723=>"110001111",
  44724=>"010000010",
  44725=>"110100110",
  44726=>"000111000",
  44727=>"011111101",
  44728=>"001111111",
  44729=>"010010110",
  44730=>"111110010",
  44731=>"000111101",
  44732=>"001100011",
  44733=>"000110001",
  44734=>"001100001",
  44735=>"100000100",
  44736=>"100110010",
  44737=>"010001111",
  44738=>"110110110",
  44739=>"111111011",
  44740=>"000010110",
  44741=>"000100001",
  44742=>"101100011",
  44743=>"110010111",
  44744=>"100010000",
  44745=>"110110100",
  44746=>"011001010",
  44747=>"100001101",
  44748=>"000100101",
  44749=>"010100101",
  44750=>"100011001",
  44751=>"011011111",
  44752=>"100110100",
  44753=>"000100000",
  44754=>"010101111",
  44755=>"001110101",
  44756=>"110100111",
  44757=>"001011001",
  44758=>"000011100",
  44759=>"010000010",
  44760=>"000010111",
  44761=>"000100010",
  44762=>"100101010",
  44763=>"000001011",
  44764=>"111100001",
  44765=>"100110011",
  44766=>"001100110",
  44767=>"100000110",
  44768=>"001001101",
  44769=>"101001111",
  44770=>"111000111",
  44771=>"000111011",
  44772=>"101110001",
  44773=>"110110101",
  44774=>"100001110",
  44775=>"010010000",
  44776=>"100000101",
  44777=>"010100000",
  44778=>"011111100",
  44779=>"011000111",
  44780=>"110011111",
  44781=>"001101010",
  44782=>"110111000",
  44783=>"111111111",
  44784=>"110010111",
  44785=>"010100100",
  44786=>"110010000",
  44787=>"101010111",
  44788=>"111011101",
  44789=>"100100000",
  44790=>"000101010",
  44791=>"111010111",
  44792=>"000000100",
  44793=>"111010100",
  44794=>"011001011",
  44795=>"000011100",
  44796=>"011011011",
  44797=>"000101110",
  44798=>"011101011",
  44799=>"001110000",
  44800=>"001101000",
  44801=>"101100001",
  44802=>"000011110",
  44803=>"010010011",
  44804=>"000001001",
  44805=>"111001110",
  44806=>"001111000",
  44807=>"101001111",
  44808=>"011000000",
  44809=>"101110100",
  44810=>"000110101",
  44811=>"000100100",
  44812=>"110010001",
  44813=>"110011110",
  44814=>"111101000",
  44815=>"111100110",
  44816=>"011101100",
  44817=>"010110100",
  44818=>"011101000",
  44819=>"101000101",
  44820=>"101001001",
  44821=>"110000110",
  44822=>"101111000",
  44823=>"111000001",
  44824=>"001101001",
  44825=>"000111001",
  44826=>"001100011",
  44827=>"101111111",
  44828=>"010110001",
  44829=>"110111010",
  44830=>"010011110",
  44831=>"001000010",
  44832=>"000000010",
  44833=>"011101110",
  44834=>"101111111",
  44835=>"011001000",
  44836=>"111101111",
  44837=>"000001001",
  44838=>"011010011",
  44839=>"010000111",
  44840=>"010011100",
  44841=>"110100011",
  44842=>"100011111",
  44843=>"011111100",
  44844=>"111110000",
  44845=>"001001011",
  44846=>"001011000",
  44847=>"010100010",
  44848=>"010111100",
  44849=>"111111100",
  44850=>"000110111",
  44851=>"000111010",
  44852=>"101100100",
  44853=>"001000111",
  44854=>"011100110",
  44855=>"110011011",
  44856=>"000110101",
  44857=>"000001010",
  44858=>"111000010",
  44859=>"110011110",
  44860=>"100000101",
  44861=>"100100001",
  44862=>"101101111",
  44863=>"000101111",
  44864=>"000111001",
  44865=>"110011111",
  44866=>"000110111",
  44867=>"100100000",
  44868=>"101111000",
  44869=>"101000011",
  44870=>"111001100",
  44871=>"000001001",
  44872=>"001001010",
  44873=>"100011100",
  44874=>"110101010",
  44875=>"111010100",
  44876=>"100110110",
  44877=>"110100000",
  44878=>"000001001",
  44879=>"000111100",
  44880=>"100100001",
  44881=>"101010000",
  44882=>"000000000",
  44883=>"110011110",
  44884=>"011101010",
  44885=>"010111010",
  44886=>"100101001",
  44887=>"101001110",
  44888=>"001111010",
  44889=>"111111000",
  44890=>"000100001",
  44891=>"000110110",
  44892=>"010011010",
  44893=>"111011011",
  44894=>"010000010",
  44895=>"001101101",
  44896=>"100110000",
  44897=>"111100101",
  44898=>"010011011",
  44899=>"101010110",
  44900=>"110010110",
  44901=>"011011101",
  44902=>"001011001",
  44903=>"011010110",
  44904=>"100011011",
  44905=>"101011011",
  44906=>"011111000",
  44907=>"111010000",
  44908=>"101000011",
  44909=>"101100101",
  44910=>"011011011",
  44911=>"010011000",
  44912=>"100101110",
  44913=>"101110111",
  44914=>"111000000",
  44915=>"000001000",
  44916=>"000111101",
  44917=>"111111111",
  44918=>"001000110",
  44919=>"101000001",
  44920=>"001011110",
  44921=>"000010111",
  44922=>"010101101",
  44923=>"010100000",
  44924=>"000111110",
  44925=>"110000101",
  44926=>"001011111",
  44927=>"100011010",
  44928=>"100001110",
  44929=>"110001001",
  44930=>"010011111",
  44931=>"111010101",
  44932=>"010110100",
  44933=>"101001000",
  44934=>"000100000",
  44935=>"010100010",
  44936=>"000101100",
  44937=>"101001011",
  44938=>"100110011",
  44939=>"110011111",
  44940=>"011001011",
  44941=>"001111011",
  44942=>"101110000",
  44943=>"101100011",
  44944=>"010101111",
  44945=>"101001000",
  44946=>"001001010",
  44947=>"101101001",
  44948=>"011101010",
  44949=>"011100010",
  44950=>"010010111",
  44951=>"111101011",
  44952=>"001110101",
  44953=>"100100010",
  44954=>"111001011",
  44955=>"000111000",
  44956=>"101111010",
  44957=>"010101000",
  44958=>"010110001",
  44959=>"011111110",
  44960=>"100111010",
  44961=>"110100111",
  44962=>"011011110",
  44963=>"000111110",
  44964=>"001001101",
  44965=>"100100011",
  44966=>"111111000",
  44967=>"111000001",
  44968=>"000100111",
  44969=>"101111011",
  44970=>"011111110",
  44971=>"111110110",
  44972=>"010000000",
  44973=>"100010010",
  44974=>"101000101",
  44975=>"100001000",
  44976=>"100111000",
  44977=>"000001101",
  44978=>"010110110",
  44979=>"101011111",
  44980=>"011011001",
  44981=>"110100111",
  44982=>"011001110",
  44983=>"100101111",
  44984=>"011011111",
  44985=>"111111011",
  44986=>"111011001",
  44987=>"111110010",
  44988=>"011000111",
  44989=>"010000101",
  44990=>"010010111",
  44991=>"011110100",
  44992=>"101111110",
  44993=>"011111000",
  44994=>"001110100",
  44995=>"101001000",
  44996=>"100101100",
  44997=>"001010011",
  44998=>"100000110",
  44999=>"111110111",
  45000=>"001101100",
  45001=>"000011011",
  45002=>"010000111",
  45003=>"010111111",
  45004=>"010010010",
  45005=>"110100101",
  45006=>"100110100",
  45007=>"111111101",
  45008=>"100100100",
  45009=>"101000111",
  45010=>"111000010",
  45011=>"110011011",
  45012=>"011101011",
  45013=>"100001110",
  45014=>"011000000",
  45015=>"111100010",
  45016=>"001110010",
  45017=>"011011101",
  45018=>"110100010",
  45019=>"111100011",
  45020=>"111010110",
  45021=>"110000101",
  45022=>"110100110",
  45023=>"100001001",
  45024=>"101110010",
  45025=>"001000101",
  45026=>"100011011",
  45027=>"001100111",
  45028=>"000011000",
  45029=>"110010110",
  45030=>"000001001",
  45031=>"010111010",
  45032=>"000000101",
  45033=>"011101110",
  45034=>"010100000",
  45035=>"101011100",
  45036=>"000000010",
  45037=>"110010111",
  45038=>"011010101",
  45039=>"101101010",
  45040=>"011111001",
  45041=>"000010110",
  45042=>"010000001",
  45043=>"100100100",
  45044=>"110010111",
  45045=>"111100011",
  45046=>"011001110",
  45047=>"000011101",
  45048=>"111111001",
  45049=>"100011110",
  45050=>"111110100",
  45051=>"100011000",
  45052=>"011001001",
  45053=>"001000010",
  45054=>"000000010",
  45055=>"011010111",
  45056=>"100101011",
  45057=>"110111110",
  45058=>"001101010",
  45059=>"101001000",
  45060=>"101110111",
  45061=>"101111101",
  45062=>"001010110",
  45063=>"101101011",
  45064=>"010001010",
  45065=>"100100000",
  45066=>"000100001",
  45067=>"000011100",
  45068=>"000100111",
  45069=>"000001001",
  45070=>"111010000",
  45071=>"010001011",
  45072=>"100010001",
  45073=>"000101101",
  45074=>"111110000",
  45075=>"110111110",
  45076=>"000011011",
  45077=>"000101001",
  45078=>"101001010",
  45079=>"110011000",
  45080=>"011110000",
  45081=>"110001011",
  45082=>"100111111",
  45083=>"001100101",
  45084=>"101100101",
  45085=>"010010010",
  45086=>"000110001",
  45087=>"011011101",
  45088=>"000110011",
  45089=>"000100111",
  45090=>"100000001",
  45091=>"100100000",
  45092=>"001011001",
  45093=>"111011100",
  45094=>"001111010",
  45095=>"101111110",
  45096=>"010100010",
  45097=>"100000100",
  45098=>"000100111",
  45099=>"011101111",
  45100=>"100011010",
  45101=>"101101110",
  45102=>"011000100",
  45103=>"001000100",
  45104=>"111111100",
  45105=>"000000000",
  45106=>"101010011",
  45107=>"110101100",
  45108=>"110001111",
  45109=>"000000100",
  45110=>"000111111",
  45111=>"000110110",
  45112=>"001001101",
  45113=>"000000100",
  45114=>"010001110",
  45115=>"010101011",
  45116=>"100001110",
  45117=>"000001100",
  45118=>"011101101",
  45119=>"000010011",
  45120=>"000000010",
  45121=>"001000011",
  45122=>"111110100",
  45123=>"011111110",
  45124=>"001100101",
  45125=>"000101011",
  45126=>"011110011",
  45127=>"101011100",
  45128=>"000111110",
  45129=>"101010000",
  45130=>"001000001",
  45131=>"100000011",
  45132=>"011100111",
  45133=>"010101010",
  45134=>"110011110",
  45135=>"000111111",
  45136=>"100110001",
  45137=>"100111000",
  45138=>"010011011",
  45139=>"010111010",
  45140=>"010001100",
  45141=>"101001111",
  45142=>"000101000",
  45143=>"001010111",
  45144=>"001101110",
  45145=>"001111100",
  45146=>"110011000",
  45147=>"010000101",
  45148=>"110010011",
  45149=>"000001111",
  45150=>"011001011",
  45151=>"101000100",
  45152=>"101100110",
  45153=>"110000001",
  45154=>"100110101",
  45155=>"011010000",
  45156=>"000101111",
  45157=>"110010000",
  45158=>"110000000",
  45159=>"111010000",
  45160=>"001000001",
  45161=>"110110010",
  45162=>"100111010",
  45163=>"100110011",
  45164=>"110100000",
  45165=>"011101100",
  45166=>"010100010",
  45167=>"001101010",
  45168=>"010000101",
  45169=>"001110011",
  45170=>"000111111",
  45171=>"101101011",
  45172=>"100010011",
  45173=>"110001001",
  45174=>"010101001",
  45175=>"010001011",
  45176=>"000011000",
  45177=>"010100101",
  45178=>"000011110",
  45179=>"111000101",
  45180=>"000110011",
  45181=>"001010011",
  45182=>"101101111",
  45183=>"111100000",
  45184=>"000110010",
  45185=>"011110111",
  45186=>"001001110",
  45187=>"001111100",
  45188=>"010000001",
  45189=>"101011010",
  45190=>"110000111",
  45191=>"000010001",
  45192=>"000010101",
  45193=>"100110100",
  45194=>"100111011",
  45195=>"001010010",
  45196=>"010000110",
  45197=>"010111110",
  45198=>"110100101",
  45199=>"101110111",
  45200=>"011010111",
  45201=>"011100110",
  45202=>"000001110",
  45203=>"010001101",
  45204=>"000011000",
  45205=>"100101001",
  45206=>"101001001",
  45207=>"001100001",
  45208=>"110100001",
  45209=>"110011111",
  45210=>"000101001",
  45211=>"100001101",
  45212=>"001010011",
  45213=>"101111001",
  45214=>"111100110",
  45215=>"110010011",
  45216=>"001000001",
  45217=>"100101110",
  45218=>"111000000",
  45219=>"010001001",
  45220=>"001000100",
  45221=>"010111110",
  45222=>"101000100",
  45223=>"001110110",
  45224=>"000000001",
  45225=>"000011110",
  45226=>"000100001",
  45227=>"001100011",
  45228=>"001010110",
  45229=>"010010111",
  45230=>"110100110",
  45231=>"110001100",
  45232=>"110000001",
  45233=>"100010010",
  45234=>"100000100",
  45235=>"000001100",
  45236=>"010110000",
  45237=>"010011001",
  45238=>"110100000",
  45239=>"001001101",
  45240=>"001101100",
  45241=>"100010110",
  45242=>"111001100",
  45243=>"110001111",
  45244=>"111111001",
  45245=>"011001111",
  45246=>"111101001",
  45247=>"100011010",
  45248=>"011000111",
  45249=>"000101001",
  45250=>"000100010",
  45251=>"000111011",
  45252=>"100001010",
  45253=>"000111111",
  45254=>"011111110",
  45255=>"011111000",
  45256=>"110011110",
  45257=>"001111110",
  45258=>"001011111",
  45259=>"100110111",
  45260=>"000001110",
  45261=>"001100011",
  45262=>"011101011",
  45263=>"000100010",
  45264=>"100001100",
  45265=>"010001111",
  45266=>"100001000",
  45267=>"000101100",
  45268=>"101000000",
  45269=>"100110111",
  45270=>"110001000",
  45271=>"010011010",
  45272=>"011101000",
  45273=>"100110001",
  45274=>"111001000",
  45275=>"010011010",
  45276=>"001101111",
  45277=>"011111001",
  45278=>"010011001",
  45279=>"011110000",
  45280=>"110110100",
  45281=>"010001000",
  45282=>"001000101",
  45283=>"111001011",
  45284=>"011011001",
  45285=>"100010101",
  45286=>"001000101",
  45287=>"101110110",
  45288=>"100111101",
  45289=>"011111101",
  45290=>"010100101",
  45291=>"111111000",
  45292=>"101111100",
  45293=>"101000000",
  45294=>"110100111",
  45295=>"010111000",
  45296=>"010101010",
  45297=>"001110111",
  45298=>"000001000",
  45299=>"011011100",
  45300=>"101111001",
  45301=>"000111100",
  45302=>"110011011",
  45303=>"101000100",
  45304=>"111100011",
  45305=>"111000010",
  45306=>"011111001",
  45307=>"111110101",
  45308=>"110110011",
  45309=>"110100110",
  45310=>"110000001",
  45311=>"110010101",
  45312=>"100001101",
  45313=>"001010011",
  45314=>"110110111",
  45315=>"001000111",
  45316=>"011011101",
  45317=>"010100111",
  45318=>"111010011",
  45319=>"110000001",
  45320=>"000100011",
  45321=>"000010100",
  45322=>"000101001",
  45323=>"001011001",
  45324=>"011100001",
  45325=>"000111101",
  45326=>"110001111",
  45327=>"100101101",
  45328=>"110101110",
  45329=>"111111110",
  45330=>"111010011",
  45331=>"001011011",
  45332=>"001100011",
  45333=>"001000100",
  45334=>"001110110",
  45335=>"101000110",
  45336=>"100100001",
  45337=>"101000001",
  45338=>"000111001",
  45339=>"011111101",
  45340=>"000100001",
  45341=>"110111010",
  45342=>"010000101",
  45343=>"110001000",
  45344=>"101100100",
  45345=>"001001100",
  45346=>"100110101",
  45347=>"001110010",
  45348=>"110011000",
  45349=>"101110000",
  45350=>"011101000",
  45351=>"110011111",
  45352=>"110110110",
  45353=>"100100001",
  45354=>"111000011",
  45355=>"100000110",
  45356=>"110110001",
  45357=>"010001110",
  45358=>"110000000",
  45359=>"010110101",
  45360=>"100110100",
  45361=>"110011000",
  45362=>"111010101",
  45363=>"101100110",
  45364=>"110100100",
  45365=>"011100011",
  45366=>"100001011",
  45367=>"011100001",
  45368=>"010001100",
  45369=>"111100001",
  45370=>"110100011",
  45371=>"111011101",
  45372=>"000111111",
  45373=>"110100110",
  45374=>"011100111",
  45375=>"001111101",
  45376=>"001000000",
  45377=>"000000101",
  45378=>"110011110",
  45379=>"111101010",
  45380=>"111110101",
  45381=>"100011111",
  45382=>"011100001",
  45383=>"010000000",
  45384=>"110010000",
  45385=>"001000101",
  45386=>"010001000",
  45387=>"110000010",
  45388=>"100111110",
  45389=>"110100100",
  45390=>"011110011",
  45391=>"010010010",
  45392=>"100101010",
  45393=>"101110010",
  45394=>"111001111",
  45395=>"011010000",
  45396=>"011100010",
  45397=>"011010011",
  45398=>"110010000",
  45399=>"001111001",
  45400=>"101111100",
  45401=>"000101001",
  45402=>"001110001",
  45403=>"011000101",
  45404=>"010110000",
  45405=>"001100000",
  45406=>"111110110",
  45407=>"110100101",
  45408=>"000111100",
  45409=>"110011011",
  45410=>"101101011",
  45411=>"010001111",
  45412=>"010101101",
  45413=>"100010001",
  45414=>"000010110",
  45415=>"111111101",
  45416=>"010111111",
  45417=>"011100000",
  45418=>"110101010",
  45419=>"010000111",
  45420=>"011101100",
  45421=>"000111010",
  45422=>"101000111",
  45423=>"101010111",
  45424=>"001000001",
  45425=>"011001000",
  45426=>"011100011",
  45427=>"110110000",
  45428=>"011000110",
  45429=>"111101111",
  45430=>"101010110",
  45431=>"100110110",
  45432=>"100001101",
  45433=>"111100010",
  45434=>"100000101",
  45435=>"011100100",
  45436=>"000110100",
  45437=>"000010000",
  45438=>"000000110",
  45439=>"001010111",
  45440=>"100011010",
  45441=>"101011100",
  45442=>"101000101",
  45443=>"100110110",
  45444=>"101010111",
  45445=>"001101000",
  45446=>"111011010",
  45447=>"110100101",
  45448=>"101010000",
  45449=>"010000000",
  45450=>"111011011",
  45451=>"000000100",
  45452=>"010100011",
  45453=>"100000101",
  45454=>"000010011",
  45455=>"010101011",
  45456=>"110001000",
  45457=>"000111101",
  45458=>"100110110",
  45459=>"111101001",
  45460=>"000011110",
  45461=>"100001111",
  45462=>"111010001",
  45463=>"110111000",
  45464=>"111000110",
  45465=>"000000111",
  45466=>"010111001",
  45467=>"111001100",
  45468=>"001000110",
  45469=>"101111010",
  45470=>"111000011",
  45471=>"010000000",
  45472=>"100100100",
  45473=>"001101000",
  45474=>"011100110",
  45475=>"101010101",
  45476=>"101110110",
  45477=>"001100101",
  45478=>"011111111",
  45479=>"101101011",
  45480=>"100111111",
  45481=>"001001000",
  45482=>"111010000",
  45483=>"011000001",
  45484=>"100110011",
  45485=>"010010001",
  45486=>"010100101",
  45487=>"000100001",
  45488=>"101001101",
  45489=>"110101010",
  45490=>"010111101",
  45491=>"010000111",
  45492=>"101100100",
  45493=>"000100101",
  45494=>"101000101",
  45495=>"001111100",
  45496=>"010100011",
  45497=>"011000111",
  45498=>"101010100",
  45499=>"110010011",
  45500=>"110010001",
  45501=>"000111101",
  45502=>"011011110",
  45503=>"101110100",
  45504=>"001101001",
  45505=>"001111110",
  45506=>"010110101",
  45507=>"011010011",
  45508=>"010101010",
  45509=>"100000001",
  45510=>"011011001",
  45511=>"000100000",
  45512=>"000100101",
  45513=>"101111110",
  45514=>"010010111",
  45515=>"101000010",
  45516=>"111111101",
  45517=>"010000100",
  45518=>"010000111",
  45519=>"111010101",
  45520=>"100010110",
  45521=>"110010010",
  45522=>"010010111",
  45523=>"010111010",
  45524=>"001000110",
  45525=>"110001000",
  45526=>"100001100",
  45527=>"000001000",
  45528=>"111010011",
  45529=>"100010011",
  45530=>"010001101",
  45531=>"010100000",
  45532=>"110010010",
  45533=>"100001111",
  45534=>"000110101",
  45535=>"001101010",
  45536=>"100110111",
  45537=>"001011110",
  45538=>"010110100",
  45539=>"000100110",
  45540=>"110001010",
  45541=>"111011110",
  45542=>"100001011",
  45543=>"101100111",
  45544=>"010111010",
  45545=>"111111010",
  45546=>"001010000",
  45547=>"000011100",
  45548=>"110111111",
  45549=>"110100110",
  45550=>"100011000",
  45551=>"010000101",
  45552=>"100010111",
  45553=>"111100011",
  45554=>"100101010",
  45555=>"000011101",
  45556=>"010111100",
  45557=>"010100111",
  45558=>"111111011",
  45559=>"100111100",
  45560=>"111001110",
  45561=>"111100011",
  45562=>"000001010",
  45563=>"011110111",
  45564=>"000001100",
  45565=>"111010101",
  45566=>"110101011",
  45567=>"110011010",
  45568=>"010001000",
  45569=>"101011011",
  45570=>"011100000",
  45571=>"110101001",
  45572=>"100110111",
  45573=>"010010100",
  45574=>"001000101",
  45575=>"010010001",
  45576=>"010010100",
  45577=>"101100111",
  45578=>"101000111",
  45579=>"110001011",
  45580=>"001101000",
  45581=>"111010111",
  45582=>"000000010",
  45583=>"110100011",
  45584=>"001011010",
  45585=>"010011011",
  45586=>"100001011",
  45587=>"010100100",
  45588=>"001010011",
  45589=>"111101101",
  45590=>"000010100",
  45591=>"001010111",
  45592=>"000100111",
  45593=>"110101001",
  45594=>"100001010",
  45595=>"011110011",
  45596=>"101000110",
  45597=>"001010101",
  45598=>"010011011",
  45599=>"000011111",
  45600=>"000010010",
  45601=>"101000010",
  45602=>"111101010",
  45603=>"000001111",
  45604=>"000001000",
  45605=>"110001100",
  45606=>"001110010",
  45607=>"101001111",
  45608=>"100001100",
  45609=>"001111011",
  45610=>"111100011",
  45611=>"111011011",
  45612=>"000111011",
  45613=>"000111111",
  45614=>"010010101",
  45615=>"001010110",
  45616=>"111011111",
  45617=>"000111010",
  45618=>"000000000",
  45619=>"001010000",
  45620=>"000110110",
  45621=>"101010100",
  45622=>"000010100",
  45623=>"000100010",
  45624=>"011010011",
  45625=>"111100101",
  45626=>"001110000",
  45627=>"000010001",
  45628=>"010110100",
  45629=>"010111100",
  45630=>"111010111",
  45631=>"100001101",
  45632=>"111010111",
  45633=>"001000000",
  45634=>"000110110",
  45635=>"100000100",
  45636=>"011100100",
  45637=>"011110111",
  45638=>"100001001",
  45639=>"100111010",
  45640=>"111000100",
  45641=>"111110001",
  45642=>"011111001",
  45643=>"011001101",
  45644=>"001001001",
  45645=>"101101100",
  45646=>"100100001",
  45647=>"100101110",
  45648=>"110011110",
  45649=>"010101010",
  45650=>"001010100",
  45651=>"100100001",
  45652=>"001010001",
  45653=>"001101111",
  45654=>"010000001",
  45655=>"010011110",
  45656=>"011111111",
  45657=>"101010111",
  45658=>"101001100",
  45659=>"000101010",
  45660=>"010001110",
  45661=>"000100100",
  45662=>"000110100",
  45663=>"010111010",
  45664=>"101100000",
  45665=>"010100111",
  45666=>"101000000",
  45667=>"001000001",
  45668=>"100011000",
  45669=>"001001010",
  45670=>"111100111",
  45671=>"101010001",
  45672=>"000110001",
  45673=>"000101000",
  45674=>"001111101",
  45675=>"111101111",
  45676=>"100101100",
  45677=>"010011001",
  45678=>"101110001",
  45679=>"010010000",
  45680=>"101010001",
  45681=>"000101010",
  45682=>"111011011",
  45683=>"101001100",
  45684=>"110111001",
  45685=>"010101001",
  45686=>"101010110",
  45687=>"100000101",
  45688=>"000111101",
  45689=>"111100000",
  45690=>"000001101",
  45691=>"111110111",
  45692=>"000001011",
  45693=>"000000111",
  45694=>"011011010",
  45695=>"000111111",
  45696=>"101001100",
  45697=>"010110100",
  45698=>"000001000",
  45699=>"000011100",
  45700=>"100001101",
  45701=>"111110001",
  45702=>"011111011",
  45703=>"111000000",
  45704=>"011011000",
  45705=>"011111100",
  45706=>"010111110",
  45707=>"101011010",
  45708=>"101010100",
  45709=>"011100101",
  45710=>"111111101",
  45711=>"001111101",
  45712=>"001001101",
  45713=>"011011001",
  45714=>"101111001",
  45715=>"111011000",
  45716=>"011100100",
  45717=>"001001100",
  45718=>"100000011",
  45719=>"011111011",
  45720=>"110101000",
  45721=>"010000011",
  45722=>"110010001",
  45723=>"101100011",
  45724=>"001001100",
  45725=>"011101101",
  45726=>"111110000",
  45727=>"110010000",
  45728=>"110010110",
  45729=>"101100101",
  45730=>"010011101",
  45731=>"001001110",
  45732=>"101110011",
  45733=>"111011000",
  45734=>"111000110",
  45735=>"001100111",
  45736=>"000000010",
  45737=>"101010101",
  45738=>"110001111",
  45739=>"111100000",
  45740=>"011000001",
  45741=>"011011010",
  45742=>"010100100",
  45743=>"101010101",
  45744=>"101111111",
  45745=>"100101100",
  45746=>"001011001",
  45747=>"011010010",
  45748=>"001100101",
  45749=>"100010110",
  45750=>"110000000",
  45751=>"101100101",
  45752=>"101111110",
  45753=>"110001001",
  45754=>"011100111",
  45755=>"111110101",
  45756=>"111111111",
  45757=>"110001001",
  45758=>"001001000",
  45759=>"010000100",
  45760=>"001011000",
  45761=>"100111110",
  45762=>"000000100",
  45763=>"001011010",
  45764=>"100001000",
  45765=>"010010100",
  45766=>"101101011",
  45767=>"111011010",
  45768=>"000001011",
  45769=>"011100000",
  45770=>"111011110",
  45771=>"101100011",
  45772=>"100110110",
  45773=>"101010111",
  45774=>"011000001",
  45775=>"000001000",
  45776=>"011111110",
  45777=>"000111100",
  45778=>"111000101",
  45779=>"010000001",
  45780=>"010111011",
  45781=>"000101011",
  45782=>"110111101",
  45783=>"111111110",
  45784=>"110011101",
  45785=>"011001011",
  45786=>"011100110",
  45787=>"010101111",
  45788=>"000001100",
  45789=>"101010000",
  45790=>"101100100",
  45791=>"110101010",
  45792=>"101110101",
  45793=>"000110011",
  45794=>"011110111",
  45795=>"110100100",
  45796=>"100111101",
  45797=>"111100010",
  45798=>"111000011",
  45799=>"100001110",
  45800=>"011010111",
  45801=>"000111111",
  45802=>"011100011",
  45803=>"100110111",
  45804=>"011001110",
  45805=>"100101101",
  45806=>"001101000",
  45807=>"110011011",
  45808=>"101000000",
  45809=>"111100000",
  45810=>"011101010",
  45811=>"100101100",
  45812=>"110110111",
  45813=>"100000100",
  45814=>"000000010",
  45815=>"001000100",
  45816=>"011111010",
  45817=>"011001101",
  45818=>"010011001",
  45819=>"101101010",
  45820=>"111100010",
  45821=>"101100110",
  45822=>"110110001",
  45823=>"000010110",
  45824=>"001100010",
  45825=>"000011101",
  45826=>"111000100",
  45827=>"101000110",
  45828=>"011001001",
  45829=>"000010000",
  45830=>"000001000",
  45831=>"000000110",
  45832=>"101011011",
  45833=>"111100001",
  45834=>"101110101",
  45835=>"110001101",
  45836=>"101010011",
  45837=>"011101100",
  45838=>"110110111",
  45839=>"111110000",
  45840=>"001000001",
  45841=>"010010100",
  45842=>"100000011",
  45843=>"011100101",
  45844=>"101011101",
  45845=>"010111101",
  45846=>"000000010",
  45847=>"001100001",
  45848=>"010100111",
  45849=>"011000101",
  45850=>"000010001",
  45851=>"011001010",
  45852=>"011001011",
  45853=>"100101010",
  45854=>"100100000",
  45855=>"010010010",
  45856=>"100111000",
  45857=>"111000000",
  45858=>"111010010",
  45859=>"110010010",
  45860=>"111111111",
  45861=>"101010101",
  45862=>"011001000",
  45863=>"000101100",
  45864=>"010110010",
  45865=>"011111110",
  45866=>"010001011",
  45867=>"011111111",
  45868=>"110011110",
  45869=>"010010110",
  45870=>"100011000",
  45871=>"111110010",
  45872=>"000111101",
  45873=>"000001110",
  45874=>"000000001",
  45875=>"111010111",
  45876=>"100010100",
  45877=>"010111011",
  45878=>"011110100",
  45879=>"111110101",
  45880=>"011100100",
  45881=>"101000101",
  45882=>"001011111",
  45883=>"111110010",
  45884=>"110101010",
  45885=>"110110100",
  45886=>"100001111",
  45887=>"011010101",
  45888=>"010010101",
  45889=>"000111111",
  45890=>"101010111",
  45891=>"100000111",
  45892=>"100100101",
  45893=>"110001110",
  45894=>"000101010",
  45895=>"011100111",
  45896=>"011101011",
  45897=>"110011010",
  45898=>"011110000",
  45899=>"111010001",
  45900=>"100101101",
  45901=>"100111001",
  45902=>"010001110",
  45903=>"111010100",
  45904=>"110101111",
  45905=>"001111000",
  45906=>"010110101",
  45907=>"010000111",
  45908=>"101000101",
  45909=>"111101100",
  45910=>"110010001",
  45911=>"100010011",
  45912=>"010001011",
  45913=>"111001111",
  45914=>"110000010",
  45915=>"111101101",
  45916=>"111101011",
  45917=>"001011010",
  45918=>"101001010",
  45919=>"000100011",
  45920=>"101110011",
  45921=>"001001100",
  45922=>"100111000",
  45923=>"011110101",
  45924=>"011010000",
  45925=>"100011011",
  45926=>"010001110",
  45927=>"001111001",
  45928=>"101101001",
  45929=>"010101001",
  45930=>"100001001",
  45931=>"010101001",
  45932=>"000111101",
  45933=>"000000101",
  45934=>"111110101",
  45935=>"010001111",
  45936=>"010011000",
  45937=>"000010111",
  45938=>"000000110",
  45939=>"100011111",
  45940=>"010000101",
  45941=>"001110001",
  45942=>"110001111",
  45943=>"100001011",
  45944=>"111011111",
  45945=>"001000101",
  45946=>"101111010",
  45947=>"101111101",
  45948=>"000001101",
  45949=>"110000101",
  45950=>"101101111",
  45951=>"101011100",
  45952=>"010000001",
  45953=>"000000100",
  45954=>"110001011",
  45955=>"101110011",
  45956=>"111000101",
  45957=>"111001110",
  45958=>"011010111",
  45959=>"001110100",
  45960=>"111111011",
  45961=>"101011010",
  45962=>"010010100",
  45963=>"010011000",
  45964=>"010001101",
  45965=>"001110000",
  45966=>"011110100",
  45967=>"100010010",
  45968=>"001110100",
  45969=>"000010100",
  45970=>"000010111",
  45971=>"100000001",
  45972=>"010011001",
  45973=>"110000000",
  45974=>"001000010",
  45975=>"110100010",
  45976=>"100110100",
  45977=>"001011010",
  45978=>"001010101",
  45979=>"000001100",
  45980=>"111011111",
  45981=>"100100010",
  45982=>"111001101",
  45983=>"101101111",
  45984=>"101001100",
  45985=>"011111101",
  45986=>"110101101",
  45987=>"000010101",
  45988=>"010001011",
  45989=>"001001110",
  45990=>"100100110",
  45991=>"101010001",
  45992=>"010011111",
  45993=>"101100011",
  45994=>"110001111",
  45995=>"111001100",
  45996=>"000001011",
  45997=>"101100101",
  45998=>"010010000",
  45999=>"101010010",
  46000=>"110100001",
  46001=>"111001100",
  46002=>"100011010",
  46003=>"000011001",
  46004=>"111011111",
  46005=>"001101001",
  46006=>"100000010",
  46007=>"100111110",
  46008=>"000111001",
  46009=>"001100111",
  46010=>"110010011",
  46011=>"001100100",
  46012=>"001010011",
  46013=>"000100010",
  46014=>"011001110",
  46015=>"010001010",
  46016=>"010100001",
  46017=>"000000000",
  46018=>"000011000",
  46019=>"111011110",
  46020=>"110000001",
  46021=>"001100110",
  46022=>"110011001",
  46023=>"110000011",
  46024=>"111100001",
  46025=>"000110001",
  46026=>"000101000",
  46027=>"000001000",
  46028=>"010100110",
  46029=>"100100110",
  46030=>"000110011",
  46031=>"111100111",
  46032=>"110101001",
  46033=>"001011000",
  46034=>"000110110",
  46035=>"010010111",
  46036=>"000110000",
  46037=>"000111111",
  46038=>"010001100",
  46039=>"001110010",
  46040=>"110101110",
  46041=>"101100010",
  46042=>"111000000",
  46043=>"001110110",
  46044=>"100001111",
  46045=>"001010101",
  46046=>"001001101",
  46047=>"000110110",
  46048=>"011000001",
  46049=>"100000011",
  46050=>"001011000",
  46051=>"000011010",
  46052=>"110110101",
  46053=>"101100100",
  46054=>"011101110",
  46055=>"100110101",
  46056=>"011011000",
  46057=>"111110001",
  46058=>"001100101",
  46059=>"100100011",
  46060=>"000011111",
  46061=>"010000011",
  46062=>"011011001",
  46063=>"101101111",
  46064=>"000100000",
  46065=>"110011110",
  46066=>"100111000",
  46067=>"001101001",
  46068=>"110011000",
  46069=>"000011100",
  46070=>"110110110",
  46071=>"001110100",
  46072=>"000110000",
  46073=>"000110110",
  46074=>"100000000",
  46075=>"111110101",
  46076=>"010011100",
  46077=>"111010000",
  46078=>"100110001",
  46079=>"000001010",
  46080=>"101011001",
  46081=>"101101011",
  46082=>"100110111",
  46083=>"011111010",
  46084=>"110001111",
  46085=>"111010001",
  46086=>"111100011",
  46087=>"101010011",
  46088=>"010000001",
  46089=>"110010010",
  46090=>"010011110",
  46091=>"000001010",
  46092=>"110100111",
  46093=>"010110011",
  46094=>"000111110",
  46095=>"100111000",
  46096=>"101011100",
  46097=>"110101011",
  46098=>"010000100",
  46099=>"111100100",
  46100=>"101100010",
  46101=>"110110101",
  46102=>"001110111",
  46103=>"001010110",
  46104=>"001101000",
  46105=>"001101001",
  46106=>"100101010",
  46107=>"111111011",
  46108=>"111010101",
  46109=>"110010101",
  46110=>"010101000",
  46111=>"100001000",
  46112=>"011011000",
  46113=>"101110111",
  46114=>"111010011",
  46115=>"100010000",
  46116=>"100001111",
  46117=>"000111110",
  46118=>"011110100",
  46119=>"000001000",
  46120=>"101010011",
  46121=>"111111000",
  46122=>"001000110",
  46123=>"011110001",
  46124=>"000011100",
  46125=>"101001010",
  46126=>"001110100",
  46127=>"100011011",
  46128=>"110000110",
  46129=>"111101110",
  46130=>"011001010",
  46131=>"110011010",
  46132=>"111111000",
  46133=>"000100110",
  46134=>"100010001",
  46135=>"011101000",
  46136=>"111110011",
  46137=>"001101101",
  46138=>"011101010",
  46139=>"000101110",
  46140=>"100111001",
  46141=>"101000000",
  46142=>"000000010",
  46143=>"101000110",
  46144=>"011110101",
  46145=>"010000101",
  46146=>"010011001",
  46147=>"010110110",
  46148=>"111111101",
  46149=>"000100000",
  46150=>"100010100",
  46151=>"110111100",
  46152=>"001101001",
  46153=>"100111011",
  46154=>"110100101",
  46155=>"011110011",
  46156=>"000010010",
  46157=>"000110111",
  46158=>"111111111",
  46159=>"000111011",
  46160=>"000101111",
  46161=>"010001001",
  46162=>"111001000",
  46163=>"100010111",
  46164=>"010001100",
  46165=>"101011111",
  46166=>"100001111",
  46167=>"110111101",
  46168=>"101110101",
  46169=>"001010000",
  46170=>"111100010",
  46171=>"000101110",
  46172=>"001111111",
  46173=>"010101000",
  46174=>"111010110",
  46175=>"000101000",
  46176=>"001001000",
  46177=>"110101100",
  46178=>"111000101",
  46179=>"011000000",
  46180=>"100000100",
  46181=>"001101100",
  46182=>"010111101",
  46183=>"111110011",
  46184=>"100110110",
  46185=>"011110100",
  46186=>"011000001",
  46187=>"011001101",
  46188=>"110101010",
  46189=>"001111010",
  46190=>"010000010",
  46191=>"101001101",
  46192=>"111011101",
  46193=>"100100100",
  46194=>"001101011",
  46195=>"101101000",
  46196=>"100011010",
  46197=>"010010100",
  46198=>"111110000",
  46199=>"101010100",
  46200=>"001000010",
  46201=>"101110111",
  46202=>"001101001",
  46203=>"110111101",
  46204=>"000010111",
  46205=>"101100010",
  46206=>"111001011",
  46207=>"100001111",
  46208=>"000100110",
  46209=>"110000101",
  46210=>"000100011",
  46211=>"010111110",
  46212=>"000000100",
  46213=>"001100000",
  46214=>"010001000",
  46215=>"000101011",
  46216=>"100101011",
  46217=>"100100001",
  46218=>"111001100",
  46219=>"011001111",
  46220=>"111111010",
  46221=>"010110110",
  46222=>"001000101",
  46223=>"110110111",
  46224=>"011001101",
  46225=>"101001100",
  46226=>"011101110",
  46227=>"010011100",
  46228=>"010101011",
  46229=>"111101010",
  46230=>"010101100",
  46231=>"010100111",
  46232=>"111111101",
  46233=>"100100110",
  46234=>"000110000",
  46235=>"000001110",
  46236=>"110000100",
  46237=>"110001111",
  46238=>"111001100",
  46239=>"001011111",
  46240=>"000000000",
  46241=>"110011000",
  46242=>"010110000",
  46243=>"110111010",
  46244=>"001011100",
  46245=>"001110100",
  46246=>"101110001",
  46247=>"001011011",
  46248=>"101010101",
  46249=>"010100010",
  46250=>"111110101",
  46251=>"001001101",
  46252=>"001111000",
  46253=>"110100101",
  46254=>"110100101",
  46255=>"001101000",
  46256=>"001010111",
  46257=>"101100110",
  46258=>"000111111",
  46259=>"000110110",
  46260=>"101001000",
  46261=>"110001100",
  46262=>"010001000",
  46263=>"110111010",
  46264=>"000110101",
  46265=>"111001001",
  46266=>"000110111",
  46267=>"111001110",
  46268=>"111101001",
  46269=>"110110010",
  46270=>"001100001",
  46271=>"001110001",
  46272=>"010110110",
  46273=>"011000101",
  46274=>"010010110",
  46275=>"001000100",
  46276=>"111101111",
  46277=>"100001001",
  46278=>"100110011",
  46279=>"101101001",
  46280=>"010011011",
  46281=>"100001110",
  46282=>"000111100",
  46283=>"111110011",
  46284=>"101101100",
  46285=>"101000001",
  46286=>"001000100",
  46287=>"010100010",
  46288=>"011001000",
  46289=>"010100110",
  46290=>"011010110",
  46291=>"111000101",
  46292=>"110111010",
  46293=>"001110000",
  46294=>"011011001",
  46295=>"100011010",
  46296=>"010001001",
  46297=>"101111111",
  46298=>"001101100",
  46299=>"011100011",
  46300=>"111001010",
  46301=>"010111101",
  46302=>"100001000",
  46303=>"101100111",
  46304=>"101000101",
  46305=>"000110110",
  46306=>"101101110",
  46307=>"001101111",
  46308=>"101001010",
  46309=>"111111011",
  46310=>"000011000",
  46311=>"111001111",
  46312=>"011101000",
  46313=>"101110010",
  46314=>"101110001",
  46315=>"110110000",
  46316=>"111010001",
  46317=>"101101001",
  46318=>"001101100",
  46319=>"100000111",
  46320=>"010111101",
  46321=>"101010101",
  46322=>"101100011",
  46323=>"010010011",
  46324=>"101000011",
  46325=>"000110110",
  46326=>"010001000",
  46327=>"111101100",
  46328=>"001110110",
  46329=>"001101101",
  46330=>"100111110",
  46331=>"011011010",
  46332=>"010011111",
  46333=>"110101111",
  46334=>"101110100",
  46335=>"100000000",
  46336=>"001010010",
  46337=>"010001100",
  46338=>"000000100",
  46339=>"011011110",
  46340=>"000001100",
  46341=>"100101111",
  46342=>"001101010",
  46343=>"000110101",
  46344=>"110100101",
  46345=>"110011010",
  46346=>"101010100",
  46347=>"100111101",
  46348=>"011101001",
  46349=>"100101111",
  46350=>"001000011",
  46351=>"010111011",
  46352=>"000011110",
  46353=>"111011011",
  46354=>"001000100",
  46355=>"000110111",
  46356=>"001000010",
  46357=>"001000100",
  46358=>"001011101",
  46359=>"010001000",
  46360=>"011010011",
  46361=>"110110001",
  46362=>"010101000",
  46363=>"100011000",
  46364=>"000110110",
  46365=>"100100110",
  46366=>"101110000",
  46367=>"100001111",
  46368=>"000000100",
  46369=>"111000000",
  46370=>"011111011",
  46371=>"011110011",
  46372=>"010000111",
  46373=>"011000001",
  46374=>"101100000",
  46375=>"001110010",
  46376=>"000100000",
  46377=>"100111111",
  46378=>"011100111",
  46379=>"011000111",
  46380=>"111001100",
  46381=>"110110010",
  46382=>"000010000",
  46383=>"010111101",
  46384=>"010011011",
  46385=>"110100001",
  46386=>"011111111",
  46387=>"001001010",
  46388=>"000010010",
  46389=>"011000100",
  46390=>"111001011",
  46391=>"100011111",
  46392=>"000110111",
  46393=>"011011010",
  46394=>"000110010",
  46395=>"101110101",
  46396=>"000110111",
  46397=>"000001001",
  46398=>"101001010",
  46399=>"001000101",
  46400=>"011111110",
  46401=>"100001101",
  46402=>"000101000",
  46403=>"100000001",
  46404=>"111000100",
  46405=>"000011100",
  46406=>"111010111",
  46407=>"111011010",
  46408=>"000011100",
  46409=>"001101100",
  46410=>"110110011",
  46411=>"001001101",
  46412=>"101010000",
  46413=>"111011001",
  46414=>"011011001",
  46415=>"010101010",
  46416=>"010100010",
  46417=>"110100101",
  46418=>"001011111",
  46419=>"000011111",
  46420=>"000000111",
  46421=>"101110100",
  46422=>"111000010",
  46423=>"010110100",
  46424=>"001010011",
  46425=>"110101100",
  46426=>"111111011",
  46427=>"001011111",
  46428=>"101111101",
  46429=>"110110110",
  46430=>"011000000",
  46431=>"010110000",
  46432=>"000010011",
  46433=>"111111110",
  46434=>"101001100",
  46435=>"111110110",
  46436=>"111100011",
  46437=>"100011111",
  46438=>"000110111",
  46439=>"100101101",
  46440=>"111101001",
  46441=>"000000001",
  46442=>"011010100",
  46443=>"000001110",
  46444=>"000100101",
  46445=>"000000011",
  46446=>"000111011",
  46447=>"000010010",
  46448=>"110001100",
  46449=>"111110111",
  46450=>"010111011",
  46451=>"010110000",
  46452=>"110001100",
  46453=>"100001100",
  46454=>"001011010",
  46455=>"110110011",
  46456=>"010110101",
  46457=>"011000111",
  46458=>"000110011",
  46459=>"011010101",
  46460=>"111011011",
  46461=>"011001000",
  46462=>"101111000",
  46463=>"110110100",
  46464=>"000001110",
  46465=>"001111111",
  46466=>"011111010",
  46467=>"010101110",
  46468=>"101001001",
  46469=>"000000000",
  46470=>"111110011",
  46471=>"100100101",
  46472=>"010010101",
  46473=>"111000000",
  46474=>"101100110",
  46475=>"000111010",
  46476=>"001101100",
  46477=>"011111000",
  46478=>"000101100",
  46479=>"101110100",
  46480=>"001100010",
  46481=>"111001100",
  46482=>"010011010",
  46483=>"101010100",
  46484=>"001011000",
  46485=>"011010001",
  46486=>"000100100",
  46487=>"100001111",
  46488=>"111001101",
  46489=>"101000110",
  46490=>"011001110",
  46491=>"001001001",
  46492=>"111011101",
  46493=>"000100011",
  46494=>"001010110",
  46495=>"011001010",
  46496=>"100000110",
  46497=>"100101000",
  46498=>"110110101",
  46499=>"001110111",
  46500=>"011111000",
  46501=>"111101011",
  46502=>"011011011",
  46503=>"000010001",
  46504=>"111101000",
  46505=>"000110100",
  46506=>"111010111",
  46507=>"000011100",
  46508=>"100011111",
  46509=>"100100100",
  46510=>"000011000",
  46511=>"011010100",
  46512=>"011010011",
  46513=>"100010010",
  46514=>"100110110",
  46515=>"000110011",
  46516=>"111101110",
  46517=>"010100001",
  46518=>"100111100",
  46519=>"001101110",
  46520=>"001001001",
  46521=>"010100001",
  46522=>"101100000",
  46523=>"000000100",
  46524=>"111011110",
  46525=>"110110100",
  46526=>"110011101",
  46527=>"001111111",
  46528=>"010101100",
  46529=>"011011101",
  46530=>"101001010",
  46531=>"101110000",
  46532=>"011010000",
  46533=>"000010101",
  46534=>"101010111",
  46535=>"110110110",
  46536=>"001001101",
  46537=>"001000110",
  46538=>"111101011",
  46539=>"000010111",
  46540=>"110011010",
  46541=>"111110110",
  46542=>"011100001",
  46543=>"001100100",
  46544=>"110101011",
  46545=>"010110110",
  46546=>"110001011",
  46547=>"010101100",
  46548=>"110101111",
  46549=>"011001111",
  46550=>"110100011",
  46551=>"111010010",
  46552=>"110011110",
  46553=>"001111001",
  46554=>"001001101",
  46555=>"000101101",
  46556=>"101100101",
  46557=>"000110101",
  46558=>"011100010",
  46559=>"100001000",
  46560=>"011011011",
  46561=>"001101001",
  46562=>"101100011",
  46563=>"111111011",
  46564=>"010001001",
  46565=>"011001110",
  46566=>"111010110",
  46567=>"000110010",
  46568=>"101001000",
  46569=>"101101001",
  46570=>"100101000",
  46571=>"000110101",
  46572=>"101100100",
  46573=>"111011110",
  46574=>"010111101",
  46575=>"101110000",
  46576=>"101110101",
  46577=>"011000110",
  46578=>"010100000",
  46579=>"001100011",
  46580=>"100000100",
  46581=>"010011110",
  46582=>"110101000",
  46583=>"001110101",
  46584=>"101001000",
  46585=>"011011100",
  46586=>"010000110",
  46587=>"100100100",
  46588=>"101101110",
  46589=>"001010101",
  46590=>"110101101",
  46591=>"001111101",
  46592=>"011100011",
  46593=>"100000110",
  46594=>"011011100",
  46595=>"111010101",
  46596=>"101111101",
  46597=>"001110010",
  46598=>"010000000",
  46599=>"101001001",
  46600=>"000001110",
  46601=>"010001110",
  46602=>"000101110",
  46603=>"011011111",
  46604=>"010010001",
  46605=>"011001101",
  46606=>"110001000",
  46607=>"001100001",
  46608=>"011011110",
  46609=>"011000001",
  46610=>"010110010",
  46611=>"000011011",
  46612=>"011000110",
  46613=>"011111011",
  46614=>"100000010",
  46615=>"001000001",
  46616=>"110001111",
  46617=>"001111100",
  46618=>"001001101",
  46619=>"110001001",
  46620=>"011101111",
  46621=>"011011001",
  46622=>"100010110",
  46623=>"101100101",
  46624=>"011010000",
  46625=>"100011010",
  46626=>"000110011",
  46627=>"010000110",
  46628=>"010010100",
  46629=>"001100111",
  46630=>"101010101",
  46631=>"101001010",
  46632=>"111111100",
  46633=>"100110001",
  46634=>"111110110",
  46635=>"001110000",
  46636=>"001000011",
  46637=>"010001010",
  46638=>"010100101",
  46639=>"000110000",
  46640=>"110110101",
  46641=>"110101110",
  46642=>"010111011",
  46643=>"101010011",
  46644=>"000110010",
  46645=>"010011111",
  46646=>"010100000",
  46647=>"010001100",
  46648=>"000001110",
  46649=>"100111111",
  46650=>"100011001",
  46651=>"101100111",
  46652=>"000111101",
  46653=>"111011001",
  46654=>"011110110",
  46655=>"110000100",
  46656=>"001000010",
  46657=>"000011000",
  46658=>"010101111",
  46659=>"001010011",
  46660=>"001110110",
  46661=>"111101111",
  46662=>"111111100",
  46663=>"100010000",
  46664=>"011001010",
  46665=>"111111000",
  46666=>"000011100",
  46667=>"100101110",
  46668=>"100101111",
  46669=>"000100011",
  46670=>"110100101",
  46671=>"101111111",
  46672=>"101001001",
  46673=>"100111100",
  46674=>"001001100",
  46675=>"001001010",
  46676=>"010010101",
  46677=>"101101001",
  46678=>"100010110",
  46679=>"111111100",
  46680=>"100111000",
  46681=>"111110011",
  46682=>"101101101",
  46683=>"110110011",
  46684=>"010010010",
  46685=>"111110101",
  46686=>"111000111",
  46687=>"000010011",
  46688=>"001101100",
  46689=>"111010001",
  46690=>"110011010",
  46691=>"001010010",
  46692=>"000000111",
  46693=>"011100010",
  46694=>"110001010",
  46695=>"001000011",
  46696=>"011111111",
  46697=>"000000011",
  46698=>"110011011",
  46699=>"000000100",
  46700=>"001100001",
  46701=>"110111100",
  46702=>"101011100",
  46703=>"011011011",
  46704=>"000100111",
  46705=>"010000000",
  46706=>"000101111",
  46707=>"001010110",
  46708=>"100111100",
  46709=>"111011011",
  46710=>"000100110",
  46711=>"101000111",
  46712=>"010111011",
  46713=>"001000111",
  46714=>"001101001",
  46715=>"111100110",
  46716=>"011000010",
  46717=>"011110110",
  46718=>"011000110",
  46719=>"001010011",
  46720=>"111100101",
  46721=>"001010100",
  46722=>"011010001",
  46723=>"000001101",
  46724=>"111110011",
  46725=>"110111011",
  46726=>"000001111",
  46727=>"001111111",
  46728=>"110000010",
  46729=>"011011000",
  46730=>"101000001",
  46731=>"101110110",
  46732=>"000011011",
  46733=>"011110111",
  46734=>"001000111",
  46735=>"011111110",
  46736=>"110111100",
  46737=>"110000000",
  46738=>"000101010",
  46739=>"011110100",
  46740=>"011000110",
  46741=>"010011110",
  46742=>"010000111",
  46743=>"000111000",
  46744=>"001101010",
  46745=>"111111001",
  46746=>"000101111",
  46747=>"100000011",
  46748=>"110101111",
  46749=>"011011111",
  46750=>"001001010",
  46751=>"010101000",
  46752=>"100000110",
  46753=>"001010001",
  46754=>"100110101",
  46755=>"111001010",
  46756=>"010001011",
  46757=>"101000001",
  46758=>"100011101",
  46759=>"111010111",
  46760=>"010100001",
  46761=>"111000001",
  46762=>"100111010",
  46763=>"000100111",
  46764=>"110111000",
  46765=>"100001110",
  46766=>"110111001",
  46767=>"101000010",
  46768=>"110001011",
  46769=>"100010111",
  46770=>"000111111",
  46771=>"110011010",
  46772=>"101100101",
  46773=>"011101100",
  46774=>"011111011",
  46775=>"100100010",
  46776=>"001011001",
  46777=>"101001000",
  46778=>"110001011",
  46779=>"111101100",
  46780=>"011100100",
  46781=>"001001001",
  46782=>"110110101",
  46783=>"110000001",
  46784=>"010101010",
  46785=>"011011101",
  46786=>"000101111",
  46787=>"011011011",
  46788=>"001001111",
  46789=>"101100100",
  46790=>"111101101",
  46791=>"000100111",
  46792=>"111010110",
  46793=>"000010000",
  46794=>"110001010",
  46795=>"101011110",
  46796=>"011010100",
  46797=>"100000010",
  46798=>"000010110",
  46799=>"000000001",
  46800=>"110111000",
  46801=>"111111111",
  46802=>"000001110",
  46803=>"111101110",
  46804=>"100101100",
  46805=>"110000111",
  46806=>"001110000",
  46807=>"000010111",
  46808=>"011101110",
  46809=>"011000010",
  46810=>"001110000",
  46811=>"101000000",
  46812=>"001000001",
  46813=>"010001010",
  46814=>"011001010",
  46815=>"001101011",
  46816=>"010110111",
  46817=>"111010101",
  46818=>"100001101",
  46819=>"111010011",
  46820=>"100001101",
  46821=>"101100101",
  46822=>"001010100",
  46823=>"011100101",
  46824=>"100010000",
  46825=>"011101011",
  46826=>"111111101",
  46827=>"000110000",
  46828=>"000000101",
  46829=>"100000001",
  46830=>"100101000",
  46831=>"100011111",
  46832=>"001000100",
  46833=>"111111110",
  46834=>"000001111",
  46835=>"001110000",
  46836=>"111011100",
  46837=>"100101110",
  46838=>"101010000",
  46839=>"010110111",
  46840=>"111101110",
  46841=>"101100110",
  46842=>"110100101",
  46843=>"011100100",
  46844=>"011010001",
  46845=>"000010011",
  46846=>"101100101",
  46847=>"111001110",
  46848=>"010110000",
  46849=>"101110101",
  46850=>"011111110",
  46851=>"011110110",
  46852=>"101111110",
  46853=>"111111111",
  46854=>"000001001",
  46855=>"001001100",
  46856=>"000001011",
  46857=>"101110101",
  46858=>"111110001",
  46859=>"111000000",
  46860=>"101100010",
  46861=>"011111101",
  46862=>"001000001",
  46863=>"010001011",
  46864=>"011101110",
  46865=>"000011111",
  46866=>"010101101",
  46867=>"000010111",
  46868=>"001011011",
  46869=>"011011001",
  46870=>"101010010",
  46871=>"101010000",
  46872=>"101001101",
  46873=>"110001010",
  46874=>"000001011",
  46875=>"110110111",
  46876=>"011000000",
  46877=>"010110110",
  46878=>"111010000",
  46879=>"001011111",
  46880=>"100000011",
  46881=>"111000001",
  46882=>"110101110",
  46883=>"000010110",
  46884=>"100101000",
  46885=>"001101100",
  46886=>"101010011",
  46887=>"001100010",
  46888=>"101010100",
  46889=>"111110111",
  46890=>"001100100",
  46891=>"100000001",
  46892=>"001111110",
  46893=>"000111001",
  46894=>"011111101",
  46895=>"101010011",
  46896=>"111100001",
  46897=>"011001111",
  46898=>"100000111",
  46899=>"010001100",
  46900=>"101010011",
  46901=>"010001001",
  46902=>"110101101",
  46903=>"100111000",
  46904=>"110101000",
  46905=>"101000100",
  46906=>"011011010",
  46907=>"111010101",
  46908=>"101100001",
  46909=>"111110110",
  46910=>"101101110",
  46911=>"001010000",
  46912=>"000101011",
  46913=>"011001100",
  46914=>"111111000",
  46915=>"111101110",
  46916=>"100000011",
  46917=>"111000100",
  46918=>"001110001",
  46919=>"101100000",
  46920=>"110101000",
  46921=>"000111101",
  46922=>"110111101",
  46923=>"100111110",
  46924=>"111111000",
  46925=>"001100011",
  46926=>"111000110",
  46927=>"110111111",
  46928=>"011100000",
  46929=>"111000011",
  46930=>"001011000",
  46931=>"111000111",
  46932=>"000111101",
  46933=>"100101100",
  46934=>"100111010",
  46935=>"010110111",
  46936=>"111010110",
  46937=>"011100111",
  46938=>"111001011",
  46939=>"111111111",
  46940=>"100011010",
  46941=>"011101101",
  46942=>"001011000",
  46943=>"011100001",
  46944=>"011011001",
  46945=>"110111101",
  46946=>"001000011",
  46947=>"010000101",
  46948=>"110001110",
  46949=>"001000110",
  46950=>"011001011",
  46951=>"110000110",
  46952=>"000011010",
  46953=>"010000011",
  46954=>"110101001",
  46955=>"101100011",
  46956=>"011001110",
  46957=>"111100001",
  46958=>"110100100",
  46959=>"000000010",
  46960=>"001000101",
  46961=>"000100001",
  46962=>"111001110",
  46963=>"111011100",
  46964=>"101001100",
  46965=>"100000100",
  46966=>"110011011",
  46967=>"111011100",
  46968=>"110111101",
  46969=>"100000000",
  46970=>"101100110",
  46971=>"001101000",
  46972=>"001010010",
  46973=>"110111111",
  46974=>"100101010",
  46975=>"000011010",
  46976=>"010000100",
  46977=>"011010000",
  46978=>"100111000",
  46979=>"101000111",
  46980=>"000011011",
  46981=>"100111011",
  46982=>"111011111",
  46983=>"010011001",
  46984=>"001110010",
  46985=>"001100001",
  46986=>"111101000",
  46987=>"110111111",
  46988=>"010010110",
  46989=>"011100110",
  46990=>"111111000",
  46991=>"000100000",
  46992=>"011100011",
  46993=>"111011111",
  46994=>"111100010",
  46995=>"011101101",
  46996=>"001010110",
  46997=>"010000001",
  46998=>"011101011",
  46999=>"011110110",
  47000=>"010111010",
  47001=>"000000001",
  47002=>"100100100",
  47003=>"110101110",
  47004=>"110001110",
  47005=>"001011110",
  47006=>"100000010",
  47007=>"010110011",
  47008=>"111101101",
  47009=>"110111111",
  47010=>"000100111",
  47011=>"011100100",
  47012=>"000010000",
  47013=>"100000110",
  47014=>"010111010",
  47015=>"100011110",
  47016=>"000110101",
  47017=>"001000110",
  47018=>"100110110",
  47019=>"011011101",
  47020=>"111111101",
  47021=>"011101111",
  47022=>"000010000",
  47023=>"011110101",
  47024=>"111111101",
  47025=>"111000000",
  47026=>"011101011",
  47027=>"011110101",
  47028=>"100010110",
  47029=>"011101011",
  47030=>"011001111",
  47031=>"101111001",
  47032=>"000100100",
  47033=>"110110000",
  47034=>"010111011",
  47035=>"001101101",
  47036=>"010101110",
  47037=>"100100111",
  47038=>"001111000",
  47039=>"100100100",
  47040=>"111001100",
  47041=>"100111110",
  47042=>"001101110",
  47043=>"011100011",
  47044=>"010101000",
  47045=>"110000100",
  47046=>"100000101",
  47047=>"000001010",
  47048=>"001110101",
  47049=>"001101110",
  47050=>"000001011",
  47051=>"101001111",
  47052=>"011110000",
  47053=>"000100110",
  47054=>"110010001",
  47055=>"110010001",
  47056=>"000110001",
  47057=>"110000010",
  47058=>"110010000",
  47059=>"110010000",
  47060=>"101000100",
  47061=>"011101000",
  47062=>"010101111",
  47063=>"110100111",
  47064=>"110010010",
  47065=>"111010011",
  47066=>"010111111",
  47067=>"101100000",
  47068=>"010010011",
  47069=>"000001101",
  47070=>"110011011",
  47071=>"010010100",
  47072=>"111110100",
  47073=>"001010000",
  47074=>"101010000",
  47075=>"001011001",
  47076=>"001000010",
  47077=>"110100100",
  47078=>"101011111",
  47079=>"101101010",
  47080=>"000111000",
  47081=>"101000101",
  47082=>"011111110",
  47083=>"100010000",
  47084=>"011111110",
  47085=>"110110011",
  47086=>"011011110",
  47087=>"111110111",
  47088=>"100001111",
  47089=>"101100011",
  47090=>"001000000",
  47091=>"010100011",
  47092=>"100000011",
  47093=>"101010001",
  47094=>"101000000",
  47095=>"100010000",
  47096=>"010101010",
  47097=>"110110011",
  47098=>"111001011",
  47099=>"000000001",
  47100=>"011000001",
  47101=>"101000000",
  47102=>"100000001",
  47103=>"011111010",
  47104=>"000001011",
  47105=>"011011101",
  47106=>"000101100",
  47107=>"100111001",
  47108=>"101000000",
  47109=>"011111100",
  47110=>"100111111",
  47111=>"011010101",
  47112=>"011110000",
  47113=>"011101111",
  47114=>"010100111",
  47115=>"100011010",
  47116=>"100101011",
  47117=>"000110010",
  47118=>"101010001",
  47119=>"000110111",
  47120=>"011100010",
  47121=>"000011001",
  47122=>"001110010",
  47123=>"001011011",
  47124=>"011111100",
  47125=>"100000000",
  47126=>"101010100",
  47127=>"110111001",
  47128=>"000000001",
  47129=>"011010010",
  47130=>"110101011",
  47131=>"000100010",
  47132=>"011011100",
  47133=>"000011110",
  47134=>"010010010",
  47135=>"110101101",
  47136=>"011110110",
  47137=>"101111101",
  47138=>"101010010",
  47139=>"011100111",
  47140=>"010001111",
  47141=>"111100010",
  47142=>"011001101",
  47143=>"110011111",
  47144=>"111010101",
  47145=>"010010110",
  47146=>"100010001",
  47147=>"001011110",
  47148=>"011110111",
  47149=>"111101001",
  47150=>"010110110",
  47151=>"100101001",
  47152=>"111110000",
  47153=>"011110001",
  47154=>"000111010",
  47155=>"000110001",
  47156=>"010111010",
  47157=>"001100001",
  47158=>"000011100",
  47159=>"011111011",
  47160=>"011101001",
  47161=>"111010101",
  47162=>"110101101",
  47163=>"000100001",
  47164=>"011110111",
  47165=>"010101110",
  47166=>"010011110",
  47167=>"100110011",
  47168=>"100100100",
  47169=>"100110101",
  47170=>"011000111",
  47171=>"100010111",
  47172=>"000110001",
  47173=>"011001000",
  47174=>"010010000",
  47175=>"111100111",
  47176=>"111101101",
  47177=>"100110111",
  47178=>"011001001",
  47179=>"011111111",
  47180=>"101011000",
  47181=>"001001010",
  47182=>"110100001",
  47183=>"010001111",
  47184=>"110111111",
  47185=>"010110000",
  47186=>"011101000",
  47187=>"000111001",
  47188=>"100100100",
  47189=>"000100000",
  47190=>"101011010",
  47191=>"111001000",
  47192=>"100110000",
  47193=>"000101101",
  47194=>"010100001",
  47195=>"100100111",
  47196=>"101010100",
  47197=>"111010000",
  47198=>"111000000",
  47199=>"110010001",
  47200=>"000101001",
  47201=>"010100000",
  47202=>"000101110",
  47203=>"000010001",
  47204=>"011101001",
  47205=>"011111111",
  47206=>"111001100",
  47207=>"110010010",
  47208=>"100011001",
  47209=>"111110100",
  47210=>"111110001",
  47211=>"011101010",
  47212=>"000111011",
  47213=>"111010110",
  47214=>"100110000",
  47215=>"110110000",
  47216=>"010000011",
  47217=>"110011110",
  47218=>"000110011",
  47219=>"110110111",
  47220=>"011100101",
  47221=>"011111001",
  47222=>"000110001",
  47223=>"000000011",
  47224=>"110000011",
  47225=>"100101000",
  47226=>"000010100",
  47227=>"000000000",
  47228=>"110110000",
  47229=>"101010000",
  47230=>"010101101",
  47231=>"110001000",
  47232=>"001010110",
  47233=>"100011001",
  47234=>"010011011",
  47235=>"101111111",
  47236=>"011011110",
  47237=>"000001001",
  47238=>"011101101",
  47239=>"100111010",
  47240=>"001001000",
  47241=>"111011111",
  47242=>"011101100",
  47243=>"111111110",
  47244=>"100111011",
  47245=>"100101110",
  47246=>"110101110",
  47247=>"111101010",
  47248=>"001100100",
  47249=>"100101100",
  47250=>"100111101",
  47251=>"111011000",
  47252=>"010111100",
  47253=>"100110110",
  47254=>"000011001",
  47255=>"001101110",
  47256=>"010000100",
  47257=>"000010100",
  47258=>"100111101",
  47259=>"011001110",
  47260=>"001101011",
  47261=>"100111000",
  47262=>"101100011",
  47263=>"101000000",
  47264=>"110010111",
  47265=>"011111000",
  47266=>"101000000",
  47267=>"001101100",
  47268=>"011001111",
  47269=>"100010011",
  47270=>"000011001",
  47271=>"100001000",
  47272=>"001111101",
  47273=>"001001011",
  47274=>"111110111",
  47275=>"111110111",
  47276=>"111000000",
  47277=>"000101001",
  47278=>"110010101",
  47279=>"101110110",
  47280=>"111010001",
  47281=>"010100100",
  47282=>"101101111",
  47283=>"110101011",
  47284=>"011110001",
  47285=>"111110000",
  47286=>"010011010",
  47287=>"011111001",
  47288=>"110111010",
  47289=>"101101101",
  47290=>"110111100",
  47291=>"011111000",
  47292=>"111001100",
  47293=>"111000000",
  47294=>"110010011",
  47295=>"111111111",
  47296=>"111001100",
  47297=>"000000100",
  47298=>"101001100",
  47299=>"010011010",
  47300=>"110011000",
  47301=>"001000010",
  47302=>"001111110",
  47303=>"110011011",
  47304=>"000010000",
  47305=>"010101010",
  47306=>"111010001",
  47307=>"111101110",
  47308=>"111011011",
  47309=>"110110111",
  47310=>"011011101",
  47311=>"000101001",
  47312=>"011011100",
  47313=>"101101100",
  47314=>"011101001",
  47315=>"010001101",
  47316=>"010010001",
  47317=>"100000100",
  47318=>"111111111",
  47319=>"111011100",
  47320=>"000100101",
  47321=>"000101010",
  47322=>"111000111",
  47323=>"000101101",
  47324=>"010000110",
  47325=>"011101001",
  47326=>"001001001",
  47327=>"100111100",
  47328=>"111000000",
  47329=>"110010000",
  47330=>"111111101",
  47331=>"111110001",
  47332=>"101001010",
  47333=>"001000000",
  47334=>"110110000",
  47335=>"110001001",
  47336=>"100011100",
  47337=>"010010011",
  47338=>"101011001",
  47339=>"110101101",
  47340=>"100101010",
  47341=>"000110101",
  47342=>"000000011",
  47343=>"111001000",
  47344=>"101101001",
  47345=>"011000001",
  47346=>"101000101",
  47347=>"111101110",
  47348=>"010011010",
  47349=>"000101111",
  47350=>"100011011",
  47351=>"000001110",
  47352=>"110101101",
  47353=>"111001011",
  47354=>"010100111",
  47355=>"001111001",
  47356=>"101110010",
  47357=>"110011111",
  47358=>"001101100",
  47359=>"001100111",
  47360=>"010000010",
  47361=>"011011110",
  47362=>"001000000",
  47363=>"010111000",
  47364=>"010101010",
  47365=>"000101011",
  47366=>"000101101",
  47367=>"100101100",
  47368=>"101111001",
  47369=>"100110101",
  47370=>"100000101",
  47371=>"110100000",
  47372=>"010011011",
  47373=>"100101111",
  47374=>"101111110",
  47375=>"101100101",
  47376=>"110001011",
  47377=>"001001001",
  47378=>"000110000",
  47379=>"111010110",
  47380=>"101100000",
  47381=>"101001111",
  47382=>"100011000",
  47383=>"001111000",
  47384=>"110001110",
  47385=>"100001100",
  47386=>"101111011",
  47387=>"100111010",
  47388=>"111100010",
  47389=>"100011110",
  47390=>"110011110",
  47391=>"100010001",
  47392=>"000101101",
  47393=>"101011001",
  47394=>"001101110",
  47395=>"111000100",
  47396=>"000011010",
  47397=>"111101110",
  47398=>"110110100",
  47399=>"111101001",
  47400=>"101000010",
  47401=>"110001001",
  47402=>"011001001",
  47403=>"100100111",
  47404=>"110011110",
  47405=>"010001100",
  47406=>"110111001",
  47407=>"111110111",
  47408=>"101110011",
  47409=>"010011110",
  47410=>"011101110",
  47411=>"000000000",
  47412=>"100001011",
  47413=>"000011011",
  47414=>"111101010",
  47415=>"000111100",
  47416=>"100101110",
  47417=>"011011000",
  47418=>"101101011",
  47419=>"111011001",
  47420=>"101101110",
  47421=>"001010010",
  47422=>"010100111",
  47423=>"010010111",
  47424=>"101110011",
  47425=>"100101000",
  47426=>"010011001",
  47427=>"000111110",
  47428=>"100110110",
  47429=>"110000000",
  47430=>"000110001",
  47431=>"100110100",
  47432=>"011101101",
  47433=>"100010010",
  47434=>"001011011",
  47435=>"010011001",
  47436=>"100101101",
  47437=>"100010111",
  47438=>"000000110",
  47439=>"010001101",
  47440=>"110011110",
  47441=>"001110000",
  47442=>"111100010",
  47443=>"100111111",
  47444=>"000001001",
  47445=>"110101110",
  47446=>"001000011",
  47447=>"010101000",
  47448=>"001110110",
  47449=>"110010000",
  47450=>"010100000",
  47451=>"101111001",
  47452=>"001100111",
  47453=>"010111111",
  47454=>"111010111",
  47455=>"100111001",
  47456=>"100000011",
  47457=>"010110110",
  47458=>"111001010",
  47459=>"111110000",
  47460=>"010011010",
  47461=>"101000111",
  47462=>"111111011",
  47463=>"011111010",
  47464=>"000101111",
  47465=>"111100010",
  47466=>"000100100",
  47467=>"101100111",
  47468=>"100001110",
  47469=>"001001110",
  47470=>"100101101",
  47471=>"001111000",
  47472=>"100100111",
  47473=>"101100000",
  47474=>"011100101",
  47475=>"100111110",
  47476=>"011100100",
  47477=>"110000001",
  47478=>"001011011",
  47479=>"001001101",
  47480=>"110000011",
  47481=>"110010110",
  47482=>"101000100",
  47483=>"101100101",
  47484=>"011101000",
  47485=>"100110010",
  47486=>"011100010",
  47487=>"000101001",
  47488=>"110001000",
  47489=>"001111111",
  47490=>"100101011",
  47491=>"100101010",
  47492=>"110101100",
  47493=>"010100001",
  47494=>"100001111",
  47495=>"111100110",
  47496=>"000000101",
  47497=>"101000110",
  47498=>"001001111",
  47499=>"011110101",
  47500=>"010111101",
  47501=>"000000011",
  47502=>"010001110",
  47503=>"010110010",
  47504=>"010110001",
  47505=>"111001001",
  47506=>"001000101",
  47507=>"001010010",
  47508=>"110101110",
  47509=>"111011100",
  47510=>"111101001",
  47511=>"111111100",
  47512=>"101101011",
  47513=>"111101011",
  47514=>"001011110",
  47515=>"001101000",
  47516=>"100011111",
  47517=>"111001011",
  47518=>"100011001",
  47519=>"111010000",
  47520=>"101101000",
  47521=>"111000011",
  47522=>"110111010",
  47523=>"101011001",
  47524=>"010001100",
  47525=>"101101100",
  47526=>"000011111",
  47527=>"001100000",
  47528=>"101000011",
  47529=>"111000000",
  47530=>"101101000",
  47531=>"111001101",
  47532=>"011000011",
  47533=>"010100000",
  47534=>"010011110",
  47535=>"011110011",
  47536=>"110001010",
  47537=>"100000101",
  47538=>"000100001",
  47539=>"001000010",
  47540=>"100110010",
  47541=>"011101010",
  47542=>"100011111",
  47543=>"010101000",
  47544=>"000101000",
  47545=>"101000111",
  47546=>"111011110",
  47547=>"011011100",
  47548=>"001110000",
  47549=>"110001111",
  47550=>"000100011",
  47551=>"001011000",
  47552=>"010100011",
  47553=>"000111010",
  47554=>"011010100",
  47555=>"110100001",
  47556=>"101100100",
  47557=>"111111111",
  47558=>"111100011",
  47559=>"101101000",
  47560=>"111000111",
  47561=>"001101111",
  47562=>"000100001",
  47563=>"011110011",
  47564=>"001100110",
  47565=>"010010001",
  47566=>"100110101",
  47567=>"010111010",
  47568=>"000001000",
  47569=>"111110110",
  47570=>"101100100",
  47571=>"101110101",
  47572=>"110101111",
  47573=>"011011000",
  47574=>"100111010",
  47575=>"110011011",
  47576=>"001100011",
  47577=>"010000110",
  47578=>"100111100",
  47579=>"001011100",
  47580=>"011010001",
  47581=>"001001001",
  47582=>"011110010",
  47583=>"001001010",
  47584=>"111010100",
  47585=>"111010011",
  47586=>"110111110",
  47587=>"001011001",
  47588=>"111111001",
  47589=>"000100000",
  47590=>"110010101",
  47591=>"000110111",
  47592=>"001000100",
  47593=>"110101100",
  47594=>"001000000",
  47595=>"011110101",
  47596=>"111100101",
  47597=>"111001100",
  47598=>"100111111",
  47599=>"001111111",
  47600=>"111111000",
  47601=>"000001010",
  47602=>"010010011",
  47603=>"100100110",
  47604=>"110110100",
  47605=>"010101101",
  47606=>"000101011",
  47607=>"011111100",
  47608=>"110100100",
  47609=>"100011101",
  47610=>"101000001",
  47611=>"010111010",
  47612=>"000101100",
  47613=>"111110001",
  47614=>"001010011",
  47615=>"001010001",
  47616=>"100011011",
  47617=>"010001111",
  47618=>"010011000",
  47619=>"101001101",
  47620=>"100111110",
  47621=>"111000001",
  47622=>"110000111",
  47623=>"011100100",
  47624=>"100111011",
  47625=>"000011110",
  47626=>"111011010",
  47627=>"000010011",
  47628=>"100000110",
  47629=>"100101101",
  47630=>"011000010",
  47631=>"111001110",
  47632=>"001110110",
  47633=>"000000011",
  47634=>"000111001",
  47635=>"001001001",
  47636=>"110111010",
  47637=>"101010101",
  47638=>"011011100",
  47639=>"000011011",
  47640=>"001011110",
  47641=>"101110000",
  47642=>"110101111",
  47643=>"100001000",
  47644=>"110111011",
  47645=>"100010111",
  47646=>"000000010",
  47647=>"010010100",
  47648=>"011011101",
  47649=>"110101101",
  47650=>"111011000",
  47651=>"101111111",
  47652=>"001101001",
  47653=>"110111111",
  47654=>"001110101",
  47655=>"101000000",
  47656=>"011110110",
  47657=>"100000000",
  47658=>"011011100",
  47659=>"111010111",
  47660=>"010000011",
  47661=>"111001101",
  47662=>"111110100",
  47663=>"110001110",
  47664=>"000110110",
  47665=>"010100100",
  47666=>"010110100",
  47667=>"000000101",
  47668=>"101111010",
  47669=>"110110110",
  47670=>"001001110",
  47671=>"100000010",
  47672=>"100011111",
  47673=>"110010101",
  47674=>"010001100",
  47675=>"001000000",
  47676=>"111111110",
  47677=>"010100010",
  47678=>"011000001",
  47679=>"000111001",
  47680=>"111110011",
  47681=>"000000110",
  47682=>"100001101",
  47683=>"100011111",
  47684=>"010101000",
  47685=>"011111100",
  47686=>"111001001",
  47687=>"001010000",
  47688=>"011001110",
  47689=>"101011111",
  47690=>"100111010",
  47691=>"101101000",
  47692=>"000000011",
  47693=>"101000101",
  47694=>"100111111",
  47695=>"000101011",
  47696=>"110111110",
  47697=>"110110111",
  47698=>"001000001",
  47699=>"011110011",
  47700=>"000001011",
  47701=>"101111010",
  47702=>"100001101",
  47703=>"010110010",
  47704=>"001110001",
  47705=>"101000001",
  47706=>"001100101",
  47707=>"101001101",
  47708=>"010011111",
  47709=>"010000101",
  47710=>"101100001",
  47711=>"000001000",
  47712=>"101001011",
  47713=>"101001001",
  47714=>"010100101",
  47715=>"111100111",
  47716=>"100111101",
  47717=>"100100100",
  47718=>"001100110",
  47719=>"111101011",
  47720=>"111111101",
  47721=>"011110010",
  47722=>"000000011",
  47723=>"011111101",
  47724=>"101001010",
  47725=>"110000111",
  47726=>"100110111",
  47727=>"001111110",
  47728=>"001111110",
  47729=>"001100101",
  47730=>"110000010",
  47731=>"101010101",
  47732=>"111110101",
  47733=>"101011001",
  47734=>"101100111",
  47735=>"101100000",
  47736=>"110011001",
  47737=>"101100011",
  47738=>"100001110",
  47739=>"010011101",
  47740=>"000100010",
  47741=>"100111011",
  47742=>"011010000",
  47743=>"010101111",
  47744=>"101001001",
  47745=>"001101100",
  47746=>"101110000",
  47747=>"100100101",
  47748=>"011010111",
  47749=>"001000000",
  47750=>"011100000",
  47751=>"110100001",
  47752=>"111100011",
  47753=>"001100101",
  47754=>"100111001",
  47755=>"010000110",
  47756=>"111100011",
  47757=>"101111110",
  47758=>"011100101",
  47759=>"101101010",
  47760=>"111011101",
  47761=>"011101011",
  47762=>"100010100",
  47763=>"110110111",
  47764=>"000111000",
  47765=>"101001011",
  47766=>"110000101",
  47767=>"110111101",
  47768=>"000010001",
  47769=>"010111000",
  47770=>"011101000",
  47771=>"000011101",
  47772=>"000111000",
  47773=>"011100111",
  47774=>"010110011",
  47775=>"101110110",
  47776=>"111000000",
  47777=>"010010101",
  47778=>"111101010",
  47779=>"110110111",
  47780=>"101010110",
  47781=>"101111100",
  47782=>"110011111",
  47783=>"101001111",
  47784=>"101111011",
  47785=>"010011011",
  47786=>"010101101",
  47787=>"010011111",
  47788=>"110010001",
  47789=>"111011001",
  47790=>"101101000",
  47791=>"101111101",
  47792=>"011100101",
  47793=>"110110100",
  47794=>"011111111",
  47795=>"001001001",
  47796=>"100111111",
  47797=>"100011110",
  47798=>"101100100",
  47799=>"001011000",
  47800=>"010000000",
  47801=>"101101110",
  47802=>"101010000",
  47803=>"010111110",
  47804=>"001011010",
  47805=>"001000010",
  47806=>"010001011",
  47807=>"011111011",
  47808=>"100111100",
  47809=>"001101011",
  47810=>"011010100",
  47811=>"100000100",
  47812=>"000010001",
  47813=>"011110111",
  47814=>"110000111",
  47815=>"101111000",
  47816=>"001100000",
  47817=>"111110111",
  47818=>"001100001",
  47819=>"001000001",
  47820=>"111111110",
  47821=>"101000100",
  47822=>"010011000",
  47823=>"010111011",
  47824=>"000000011",
  47825=>"011110111",
  47826=>"010000100",
  47827=>"011011000",
  47828=>"100111001",
  47829=>"000000110",
  47830=>"011010101",
  47831=>"110100010",
  47832=>"110000101",
  47833=>"101100000",
  47834=>"000011010",
  47835=>"010000110",
  47836=>"101001100",
  47837=>"010001100",
  47838=>"110101010",
  47839=>"010001101",
  47840=>"101100011",
  47841=>"100101000",
  47842=>"101000011",
  47843=>"101100011",
  47844=>"100111111",
  47845=>"011010000",
  47846=>"110001001",
  47847=>"000101000",
  47848=>"110101100",
  47849=>"101010001",
  47850=>"101000000",
  47851=>"101011011",
  47852=>"100100000",
  47853=>"011111101",
  47854=>"101101101",
  47855=>"011111001",
  47856=>"000110011",
  47857=>"101110110",
  47858=>"101101000",
  47859=>"101110011",
  47860=>"011011010",
  47861=>"000010110",
  47862=>"100101111",
  47863=>"000010110",
  47864=>"111001011",
  47865=>"010100010",
  47866=>"011110010",
  47867=>"010000000",
  47868=>"001010101",
  47869=>"100010001",
  47870=>"011110101",
  47871=>"100010010",
  47872=>"110011110",
  47873=>"111100011",
  47874=>"111000111",
  47875=>"001101010",
  47876=>"100000110",
  47877=>"100110101",
  47878=>"111010011",
  47879=>"010111011",
  47880=>"011011001",
  47881=>"110110001",
  47882=>"110010010",
  47883=>"011111100",
  47884=>"101101101",
  47885=>"011100000",
  47886=>"110110111",
  47887=>"000111011",
  47888=>"101010000",
  47889=>"001111110",
  47890=>"110110110",
  47891=>"101000001",
  47892=>"110011010",
  47893=>"100000010",
  47894=>"110100110",
  47895=>"001110001",
  47896=>"101001001",
  47897=>"101011101",
  47898=>"101101000",
  47899=>"110111111",
  47900=>"101101000",
  47901=>"111111100",
  47902=>"000111001",
  47903=>"111011101",
  47904=>"010110111",
  47905=>"110100110",
  47906=>"010000101",
  47907=>"100111000",
  47908=>"011011101",
  47909=>"010100101",
  47910=>"100100111",
  47911=>"011101010",
  47912=>"101011101",
  47913=>"000111110",
  47914=>"011110100",
  47915=>"101100101",
  47916=>"000100000",
  47917=>"101000100",
  47918=>"110001101",
  47919=>"110110111",
  47920=>"000010111",
  47921=>"011011101",
  47922=>"000000010",
  47923=>"111111111",
  47924=>"111110011",
  47925=>"110110000",
  47926=>"010011001",
  47927=>"010100011",
  47928=>"101100110",
  47929=>"111000001",
  47930=>"001100001",
  47931=>"011011010",
  47932=>"101101001",
  47933=>"110001100",
  47934=>"000010110",
  47935=>"110100100",
  47936=>"111101110",
  47937=>"000111000",
  47938=>"010110110",
  47939=>"011100001",
  47940=>"000111111",
  47941=>"011101110",
  47942=>"100010101",
  47943=>"111001011",
  47944=>"000110000",
  47945=>"011100000",
  47946=>"001100110",
  47947=>"100000101",
  47948=>"100111110",
  47949=>"000000100",
  47950=>"110100001",
  47951=>"100110100",
  47952=>"100000000",
  47953=>"101000110",
  47954=>"001001011",
  47955=>"110111000",
  47956=>"001100011",
  47957=>"111000100",
  47958=>"110100101",
  47959=>"001000000",
  47960=>"110111011",
  47961=>"000001111",
  47962=>"110010001",
  47963=>"010000011",
  47964=>"000101010",
  47965=>"101000111",
  47966=>"001101000",
  47967=>"001101010",
  47968=>"111100100",
  47969=>"011101010",
  47970=>"001000001",
  47971=>"101001000",
  47972=>"011100110",
  47973=>"011101101",
  47974=>"101100001",
  47975=>"100010100",
  47976=>"110000000",
  47977=>"100101011",
  47978=>"110011100",
  47979=>"011111101",
  47980=>"110101011",
  47981=>"101001101",
  47982=>"001101101",
  47983=>"001110011",
  47984=>"111110101",
  47985=>"001000001",
  47986=>"011111101",
  47987=>"011001000",
  47988=>"111001010",
  47989=>"101001100",
  47990=>"101100011",
  47991=>"101011100",
  47992=>"101111110",
  47993=>"110000001",
  47994=>"111001010",
  47995=>"110001110",
  47996=>"111011111",
  47997=>"101000001",
  47998=>"111001101",
  47999=>"011100001",
  48000=>"111111001",
  48001=>"101110111",
  48002=>"001100010",
  48003=>"011100101",
  48004=>"011100111",
  48005=>"101110111",
  48006=>"101000100",
  48007=>"010101111",
  48008=>"101100111",
  48009=>"011111010",
  48010=>"110100000",
  48011=>"101110011",
  48012=>"100110001",
  48013=>"111010011",
  48014=>"000100110",
  48015=>"001100111",
  48016=>"010011111",
  48017=>"000111111",
  48018=>"011010101",
  48019=>"000110010",
  48020=>"010110110",
  48021=>"101101000",
  48022=>"101001101",
  48023=>"100101010",
  48024=>"011100111",
  48025=>"000001000",
  48026=>"100010011",
  48027=>"011100101",
  48028=>"110110000",
  48029=>"101101001",
  48030=>"101001111",
  48031=>"000101001",
  48032=>"111111100",
  48033=>"111111100",
  48034=>"101101100",
  48035=>"101111110",
  48036=>"000011001",
  48037=>"001011000",
  48038=>"111001111",
  48039=>"110010010",
  48040=>"010110011",
  48041=>"110101100",
  48042=>"110011011",
  48043=>"100101101",
  48044=>"010101100",
  48045=>"110001001",
  48046=>"101101111",
  48047=>"110011001",
  48048=>"010111111",
  48049=>"100101111",
  48050=>"001000110",
  48051=>"011001010",
  48052=>"111100010",
  48053=>"111101111",
  48054=>"100001101",
  48055=>"101100011",
  48056=>"110111001",
  48057=>"110011011",
  48058=>"110100110",
  48059=>"100010111",
  48060=>"000010100",
  48061=>"000100100",
  48062=>"000111100",
  48063=>"001001111",
  48064=>"111010010",
  48065=>"010110110",
  48066=>"011111010",
  48067=>"000101100",
  48068=>"010001111",
  48069=>"010111011",
  48070=>"001101100",
  48071=>"000100110",
  48072=>"100011000",
  48073=>"010100010",
  48074=>"011011110",
  48075=>"101010000",
  48076=>"110001000",
  48077=>"101111110",
  48078=>"001000000",
  48079=>"101110100",
  48080=>"100011110",
  48081=>"000100110",
  48082=>"011001101",
  48083=>"101010000",
  48084=>"000010010",
  48085=>"110000101",
  48086=>"101111111",
  48087=>"101000010",
  48088=>"100000000",
  48089=>"000000110",
  48090=>"000010101",
  48091=>"000111011",
  48092=>"000101101",
  48093=>"000110100",
  48094=>"010101000",
  48095=>"010100011",
  48096=>"110001100",
  48097=>"111101101",
  48098=>"111111110",
  48099=>"110010010",
  48100=>"100000111",
  48101=>"011100110",
  48102=>"111101111",
  48103=>"100001100",
  48104=>"101111011",
  48105=>"001000011",
  48106=>"011111011",
  48107=>"010011000",
  48108=>"101110100",
  48109=>"010010111",
  48110=>"101110111",
  48111=>"000100000",
  48112=>"110001011",
  48113=>"000001110",
  48114=>"001010000",
  48115=>"010100101",
  48116=>"110000101",
  48117=>"011000001",
  48118=>"000011100",
  48119=>"011100100",
  48120=>"001001101",
  48121=>"101111111",
  48122=>"111011100",
  48123=>"001010010",
  48124=>"001001110",
  48125=>"110000110",
  48126=>"101101111",
  48127=>"110111111",
  48128=>"000101000",
  48129=>"001110011",
  48130=>"011101100",
  48131=>"111000100",
  48132=>"011101011",
  48133=>"101000011",
  48134=>"010100111",
  48135=>"001111000",
  48136=>"010000010",
  48137=>"000010011",
  48138=>"001111101",
  48139=>"111101011",
  48140=>"011101011",
  48141=>"110001100",
  48142=>"100010010",
  48143=>"111000010",
  48144=>"010000100",
  48145=>"000101010",
  48146=>"000010100",
  48147=>"111100010",
  48148=>"111100010",
  48149=>"101000010",
  48150=>"010001001",
  48151=>"011101001",
  48152=>"101101000",
  48153=>"011010000",
  48154=>"101011011",
  48155=>"101110000",
  48156=>"110101011",
  48157=>"011100100",
  48158=>"000011000",
  48159=>"011000011",
  48160=>"101011001",
  48161=>"001110011",
  48162=>"110010101",
  48163=>"010000010",
  48164=>"110100001",
  48165=>"110110110",
  48166=>"100010101",
  48167=>"010001111",
  48168=>"110110000",
  48169=>"110111010",
  48170=>"111011111",
  48171=>"011000000",
  48172=>"100010001",
  48173=>"101011101",
  48174=>"111110110",
  48175=>"100111010",
  48176=>"011100011",
  48177=>"011110000",
  48178=>"111110011",
  48179=>"011000010",
  48180=>"001001000",
  48181=>"101100101",
  48182=>"100110100",
  48183=>"110010100",
  48184=>"001110111",
  48185=>"001000001",
  48186=>"110011000",
  48187=>"101000100",
  48188=>"000110111",
  48189=>"000000000",
  48190=>"010011010",
  48191=>"111011011",
  48192=>"011011000",
  48193=>"000010110",
  48194=>"010001111",
  48195=>"100001101",
  48196=>"100110000",
  48197=>"001111110",
  48198=>"011001010",
  48199=>"010001101",
  48200=>"100100111",
  48201=>"111100101",
  48202=>"110111001",
  48203=>"100000101",
  48204=>"000110010",
  48205=>"000011011",
  48206=>"110110101",
  48207=>"000100010",
  48208=>"001011101",
  48209=>"111100000",
  48210=>"010000011",
  48211=>"010011001",
  48212=>"101110010",
  48213=>"100100110",
  48214=>"111011001",
  48215=>"100000100",
  48216=>"101001000",
  48217=>"100010000",
  48218=>"110011011",
  48219=>"111100011",
  48220=>"001110000",
  48221=>"101011101",
  48222=>"010000011",
  48223=>"101111111",
  48224=>"010101111",
  48225=>"010111011",
  48226=>"010100011",
  48227=>"000010011",
  48228=>"100101101",
  48229=>"111011000",
  48230=>"010010110",
  48231=>"110111001",
  48232=>"010100100",
  48233=>"011101111",
  48234=>"101001001",
  48235=>"000001000",
  48236=>"111001100",
  48237=>"001010101",
  48238=>"111011000",
  48239=>"010100100",
  48240=>"111001111",
  48241=>"011111001",
  48242=>"111111110",
  48243=>"100101101",
  48244=>"000001110",
  48245=>"100001011",
  48246=>"101000000",
  48247=>"010001101",
  48248=>"101010000",
  48249=>"000000100",
  48250=>"000000110",
  48251=>"010001100",
  48252=>"110000010",
  48253=>"101011110",
  48254=>"011100000",
  48255=>"011010111",
  48256=>"100111000",
  48257=>"110001110",
  48258=>"110000111",
  48259=>"001010111",
  48260=>"001001111",
  48261=>"100100100",
  48262=>"101110101",
  48263=>"001001010",
  48264=>"000110100",
  48265=>"001000000",
  48266=>"010001110",
  48267=>"110110100",
  48268=>"001101100",
  48269=>"010011111",
  48270=>"011000011",
  48271=>"110000110",
  48272=>"111110100",
  48273=>"110101111",
  48274=>"101101000",
  48275=>"110001101",
  48276=>"011101111",
  48277=>"000101011",
  48278=>"001111100",
  48279=>"110110101",
  48280=>"101011110",
  48281=>"101001111",
  48282=>"111101100",
  48283=>"111111101",
  48284=>"011001101",
  48285=>"111000101",
  48286=>"001000011",
  48287=>"101011111",
  48288=>"111101000",
  48289=>"001100111",
  48290=>"000010000",
  48291=>"100111010",
  48292=>"010000101",
  48293=>"010100110",
  48294=>"000100010",
  48295=>"101001011",
  48296=>"100001100",
  48297=>"110100011",
  48298=>"010111010",
  48299=>"101111100",
  48300=>"110110000",
  48301=>"110000110",
  48302=>"101000110",
  48303=>"010110011",
  48304=>"010110110",
  48305=>"110111111",
  48306=>"011001110",
  48307=>"001101010",
  48308=>"011001000",
  48309=>"000001001",
  48310=>"011101111",
  48311=>"001101110",
  48312=>"011110101",
  48313=>"011111101",
  48314=>"011000111",
  48315=>"000111000",
  48316=>"001010110",
  48317=>"100000101",
  48318=>"000111011",
  48319=>"010110011",
  48320=>"111111011",
  48321=>"100011111",
  48322=>"100100101",
  48323=>"100001100",
  48324=>"000001111",
  48325=>"110011001",
  48326=>"101000000",
  48327=>"111100100",
  48328=>"100010110",
  48329=>"111001111",
  48330=>"101001111",
  48331=>"000110000",
  48332=>"001101000",
  48333=>"111111001",
  48334=>"000100010",
  48335=>"110100110",
  48336=>"111100110",
  48337=>"101001101",
  48338=>"000000000",
  48339=>"010111001",
  48340=>"010001100",
  48341=>"100011110",
  48342=>"110000101",
  48343=>"011111100",
  48344=>"010000110",
  48345=>"101101011",
  48346=>"000000001",
  48347=>"111001000",
  48348=>"001000100",
  48349=>"110110111",
  48350=>"111111111",
  48351=>"101101101",
  48352=>"001100111",
  48353=>"011111100",
  48354=>"010010101",
  48355=>"010010110",
  48356=>"000011110",
  48357=>"111111000",
  48358=>"010000000",
  48359=>"100000100",
  48360=>"101010110",
  48361=>"010100011",
  48362=>"101100110",
  48363=>"000011010",
  48364=>"111101010",
  48365=>"111001000",
  48366=>"101100011",
  48367=>"011001011",
  48368=>"000000111",
  48369=>"101111110",
  48370=>"100111101",
  48371=>"111111111",
  48372=>"011101101",
  48373=>"001000111",
  48374=>"000111010",
  48375=>"000110111",
  48376=>"101011001",
  48377=>"111011011",
  48378=>"000001010",
  48379=>"110000101",
  48380=>"010001111",
  48381=>"000000000",
  48382=>"011100100",
  48383=>"001010011",
  48384=>"110000001",
  48385=>"110011110",
  48386=>"000111010",
  48387=>"110011100",
  48388=>"001110100",
  48389=>"101111010",
  48390=>"111100001",
  48391=>"010110000",
  48392=>"101101010",
  48393=>"100010111",
  48394=>"011100001",
  48395=>"100110110",
  48396=>"111111010",
  48397=>"011111110",
  48398=>"110101001",
  48399=>"110010111",
  48400=>"111011110",
  48401=>"101100011",
  48402=>"100010101",
  48403=>"100111111",
  48404=>"010001001",
  48405=>"100111100",
  48406=>"010011000",
  48407=>"011011011",
  48408=>"011100011",
  48409=>"100100001",
  48410=>"111101100",
  48411=>"111010000",
  48412=>"111100110",
  48413=>"101000001",
  48414=>"001111111",
  48415=>"011100000",
  48416=>"000011101",
  48417=>"011111101",
  48418=>"001101011",
  48419=>"010000001",
  48420=>"101001000",
  48421=>"111011001",
  48422=>"101110101",
  48423=>"010000111",
  48424=>"011110000",
  48425=>"001011000",
  48426=>"100011111",
  48427=>"101011110",
  48428=>"000011010",
  48429=>"010000101",
  48430=>"111111111",
  48431=>"001111000",
  48432=>"110000110",
  48433=>"111100001",
  48434=>"100111010",
  48435=>"111010111",
  48436=>"001100010",
  48437=>"100111110",
  48438=>"110101010",
  48439=>"100010111",
  48440=>"101101011",
  48441=>"000111010",
  48442=>"000010000",
  48443=>"110100100",
  48444=>"011000110",
  48445=>"111011011",
  48446=>"001000011",
  48447=>"010100000",
  48448=>"100001000",
  48449=>"101001000",
  48450=>"110111101",
  48451=>"010010010",
  48452=>"011110011",
  48453=>"011110101",
  48454=>"001101100",
  48455=>"000110000",
  48456=>"011100111",
  48457=>"100000011",
  48458=>"111110000",
  48459=>"010000101",
  48460=>"011001101",
  48461=>"100110111",
  48462=>"100010110",
  48463=>"010111001",
  48464=>"110001111",
  48465=>"001101010",
  48466=>"101101101",
  48467=>"111100011",
  48468=>"011010010",
  48469=>"111111100",
  48470=>"000001010",
  48471=>"110010001",
  48472=>"001111111",
  48473=>"101110000",
  48474=>"000100101",
  48475=>"111111001",
  48476=>"001111111",
  48477=>"001000111",
  48478=>"101010001",
  48479=>"111000001",
  48480=>"101101111",
  48481=>"011001011",
  48482=>"101110111",
  48483=>"000101000",
  48484=>"010011100",
  48485=>"100010110",
  48486=>"011100111",
  48487=>"101110111",
  48488=>"101110001",
  48489=>"000110011",
  48490=>"001111000",
  48491=>"101010101",
  48492=>"110111001",
  48493=>"110011110",
  48494=>"001001000",
  48495=>"111111101",
  48496=>"001110000",
  48497=>"111101110",
  48498=>"101010111",
  48499=>"100011111",
  48500=>"010010010",
  48501=>"000010011",
  48502=>"101100100",
  48503=>"100111101",
  48504=>"100000010",
  48505=>"100101011",
  48506=>"110000001",
  48507=>"001100100",
  48508=>"100000010",
  48509=>"100101100",
  48510=>"000011001",
  48511=>"011110110",
  48512=>"000110110",
  48513=>"000001100",
  48514=>"000111101",
  48515=>"001000010",
  48516=>"101000110",
  48517=>"000011010",
  48518=>"010110011",
  48519=>"101000100",
  48520=>"111000111",
  48521=>"010101110",
  48522=>"000011111",
  48523=>"010010000",
  48524=>"010100010",
  48525=>"000100100",
  48526=>"000000001",
  48527=>"001010010",
  48528=>"100001111",
  48529=>"100010010",
  48530=>"000010101",
  48531=>"001011011",
  48532=>"111100100",
  48533=>"010010111",
  48534=>"010001001",
  48535=>"101000000",
  48536=>"001100110",
  48537=>"001001001",
  48538=>"100001010",
  48539=>"111111000",
  48540=>"011011011",
  48541=>"101100110",
  48542=>"011111010",
  48543=>"000100001",
  48544=>"010110011",
  48545=>"111010110",
  48546=>"001100110",
  48547=>"111100111",
  48548=>"000001101",
  48549=>"110100110",
  48550=>"111101111",
  48551=>"010101011",
  48552=>"001011110",
  48553=>"100100101",
  48554=>"100110111",
  48555=>"010000100",
  48556=>"010010111",
  48557=>"011110101",
  48558=>"010100010",
  48559=>"101011011",
  48560=>"000001100",
  48561=>"110010011",
  48562=>"101011100",
  48563=>"100010011",
  48564=>"111101101",
  48565=>"100110010",
  48566=>"011111110",
  48567=>"010111110",
  48568=>"000100110",
  48569=>"100011100",
  48570=>"000001100",
  48571=>"010000100",
  48572=>"010111110",
  48573=>"111001011",
  48574=>"101001110",
  48575=>"100101000",
  48576=>"111000101",
  48577=>"010000110",
  48578=>"101110011",
  48579=>"001010010",
  48580=>"100001010",
  48581=>"011000000",
  48582=>"101100111",
  48583=>"101111000",
  48584=>"111011000",
  48585=>"111111011",
  48586=>"110111001",
  48587=>"110101110",
  48588=>"011000011",
  48589=>"000010101",
  48590=>"001111111",
  48591=>"001101011",
  48592=>"000111010",
  48593=>"000001000",
  48594=>"000011001",
  48595=>"100011010",
  48596=>"100001101",
  48597=>"011100101",
  48598=>"110001111",
  48599=>"011011010",
  48600=>"000101100",
  48601=>"101100011",
  48602=>"011000101",
  48603=>"111001010",
  48604=>"011111000",
  48605=>"111111010",
  48606=>"111001001",
  48607=>"111000011",
  48608=>"000011010",
  48609=>"111101111",
  48610=>"010000000",
  48611=>"101001110",
  48612=>"010101100",
  48613=>"011000101",
  48614=>"011111000",
  48615=>"101011110",
  48616=>"000010110",
  48617=>"000010111",
  48618=>"100001000",
  48619=>"100101010",
  48620=>"010001100",
  48621=>"100110010",
  48622=>"010110101",
  48623=>"100110100",
  48624=>"010110000",
  48625=>"111111011",
  48626=>"010101010",
  48627=>"011000111",
  48628=>"111100100",
  48629=>"101000001",
  48630=>"101110010",
  48631=>"100110011",
  48632=>"000110000",
  48633=>"000111010",
  48634=>"000010010",
  48635=>"011100100",
  48636=>"000010100",
  48637=>"111000110",
  48638=>"101001100",
  48639=>"000011001",
  48640=>"101001000",
  48641=>"011010010",
  48642=>"111011001",
  48643=>"010111011",
  48644=>"010000010",
  48645=>"001101001",
  48646=>"001111000",
  48647=>"010000011",
  48648=>"110100100",
  48649=>"011000101",
  48650=>"111101101",
  48651=>"010100100",
  48652=>"010100010",
  48653=>"011100110",
  48654=>"000010000",
  48655=>"101101000",
  48656=>"011010110",
  48657=>"010100011",
  48658=>"010101101",
  48659=>"001100010",
  48660=>"000110010",
  48661=>"001011100",
  48662=>"000111110",
  48663=>"101011011",
  48664=>"010101000",
  48665=>"100110001",
  48666=>"111111011",
  48667=>"000110101",
  48668=>"011111110",
  48669=>"001101110",
  48670=>"100000101",
  48671=>"010111011",
  48672=>"001000000",
  48673=>"100011100",
  48674=>"110000111",
  48675=>"001101010",
  48676=>"001000101",
  48677=>"010010110",
  48678=>"111110110",
  48679=>"100000110",
  48680=>"011111001",
  48681=>"000011001",
  48682=>"010111111",
  48683=>"000101101",
  48684=>"010001110",
  48685=>"010010101",
  48686=>"000101000",
  48687=>"011100001",
  48688=>"101110010",
  48689=>"101101110",
  48690=>"101000010",
  48691=>"001010111",
  48692=>"101110110",
  48693=>"100100000",
  48694=>"100010100",
  48695=>"000111011",
  48696=>"000111111",
  48697=>"000011111",
  48698=>"010100110",
  48699=>"111100101",
  48700=>"011000000",
  48701=>"001111001",
  48702=>"011000001",
  48703=>"000010011",
  48704=>"000000000",
  48705=>"011011110",
  48706=>"000111101",
  48707=>"010111110",
  48708=>"110100001",
  48709=>"000011111",
  48710=>"000100010",
  48711=>"111101010",
  48712=>"001000111",
  48713=>"101001101",
  48714=>"000101000",
  48715=>"011001100",
  48716=>"100110000",
  48717=>"000101010",
  48718=>"001010010",
  48719=>"111010110",
  48720=>"010010101",
  48721=>"111010001",
  48722=>"000010010",
  48723=>"111111000",
  48724=>"000001101",
  48725=>"110001101",
  48726=>"010010011",
  48727=>"100010110",
  48728=>"111100111",
  48729=>"110010100",
  48730=>"010100001",
  48731=>"000010010",
  48732=>"100110101",
  48733=>"101001000",
  48734=>"101110001",
  48735=>"011101101",
  48736=>"110001011",
  48737=>"010111001",
  48738=>"010010010",
  48739=>"100011010",
  48740=>"111101000",
  48741=>"011100011",
  48742=>"010001111",
  48743=>"111110011",
  48744=>"011011101",
  48745=>"110111001",
  48746=>"000110001",
  48747=>"010100110",
  48748=>"110011000",
  48749=>"111011010",
  48750=>"001011111",
  48751=>"010101100",
  48752=>"001110000",
  48753=>"001000110",
  48754=>"100011100",
  48755=>"101111101",
  48756=>"011110001",
  48757=>"110011110",
  48758=>"111101000",
  48759=>"100101010",
  48760=>"000100010",
  48761=>"100111010",
  48762=>"011010001",
  48763=>"011101001",
  48764=>"000011001",
  48765=>"000100001",
  48766=>"110101001",
  48767=>"010110001",
  48768=>"010000001",
  48769=>"100111001",
  48770=>"111110110",
  48771=>"000100010",
  48772=>"001100101",
  48773=>"100100100",
  48774=>"000101100",
  48775=>"010010011",
  48776=>"010000110",
  48777=>"100101001",
  48778=>"100000011",
  48779=>"111110101",
  48780=>"101000101",
  48781=>"100100100",
  48782=>"101100000",
  48783=>"110010001",
  48784=>"100111101",
  48785=>"101100011",
  48786=>"101111010",
  48787=>"111001110",
  48788=>"101101101",
  48789=>"000011111",
  48790=>"000111000",
  48791=>"111100011",
  48792=>"110101111",
  48793=>"100010001",
  48794=>"110001011",
  48795=>"011111000",
  48796=>"001110110",
  48797=>"001000010",
  48798=>"010000101",
  48799=>"111111111",
  48800=>"100110011",
  48801=>"100000110",
  48802=>"100100111",
  48803=>"000101000",
  48804=>"110010001",
  48805=>"010101111",
  48806=>"111110111",
  48807=>"000000100",
  48808=>"001110010",
  48809=>"000001111",
  48810=>"000110101",
  48811=>"110010111",
  48812=>"010001001",
  48813=>"110001010",
  48814=>"111000001",
  48815=>"101101111",
  48816=>"001101011",
  48817=>"001110001",
  48818=>"001000110",
  48819=>"011010111",
  48820=>"101001000",
  48821=>"111000000",
  48822=>"001111101",
  48823=>"010011000",
  48824=>"001100010",
  48825=>"001000000",
  48826=>"110110111",
  48827=>"101110011",
  48828=>"110000001",
  48829=>"110111100",
  48830=>"100111100",
  48831=>"010110100",
  48832=>"001001011",
  48833=>"100000100",
  48834=>"011011010",
  48835=>"011110010",
  48836=>"100011000",
  48837=>"100110010",
  48838=>"111001110",
  48839=>"100110110",
  48840=>"101001111",
  48841=>"100101100",
  48842=>"001100111",
  48843=>"111101101",
  48844=>"010101101",
  48845=>"100011101",
  48846=>"100100001",
  48847=>"100110011",
  48848=>"100101010",
  48849=>"000000011",
  48850=>"011010001",
  48851=>"010011000",
  48852=>"100001000",
  48853=>"111110010",
  48854=>"001010011",
  48855=>"110111011",
  48856=>"000111011",
  48857=>"111110011",
  48858=>"001000100",
  48859=>"100100000",
  48860=>"000100110",
  48861=>"100011011",
  48862=>"010101111",
  48863=>"001100000",
  48864=>"010110110",
  48865=>"100000110",
  48866=>"010010100",
  48867=>"011100111",
  48868=>"011001100",
  48869=>"101010110",
  48870=>"110011101",
  48871=>"001000111",
  48872=>"100100001",
  48873=>"001001000",
  48874=>"000011011",
  48875=>"100001010",
  48876=>"001111011",
  48877=>"100011100",
  48878=>"000000101",
  48879=>"010001100",
  48880=>"100001001",
  48881=>"001100110",
  48882=>"001100011",
  48883=>"111010101",
  48884=>"111000011",
  48885=>"110111111",
  48886=>"111110100",
  48887=>"110001001",
  48888=>"001110110",
  48889=>"101100011",
  48890=>"101110101",
  48891=>"000000000",
  48892=>"011000100",
  48893=>"100110010",
  48894=>"101011000",
  48895=>"000000010",
  48896=>"011101111",
  48897=>"000111000",
  48898=>"111111100",
  48899=>"000101011",
  48900=>"111000010",
  48901=>"100000100",
  48902=>"101000011",
  48903=>"111100100",
  48904=>"101101000",
  48905=>"000100101",
  48906=>"110000101",
  48907=>"010110010",
  48908=>"011100001",
  48909=>"101100111",
  48910=>"001101001",
  48911=>"000101111",
  48912=>"100111000",
  48913=>"100000000",
  48914=>"010101100",
  48915=>"110000110",
  48916=>"101111111",
  48917=>"010101001",
  48918=>"111011001",
  48919=>"011001110",
  48920=>"100100110",
  48921=>"000000000",
  48922=>"100111010",
  48923=>"010100001",
  48924=>"000011110",
  48925=>"000011110",
  48926=>"000101000",
  48927=>"101000000",
  48928=>"110000010",
  48929=>"101001010",
  48930=>"010111101",
  48931=>"001001001",
  48932=>"111100110",
  48933=>"010101101",
  48934=>"111011101",
  48935=>"111100001",
  48936=>"000011000",
  48937=>"000000100",
  48938=>"100010000",
  48939=>"100010101",
  48940=>"110100000",
  48941=>"000010100",
  48942=>"110010101",
  48943=>"100110010",
  48944=>"111101001",
  48945=>"101111000",
  48946=>"011011001",
  48947=>"010101110",
  48948=>"101111011",
  48949=>"111001000",
  48950=>"011110111",
  48951=>"110111101",
  48952=>"100100110",
  48953=>"011111000",
  48954=>"101010111",
  48955=>"101000000",
  48956=>"111101100",
  48957=>"001101111",
  48958=>"111111111",
  48959=>"001010011",
  48960=>"001100100",
  48961=>"011011010",
  48962=>"011001101",
  48963=>"010111111",
  48964=>"101110000",
  48965=>"001110010",
  48966=>"110010111",
  48967=>"110001010",
  48968=>"100110001",
  48969=>"111111001",
  48970=>"110001101",
  48971=>"010101010",
  48972=>"001110010",
  48973=>"000110000",
  48974=>"111100010",
  48975=>"110111010",
  48976=>"110111010",
  48977=>"110101001",
  48978=>"100100000",
  48979=>"000011000",
  48980=>"010001110",
  48981=>"100111011",
  48982=>"111111110",
  48983=>"101101011",
  48984=>"011001000",
  48985=>"110001000",
  48986=>"101110111",
  48987=>"000001111",
  48988=>"010111001",
  48989=>"100001011",
  48990=>"100001101",
  48991=>"010000001",
  48992=>"100101011",
  48993=>"010100010",
  48994=>"101001100",
  48995=>"000110101",
  48996=>"110000010",
  48997=>"101010101",
  48998=>"101101101",
  48999=>"000111011",
  49000=>"101110110",
  49001=>"111100111",
  49002=>"011010110",
  49003=>"001010010",
  49004=>"000001110",
  49005=>"100101000",
  49006=>"001011011",
  49007=>"111010010",
  49008=>"011100111",
  49009=>"000011100",
  49010=>"111010010",
  49011=>"000011001",
  49012=>"010000001",
  49013=>"100100101",
  49014=>"000010101",
  49015=>"111111110",
  49016=>"101010011",
  49017=>"010011001",
  49018=>"001111110",
  49019=>"111101011",
  49020=>"000000000",
  49021=>"010110110",
  49022=>"010011000",
  49023=>"101111011",
  49024=>"001100000",
  49025=>"111001011",
  49026=>"011011101",
  49027=>"111001010",
  49028=>"100111000",
  49029=>"001101000",
  49030=>"011110010",
  49031=>"100010010",
  49032=>"000001100",
  49033=>"001110000",
  49034=>"000000000",
  49035=>"110110111",
  49036=>"100111000",
  49037=>"011111010",
  49038=>"100001000",
  49039=>"011101010",
  49040=>"010001000",
  49041=>"001001101",
  49042=>"000011000",
  49043=>"100110100",
  49044=>"000001110",
  49045=>"000011000",
  49046=>"101000011",
  49047=>"001110001",
  49048=>"110111010",
  49049=>"101011101",
  49050=>"111110001",
  49051=>"101001101",
  49052=>"101001101",
  49053=>"101110000",
  49054=>"011000000",
  49055=>"100111000",
  49056=>"110101001",
  49057=>"100011110",
  49058=>"110010100",
  49059=>"101100110",
  49060=>"000101110",
  49061=>"110000111",
  49062=>"001100000",
  49063=>"010010000",
  49064=>"001000000",
  49065=>"101110110",
  49066=>"110001000",
  49067=>"111001111",
  49068=>"100000110",
  49069=>"111010000",
  49070=>"101101001",
  49071=>"111010010",
  49072=>"111111110",
  49073=>"010111001",
  49074=>"001001100",
  49075=>"110000100",
  49076=>"101101010",
  49077=>"101111110",
  49078=>"111010111",
  49079=>"010011011",
  49080=>"111001100",
  49081=>"100111111",
  49082=>"110100101",
  49083=>"001100001",
  49084=>"100010110",
  49085=>"100000110",
  49086=>"010101000",
  49087=>"000100000",
  49088=>"101100111",
  49089=>"010010111",
  49090=>"000101010",
  49091=>"010101001",
  49092=>"000101000",
  49093=>"000111011",
  49094=>"011010001",
  49095=>"010010111",
  49096=>"010110000",
  49097=>"111010100",
  49098=>"011010010",
  49099=>"101111110",
  49100=>"011001111",
  49101=>"011000101",
  49102=>"010001010",
  49103=>"110101000",
  49104=>"010111101",
  49105=>"111110100",
  49106=>"000010100",
  49107=>"111000001",
  49108=>"110011001",
  49109=>"010110111",
  49110=>"100011111",
  49111=>"101101110",
  49112=>"111101111",
  49113=>"100101101",
  49114=>"111011101",
  49115=>"000010111",
  49116=>"001000110",
  49117=>"000110011",
  49118=>"010110000",
  49119=>"111100110",
  49120=>"111000110",
  49121=>"111110100",
  49122=>"011100111",
  49123=>"101111101",
  49124=>"111010010",
  49125=>"101010100",
  49126=>"101011011",
  49127=>"111100101",
  49128=>"001101011",
  49129=>"100000110",
  49130=>"111111000",
  49131=>"001101010",
  49132=>"100010011",
  49133=>"011011000",
  49134=>"101100101",
  49135=>"100111011",
  49136=>"100010010",
  49137=>"100111111",
  49138=>"100000110",
  49139=>"100010111",
  49140=>"000011010",
  49141=>"100100110",
  49142=>"000000101",
  49143=>"001101011",
  49144=>"110011110",
  49145=>"010001011",
  49146=>"110010101",
  49147=>"110000110",
  49148=>"011001101",
  49149=>"010000101",
  49150=>"000111110",
  49151=>"110110110",
  49152=>"000011110",
  49153=>"110010010",
  49154=>"001010110",
  49155=>"000101001",
  49156=>"001010000",
  49157=>"111111100",
  49158=>"010111001",
  49159=>"000100010",
  49160=>"100100010",
  49161=>"010100011",
  49162=>"100101100",
  49163=>"011000110",
  49164=>"100111110",
  49165=>"001101100",
  49166=>"001000011",
  49167=>"010101100",
  49168=>"101100100",
  49169=>"101101010",
  49170=>"001011100",
  49171=>"000010011",
  49172=>"001111010",
  49173=>"011010001",
  49174=>"110110010",
  49175=>"101010100",
  49176=>"111110110",
  49177=>"000001001",
  49178=>"010001000",
  49179=>"001010100",
  49180=>"011010001",
  49181=>"001000011",
  49182=>"011011001",
  49183=>"101100110",
  49184=>"110110001",
  49185=>"101010000",
  49186=>"100111011",
  49187=>"100010100",
  49188=>"100101000",
  49189=>"100101011",
  49190=>"100101000",
  49191=>"110101000",
  49192=>"110101010",
  49193=>"101000100",
  49194=>"100111010",
  49195=>"111011101",
  49196=>"111101011",
  49197=>"111110110",
  49198=>"100011010",
  49199=>"101010101",
  49200=>"000001001",
  49201=>"111001010",
  49202=>"100011101",
  49203=>"000111001",
  49204=>"010001100",
  49205=>"110000010",
  49206=>"111010011",
  49207=>"100001111",
  49208=>"000001000",
  49209=>"111100000",
  49210=>"000000001",
  49211=>"000011001",
  49212=>"000001010",
  49213=>"000111001",
  49214=>"011010100",
  49215=>"100111111",
  49216=>"111101000",
  49217=>"100010000",
  49218=>"010111100",
  49219=>"010001100",
  49220=>"000111101",
  49221=>"001000001",
  49222=>"111001000",
  49223=>"100011101",
  49224=>"000000111",
  49225=>"011011010",
  49226=>"111011111",
  49227=>"111001000",
  49228=>"111011010",
  49229=>"101010110",
  49230=>"100001101",
  49231=>"111011100",
  49232=>"000000000",
  49233=>"111110111",
  49234=>"000100111",
  49235=>"011111101",
  49236=>"100111110",
  49237=>"111000001",
  49238=>"011110000",
  49239=>"011011011",
  49240=>"010000100",
  49241=>"111100001",
  49242=>"000010111",
  49243=>"101000111",
  49244=>"100000011",
  49245=>"101110101",
  49246=>"101110001",
  49247=>"100011001",
  49248=>"111110001",
  49249=>"111101111",
  49250=>"010010100",
  49251=>"000000011",
  49252=>"011000001",
  49253=>"011101100",
  49254=>"110001101",
  49255=>"111010001",
  49256=>"000001111",
  49257=>"010010110",
  49258=>"001100000",
  49259=>"111101101",
  49260=>"001010010",
  49261=>"010110111",
  49262=>"010111000",
  49263=>"001000011",
  49264=>"010100111",
  49265=>"000110101",
  49266=>"111100011",
  49267=>"010010100",
  49268=>"100001111",
  49269=>"011000100",
  49270=>"010100001",
  49271=>"010010010",
  49272=>"000100001",
  49273=>"101001001",
  49274=>"011001000",
  49275=>"010111101",
  49276=>"010111001",
  49277=>"101111011",
  49278=>"100111000",
  49279=>"101100010",
  49280=>"001000111",
  49281=>"101111101",
  49282=>"001101001",
  49283=>"100110011",
  49284=>"100000011",
  49285=>"010101001",
  49286=>"111001101",
  49287=>"111001010",
  49288=>"100001101",
  49289=>"000010100",
  49290=>"111000011",
  49291=>"101010000",
  49292=>"111101101",
  49293=>"001100010",
  49294=>"001000001",
  49295=>"010110000",
  49296=>"111111010",
  49297=>"101111100",
  49298=>"101101000",
  49299=>"001001111",
  49300=>"001101111",
  49301=>"001001000",
  49302=>"100001011",
  49303=>"111101011",
  49304=>"011110101",
  49305=>"010100011",
  49306=>"001011101",
  49307=>"111110010",
  49308=>"101000001",
  49309=>"011110000",
  49310=>"010100000",
  49311=>"111001101",
  49312=>"101100110",
  49313=>"101100001",
  49314=>"010110010",
  49315=>"000101111",
  49316=>"000001001",
  49317=>"100111100",
  49318=>"111111011",
  49319=>"100000100",
  49320=>"100101111",
  49321=>"001101000",
  49322=>"001001010",
  49323=>"010001111",
  49324=>"101010000",
  49325=>"011100010",
  49326=>"110101010",
  49327=>"111100001",
  49328=>"000110111",
  49329=>"000110100",
  49330=>"111100101",
  49331=>"111100000",
  49332=>"011010110",
  49333=>"011111000",
  49334=>"100000000",
  49335=>"101100110",
  49336=>"100100011",
  49337=>"110110111",
  49338=>"100011111",
  49339=>"000010010",
  49340=>"100110011",
  49341=>"001011011",
  49342=>"111101111",
  49343=>"011101101",
  49344=>"100111000",
  49345=>"000101011",
  49346=>"001101000",
  49347=>"111011010",
  49348=>"011001100",
  49349=>"101010111",
  49350=>"011101011",
  49351=>"000100011",
  49352=>"011010111",
  49353=>"110000001",
  49354=>"101101110",
  49355=>"100001101",
  49356=>"001110000",
  49357=>"101101010",
  49358=>"000000111",
  49359=>"101001101",
  49360=>"111000111",
  49361=>"010101111",
  49362=>"001110010",
  49363=>"101101111",
  49364=>"101101101",
  49365=>"000110101",
  49366=>"111011100",
  49367=>"010011000",
  49368=>"000101000",
  49369=>"000000001",
  49370=>"000111010",
  49371=>"101111000",
  49372=>"010111010",
  49373=>"001010011",
  49374=>"111010011",
  49375=>"101000010",
  49376=>"011000100",
  49377=>"110110111",
  49378=>"111111010",
  49379=>"111101000",
  49380=>"011000000",
  49381=>"111001101",
  49382=>"100111111",
  49383=>"100001010",
  49384=>"100011110",
  49385=>"110100000",
  49386=>"100101001",
  49387=>"101100010",
  49388=>"111111011",
  49389=>"110000000",
  49390=>"000000111",
  49391=>"010010000",
  49392=>"110011000",
  49393=>"111001101",
  49394=>"101001111",
  49395=>"010000011",
  49396=>"001110001",
  49397=>"010110011",
  49398=>"010101000",
  49399=>"001111001",
  49400=>"111010001",
  49401=>"000000100",
  49402=>"101111000",
  49403=>"000101001",
  49404=>"011001110",
  49405=>"000011100",
  49406=>"001110011",
  49407=>"000110111",
  49408=>"110011001",
  49409=>"011100000",
  49410=>"100010010",
  49411=>"101101000",
  49412=>"110100111",
  49413=>"101110101",
  49414=>"011001011",
  49415=>"100011001",
  49416=>"010101101",
  49417=>"000001110",
  49418=>"110110110",
  49419=>"100100001",
  49420=>"110000011",
  49421=>"010010000",
  49422=>"001100011",
  49423=>"000000010",
  49424=>"000100011",
  49425=>"010001011",
  49426=>"000001100",
  49427=>"110000100",
  49428=>"000011010",
  49429=>"000011000",
  49430=>"111010100",
  49431=>"001000001",
  49432=>"001000111",
  49433=>"110111000",
  49434=>"101101110",
  49435=>"001011000",
  49436=>"001011110",
  49437=>"000100111",
  49438=>"100011111",
  49439=>"100100111",
  49440=>"010000101",
  49441=>"010010011",
  49442=>"011101000",
  49443=>"011011111",
  49444=>"111011111",
  49445=>"000000100",
  49446=>"100011000",
  49447=>"110100110",
  49448=>"001110010",
  49449=>"011101011",
  49450=>"010110110",
  49451=>"001010001",
  49452=>"010000111",
  49453=>"110010111",
  49454=>"000001010",
  49455=>"110111101",
  49456=>"001111111",
  49457=>"100101110",
  49458=>"011010000",
  49459=>"000100010",
  49460=>"111000000",
  49461=>"111111101",
  49462=>"011000110",
  49463=>"001000011",
  49464=>"001101100",
  49465=>"011010001",
  49466=>"111011101",
  49467=>"100000000",
  49468=>"011001100",
  49469=>"110010110",
  49470=>"110101001",
  49471=>"011111101",
  49472=>"000110011",
  49473=>"011010100",
  49474=>"111000110",
  49475=>"110011111",
  49476=>"110101010",
  49477=>"101001101",
  49478=>"000010000",
  49479=>"111111011",
  49480=>"110010111",
  49481=>"111001011",
  49482=>"011011100",
  49483=>"001001001",
  49484=>"100110001",
  49485=>"000110001",
  49486=>"000111111",
  49487=>"100110000",
  49488=>"111000101",
  49489=>"110100110",
  49490=>"101111111",
  49491=>"000100000",
  49492=>"000010100",
  49493=>"010101110",
  49494=>"010100011",
  49495=>"101110110",
  49496=>"111100110",
  49497=>"000101111",
  49498=>"001111110",
  49499=>"100111000",
  49500=>"111101011",
  49501=>"111110001",
  49502=>"000010000",
  49503=>"000010010",
  49504=>"001110100",
  49505=>"111111101",
  49506=>"011001111",
  49507=>"001001001",
  49508=>"101110000",
  49509=>"000100000",
  49510=>"100000110",
  49511=>"011101100",
  49512=>"011111110",
  49513=>"011011000",
  49514=>"011100001",
  49515=>"000001011",
  49516=>"010010001",
  49517=>"001001010",
  49518=>"101101111",
  49519=>"011001001",
  49520=>"101100010",
  49521=>"010110011",
  49522=>"101110100",
  49523=>"011100011",
  49524=>"000101111",
  49525=>"111100000",
  49526=>"010011110",
  49527=>"010100010",
  49528=>"101101010",
  49529=>"100010010",
  49530=>"001110010",
  49531=>"101000011",
  49532=>"101101000",
  49533=>"010001011",
  49534=>"100111101",
  49535=>"000011110",
  49536=>"000101011",
  49537=>"111111111",
  49538=>"011001101",
  49539=>"001010111",
  49540=>"011001110",
  49541=>"010010110",
  49542=>"101011100",
  49543=>"011000000",
  49544=>"000101001",
  49545=>"101110100",
  49546=>"001100111",
  49547=>"001011000",
  49548=>"001110110",
  49549=>"101011100",
  49550=>"011011100",
  49551=>"000011000",
  49552=>"000010111",
  49553=>"100001111",
  49554=>"001000111",
  49555=>"100100010",
  49556=>"110101111",
  49557=>"000001010",
  49558=>"111100001",
  49559=>"100110000",
  49560=>"001111011",
  49561=>"101101100",
  49562=>"100010000",
  49563=>"110001000",
  49564=>"100000111",
  49565=>"111100111",
  49566=>"000000101",
  49567=>"111110101",
  49568=>"110100100",
  49569=>"100001111",
  49570=>"110000010",
  49571=>"001101010",
  49572=>"011110101",
  49573=>"111010000",
  49574=>"110111011",
  49575=>"111110100",
  49576=>"100101011",
  49577=>"011100101",
  49578=>"001000101",
  49579=>"110100101",
  49580=>"101000001",
  49581=>"001000000",
  49582=>"100110101",
  49583=>"001001010",
  49584=>"111101000",
  49585=>"010000110",
  49586=>"111010010",
  49587=>"111100011",
  49588=>"101010101",
  49589=>"100010100",
  49590=>"110011000",
  49591=>"110110011",
  49592=>"100000100",
  49593=>"100111001",
  49594=>"000101000",
  49595=>"011000000",
  49596=>"110010110",
  49597=>"111110101",
  49598=>"000100000",
  49599=>"101111000",
  49600=>"110110001",
  49601=>"110010100",
  49602=>"001010001",
  49603=>"100010111",
  49604=>"101010000",
  49605=>"011110001",
  49606=>"110110110",
  49607=>"000000001",
  49608=>"101001011",
  49609=>"000001010",
  49610=>"011110000",
  49611=>"100100101",
  49612=>"100011111",
  49613=>"001111001",
  49614=>"100000010",
  49615=>"111000110",
  49616=>"101010101",
  49617=>"010111011",
  49618=>"110000110",
  49619=>"001010011",
  49620=>"000111111",
  49621=>"010111011",
  49622=>"000001000",
  49623=>"111010011",
  49624=>"011010111",
  49625=>"000010101",
  49626=>"010101000",
  49627=>"111110000",
  49628=>"100110101",
  49629=>"011101111",
  49630=>"001111011",
  49631=>"011111101",
  49632=>"001101111",
  49633=>"011001111",
  49634=>"111001000",
  49635=>"111110010",
  49636=>"011100101",
  49637=>"100110011",
  49638=>"111010110",
  49639=>"010111111",
  49640=>"011100011",
  49641=>"011111010",
  49642=>"111011011",
  49643=>"001010100",
  49644=>"100010001",
  49645=>"101000000",
  49646=>"011110011",
  49647=>"110111010",
  49648=>"011101110",
  49649=>"001001111",
  49650=>"000110011",
  49651=>"010101000",
  49652=>"010010110",
  49653=>"110011111",
  49654=>"000000110",
  49655=>"010110100",
  49656=>"111001000",
  49657=>"110001101",
  49658=>"001100010",
  49659=>"011010010",
  49660=>"111001110",
  49661=>"001011000",
  49662=>"111011110",
  49663=>"100010001",
  49664=>"100101001",
  49665=>"010011010",
  49666=>"110100010",
  49667=>"111011000",
  49668=>"111011010",
  49669=>"011010111",
  49670=>"010100001",
  49671=>"001000010",
  49672=>"000000001",
  49673=>"010111001",
  49674=>"011110001",
  49675=>"100101100",
  49676=>"100110110",
  49677=>"000011001",
  49678=>"111000111",
  49679=>"000100010",
  49680=>"011000100",
  49681=>"111111011",
  49682=>"000001010",
  49683=>"100101111",
  49684=>"111100001",
  49685=>"110110000",
  49686=>"110010001",
  49687=>"011110000",
  49688=>"101010010",
  49689=>"000111011",
  49690=>"010010111",
  49691=>"110001111",
  49692=>"110101010",
  49693=>"010111111",
  49694=>"111111011",
  49695=>"100001001",
  49696=>"011001111",
  49697=>"011010101",
  49698=>"010101010",
  49699=>"101100101",
  49700=>"010000110",
  49701=>"000100101",
  49702=>"001101100",
  49703=>"111000101",
  49704=>"000000001",
  49705=>"011000010",
  49706=>"000000110",
  49707=>"011110101",
  49708=>"000111110",
  49709=>"100101011",
  49710=>"000111100",
  49711=>"100011010",
  49712=>"000000101",
  49713=>"000101100",
  49714=>"010111010",
  49715=>"111110100",
  49716=>"000100010",
  49717=>"110111100",
  49718=>"100101111",
  49719=>"010010010",
  49720=>"011000001",
  49721=>"000110000",
  49722=>"000111101",
  49723=>"100100111",
  49724=>"111101100",
  49725=>"000001100",
  49726=>"010011101",
  49727=>"100110111",
  49728=>"001111110",
  49729=>"101100001",
  49730=>"100000110",
  49731=>"001100001",
  49732=>"010100000",
  49733=>"001001111",
  49734=>"011101011",
  49735=>"001011111",
  49736=>"011000011",
  49737=>"110100010",
  49738=>"000011011",
  49739=>"010100011",
  49740=>"010110011",
  49741=>"110100000",
  49742=>"100101110",
  49743=>"111111000",
  49744=>"111101110",
  49745=>"010000111",
  49746=>"111111111",
  49747=>"000111100",
  49748=>"111100000",
  49749=>"100011000",
  49750=>"000000000",
  49751=>"011011001",
  49752=>"000110101",
  49753=>"100010001",
  49754=>"110000001",
  49755=>"010110100",
  49756=>"001000010",
  49757=>"110100110",
  49758=>"100110101",
  49759=>"000001000",
  49760=>"011111000",
  49761=>"101000011",
  49762=>"100111111",
  49763=>"100000100",
  49764=>"001010010",
  49765=>"111110111",
  49766=>"100000101",
  49767=>"000000100",
  49768=>"100001010",
  49769=>"111110010",
  49770=>"101101110",
  49771=>"010111110",
  49772=>"110101110",
  49773=>"111010101",
  49774=>"110011001",
  49775=>"000110110",
  49776=>"000000011",
  49777=>"011000000",
  49778=>"011111001",
  49779=>"110111110",
  49780=>"110011010",
  49781=>"000110110",
  49782=>"111000110",
  49783=>"001101101",
  49784=>"001011110",
  49785=>"001001101",
  49786=>"010000111",
  49787=>"000010110",
  49788=>"110011000",
  49789=>"101000101",
  49790=>"001111111",
  49791=>"010110010",
  49792=>"001011100",
  49793=>"011111010",
  49794=>"000000001",
  49795=>"101001110",
  49796=>"100110010",
  49797=>"001100111",
  49798=>"101101010",
  49799=>"110001100",
  49800=>"111111101",
  49801=>"000010111",
  49802=>"110011000",
  49803=>"110111111",
  49804=>"101111101",
  49805=>"000100100",
  49806=>"110101101",
  49807=>"110000010",
  49808=>"111101010",
  49809=>"110110000",
  49810=>"001110101",
  49811=>"101101011",
  49812=>"000010010",
  49813=>"110111000",
  49814=>"001111111",
  49815=>"011111001",
  49816=>"100110010",
  49817=>"101001001",
  49818=>"110111011",
  49819=>"100011111",
  49820=>"101100111",
  49821=>"010010000",
  49822=>"101101111",
  49823=>"001001001",
  49824=>"011010101",
  49825=>"101111110",
  49826=>"011000111",
  49827=>"001101000",
  49828=>"010001101",
  49829=>"111101101",
  49830=>"100011001",
  49831=>"110000101",
  49832=>"001001001",
  49833=>"110110101",
  49834=>"100101010",
  49835=>"001101100",
  49836=>"010010001",
  49837=>"000010101",
  49838=>"010010111",
  49839=>"101010010",
  49840=>"011001000",
  49841=>"010100110",
  49842=>"010101100",
  49843=>"000101011",
  49844=>"010111110",
  49845=>"011100111",
  49846=>"000010011",
  49847=>"000001011",
  49848=>"011010010",
  49849=>"101110101",
  49850=>"111101101",
  49851=>"111001111",
  49852=>"000101110",
  49853=>"000001110",
  49854=>"110100101",
  49855=>"111110100",
  49856=>"011111100",
  49857=>"110111001",
  49858=>"110011000",
  49859=>"011010101",
  49860=>"111101110",
  49861=>"111001100",
  49862=>"110111111",
  49863=>"001101101",
  49864=>"110000000",
  49865=>"111100111",
  49866=>"110011000",
  49867=>"100000011",
  49868=>"011100011",
  49869=>"000001110",
  49870=>"101100010",
  49871=>"001010111",
  49872=>"000111010",
  49873=>"101000100",
  49874=>"001010010",
  49875=>"110100000",
  49876=>"001000000",
  49877=>"001101011",
  49878=>"111010010",
  49879=>"010010000",
  49880=>"010101011",
  49881=>"010110010",
  49882=>"011101110",
  49883=>"010000010",
  49884=>"101101010",
  49885=>"101111101",
  49886=>"010000111",
  49887=>"010010000",
  49888=>"110001000",
  49889=>"110010001",
  49890=>"000000111",
  49891=>"010001000",
  49892=>"100001010",
  49893=>"111001101",
  49894=>"010011010",
  49895=>"011010011",
  49896=>"110010010",
  49897=>"100110010",
  49898=>"101000001",
  49899=>"101000000",
  49900=>"000000000",
  49901=>"001000000",
  49902=>"100010100",
  49903=>"010010111",
  49904=>"101010010",
  49905=>"010011101",
  49906=>"101001110",
  49907=>"000100111",
  49908=>"111111000",
  49909=>"110100101",
  49910=>"011111010",
  49911=>"011011111",
  49912=>"011110001",
  49913=>"110001110",
  49914=>"100000011",
  49915=>"100001011",
  49916=>"001011001",
  49917=>"001110101",
  49918=>"000101111",
  49919=>"111000001",
  49920=>"111111011",
  49921=>"000101000",
  49922=>"011100100",
  49923=>"110111101",
  49924=>"001010011",
  49925=>"001000100",
  49926=>"111010001",
  49927=>"110111011",
  49928=>"101001001",
  49929=>"101101111",
  49930=>"111111000",
  49931=>"101111000",
  49932=>"110100001",
  49933=>"010110100",
  49934=>"000000000",
  49935=>"011000111",
  49936=>"000001101",
  49937=>"011000000",
  49938=>"111000111",
  49939=>"010111001",
  49940=>"010100000",
  49941=>"010110010",
  49942=>"111010010",
  49943=>"000000010",
  49944=>"111111100",
  49945=>"101011001",
  49946=>"011111111",
  49947=>"100010101",
  49948=>"000000000",
  49949=>"001110000",
  49950=>"000110001",
  49951=>"110000100",
  49952=>"000010100",
  49953=>"001001011",
  49954=>"000000010",
  49955=>"101101011",
  49956=>"110100001",
  49957=>"110001100",
  49958=>"011100111",
  49959=>"001011011",
  49960=>"110011100",
  49961=>"011000001",
  49962=>"011001001",
  49963=>"110000111",
  49964=>"000110110",
  49965=>"000110110",
  49966=>"001111101",
  49967=>"000011010",
  49968=>"101111100",
  49969=>"100010100",
  49970=>"000110010",
  49971=>"011101111",
  49972=>"111111111",
  49973=>"101100001",
  49974=>"100000110",
  49975=>"110001110",
  49976=>"101000001",
  49977=>"111000111",
  49978=>"101000001",
  49979=>"111010111",
  49980=>"000111110",
  49981=>"101001101",
  49982=>"001000000",
  49983=>"110010011",
  49984=>"110010110",
  49985=>"011100101",
  49986=>"010101100",
  49987=>"100000100",
  49988=>"000111000",
  49989=>"101010101",
  49990=>"011111100",
  49991=>"111100011",
  49992=>"000011000",
  49993=>"010100000",
  49994=>"100110010",
  49995=>"111000111",
  49996=>"000010110",
  49997=>"101111000",
  49998=>"010000010",
  49999=>"000001011",
  50000=>"101001111",
  50001=>"000101010",
  50002=>"000111111",
  50003=>"110011101",
  50004=>"110101100",
  50005=>"100110111",
  50006=>"000010000",
  50007=>"100011101",
  50008=>"010000001",
  50009=>"100001001",
  50010=>"011001011",
  50011=>"000001010",
  50012=>"000011100",
  50013=>"011010101",
  50014=>"110111110",
  50015=>"000000110",
  50016=>"101110011",
  50017=>"001000100",
  50018=>"010100111",
  50019=>"011001011",
  50020=>"010001000",
  50021=>"110100010",
  50022=>"001010101",
  50023=>"000011111",
  50024=>"101111011",
  50025=>"010001100",
  50026=>"000110100",
  50027=>"111000010",
  50028=>"101001111",
  50029=>"000010000",
  50030=>"100110111",
  50031=>"010010000",
  50032=>"111100100",
  50033=>"010111100",
  50034=>"100000011",
  50035=>"000001100",
  50036=>"001000110",
  50037=>"000111010",
  50038=>"000011010",
  50039=>"000010111",
  50040=>"011110011",
  50041=>"011001110",
  50042=>"011100110",
  50043=>"011101011",
  50044=>"011011100",
  50045=>"010101110",
  50046=>"010111101",
  50047=>"111111011",
  50048=>"111011011",
  50049=>"011111110",
  50050=>"001001110",
  50051=>"101000000",
  50052=>"110011001",
  50053=>"110101101",
  50054=>"001010100",
  50055=>"000010101",
  50056=>"000110110",
  50057=>"000000010",
  50058=>"001111101",
  50059=>"110101010",
  50060=>"010001110",
  50061=>"011111100",
  50062=>"100110010",
  50063=>"100001111",
  50064=>"000100110",
  50065=>"010010110",
  50066=>"111000011",
  50067=>"100100101",
  50068=>"110111111",
  50069=>"001000101",
  50070=>"110010011",
  50071=>"011100000",
  50072=>"011111100",
  50073=>"000111110",
  50074=>"101011000",
  50075=>"110011111",
  50076=>"110110001",
  50077=>"001101011",
  50078=>"100111101",
  50079=>"110101010",
  50080=>"011010000",
  50081=>"010100100",
  50082=>"000001101",
  50083=>"000000010",
  50084=>"000001100",
  50085=>"011011000",
  50086=>"000111000",
  50087=>"000000000",
  50088=>"000101111",
  50089=>"011111011",
  50090=>"111000111",
  50091=>"100000111",
  50092=>"000000011",
  50093=>"101111111",
  50094=>"000010101",
  50095=>"011000110",
  50096=>"100010100",
  50097=>"011100110",
  50098=>"000111110",
  50099=>"110100111",
  50100=>"000011101",
  50101=>"011000001",
  50102=>"011000100",
  50103=>"111011100",
  50104=>"111100101",
  50105=>"111110111",
  50106=>"001111001",
  50107=>"001111001",
  50108=>"000011111",
  50109=>"101111111",
  50110=>"000010110",
  50111=>"000011001",
  50112=>"111001000",
  50113=>"011100101",
  50114=>"001111101",
  50115=>"000111001",
  50116=>"011110101",
  50117=>"000010101",
  50118=>"111001110",
  50119=>"010100100",
  50120=>"001001111",
  50121=>"100110110",
  50122=>"000100001",
  50123=>"000010100",
  50124=>"100100111",
  50125=>"011001110",
  50126=>"001000010",
  50127=>"111011001",
  50128=>"101001111",
  50129=>"110110111",
  50130=>"101010100",
  50131=>"110000001",
  50132=>"100010111",
  50133=>"101101100",
  50134=>"101110001",
  50135=>"101010111",
  50136=>"000100001",
  50137=>"110010010",
  50138=>"010100110",
  50139=>"100011111",
  50140=>"000111000",
  50141=>"101111110",
  50142=>"000100100",
  50143=>"000000000",
  50144=>"000101111",
  50145=>"000001111",
  50146=>"010011100",
  50147=>"101010100",
  50148=>"011001111",
  50149=>"000000100",
  50150=>"100101000",
  50151=>"010100100",
  50152=>"011110010",
  50153=>"111111001",
  50154=>"111100011",
  50155=>"001000000",
  50156=>"110101100",
  50157=>"110001010",
  50158=>"011110111",
  50159=>"111100101",
  50160=>"000111011",
  50161=>"011001001",
  50162=>"001101101",
  50163=>"000000001",
  50164=>"010000010",
  50165=>"111000001",
  50166=>"110110001",
  50167=>"000000000",
  50168=>"001000101",
  50169=>"101101100",
  50170=>"000100100",
  50171=>"111111110",
  50172=>"100101001",
  50173=>"101001100",
  50174=>"111010100",
  50175=>"011000000",
  50176=>"011101111",
  50177=>"101101100",
  50178=>"001000101",
  50179=>"011110011",
  50180=>"100001011",
  50181=>"100000111",
  50182=>"011011101",
  50183=>"000111101",
  50184=>"000001000",
  50185=>"101000100",
  50186=>"010010000",
  50187=>"001111001",
  50188=>"011110111",
  50189=>"011001100",
  50190=>"011110010",
  50191=>"001111110",
  50192=>"111111101",
  50193=>"010101001",
  50194=>"101100001",
  50195=>"100000011",
  50196=>"001101110",
  50197=>"100111011",
  50198=>"110011110",
  50199=>"100110011",
  50200=>"000101110",
  50201=>"000010000",
  50202=>"000110010",
  50203=>"101010100",
  50204=>"000001010",
  50205=>"001111111",
  50206=>"100000101",
  50207=>"100010001",
  50208=>"000011100",
  50209=>"001010100",
  50210=>"011010011",
  50211=>"110000110",
  50212=>"000100111",
  50213=>"000110011",
  50214=>"111111111",
  50215=>"010000100",
  50216=>"010111000",
  50217=>"001101010",
  50218=>"110111110",
  50219=>"000110111",
  50220=>"000101110",
  50221=>"110101011",
  50222=>"000000100",
  50223=>"110100100",
  50224=>"110011010",
  50225=>"111111100",
  50226=>"000010111",
  50227=>"001001100",
  50228=>"001001111",
  50229=>"111001111",
  50230=>"010011011",
  50231=>"101110010",
  50232=>"110111000",
  50233=>"001100001",
  50234=>"001000011",
  50235=>"011001101",
  50236=>"101110111",
  50237=>"110100011",
  50238=>"110011001",
  50239=>"000001101",
  50240=>"011000011",
  50241=>"000000001",
  50242=>"000011000",
  50243=>"110100000",
  50244=>"100110010",
  50245=>"000001000",
  50246=>"000110100",
  50247=>"110001101",
  50248=>"000010011",
  50249=>"000000011",
  50250=>"010111100",
  50251=>"010010000",
  50252=>"101100100",
  50253=>"010000000",
  50254=>"000010010",
  50255=>"100110111",
  50256=>"100001100",
  50257=>"110110011",
  50258=>"101111110",
  50259=>"001011000",
  50260=>"110001000",
  50261=>"010000000",
  50262=>"101011111",
  50263=>"101100001",
  50264=>"100010011",
  50265=>"001111010",
  50266=>"011010000",
  50267=>"001001110",
  50268=>"010100111",
  50269=>"100110111",
  50270=>"110100101",
  50271=>"010110000",
  50272=>"010010111",
  50273=>"001101100",
  50274=>"110000000",
  50275=>"001100001",
  50276=>"100101101",
  50277=>"001111010",
  50278=>"010001110",
  50279=>"011100001",
  50280=>"110100101",
  50281=>"000110000",
  50282=>"100001101",
  50283=>"000000010",
  50284=>"101111011",
  50285=>"011101011",
  50286=>"011100111",
  50287=>"111100100",
  50288=>"101101000",
  50289=>"100111000",
  50290=>"101000011",
  50291=>"001000010",
  50292=>"111011001",
  50293=>"010000010",
  50294=>"111000011",
  50295=>"010111110",
  50296=>"010101100",
  50297=>"010110110",
  50298=>"001101100",
  50299=>"110000100",
  50300=>"101010000",
  50301=>"000100110",
  50302=>"111111111",
  50303=>"010000101",
  50304=>"010000010",
  50305=>"100010011",
  50306=>"111101001",
  50307=>"000001011",
  50308=>"001100001",
  50309=>"001001001",
  50310=>"000000111",
  50311=>"111011111",
  50312=>"110100101",
  50313=>"001000101",
  50314=>"000101011",
  50315=>"111110111",
  50316=>"001100110",
  50317=>"101101100",
  50318=>"100100011",
  50319=>"011100000",
  50320=>"111110111",
  50321=>"011101110",
  50322=>"111100111",
  50323=>"100011110",
  50324=>"000101010",
  50325=>"011110110",
  50326=>"100100100",
  50327=>"100001100",
  50328=>"100111001",
  50329=>"110000011",
  50330=>"011101010",
  50331=>"100011010",
  50332=>"010111010",
  50333=>"101010111",
  50334=>"100001000",
  50335=>"011011100",
  50336=>"101110010",
  50337=>"111110111",
  50338=>"101100111",
  50339=>"100100110",
  50340=>"000100011",
  50341=>"111101110",
  50342=>"111100000",
  50343=>"011000111",
  50344=>"110001111",
  50345=>"101100100",
  50346=>"001011101",
  50347=>"111010001",
  50348=>"001100110",
  50349=>"100111101",
  50350=>"111110110",
  50351=>"000101001",
  50352=>"001101000",
  50353=>"000010001",
  50354=>"101100010",
  50355=>"100100000",
  50356=>"001010100",
  50357=>"010011111",
  50358=>"001110111",
  50359=>"100100010",
  50360=>"100110000",
  50361=>"001101001",
  50362=>"101011110",
  50363=>"101010111",
  50364=>"100101101",
  50365=>"110111000",
  50366=>"010010010",
  50367=>"000100000",
  50368=>"110010110",
  50369=>"110000001",
  50370=>"111000010",
  50371=>"100100011",
  50372=>"110100000",
  50373=>"001000100",
  50374=>"000111101",
  50375=>"110100000",
  50376=>"001100100",
  50377=>"011111111",
  50378=>"001011001",
  50379=>"111111010",
  50380=>"001100011",
  50381=>"100111010",
  50382=>"001110111",
  50383=>"010100001",
  50384=>"110001000",
  50385=>"011010011",
  50386=>"000010101",
  50387=>"011000010",
  50388=>"000000010",
  50389=>"011000101",
  50390=>"100110111",
  50391=>"100101010",
  50392=>"100010001",
  50393=>"010010101",
  50394=>"111111001",
  50395=>"111101101",
  50396=>"011011010",
  50397=>"100100011",
  50398=>"110001001",
  50399=>"000101101",
  50400=>"010011101",
  50401=>"000100010",
  50402=>"101100001",
  50403=>"010100011",
  50404=>"000101000",
  50405=>"100100100",
  50406=>"111000100",
  50407=>"111111011",
  50408=>"111011010",
  50409=>"001101011",
  50410=>"101010001",
  50411=>"110111010",
  50412=>"111000101",
  50413=>"000101110",
  50414=>"101110101",
  50415=>"100001000",
  50416=>"100001100",
  50417=>"010000000",
  50418=>"000100000",
  50419=>"111001000",
  50420=>"001111110",
  50421=>"111010001",
  50422=>"110110011",
  50423=>"000100011",
  50424=>"100000111",
  50425=>"001000111",
  50426=>"001111100",
  50427=>"000110011",
  50428=>"011001101",
  50429=>"011001100",
  50430=>"101101001",
  50431=>"111111001",
  50432=>"000000000",
  50433=>"001000001",
  50434=>"101110000",
  50435=>"101101110",
  50436=>"011000001",
  50437=>"111101111",
  50438=>"011010100",
  50439=>"100000010",
  50440=>"011000100",
  50441=>"110000001",
  50442=>"000100000",
  50443=>"101101010",
  50444=>"011101011",
  50445=>"001000000",
  50446=>"000011000",
  50447=>"010000011",
  50448=>"010001101",
  50449=>"001010101",
  50450=>"010111111",
  50451=>"001011011",
  50452=>"110110101",
  50453=>"110011100",
  50454=>"000001001",
  50455=>"101100110",
  50456=>"000000010",
  50457=>"101011111",
  50458=>"011010110",
  50459=>"000011110",
  50460=>"000011110",
  50461=>"001111101",
  50462=>"010111001",
  50463=>"001001111",
  50464=>"000000000",
  50465=>"100100011",
  50466=>"100101001",
  50467=>"010101000",
  50468=>"111110001",
  50469=>"001001011",
  50470=>"100110000",
  50471=>"111110111",
  50472=>"010110000",
  50473=>"110100110",
  50474=>"011000000",
  50475=>"011011010",
  50476=>"100011010",
  50477=>"000010101",
  50478=>"000000011",
  50479=>"100010110",
  50480=>"100101100",
  50481=>"001101100",
  50482=>"011100001",
  50483=>"101101111",
  50484=>"100001101",
  50485=>"010000011",
  50486=>"000010000",
  50487=>"000000001",
  50488=>"101110111",
  50489=>"001111110",
  50490=>"101100100",
  50491=>"101011100",
  50492=>"011000011",
  50493=>"110011100",
  50494=>"001011111",
  50495=>"110100010",
  50496=>"010011111",
  50497=>"100100110",
  50498=>"011000011",
  50499=>"000100110",
  50500=>"110101101",
  50501=>"110100100",
  50502=>"010100000",
  50503=>"001110000",
  50504=>"100000100",
  50505=>"111011000",
  50506=>"110000110",
  50507=>"010001111",
  50508=>"111011010",
  50509=>"100101001",
  50510=>"001001110",
  50511=>"010000010",
  50512=>"010001000",
  50513=>"011010101",
  50514=>"011101000",
  50515=>"000111001",
  50516=>"000111011",
  50517=>"001000000",
  50518=>"101111101",
  50519=>"111101111",
  50520=>"000100011",
  50521=>"101111011",
  50522=>"101001010",
  50523=>"001111100",
  50524=>"010110101",
  50525=>"000101111",
  50526=>"101101111",
  50527=>"001111011",
  50528=>"001010111",
  50529=>"000000111",
  50530=>"101010001",
  50531=>"000011100",
  50532=>"010011101",
  50533=>"011110111",
  50534=>"110000011",
  50535=>"010101001",
  50536=>"111100011",
  50537=>"001010101",
  50538=>"101011011",
  50539=>"000110100",
  50540=>"100111010",
  50541=>"001001011",
  50542=>"110111111",
  50543=>"001110111",
  50544=>"010001110",
  50545=>"100011101",
  50546=>"100011100",
  50547=>"010111100",
  50548=>"100110100",
  50549=>"010100111",
  50550=>"101001000",
  50551=>"010100010",
  50552=>"100111110",
  50553=>"001000011",
  50554=>"100000001",
  50555=>"111101111",
  50556=>"111111000",
  50557=>"101010000",
  50558=>"010111000",
  50559=>"010011111",
  50560=>"111110100",
  50561=>"110100110",
  50562=>"101011010",
  50563=>"011101110",
  50564=>"100100010",
  50565=>"000100110",
  50566=>"011111010",
  50567=>"100100001",
  50568=>"001000100",
  50569=>"000001011",
  50570=>"000011110",
  50571=>"010011000",
  50572=>"100100110",
  50573=>"100000101",
  50574=>"001111011",
  50575=>"101001010",
  50576=>"001101110",
  50577=>"111111000",
  50578=>"001100010",
  50579=>"001011100",
  50580=>"111010011",
  50581=>"100001000",
  50582=>"000001010",
  50583=>"110010000",
  50584=>"001000000",
  50585=>"000001000",
  50586=>"100000111",
  50587=>"101001100",
  50588=>"100001111",
  50589=>"110001010",
  50590=>"101001000",
  50591=>"110010100",
  50592=>"111010101",
  50593=>"000100010",
  50594=>"001101001",
  50595=>"001001001",
  50596=>"101010111",
  50597=>"101001100",
  50598=>"001010101",
  50599=>"101010101",
  50600=>"001111010",
  50601=>"110001100",
  50602=>"100001000",
  50603=>"111011100",
  50604=>"110110100",
  50605=>"111110011",
  50606=>"000010000",
  50607=>"001111100",
  50608=>"000010101",
  50609=>"000111001",
  50610=>"101011010",
  50611=>"100011010",
  50612=>"110101010",
  50613=>"000101001",
  50614=>"011101011",
  50615=>"001101111",
  50616=>"011111000",
  50617=>"010111111",
  50618=>"111111101",
  50619=>"101100000",
  50620=>"001100100",
  50621=>"111011110",
  50622=>"101101011",
  50623=>"101100110",
  50624=>"010111110",
  50625=>"011000100",
  50626=>"001011010",
  50627=>"000111001",
  50628=>"111111111",
  50629=>"001010000",
  50630=>"011000100",
  50631=>"000110010",
  50632=>"101001011",
  50633=>"000000011",
  50634=>"101111111",
  50635=>"011011010",
  50636=>"110100101",
  50637=>"000010001",
  50638=>"100110010",
  50639=>"011011111",
  50640=>"110110100",
  50641=>"011100001",
  50642=>"110111101",
  50643=>"111110101",
  50644=>"010111010",
  50645=>"001110001",
  50646=>"100000111",
  50647=>"101010000",
  50648=>"000111010",
  50649=>"000000010",
  50650=>"010001010",
  50651=>"101010110",
  50652=>"011101110",
  50653=>"001110110",
  50654=>"100111001",
  50655=>"100110011",
  50656=>"000101110",
  50657=>"110110100",
  50658=>"110001010",
  50659=>"100011101",
  50660=>"011010101",
  50661=>"000011110",
  50662=>"001000000",
  50663=>"100010110",
  50664=>"000010001",
  50665=>"101001110",
  50666=>"010000010",
  50667=>"110101000",
  50668=>"010000101",
  50669=>"111111111",
  50670=>"111001101",
  50671=>"000111000",
  50672=>"000011010",
  50673=>"010001010",
  50674=>"011101011",
  50675=>"011001011",
  50676=>"111000111",
  50677=>"010001010",
  50678=>"001000111",
  50679=>"100101001",
  50680=>"010110010",
  50681=>"000000111",
  50682=>"110010100",
  50683=>"001010111",
  50684=>"011111110",
  50685=>"010100011",
  50686=>"001110110",
  50687=>"000000000",
  50688=>"011000111",
  50689=>"110101110",
  50690=>"000011100",
  50691=>"000010100",
  50692=>"110111010",
  50693=>"101000001",
  50694=>"000001110",
  50695=>"010100111",
  50696=>"111111010",
  50697=>"001000011",
  50698=>"110111001",
  50699=>"010000000",
  50700=>"011111100",
  50701=>"101001100",
  50702=>"001001100",
  50703=>"001011001",
  50704=>"001000010",
  50705=>"111011101",
  50706=>"101100001",
  50707=>"001100110",
  50708=>"100011111",
  50709=>"111001000",
  50710=>"101100101",
  50711=>"100001000",
  50712=>"000101000",
  50713=>"011001100",
  50714=>"110000110",
  50715=>"011111101",
  50716=>"000010101",
  50717=>"011001010",
  50718=>"011101000",
  50719=>"010001101",
  50720=>"011101110",
  50721=>"010100011",
  50722=>"100000011",
  50723=>"001101100",
  50724=>"110000010",
  50725=>"011001000",
  50726=>"011110111",
  50727=>"111010010",
  50728=>"001110111",
  50729=>"000001000",
  50730=>"011110010",
  50731=>"010100100",
  50732=>"001100011",
  50733=>"110000110",
  50734=>"010011000",
  50735=>"000100101",
  50736=>"011101111",
  50737=>"010110111",
  50738=>"000100101",
  50739=>"111110011",
  50740=>"110011000",
  50741=>"101011101",
  50742=>"101001100",
  50743=>"010101100",
  50744=>"001011110",
  50745=>"001010000",
  50746=>"111000011",
  50747=>"011011011",
  50748=>"110000110",
  50749=>"011100000",
  50750=>"010011100",
  50751=>"100010000",
  50752=>"111000111",
  50753=>"101001000",
  50754=>"001001111",
  50755=>"100101100",
  50756=>"110110001",
  50757=>"010110011",
  50758=>"000001001",
  50759=>"010010001",
  50760=>"111010001",
  50761=>"111101101",
  50762=>"110011101",
  50763=>"110101010",
  50764=>"100101111",
  50765=>"000001011",
  50766=>"001101100",
  50767=>"001011011",
  50768=>"000011011",
  50769=>"011110101",
  50770=>"101010001",
  50771=>"101001000",
  50772=>"010111000",
  50773=>"100010100",
  50774=>"010011110",
  50775=>"101000100",
  50776=>"110110010",
  50777=>"110010001",
  50778=>"011101010",
  50779=>"001111101",
  50780=>"110000000",
  50781=>"010000110",
  50782=>"111010101",
  50783=>"100010100",
  50784=>"101111011",
  50785=>"001000001",
  50786=>"101110010",
  50787=>"000101001",
  50788=>"100101011",
  50789=>"000010001",
  50790=>"011001010",
  50791=>"000010000",
  50792=>"000101111",
  50793=>"000011100",
  50794=>"110110100",
  50795=>"000001000",
  50796=>"010101000",
  50797=>"111000011",
  50798=>"111100011",
  50799=>"001000000",
  50800=>"100101001",
  50801=>"011100101",
  50802=>"100111011",
  50803=>"001111000",
  50804=>"000101010",
  50805=>"110001110",
  50806=>"000110011",
  50807=>"011011010",
  50808=>"110111000",
  50809=>"010010001",
  50810=>"101100010",
  50811=>"001011010",
  50812=>"100001011",
  50813=>"100100011",
  50814=>"010000000",
  50815=>"101101110",
  50816=>"100001101",
  50817=>"000110000",
  50818=>"000101101",
  50819=>"001000000",
  50820=>"101001001",
  50821=>"001110000",
  50822=>"010100100",
  50823=>"101111000",
  50824=>"111010101",
  50825=>"101000111",
  50826=>"011110011",
  50827=>"000110011",
  50828=>"010001000",
  50829=>"100111101",
  50830=>"100001111",
  50831=>"111110111",
  50832=>"000001000",
  50833=>"010100111",
  50834=>"001110010",
  50835=>"100011111",
  50836=>"000001100",
  50837=>"011000101",
  50838=>"110100111",
  50839=>"111101110",
  50840=>"010100101",
  50841=>"111011110",
  50842=>"010101011",
  50843=>"101110001",
  50844=>"101011000",
  50845=>"000101110",
  50846=>"001110011",
  50847=>"110010001",
  50848=>"010110000",
  50849=>"010100010",
  50850=>"011011010",
  50851=>"001011111",
  50852=>"110011001",
  50853=>"101111111",
  50854=>"111010101",
  50855=>"110011111",
  50856=>"001000010",
  50857=>"101101011",
  50858=>"011101110",
  50859=>"101101001",
  50860=>"011101111",
  50861=>"010110100",
  50862=>"000100011",
  50863=>"111111110",
  50864=>"001000101",
  50865=>"110001100",
  50866=>"000100010",
  50867=>"010001111",
  50868=>"001101011",
  50869=>"101000010",
  50870=>"100001111",
  50871=>"001001000",
  50872=>"100001001",
  50873=>"011111110",
  50874=>"101110111",
  50875=>"101110000",
  50876=>"000111000",
  50877=>"001010001",
  50878=>"001001001",
  50879=>"100110101",
  50880=>"010000110",
  50881=>"111100001",
  50882=>"011101010",
  50883=>"001011111",
  50884=>"000000111",
  50885=>"101010101",
  50886=>"100011000",
  50887=>"110010001",
  50888=>"111101111",
  50889=>"111010000",
  50890=>"101000111",
  50891=>"000101010",
  50892=>"000111101",
  50893=>"101001000",
  50894=>"111110110",
  50895=>"100100110",
  50896=>"100001100",
  50897=>"111101101",
  50898=>"100000001",
  50899=>"111101011",
  50900=>"000010110",
  50901=>"001100010",
  50902=>"101011100",
  50903=>"011010001",
  50904=>"111100101",
  50905=>"100000101",
  50906=>"100100000",
  50907=>"000011010",
  50908=>"000111101",
  50909=>"000010001",
  50910=>"110101110",
  50911=>"110100010",
  50912=>"110000000",
  50913=>"111000011",
  50914=>"011000100",
  50915=>"100010100",
  50916=>"010001000",
  50917=>"110011000",
  50918=>"110111000",
  50919=>"010110100",
  50920=>"111110110",
  50921=>"101011010",
  50922=>"111000110",
  50923=>"100101111",
  50924=>"111110111",
  50925=>"111011111",
  50926=>"100111001",
  50927=>"011111101",
  50928=>"110100001",
  50929=>"111101000",
  50930=>"000001000",
  50931=>"110001010",
  50932=>"001000101",
  50933=>"001110100",
  50934=>"101011110",
  50935=>"000100011",
  50936=>"101110110",
  50937=>"111010011",
  50938=>"100010010",
  50939=>"101010001",
  50940=>"111000010",
  50941=>"011111001",
  50942=>"111111000",
  50943=>"111111011",
  50944=>"010000000",
  50945=>"000001000",
  50946=>"100001110",
  50947=>"010000110",
  50948=>"010101101",
  50949=>"000001010",
  50950=>"001011101",
  50951=>"110000000",
  50952=>"001010001",
  50953=>"110111101",
  50954=>"010111001",
  50955=>"110001100",
  50956=>"100111011",
  50957=>"001101000",
  50958=>"111101001",
  50959=>"100001010",
  50960=>"010010010",
  50961=>"111010010",
  50962=>"111111100",
  50963=>"011011101",
  50964=>"000110001",
  50965=>"111001100",
  50966=>"111100101",
  50967=>"001101001",
  50968=>"000001110",
  50969=>"000101001",
  50970=>"000110111",
  50971=>"011001001",
  50972=>"001111100",
  50973=>"110111111",
  50974=>"000110100",
  50975=>"010010111",
  50976=>"100111101",
  50977=>"010011000",
  50978=>"100110000",
  50979=>"001010100",
  50980=>"010110010",
  50981=>"101011000",
  50982=>"101011100",
  50983=>"001111010",
  50984=>"111111011",
  50985=>"111101010",
  50986=>"101011000",
  50987=>"100111111",
  50988=>"000010001",
  50989=>"000100010",
  50990=>"010100100",
  50991=>"101011010",
  50992=>"100001000",
  50993=>"111000100",
  50994=>"000000101",
  50995=>"001101010",
  50996=>"001000000",
  50997=>"010010010",
  50998=>"101110010",
  50999=>"000110101",
  51000=>"011010011",
  51001=>"100010111",
  51002=>"000011000",
  51003=>"110010101",
  51004=>"101001101",
  51005=>"111111010",
  51006=>"001010100",
  51007=>"101100000",
  51008=>"101101010",
  51009=>"111100110",
  51010=>"100000111",
  51011=>"100010010",
  51012=>"011101100",
  51013=>"111010101",
  51014=>"010111110",
  51015=>"110001000",
  51016=>"111100100",
  51017=>"111110011",
  51018=>"101000001",
  51019=>"101000101",
  51020=>"110010100",
  51021=>"111100001",
  51022=>"111111011",
  51023=>"100101111",
  51024=>"000001000",
  51025=>"011101110",
  51026=>"000101111",
  51027=>"110011011",
  51028=>"111000111",
  51029=>"111010000",
  51030=>"000001110",
  51031=>"100000011",
  51032=>"101000101",
  51033=>"110001001",
  51034=>"000111010",
  51035=>"001001110",
  51036=>"110110110",
  51037=>"000001110",
  51038=>"100010011",
  51039=>"110110000",
  51040=>"000010001",
  51041=>"111011111",
  51042=>"100000011",
  51043=>"011000011",
  51044=>"010110101",
  51045=>"001010110",
  51046=>"100110011",
  51047=>"100100100",
  51048=>"100011000",
  51049=>"100011111",
  51050=>"001101010",
  51051=>"000101000",
  51052=>"101101011",
  51053=>"000000100",
  51054=>"100111010",
  51055=>"000111000",
  51056=>"000101000",
  51057=>"111011100",
  51058=>"111110001",
  51059=>"111000101",
  51060=>"001001110",
  51061=>"101101111",
  51062=>"111111101",
  51063=>"011110000",
  51064=>"000000001",
  51065=>"001001011",
  51066=>"100101001",
  51067=>"010100111",
  51068=>"000000011",
  51069=>"111110101",
  51070=>"110111100",
  51071=>"111000001",
  51072=>"110110001",
  51073=>"010000010",
  51074=>"010110010",
  51075=>"101001011",
  51076=>"000001110",
  51077=>"110000110",
  51078=>"111110110",
  51079=>"001101110",
  51080=>"101011000",
  51081=>"011111100",
  51082=>"000100101",
  51083=>"010110110",
  51084=>"010100010",
  51085=>"001110011",
  51086=>"001101000",
  51087=>"110110000",
  51088=>"111001111",
  51089=>"111001000",
  51090=>"000000001",
  51091=>"011001001",
  51092=>"001001111",
  51093=>"101010011",
  51094=>"000011010",
  51095=>"010101011",
  51096=>"101100111",
  51097=>"000010000",
  51098=>"010110110",
  51099=>"010101001",
  51100=>"000011101",
  51101=>"110010001",
  51102=>"000100011",
  51103=>"001001000",
  51104=>"011000111",
  51105=>"000010110",
  51106=>"010110110",
  51107=>"001011010",
  51108=>"000010011",
  51109=>"000000110",
  51110=>"001110101",
  51111=>"101111111",
  51112=>"010100111",
  51113=>"010010001",
  51114=>"101110001",
  51115=>"100100100",
  51116=>"010101101",
  51117=>"010000111",
  51118=>"110110101",
  51119=>"001001111",
  51120=>"110001100",
  51121=>"101011110",
  51122=>"001101011",
  51123=>"111101101",
  51124=>"110110000",
  51125=>"111000111",
  51126=>"101100011",
  51127=>"110101010",
  51128=>"101101001",
  51129=>"101011001",
  51130=>"001100111",
  51131=>"101110011",
  51132=>"011100010",
  51133=>"011001100",
  51134=>"000000000",
  51135=>"010110110",
  51136=>"000011111",
  51137=>"110100110",
  51138=>"111111011",
  51139=>"010111111",
  51140=>"111101011",
  51141=>"010110100",
  51142=>"101011110",
  51143=>"111011010",
  51144=>"111100000",
  51145=>"010000000",
  51146=>"100100111",
  51147=>"000110111",
  51148=>"111101010",
  51149=>"111111011",
  51150=>"000011100",
  51151=>"011101101",
  51152=>"110001110",
  51153=>"001101010",
  51154=>"110011110",
  51155=>"000001000",
  51156=>"100010010",
  51157=>"110011011",
  51158=>"010010100",
  51159=>"001100111",
  51160=>"011110011",
  51161=>"111101111",
  51162=>"001110111",
  51163=>"100111011",
  51164=>"011011011",
  51165=>"000011100",
  51166=>"001100011",
  51167=>"010101000",
  51168=>"001011010",
  51169=>"011100000",
  51170=>"001011101",
  51171=>"011100000",
  51172=>"100001010",
  51173=>"000010011",
  51174=>"100100000",
  51175=>"101100110",
  51176=>"111001000",
  51177=>"011111100",
  51178=>"000101100",
  51179=>"111011101",
  51180=>"000101011",
  51181=>"101011001",
  51182=>"001011001",
  51183=>"110000101",
  51184=>"110010010",
  51185=>"100101100",
  51186=>"111011101",
  51187=>"110011111",
  51188=>"000000111",
  51189=>"110101000",
  51190=>"011101010",
  51191=>"101111011",
  51192=>"001000010",
  51193=>"001100101",
  51194=>"000111010",
  51195=>"110001101",
  51196=>"011010010",
  51197=>"101110000",
  51198=>"110100010",
  51199=>"101111111",
  51200=>"100011000",
  51201=>"100001100",
  51202=>"101010111",
  51203=>"001111101",
  51204=>"110001011",
  51205=>"101001001",
  51206=>"101101001",
  51207=>"100011011",
  51208=>"101001001",
  51209=>"010010001",
  51210=>"101101100",
  51211=>"011011100",
  51212=>"000010101",
  51213=>"100001011",
  51214=>"110111001",
  51215=>"110001011",
  51216=>"101001101",
  51217=>"001000000",
  51218=>"010111010",
  51219=>"001111101",
  51220=>"011011101",
  51221=>"011011010",
  51222=>"010001000",
  51223=>"110101011",
  51224=>"111110000",
  51225=>"111011100",
  51226=>"010000100",
  51227=>"111011011",
  51228=>"111110100",
  51229=>"100101010",
  51230=>"000000001",
  51231=>"010000100",
  51232=>"011001100",
  51233=>"101101011",
  51234=>"100001110",
  51235=>"110011110",
  51236=>"110100111",
  51237=>"010100001",
  51238=>"111100110",
  51239=>"100101111",
  51240=>"001110110",
  51241=>"010110111",
  51242=>"110101001",
  51243=>"100101111",
  51244=>"111010111",
  51245=>"101100100",
  51246=>"101001100",
  51247=>"001001000",
  51248=>"100011010",
  51249=>"010111100",
  51250=>"110100101",
  51251=>"011100011",
  51252=>"111111011",
  51253=>"100001010",
  51254=>"111111110",
  51255=>"101100010",
  51256=>"011001010",
  51257=>"010011110",
  51258=>"101101111",
  51259=>"101111010",
  51260=>"001001110",
  51261=>"001111010",
  51262=>"100100110",
  51263=>"111010011",
  51264=>"000111010",
  51265=>"000110010",
  51266=>"110111111",
  51267=>"100000011",
  51268=>"011001010",
  51269=>"111111000",
  51270=>"100000010",
  51271=>"100000001",
  51272=>"110000001",
  51273=>"000001111",
  51274=>"000100111",
  51275=>"010110111",
  51276=>"000001010",
  51277=>"011110000",
  51278=>"101101100",
  51279=>"000110011",
  51280=>"101100101",
  51281=>"111101100",
  51282=>"001000001",
  51283=>"100100101",
  51284=>"101100010",
  51285=>"111101101",
  51286=>"111110011",
  51287=>"101101111",
  51288=>"110000100",
  51289=>"101101011",
  51290=>"110100010",
  51291=>"101101110",
  51292=>"001001101",
  51293=>"111111100",
  51294=>"100010010",
  51295=>"111010110",
  51296=>"111000101",
  51297=>"110111010",
  51298=>"001101000",
  51299=>"000100010",
  51300=>"011000100",
  51301=>"001010000",
  51302=>"111001000",
  51303=>"100111010",
  51304=>"101101111",
  51305=>"111010011",
  51306=>"010000001",
  51307=>"010101000",
  51308=>"111011010",
  51309=>"100001010",
  51310=>"111000111",
  51311=>"111111110",
  51312=>"011100100",
  51313=>"111001101",
  51314=>"111110101",
  51315=>"011100001",
  51316=>"010110110",
  51317=>"000000011",
  51318=>"101111011",
  51319=>"100011111",
  51320=>"000101001",
  51321=>"101111100",
  51322=>"000001000",
  51323=>"011100011",
  51324=>"100100010",
  51325=>"010001011",
  51326=>"000111100",
  51327=>"110000000",
  51328=>"101100011",
  51329=>"000100011",
  51330=>"010001011",
  51331=>"101111010",
  51332=>"010111010",
  51333=>"110011100",
  51334=>"101000111",
  51335=>"111100000",
  51336=>"101011001",
  51337=>"011000011",
  51338=>"000011110",
  51339=>"000001110",
  51340=>"110100111",
  51341=>"100111110",
  51342=>"001010110",
  51343=>"011001011",
  51344=>"100110100",
  51345=>"111000111",
  51346=>"111010011",
  51347=>"011101101",
  51348=>"001011110",
  51349=>"110111011",
  51350=>"000000001",
  51351=>"001100110",
  51352=>"000011010",
  51353=>"010101000",
  51354=>"000110000",
  51355=>"100000000",
  51356=>"101010101",
  51357=>"000010111",
  51358=>"000001001",
  51359=>"010011010",
  51360=>"110001110",
  51361=>"101110001",
  51362=>"110111101",
  51363=>"001010110",
  51364=>"011101101",
  51365=>"100111011",
  51366=>"001110011",
  51367=>"001011111",
  51368=>"011111011",
  51369=>"110011000",
  51370=>"010011101",
  51371=>"000010001",
  51372=>"101000110",
  51373=>"111111110",
  51374=>"010001000",
  51375=>"001000110",
  51376=>"010101011",
  51377=>"111001101",
  51378=>"010101001",
  51379=>"101101011",
  51380=>"101100001",
  51381=>"010000010",
  51382=>"100111110",
  51383=>"011100111",
  51384=>"001011010",
  51385=>"110110010",
  51386=>"000001001",
  51387=>"011111110",
  51388=>"101101111",
  51389=>"000100100",
  51390=>"111000000",
  51391=>"010011001",
  51392=>"101001110",
  51393=>"101110000",
  51394=>"111011001",
  51395=>"000110101",
  51396=>"010111001",
  51397=>"111001101",
  51398=>"111111111",
  51399=>"101011100",
  51400=>"101010000",
  51401=>"011110000",
  51402=>"000101111",
  51403=>"101000001",
  51404=>"011111000",
  51405=>"111111111",
  51406=>"000101101",
  51407=>"000011111",
  51408=>"010011101",
  51409=>"111000110",
  51410=>"111100010",
  51411=>"101111101",
  51412=>"000010110",
  51413=>"100110110",
  51414=>"110010111",
  51415=>"001010001",
  51416=>"010000100",
  51417=>"100000001",
  51418=>"110101100",
  51419=>"100000011",
  51420=>"000100110",
  51421=>"010010110",
  51422=>"001101000",
  51423=>"011100011",
  51424=>"100110101",
  51425=>"101111000",
  51426=>"111110110",
  51427=>"111111100",
  51428=>"110110001",
  51429=>"001000110",
  51430=>"010100010",
  51431=>"011010110",
  51432=>"110101101",
  51433=>"001110101",
  51434=>"100010110",
  51435=>"001101111",
  51436=>"010010101",
  51437=>"010111011",
  51438=>"110000111",
  51439=>"111000001",
  51440=>"110100111",
  51441=>"001100101",
  51442=>"010010101",
  51443=>"101101011",
  51444=>"000001101",
  51445=>"001011110",
  51446=>"000001000",
  51447=>"100100001",
  51448=>"001101110",
  51449=>"100010101",
  51450=>"101101100",
  51451=>"000001100",
  51452=>"001000100",
  51453=>"011110000",
  51454=>"000011110",
  51455=>"111011001",
  51456=>"001001110",
  51457=>"101011111",
  51458=>"010001110",
  51459=>"010000111",
  51460=>"101100101",
  51461=>"111100001",
  51462=>"110000000",
  51463=>"100111111",
  51464=>"100110011",
  51465=>"101001001",
  51466=>"001101110",
  51467=>"101101111",
  51468=>"001111001",
  51469=>"000101101",
  51470=>"011000010",
  51471=>"010001111",
  51472=>"001011110",
  51473=>"010100101",
  51474=>"111100101",
  51475=>"010101000",
  51476=>"111011111",
  51477=>"110000010",
  51478=>"010110010",
  51479=>"111011100",
  51480=>"010001010",
  51481=>"110101011",
  51482=>"001010101",
  51483=>"010101111",
  51484=>"000110010",
  51485=>"010000110",
  51486=>"100010001",
  51487=>"101011100",
  51488=>"001001101",
  51489=>"010111011",
  51490=>"110110110",
  51491=>"010110100",
  51492=>"010010110",
  51493=>"110100100",
  51494=>"010101101",
  51495=>"111011101",
  51496=>"010011000",
  51497=>"100110101",
  51498=>"111001000",
  51499=>"100000001",
  51500=>"010100111",
  51501=>"111111000",
  51502=>"101001010",
  51503=>"111101110",
  51504=>"001011000",
  51505=>"010011010",
  51506=>"001010100",
  51507=>"101100111",
  51508=>"010110011",
  51509=>"001000100",
  51510=>"010110101",
  51511=>"110100011",
  51512=>"000010011",
  51513=>"011011110",
  51514=>"000010110",
  51515=>"111001101",
  51516=>"101010011",
  51517=>"000011101",
  51518=>"010000010",
  51519=>"010101110",
  51520=>"010111100",
  51521=>"010000000",
  51522=>"110111001",
  51523=>"000110101",
  51524=>"011001101",
  51525=>"110011001",
  51526=>"110110001",
  51527=>"010110101",
  51528=>"111011101",
  51529=>"101000000",
  51530=>"000000011",
  51531=>"101011111",
  51532=>"100011100",
  51533=>"010100001",
  51534=>"010001101",
  51535=>"001110011",
  51536=>"010000000",
  51537=>"101110110",
  51538=>"000110110",
  51539=>"010100000",
  51540=>"000101110",
  51541=>"011100001",
  51542=>"011111111",
  51543=>"001110010",
  51544=>"000000000",
  51545=>"000110000",
  51546=>"010100000",
  51547=>"010011110",
  51548=>"101110001",
  51549=>"111111111",
  51550=>"010001101",
  51551=>"100110111",
  51552=>"110010000",
  51553=>"101001001",
  51554=>"000110110",
  51555=>"000000110",
  51556=>"100100100",
  51557=>"011111011",
  51558=>"111111000",
  51559=>"010011001",
  51560=>"110001111",
  51561=>"101100000",
  51562=>"010010101",
  51563=>"110000100",
  51564=>"010010101",
  51565=>"001110110",
  51566=>"010110111",
  51567=>"101110010",
  51568=>"011000111",
  51569=>"011001000",
  51570=>"110010010",
  51571=>"110100100",
  51572=>"101101100",
  51573=>"010100011",
  51574=>"111000000",
  51575=>"011011011",
  51576=>"111100011",
  51577=>"000001100",
  51578=>"111010110",
  51579=>"101000001",
  51580=>"101111111",
  51581=>"100111001",
  51582=>"000110001",
  51583=>"111000011",
  51584=>"111101111",
  51585=>"101101100",
  51586=>"011000010",
  51587=>"110111001",
  51588=>"101001000",
  51589=>"010111001",
  51590=>"001010101",
  51591=>"000000111",
  51592=>"100001010",
  51593=>"011111001",
  51594=>"110001100",
  51595=>"001000000",
  51596=>"000001101",
  51597=>"111100110",
  51598=>"111111111",
  51599=>"110010011",
  51600=>"110011111",
  51601=>"011100010",
  51602=>"000011011",
  51603=>"010010010",
  51604=>"110110100",
  51605=>"000000000",
  51606=>"000110011",
  51607=>"001101010",
  51608=>"010110001",
  51609=>"000001100",
  51610=>"000011000",
  51611=>"111110111",
  51612=>"111100100",
  51613=>"000001100",
  51614=>"000111111",
  51615=>"011010001",
  51616=>"111101011",
  51617=>"010000100",
  51618=>"110001100",
  51619=>"001101111",
  51620=>"001010010",
  51621=>"100000010",
  51622=>"011100000",
  51623=>"110000101",
  51624=>"011110011",
  51625=>"000100000",
  51626=>"100000010",
  51627=>"100100001",
  51628=>"100001110",
  51629=>"111100100",
  51630=>"110011100",
  51631=>"011110000",
  51632=>"000101000",
  51633=>"001000000",
  51634=>"001111000",
  51635=>"111101110",
  51636=>"111101001",
  51637=>"110111111",
  51638=>"111101101",
  51639=>"000010111",
  51640=>"110011101",
  51641=>"100010111",
  51642=>"101111110",
  51643=>"011101010",
  51644=>"110101000",
  51645=>"000111000",
  51646=>"000101000",
  51647=>"001101111",
  51648=>"010100110",
  51649=>"000000001",
  51650=>"011011010",
  51651=>"111000000",
  51652=>"111110101",
  51653=>"111111000",
  51654=>"000001011",
  51655=>"100111111",
  51656=>"000111100",
  51657=>"011000100",
  51658=>"111001011",
  51659=>"001011001",
  51660=>"000100010",
  51661=>"101010001",
  51662=>"011101010",
  51663=>"011010010",
  51664=>"110110010",
  51665=>"110011010",
  51666=>"101111111",
  51667=>"100010000",
  51668=>"111111111",
  51669=>"110110001",
  51670=>"010100001",
  51671=>"100001010",
  51672=>"011001010",
  51673=>"101100100",
  51674=>"011000000",
  51675=>"010011000",
  51676=>"111010001",
  51677=>"101001110",
  51678=>"110011011",
  51679=>"111111101",
  51680=>"111101000",
  51681=>"011010111",
  51682=>"011011010",
  51683=>"101000011",
  51684=>"000110011",
  51685=>"101111011",
  51686=>"101010011",
  51687=>"111101100",
  51688=>"100110000",
  51689=>"000110000",
  51690=>"101101011",
  51691=>"100000110",
  51692=>"100010110",
  51693=>"100001100",
  51694=>"100001101",
  51695=>"011010101",
  51696=>"110011110",
  51697=>"110100111",
  51698=>"100010010",
  51699=>"000000101",
  51700=>"100100001",
  51701=>"100111101",
  51702=>"100111000",
  51703=>"011100001",
  51704=>"110101010",
  51705=>"111000011",
  51706=>"001001100",
  51707=>"011110111",
  51708=>"111011110",
  51709=>"110100100",
  51710=>"000100001",
  51711=>"011101000",
  51712=>"011011011",
  51713=>"100110000",
  51714=>"011010110",
  51715=>"100110111",
  51716=>"001010001",
  51717=>"010000111",
  51718=>"101001100",
  51719=>"110101010",
  51720=>"001011110",
  51721=>"111111011",
  51722=>"001101111",
  51723=>"001101110",
  51724=>"111111111",
  51725=>"110101111",
  51726=>"011011111",
  51727=>"000111001",
  51728=>"010110000",
  51729=>"111101001",
  51730=>"010000000",
  51731=>"110110101",
  51732=>"110100000",
  51733=>"000010011",
  51734=>"101100010",
  51735=>"000010101",
  51736=>"111001101",
  51737=>"100101001",
  51738=>"100111101",
  51739=>"110110100",
  51740=>"010000000",
  51741=>"011100111",
  51742=>"000100111",
  51743=>"110101011",
  51744=>"001000101",
  51745=>"100111101",
  51746=>"111110100",
  51747=>"111101100",
  51748=>"100101110",
  51749=>"010101101",
  51750=>"100011011",
  51751=>"000010010",
  51752=>"001001000",
  51753=>"010110100",
  51754=>"111111101",
  51755=>"110010011",
  51756=>"100100010",
  51757=>"110111001",
  51758=>"011110010",
  51759=>"001001100",
  51760=>"000111111",
  51761=>"111010111",
  51762=>"111000011",
  51763=>"011011111",
  51764=>"000100000",
  51765=>"101111010",
  51766=>"100001010",
  51767=>"010101011",
  51768=>"100101100",
  51769=>"111111011",
  51770=>"110010010",
  51771=>"100011110",
  51772=>"111000111",
  51773=>"111101001",
  51774=>"000000110",
  51775=>"110011100",
  51776=>"101010001",
  51777=>"001110101",
  51778=>"001100101",
  51779=>"110110101",
  51780=>"000110111",
  51781=>"010100010",
  51782=>"111100111",
  51783=>"100110100",
  51784=>"000011011",
  51785=>"101000110",
  51786=>"011010000",
  51787=>"100000001",
  51788=>"010100010",
  51789=>"110010110",
  51790=>"101000100",
  51791=>"001111010",
  51792=>"111000101",
  51793=>"111010101",
  51794=>"110011011",
  51795=>"101100100",
  51796=>"110110100",
  51797=>"001110100",
  51798=>"110000100",
  51799=>"111001000",
  51800=>"011111011",
  51801=>"111100101",
  51802=>"001100101",
  51803=>"011101010",
  51804=>"010101111",
  51805=>"010101111",
  51806=>"010111110",
  51807=>"001011111",
  51808=>"111010111",
  51809=>"111110110",
  51810=>"001111000",
  51811=>"011011110",
  51812=>"010001111",
  51813=>"010011011",
  51814=>"111101100",
  51815=>"000110101",
  51816=>"111111101",
  51817=>"000100111",
  51818=>"111010110",
  51819=>"110000110",
  51820=>"100001101",
  51821=>"001110100",
  51822=>"011000111",
  51823=>"110100011",
  51824=>"110101010",
  51825=>"110111100",
  51826=>"010111110",
  51827=>"010011100",
  51828=>"010111001",
  51829=>"100000011",
  51830=>"010000010",
  51831=>"001010000",
  51832=>"010011011",
  51833=>"101011111",
  51834=>"000010101",
  51835=>"110100111",
  51836=>"000001010",
  51837=>"000001111",
  51838=>"011101010",
  51839=>"011101010",
  51840=>"011000011",
  51841=>"011110111",
  51842=>"000000000",
  51843=>"111100101",
  51844=>"110101010",
  51845=>"000111001",
  51846=>"110000100",
  51847=>"001111111",
  51848=>"111110110",
  51849=>"000110000",
  51850=>"100100010",
  51851=>"011110100",
  51852=>"101000001",
  51853=>"010100101",
  51854=>"100010111",
  51855=>"100100111",
  51856=>"101000100",
  51857=>"000100001",
  51858=>"011000100",
  51859=>"110010001",
  51860=>"001001000",
  51861=>"000011111",
  51862=>"101001000",
  51863=>"101010011",
  51864=>"000011000",
  51865=>"000101100",
  51866=>"110000000",
  51867=>"000100000",
  51868=>"111001001",
  51869=>"010001101",
  51870=>"000110101",
  51871=>"010100010",
  51872=>"101100100",
  51873=>"010001010",
  51874=>"110101000",
  51875=>"100000001",
  51876=>"111101111",
  51877=>"111010010",
  51878=>"001110110",
  51879=>"110100111",
  51880=>"010000100",
  51881=>"011101110",
  51882=>"100011111",
  51883=>"110110100",
  51884=>"111101001",
  51885=>"010110010",
  51886=>"000001110",
  51887=>"100000000",
  51888=>"101111000",
  51889=>"111110000",
  51890=>"100000100",
  51891=>"010111100",
  51892=>"010000000",
  51893=>"101010000",
  51894=>"101100001",
  51895=>"110101000",
  51896=>"110100000",
  51897=>"000100011",
  51898=>"100111010",
  51899=>"111100011",
  51900=>"000110011",
  51901=>"101111111",
  51902=>"101101011",
  51903=>"111000010",
  51904=>"011101101",
  51905=>"010101110",
  51906=>"101000110",
  51907=>"001001010",
  51908=>"101010011",
  51909=>"011000100",
  51910=>"000010010",
  51911=>"010111010",
  51912=>"100100110",
  51913=>"000000011",
  51914=>"110100011",
  51915=>"111010011",
  51916=>"000111010",
  51917=>"001111011",
  51918=>"111110110",
  51919=>"111101110",
  51920=>"010101101",
  51921=>"111001110",
  51922=>"011011000",
  51923=>"111001101",
  51924=>"111101101",
  51925=>"011101010",
  51926=>"100000101",
  51927=>"001001001",
  51928=>"111001001",
  51929=>"111111010",
  51930=>"111001111",
  51931=>"110010010",
  51932=>"001110000",
  51933=>"111100100",
  51934=>"011011010",
  51935=>"100101001",
  51936=>"100110110",
  51937=>"010000011",
  51938=>"001011101",
  51939=>"101110111",
  51940=>"011010001",
  51941=>"100111000",
  51942=>"101111001",
  51943=>"101100111",
  51944=>"000111000",
  51945=>"100100111",
  51946=>"010000000",
  51947=>"011011001",
  51948=>"111111111",
  51949=>"000110011",
  51950=>"001010000",
  51951=>"001101100",
  51952=>"000101001",
  51953=>"100001011",
  51954=>"110111000",
  51955=>"000000110",
  51956=>"100110001",
  51957=>"100000110",
  51958=>"101011010",
  51959=>"100100100",
  51960=>"101101001",
  51961=>"001100000",
  51962=>"010000001",
  51963=>"101101100",
  51964=>"010011011",
  51965=>"000101111",
  51966=>"011110111",
  51967=>"110001111",
  51968=>"110110111",
  51969=>"000000011",
  51970=>"000000110",
  51971=>"010001011",
  51972=>"000010001",
  51973=>"100111110",
  51974=>"001111110",
  51975=>"101110100",
  51976=>"010100000",
  51977=>"001001000",
  51978=>"100111110",
  51979=>"000010000",
  51980=>"100000011",
  51981=>"011101001",
  51982=>"010111000",
  51983=>"011101010",
  51984=>"111001001",
  51985=>"001101000",
  51986=>"101110001",
  51987=>"010001010",
  51988=>"110011010",
  51989=>"010110011",
  51990=>"010101000",
  51991=>"111001111",
  51992=>"001100111",
  51993=>"101110110",
  51994=>"111110110",
  51995=>"000100010",
  51996=>"110111000",
  51997=>"011111011",
  51998=>"101001100",
  51999=>"100000111",
  52000=>"010000010",
  52001=>"101111000",
  52002=>"111110000",
  52003=>"000110001",
  52004=>"000011001",
  52005=>"111001111",
  52006=>"100010101",
  52007=>"100110000",
  52008=>"100101100",
  52009=>"100000110",
  52010=>"001000011",
  52011=>"110111001",
  52012=>"001011111",
  52013=>"001001110",
  52014=>"101100011",
  52015=>"100000010",
  52016=>"101111010",
  52017=>"010011101",
  52018=>"011001100",
  52019=>"000011110",
  52020=>"100101011",
  52021=>"010011100",
  52022=>"110001001",
  52023=>"000101010",
  52024=>"000101101",
  52025=>"100000100",
  52026=>"010001001",
  52027=>"101111000",
  52028=>"101101101",
  52029=>"000001000",
  52030=>"000100111",
  52031=>"110111001",
  52032=>"010010010",
  52033=>"001011001",
  52034=>"000110100",
  52035=>"111010111",
  52036=>"000001101",
  52037=>"110000111",
  52038=>"111101011",
  52039=>"000100011",
  52040=>"000011000",
  52041=>"001011011",
  52042=>"110001000",
  52043=>"101010110",
  52044=>"000001000",
  52045=>"110110010",
  52046=>"100110010",
  52047=>"000000100",
  52048=>"111111100",
  52049=>"001111010",
  52050=>"100110110",
  52051=>"011100011",
  52052=>"101010011",
  52053=>"011011100",
  52054=>"110011100",
  52055=>"011000111",
  52056=>"101101010",
  52057=>"010001001",
  52058=>"001000010",
  52059=>"000001101",
  52060=>"111110100",
  52061=>"000010000",
  52062=>"001110010",
  52063=>"111101011",
  52064=>"111000011",
  52065=>"011110110",
  52066=>"100111010",
  52067=>"001110001",
  52068=>"000101101",
  52069=>"001001010",
  52070=>"000000110",
  52071=>"110011010",
  52072=>"011000100",
  52073=>"100000001",
  52074=>"000111010",
  52075=>"000010111",
  52076=>"101011111",
  52077=>"100000101",
  52078=>"101000011",
  52079=>"110110010",
  52080=>"100100010",
  52081=>"011001010",
  52082=>"011100110",
  52083=>"001000110",
  52084=>"110100100",
  52085=>"111110101",
  52086=>"011010001",
  52087=>"111000001",
  52088=>"010001000",
  52089=>"100111001",
  52090=>"101000101",
  52091=>"001111000",
  52092=>"011111000",
  52093=>"111100110",
  52094=>"110101101",
  52095=>"000100011",
  52096=>"100101010",
  52097=>"001101011",
  52098=>"001100110",
  52099=>"110010100",
  52100=>"100110110",
  52101=>"111010011",
  52102=>"100101011",
  52103=>"111000010",
  52104=>"111001011",
  52105=>"001111111",
  52106=>"111010010",
  52107=>"000100100",
  52108=>"010010001",
  52109=>"000110000",
  52110=>"010101001",
  52111=>"010001101",
  52112=>"111111010",
  52113=>"101110010",
  52114=>"110110100",
  52115=>"011011111",
  52116=>"001111111",
  52117=>"010001110",
  52118=>"111000000",
  52119=>"010100100",
  52120=>"110000011",
  52121=>"001010101",
  52122=>"111111100",
  52123=>"000110100",
  52124=>"001001011",
  52125=>"110101100",
  52126=>"001000010",
  52127=>"000100001",
  52128=>"011011001",
  52129=>"100010011",
  52130=>"101111001",
  52131=>"101100000",
  52132=>"010000011",
  52133=>"110101000",
  52134=>"110010101",
  52135=>"001000001",
  52136=>"011000111",
  52137=>"000000000",
  52138=>"101111001",
  52139=>"001100001",
  52140=>"101001111",
  52141=>"111001111",
  52142=>"001110111",
  52143=>"011110010",
  52144=>"110000000",
  52145=>"101101100",
  52146=>"101000001",
  52147=>"011100101",
  52148=>"000110011",
  52149=>"000000101",
  52150=>"110101010",
  52151=>"111001100",
  52152=>"010011001",
  52153=>"100010100",
  52154=>"000110001",
  52155=>"111001100",
  52156=>"010100011",
  52157=>"011011001",
  52158=>"110001110",
  52159=>"000100001",
  52160=>"000101011",
  52161=>"000011010",
  52162=>"011011110",
  52163=>"110011111",
  52164=>"010001110",
  52165=>"111100001",
  52166=>"111100000",
  52167=>"101011001",
  52168=>"110101010",
  52169=>"000110011",
  52170=>"010000000",
  52171=>"101111011",
  52172=>"001110110",
  52173=>"011111010",
  52174=>"000100100",
  52175=>"001011111",
  52176=>"010111011",
  52177=>"000011010",
  52178=>"100000101",
  52179=>"101111101",
  52180=>"111101101",
  52181=>"111110111",
  52182=>"010011100",
  52183=>"111110001",
  52184=>"001110100",
  52185=>"111100100",
  52186=>"000111000",
  52187=>"011000101",
  52188=>"000010000",
  52189=>"100111000",
  52190=>"111010011",
  52191=>"010000000",
  52192=>"001100011",
  52193=>"100011111",
  52194=>"011100000",
  52195=>"000011100",
  52196=>"100100101",
  52197=>"011100101",
  52198=>"001100110",
  52199=>"101101101",
  52200=>"100000100",
  52201=>"000000111",
  52202=>"000010111",
  52203=>"001010001",
  52204=>"100100000",
  52205=>"000000000",
  52206=>"101111001",
  52207=>"111101000",
  52208=>"101010010",
  52209=>"100000111",
  52210=>"101000111",
  52211=>"101011110",
  52212=>"010010100",
  52213=>"110100000",
  52214=>"111101100",
  52215=>"001101000",
  52216=>"101000011",
  52217=>"000101011",
  52218=>"001000110",
  52219=>"101111111",
  52220=>"010001101",
  52221=>"011001100",
  52222=>"101011111",
  52223=>"111101000",
  52224=>"010100100",
  52225=>"100101101",
  52226=>"110110000",
  52227=>"011010100",
  52228=>"101001101",
  52229=>"111111000",
  52230=>"011110011",
  52231=>"010101000",
  52232=>"101101010",
  52233=>"110010101",
  52234=>"011111011",
  52235=>"110011001",
  52236=>"110101011",
  52237=>"000011001",
  52238=>"100000001",
  52239=>"000011110",
  52240=>"110001000",
  52241=>"000001101",
  52242=>"100011111",
  52243=>"110010000",
  52244=>"111111001",
  52245=>"100111100",
  52246=>"111011111",
  52247=>"100111010",
  52248=>"001001111",
  52249=>"011101110",
  52250=>"100110100",
  52251=>"011001001",
  52252=>"111101011",
  52253=>"010010100",
  52254=>"011010010",
  52255=>"011000101",
  52256=>"001010111",
  52257=>"011011000",
  52258=>"101010111",
  52259=>"011110010",
  52260=>"010010010",
  52261=>"000011010",
  52262=>"001000101",
  52263=>"111100101",
  52264=>"000010010",
  52265=>"010001000",
  52266=>"000001011",
  52267=>"010011000",
  52268=>"001111100",
  52269=>"000001111",
  52270=>"110100101",
  52271=>"110101010",
  52272=>"010111101",
  52273=>"111101011",
  52274=>"010001010",
  52275=>"100010100",
  52276=>"000000100",
  52277=>"110011111",
  52278=>"100111101",
  52279=>"011000100",
  52280=>"101011011",
  52281=>"100010100",
  52282=>"110010001",
  52283=>"011111110",
  52284=>"011001111",
  52285=>"110001001",
  52286=>"101011101",
  52287=>"110110001",
  52288=>"111110100",
  52289=>"111111010",
  52290=>"011101101",
  52291=>"000111001",
  52292=>"100100010",
  52293=>"001100110",
  52294=>"111111101",
  52295=>"011000011",
  52296=>"101111101",
  52297=>"101010111",
  52298=>"001110100",
  52299=>"000101010",
  52300=>"001001100",
  52301=>"100000000",
  52302=>"010111011",
  52303=>"001000000",
  52304=>"101110100",
  52305=>"001010110",
  52306=>"011010000",
  52307=>"001001011",
  52308=>"010101000",
  52309=>"101111100",
  52310=>"100010100",
  52311=>"000110000",
  52312=>"111101100",
  52313=>"111010010",
  52314=>"100001000",
  52315=>"011110011",
  52316=>"010101111",
  52317=>"100111110",
  52318=>"101001111",
  52319=>"111110111",
  52320=>"000110011",
  52321=>"011001100",
  52322=>"100110000",
  52323=>"011101001",
  52324=>"000000111",
  52325=>"100101101",
  52326=>"000011110",
  52327=>"110100011",
  52328=>"001110011",
  52329=>"011111011",
  52330=>"010000000",
  52331=>"001100110",
  52332=>"011110010",
  52333=>"101001100",
  52334=>"110000110",
  52335=>"110010110",
  52336=>"011000010",
  52337=>"111110010",
  52338=>"110011010",
  52339=>"001011111",
  52340=>"110110011",
  52341=>"011010001",
  52342=>"111001011",
  52343=>"110000110",
  52344=>"011011100",
  52345=>"000001001",
  52346=>"110000111",
  52347=>"100010000",
  52348=>"011101110",
  52349=>"001011111",
  52350=>"011110011",
  52351=>"110001110",
  52352=>"100010100",
  52353=>"110011111",
  52354=>"010100010",
  52355=>"000111111",
  52356=>"111101011",
  52357=>"110010101",
  52358=>"110010000",
  52359=>"100011000",
  52360=>"111101110",
  52361=>"101000001",
  52362=>"010100000",
  52363=>"100111101",
  52364=>"000011111",
  52365=>"000011000",
  52366=>"110101111",
  52367=>"001000011",
  52368=>"011011011",
  52369=>"101010100",
  52370=>"010101100",
  52371=>"101100000",
  52372=>"010101110",
  52373=>"000111011",
  52374=>"000000100",
  52375=>"011110111",
  52376=>"110001010",
  52377=>"001100011",
  52378=>"011110101",
  52379=>"111111111",
  52380=>"001001001",
  52381=>"100010011",
  52382=>"011111010",
  52383=>"100001111",
  52384=>"110110111",
  52385=>"110101110",
  52386=>"000111100",
  52387=>"011001010",
  52388=>"011011001",
  52389=>"001101010",
  52390=>"010100001",
  52391=>"011010001",
  52392=>"010110110",
  52393=>"000100010",
  52394=>"000001111",
  52395=>"101001000",
  52396=>"010110001",
  52397=>"000011110",
  52398=>"111000010",
  52399=>"100011000",
  52400=>"111100110",
  52401=>"000010001",
  52402=>"101111100",
  52403=>"111011011",
  52404=>"101101111",
  52405=>"001011001",
  52406=>"100001101",
  52407=>"010000100",
  52408=>"010000100",
  52409=>"110011111",
  52410=>"010101000",
  52411=>"000001110",
  52412=>"000000110",
  52413=>"100111111",
  52414=>"000010001",
  52415=>"000001000",
  52416=>"001111101",
  52417=>"111000100",
  52418=>"100100011",
  52419=>"110000111",
  52420=>"000001001",
  52421=>"001101011",
  52422=>"111011010",
  52423=>"100101100",
  52424=>"101011110",
  52425=>"011001011",
  52426=>"010011000",
  52427=>"010001011",
  52428=>"110010000",
  52429=>"111011000",
  52430=>"110101001",
  52431=>"100101011",
  52432=>"010101011",
  52433=>"001011011",
  52434=>"010011110",
  52435=>"111011110",
  52436=>"011100110",
  52437=>"111110101",
  52438=>"110001011",
  52439=>"100100111",
  52440=>"001111001",
  52441=>"111001111",
  52442=>"110100101",
  52443=>"010100100",
  52444=>"011000101",
  52445=>"100000110",
  52446=>"011010011",
  52447=>"101100100",
  52448=>"111100010",
  52449=>"001110010",
  52450=>"010000011",
  52451=>"101001000",
  52452=>"100101100",
  52453=>"000011000",
  52454=>"110100001",
  52455=>"000010111",
  52456=>"101100000",
  52457=>"101010011",
  52458=>"011000100",
  52459=>"101100100",
  52460=>"110011111",
  52461=>"110100110",
  52462=>"101001001",
  52463=>"010111011",
  52464=>"100001110",
  52465=>"101000000",
  52466=>"000110001",
  52467=>"011101111",
  52468=>"111011010",
  52469=>"011111011",
  52470=>"011010101",
  52471=>"001100001",
  52472=>"001001100",
  52473=>"001111010",
  52474=>"000011000",
  52475=>"010111100",
  52476=>"110101110",
  52477=>"011001101",
  52478=>"100101001",
  52479=>"111010000",
  52480=>"000010111",
  52481=>"111111010",
  52482=>"111011010",
  52483=>"101010011",
  52484=>"011110111",
  52485=>"111000110",
  52486=>"000111010",
  52487=>"010011011",
  52488=>"110100001",
  52489=>"101111011",
  52490=>"100111111",
  52491=>"101010111",
  52492=>"101010111",
  52493=>"111011000",
  52494=>"011010010",
  52495=>"000000010",
  52496=>"000001100",
  52497=>"111110111",
  52498=>"011001000",
  52499=>"011110110",
  52500=>"111010011",
  52501=>"101111001",
  52502=>"010011100",
  52503=>"011101001",
  52504=>"011111001",
  52505=>"001111010",
  52506=>"010100111",
  52507=>"110110011",
  52508=>"101101100",
  52509=>"110010000",
  52510=>"001100010",
  52511=>"011111000",
  52512=>"111010001",
  52513=>"001011111",
  52514=>"011010010",
  52515=>"110010110",
  52516=>"100011000",
  52517=>"010001101",
  52518=>"000000110",
  52519=>"000110101",
  52520=>"001001000",
  52521=>"001110001",
  52522=>"110000010",
  52523=>"110101001",
  52524=>"000111011",
  52525=>"000000001",
  52526=>"111100111",
  52527=>"001010111",
  52528=>"101011111",
  52529=>"000101010",
  52530=>"101010100",
  52531=>"010110011",
  52532=>"101100001",
  52533=>"100000010",
  52534=>"000100101",
  52535=>"100100001",
  52536=>"101101101",
  52537=>"000010111",
  52538=>"101000101",
  52539=>"011100111",
  52540=>"001110000",
  52541=>"011110101",
  52542=>"100000000",
  52543=>"101110011",
  52544=>"100111111",
  52545=>"000100101",
  52546=>"010011110",
  52547=>"100111110",
  52548=>"110111111",
  52549=>"010000011",
  52550=>"001001101",
  52551=>"010110001",
  52552=>"010001000",
  52553=>"011010110",
  52554=>"110110010",
  52555=>"110000110",
  52556=>"110101001",
  52557=>"001100010",
  52558=>"100100000",
  52559=>"111101111",
  52560=>"100111001",
  52561=>"111100000",
  52562=>"001110000",
  52563=>"001111010",
  52564=>"001110111",
  52565=>"111010001",
  52566=>"011001001",
  52567=>"000100000",
  52568=>"111111111",
  52569=>"100010010",
  52570=>"100100011",
  52571=>"111111100",
  52572=>"011111111",
  52573=>"010010000",
  52574=>"010111111",
  52575=>"001101111",
  52576=>"111101000",
  52577=>"011110110",
  52578=>"101010101",
  52579=>"011100000",
  52580=>"101111000",
  52581=>"100101010",
  52582=>"000111010",
  52583=>"000111110",
  52584=>"011100101",
  52585=>"100001101",
  52586=>"010011101",
  52587=>"111100110",
  52588=>"011111011",
  52589=>"001111000",
  52590=>"101001101",
  52591=>"100100111",
  52592=>"101000011",
  52593=>"000110001",
  52594=>"110010100",
  52595=>"101101111",
  52596=>"101011011",
  52597=>"111111110",
  52598=>"111001101",
  52599=>"000011001",
  52600=>"100110001",
  52601=>"101000011",
  52602=>"101110000",
  52603=>"001101010",
  52604=>"011111000",
  52605=>"001110010",
  52606=>"001001111",
  52607=>"101101100",
  52608=>"100110010",
  52609=>"010100010",
  52610=>"110100111",
  52611=>"101011000",
  52612=>"110101110",
  52613=>"100001111",
  52614=>"101000110",
  52615=>"110000001",
  52616=>"010110101",
  52617=>"111100010",
  52618=>"011001000",
  52619=>"000111111",
  52620=>"001100110",
  52621=>"100000011",
  52622=>"010000100",
  52623=>"011110010",
  52624=>"000101101",
  52625=>"100000010",
  52626=>"111011010",
  52627=>"011110100",
  52628=>"101010111",
  52629=>"101111101",
  52630=>"100001110",
  52631=>"011111011",
  52632=>"110001010",
  52633=>"100011010",
  52634=>"110000011",
  52635=>"110101110",
  52636=>"100011101",
  52637=>"100111110",
  52638=>"001110011",
  52639=>"001001101",
  52640=>"001011111",
  52641=>"011001001",
  52642=>"100001111",
  52643=>"110010001",
  52644=>"000111000",
  52645=>"001011100",
  52646=>"000011000",
  52647=>"100100001",
  52648=>"000011011",
  52649=>"010000100",
  52650=>"010111111",
  52651=>"111111110",
  52652=>"110011101",
  52653=>"111111011",
  52654=>"101111100",
  52655=>"101110101",
  52656=>"011111101",
  52657=>"000000010",
  52658=>"111000100",
  52659=>"010000001",
  52660=>"111111110",
  52661=>"000111110",
  52662=>"110110000",
  52663=>"111100111",
  52664=>"001011011",
  52665=>"001010011",
  52666=>"001110001",
  52667=>"010011000",
  52668=>"010011111",
  52669=>"011001100",
  52670=>"000111101",
  52671=>"001001100",
  52672=>"000111010",
  52673=>"110011000",
  52674=>"011110101",
  52675=>"010100101",
  52676=>"111100011",
  52677=>"100001100",
  52678=>"000100100",
  52679=>"111100001",
  52680=>"111000111",
  52681=>"011111100",
  52682=>"110011110",
  52683=>"001010101",
  52684=>"011110000",
  52685=>"001001100",
  52686=>"110110111",
  52687=>"011010100",
  52688=>"011011001",
  52689=>"110101011",
  52690=>"011010110",
  52691=>"101111101",
  52692=>"101110110",
  52693=>"111011111",
  52694=>"011101111",
  52695=>"011111000",
  52696=>"110011001",
  52697=>"000100001",
  52698=>"010100100",
  52699=>"001101100",
  52700=>"010111011",
  52701=>"110100100",
  52702=>"110001100",
  52703=>"010001001",
  52704=>"110000110",
  52705=>"001110010",
  52706=>"000010100",
  52707=>"001010001",
  52708=>"010000100",
  52709=>"101000110",
  52710=>"000011011",
  52711=>"011001010",
  52712=>"100101110",
  52713=>"010011101",
  52714=>"000110100",
  52715=>"111100101",
  52716=>"100101001",
  52717=>"111101101",
  52718=>"010011001",
  52719=>"000010011",
  52720=>"010100010",
  52721=>"011011000",
  52722=>"100110011",
  52723=>"000010000",
  52724=>"110101001",
  52725=>"000001100",
  52726=>"000011010",
  52727=>"100100100",
  52728=>"101011101",
  52729=>"100001100",
  52730=>"010000101",
  52731=>"100000001",
  52732=>"000101100",
  52733=>"101111010",
  52734=>"101100110",
  52735=>"110101010",
  52736=>"010000111",
  52737=>"100101011",
  52738=>"010110110",
  52739=>"011001001",
  52740=>"001011001",
  52741=>"101000111",
  52742=>"110000100",
  52743=>"111010111",
  52744=>"101110001",
  52745=>"001010110",
  52746=>"110001111",
  52747=>"001111001",
  52748=>"100010110",
  52749=>"100100001",
  52750=>"100000010",
  52751=>"000101101",
  52752=>"100101001",
  52753=>"000100110",
  52754=>"010011110",
  52755=>"111100100",
  52756=>"000000000",
  52757=>"100000001",
  52758=>"101101111",
  52759=>"000100110",
  52760=>"001110010",
  52761=>"111000110",
  52762=>"101110100",
  52763=>"101011111",
  52764=>"111000110",
  52765=>"100000110",
  52766=>"010101000",
  52767=>"001011000",
  52768=>"110110110",
  52769=>"011110101",
  52770=>"111000100",
  52771=>"110101000",
  52772=>"000111101",
  52773=>"001110111",
  52774=>"111111110",
  52775=>"111011101",
  52776=>"101001001",
  52777=>"100011010",
  52778=>"111011100",
  52779=>"011011111",
  52780=>"100010000",
  52781=>"000101101",
  52782=>"011111000",
  52783=>"010000010",
  52784=>"110101110",
  52785=>"110100011",
  52786=>"011000111",
  52787=>"000011110",
  52788=>"100101111",
  52789=>"111100011",
  52790=>"001111011",
  52791=>"011000010",
  52792=>"011101111",
  52793=>"111110011",
  52794=>"011110101",
  52795=>"010010010",
  52796=>"101100100",
  52797=>"111001001",
  52798=>"111010100",
  52799=>"100101101",
  52800=>"010001011",
  52801=>"110101111",
  52802=>"010100101",
  52803=>"011110101",
  52804=>"100110111",
  52805=>"101110101",
  52806=>"011111111",
  52807=>"101101011",
  52808=>"000000010",
  52809=>"111010111",
  52810=>"100101011",
  52811=>"001000001",
  52812=>"010000001",
  52813=>"000000100",
  52814=>"110101001",
  52815=>"110111010",
  52816=>"000000001",
  52817=>"000110010",
  52818=>"101100000",
  52819=>"110001101",
  52820=>"111110111",
  52821=>"011111000",
  52822=>"000100100",
  52823=>"010110100",
  52824=>"111111010",
  52825=>"100111010",
  52826=>"111110011",
  52827=>"011111001",
  52828=>"101000111",
  52829=>"001010001",
  52830=>"001010101",
  52831=>"010001111",
  52832=>"010001110",
  52833=>"111100011",
  52834=>"101000001",
  52835=>"100001100",
  52836=>"101101010",
  52837=>"001001010",
  52838=>"100001100",
  52839=>"001111101",
  52840=>"001111010",
  52841=>"100110001",
  52842=>"010000001",
  52843=>"111100110",
  52844=>"000110111",
  52845=>"000001010",
  52846=>"100111110",
  52847=>"100000000",
  52848=>"011000000",
  52849=>"011001000",
  52850=>"010011010",
  52851=>"110110000",
  52852=>"101100101",
  52853=>"011000101",
  52854=>"111100000",
  52855=>"010001100",
  52856=>"101101011",
  52857=>"010000101",
  52858=>"011011111",
  52859=>"011011100",
  52860=>"101011010",
  52861=>"110011010",
  52862=>"100000011",
  52863=>"011100111",
  52864=>"101010101",
  52865=>"001111101",
  52866=>"111100111",
  52867=>"100110000",
  52868=>"110001111",
  52869=>"111011001",
  52870=>"101010110",
  52871=>"000010100",
  52872=>"000100101",
  52873=>"010000111",
  52874=>"010010101",
  52875=>"010111011",
  52876=>"010001101",
  52877=>"110001011",
  52878=>"101111100",
  52879=>"101111101",
  52880=>"010111010",
  52881=>"001110111",
  52882=>"111000110",
  52883=>"100110111",
  52884=>"001001011",
  52885=>"111100101",
  52886=>"000110110",
  52887=>"101001000",
  52888=>"110100101",
  52889=>"110000010",
  52890=>"101101110",
  52891=>"111110110",
  52892=>"000100111",
  52893=>"010011001",
  52894=>"000000000",
  52895=>"011100010",
  52896=>"111111101",
  52897=>"111111001",
  52898=>"101111101",
  52899=>"101000100",
  52900=>"111010001",
  52901=>"000001000",
  52902=>"110111010",
  52903=>"110100100",
  52904=>"000101100",
  52905=>"000100111",
  52906=>"110000101",
  52907=>"100101000",
  52908=>"001010101",
  52909=>"100000101",
  52910=>"010111011",
  52911=>"110100001",
  52912=>"100010000",
  52913=>"110110110",
  52914=>"011011011",
  52915=>"000010010",
  52916=>"101110000",
  52917=>"101111100",
  52918=>"111101101",
  52919=>"001111011",
  52920=>"100010111",
  52921=>"111000010",
  52922=>"000111000",
  52923=>"010010010",
  52924=>"111100011",
  52925=>"001110010",
  52926=>"110000100",
  52927=>"001001010",
  52928=>"101000000",
  52929=>"101101011",
  52930=>"111110110",
  52931=>"100110011",
  52932=>"011100011",
  52933=>"000001000",
  52934=>"111101010",
  52935=>"011101111",
  52936=>"011111101",
  52937=>"100010010",
  52938=>"100000000",
  52939=>"000100111",
  52940=>"011010010",
  52941=>"001000010",
  52942=>"111011010",
  52943=>"000010111",
  52944=>"100011001",
  52945=>"010001001",
  52946=>"011000101",
  52947=>"101000000",
  52948=>"000101010",
  52949=>"111101001",
  52950=>"010000110",
  52951=>"001001000",
  52952=>"001001011",
  52953=>"000110010",
  52954=>"011110000",
  52955=>"001001011",
  52956=>"001000101",
  52957=>"101010000",
  52958=>"011001110",
  52959=>"110100011",
  52960=>"001011101",
  52961=>"000100010",
  52962=>"111000011",
  52963=>"001001101",
  52964=>"101001101",
  52965=>"101100100",
  52966=>"000010101",
  52967=>"110010000",
  52968=>"101111011",
  52969=>"101100010",
  52970=>"000110100",
  52971=>"001101011",
  52972=>"100010001",
  52973=>"100010110",
  52974=>"110011111",
  52975=>"000011000",
  52976=>"010111111",
  52977=>"000101111",
  52978=>"110001100",
  52979=>"110010011",
  52980=>"111000010",
  52981=>"010101011",
  52982=>"100111101",
  52983=>"001010101",
  52984=>"110010110",
  52985=>"011010110",
  52986=>"000010110",
  52987=>"010111011",
  52988=>"001111001",
  52989=>"110100000",
  52990=>"111101010",
  52991=>"000101111",
  52992=>"001000100",
  52993=>"000010011",
  52994=>"111111111",
  52995=>"001000100",
  52996=>"010111011",
  52997=>"100011101",
  52998=>"011000100",
  52999=>"000000111",
  53000=>"111110011",
  53001=>"010111010",
  53002=>"111100101",
  53003=>"001000101",
  53004=>"100110011",
  53005=>"001011101",
  53006=>"000100101",
  53007=>"001001100",
  53008=>"100001010",
  53009=>"010110001",
  53010=>"000100110",
  53011=>"001011110",
  53012=>"010101100",
  53013=>"001000101",
  53014=>"110100000",
  53015=>"111001010",
  53016=>"110100111",
  53017=>"001001011",
  53018=>"000111110",
  53019=>"101110100",
  53020=>"110100101",
  53021=>"110101111",
  53022=>"111101010",
  53023=>"101001100",
  53024=>"011101111",
  53025=>"110010100",
  53026=>"111100111",
  53027=>"101000111",
  53028=>"011110011",
  53029=>"010100101",
  53030=>"100110010",
  53031=>"010000101",
  53032=>"101000111",
  53033=>"001100001",
  53034=>"011111010",
  53035=>"110011001",
  53036=>"110011010",
  53037=>"010010011",
  53038=>"101100011",
  53039=>"111111011",
  53040=>"010001101",
  53041=>"101101100",
  53042=>"100101010",
  53043=>"110011101",
  53044=>"000110001",
  53045=>"000110100",
  53046=>"111011010",
  53047=>"101101011",
  53048=>"100100110",
  53049=>"010000001",
  53050=>"101001101",
  53051=>"100000110",
  53052=>"110111001",
  53053=>"001110010",
  53054=>"010100101",
  53055=>"101010000",
  53056=>"000100110",
  53057=>"100101000",
  53058=>"111111010",
  53059=>"100010111",
  53060=>"101101100",
  53061=>"110001010",
  53062=>"110001000",
  53063=>"011110000",
  53064=>"010011011",
  53065=>"001010001",
  53066=>"010010111",
  53067=>"001010111",
  53068=>"111001101",
  53069=>"001100010",
  53070=>"011011101",
  53071=>"010101011",
  53072=>"011110011",
  53073=>"010000011",
  53074=>"000101000",
  53075=>"101101001",
  53076=>"110100011",
  53077=>"100011001",
  53078=>"001101010",
  53079=>"001100001",
  53080=>"101010001",
  53081=>"001010000",
  53082=>"110111000",
  53083=>"010001111",
  53084=>"000100111",
  53085=>"100001010",
  53086=>"001011111",
  53087=>"000101000",
  53088=>"001000000",
  53089=>"110001000",
  53090=>"001000101",
  53091=>"110100001",
  53092=>"011111110",
  53093=>"001011010",
  53094=>"111101111",
  53095=>"000101111",
  53096=>"100110011",
  53097=>"111101001",
  53098=>"111101110",
  53099=>"111000001",
  53100=>"000101101",
  53101=>"000001110",
  53102=>"110111110",
  53103=>"101100001",
  53104=>"001010100",
  53105=>"010000001",
  53106=>"101010000",
  53107=>"010101010",
  53108=>"001110001",
  53109=>"000011010",
  53110=>"011011001",
  53111=>"111000101",
  53112=>"100110010",
  53113=>"010100101",
  53114=>"000001100",
  53115=>"010110011",
  53116=>"010000001",
  53117=>"010001000",
  53118=>"000100100",
  53119=>"110100001",
  53120=>"111010000",
  53121=>"111010101",
  53122=>"111110111",
  53123=>"101000110",
  53124=>"010101001",
  53125=>"100011001",
  53126=>"011011110",
  53127=>"111100011",
  53128=>"000000000",
  53129=>"000110100",
  53130=>"100111000",
  53131=>"111110111",
  53132=>"111110010",
  53133=>"100010001",
  53134=>"010011000",
  53135=>"111000100",
  53136=>"101010000",
  53137=>"111111111",
  53138=>"110000101",
  53139=>"001000000",
  53140=>"110111000",
  53141=>"000000011",
  53142=>"110110100",
  53143=>"001010110",
  53144=>"000010110",
  53145=>"000110000",
  53146=>"110010110",
  53147=>"001011100",
  53148=>"110001100",
  53149=>"000000000",
  53150=>"000000011",
  53151=>"111011110",
  53152=>"010011101",
  53153=>"101111110",
  53154=>"010010000",
  53155=>"110011001",
  53156=>"010111110",
  53157=>"110110110",
  53158=>"010111111",
  53159=>"100010101",
  53160=>"110001101",
  53161=>"100010010",
  53162=>"001110111",
  53163=>"011111010",
  53164=>"010111011",
  53165=>"010000011",
  53166=>"111011110",
  53167=>"010101010",
  53168=>"111000100",
  53169=>"010001100",
  53170=>"110110110",
  53171=>"000001000",
  53172=>"111011100",
  53173=>"001110111",
  53174=>"101110101",
  53175=>"101011100",
  53176=>"110101010",
  53177=>"011001101",
  53178=>"000101001",
  53179=>"101011101",
  53180=>"111100111",
  53181=>"001100000",
  53182=>"101111001",
  53183=>"111101110",
  53184=>"100010011",
  53185=>"011011101",
  53186=>"001100001",
  53187=>"111111011",
  53188=>"010100101",
  53189=>"100011000",
  53190=>"101110001",
  53191=>"001111111",
  53192=>"101000000",
  53193=>"110000111",
  53194=>"000001110",
  53195=>"011111101",
  53196=>"111000011",
  53197=>"100100111",
  53198=>"001110011",
  53199=>"000101010",
  53200=>"111000111",
  53201=>"000010110",
  53202=>"010011011",
  53203=>"001100000",
  53204=>"000011111",
  53205=>"010010011",
  53206=>"111010000",
  53207=>"001110001",
  53208=>"111100000",
  53209=>"010000110",
  53210=>"101011101",
  53211=>"001101011",
  53212=>"100100101",
  53213=>"101101101",
  53214=>"101001000",
  53215=>"100100110",
  53216=>"100001110",
  53217=>"010101101",
  53218=>"100100100",
  53219=>"110011001",
  53220=>"100100000",
  53221=>"010101100",
  53222=>"010110101",
  53223=>"100100000",
  53224=>"000000100",
  53225=>"101111010",
  53226=>"000100010",
  53227=>"001000111",
  53228=>"111010100",
  53229=>"001000000",
  53230=>"100011011",
  53231=>"011101101",
  53232=>"000000001",
  53233=>"010011100",
  53234=>"000001100",
  53235=>"010010000",
  53236=>"011101000",
  53237=>"110011000",
  53238=>"010000110",
  53239=>"101001101",
  53240=>"000101101",
  53241=>"111111100",
  53242=>"000010111",
  53243=>"111101110",
  53244=>"110100110",
  53245=>"110101100",
  53246=>"111011001",
  53247=>"010011100",
  53248=>"100110000",
  53249=>"101101110",
  53250=>"010110001",
  53251=>"111010110",
  53252=>"001111010",
  53253=>"101111000",
  53254=>"001000110",
  53255=>"111100101",
  53256=>"110101000",
  53257=>"010100001",
  53258=>"001111110",
  53259=>"111110011",
  53260=>"010110100",
  53261=>"001001111",
  53262=>"010011101",
  53263=>"000111001",
  53264=>"101100010",
  53265=>"110001111",
  53266=>"011110111",
  53267=>"111001010",
  53268=>"100011101",
  53269=>"111000101",
  53270=>"000110100",
  53271=>"010010000",
  53272=>"011001001",
  53273=>"001010100",
  53274=>"100010111",
  53275=>"001101000",
  53276=>"011101111",
  53277=>"101101011",
  53278=>"000010001",
  53279=>"001001111",
  53280=>"111011011",
  53281=>"000100101",
  53282=>"010000000",
  53283=>"100111001",
  53284=>"000000111",
  53285=>"110101111",
  53286=>"110110000",
  53287=>"010110111",
  53288=>"011011000",
  53289=>"001011000",
  53290=>"011010100",
  53291=>"000011110",
  53292=>"110100101",
  53293=>"000110000",
  53294=>"101101101",
  53295=>"000110110",
  53296=>"010000000",
  53297=>"001011110",
  53298=>"101111001",
  53299=>"001011010",
  53300=>"100101000",
  53301=>"001010111",
  53302=>"011011110",
  53303=>"100111111",
  53304=>"000100011",
  53305=>"000000100",
  53306=>"101011111",
  53307=>"001100000",
  53308=>"001100000",
  53309=>"010011011",
  53310=>"000110111",
  53311=>"111100110",
  53312=>"010000011",
  53313=>"001100001",
  53314=>"101010011",
  53315=>"000110011",
  53316=>"010001101",
  53317=>"100111001",
  53318=>"000101000",
  53319=>"101011101",
  53320=>"011010101",
  53321=>"011110011",
  53322=>"100001001",
  53323=>"001011010",
  53324=>"001110100",
  53325=>"110111101",
  53326=>"110011010",
  53327=>"011000111",
  53328=>"010101001",
  53329=>"110110011",
  53330=>"011011011",
  53331=>"101010011",
  53332=>"011101001",
  53333=>"011010001",
  53334=>"111100111",
  53335=>"101100001",
  53336=>"010101111",
  53337=>"111111111",
  53338=>"010000111",
  53339=>"001010010",
  53340=>"001000010",
  53341=>"101100111",
  53342=>"011101111",
  53343=>"111101101",
  53344=>"001011100",
  53345=>"010100110",
  53346=>"011001101",
  53347=>"111011000",
  53348=>"101001101",
  53349=>"111000101",
  53350=>"000110010",
  53351=>"011111000",
  53352=>"100101000",
  53353=>"100011111",
  53354=>"110011111",
  53355=>"111110000",
  53356=>"011010110",
  53357=>"010100010",
  53358=>"111101100",
  53359=>"101011010",
  53360=>"110100011",
  53361=>"110011011",
  53362=>"101000001",
  53363=>"111000001",
  53364=>"011110010",
  53365=>"100110000",
  53366=>"111001000",
  53367=>"110000111",
  53368=>"001111101",
  53369=>"001111001",
  53370=>"101011001",
  53371=>"101011101",
  53372=>"001001001",
  53373=>"011010010",
  53374=>"100010101",
  53375=>"010111110",
  53376=>"110001000",
  53377=>"000100001",
  53378=>"001011110",
  53379=>"000011100",
  53380=>"100001000",
  53381=>"101111111",
  53382=>"000111101",
  53383=>"111110000",
  53384=>"010000110",
  53385=>"000111010",
  53386=>"111001000",
  53387=>"111110001",
  53388=>"010001101",
  53389=>"100001110",
  53390=>"011000110",
  53391=>"010101000",
  53392=>"100011111",
  53393=>"110010111",
  53394=>"110110010",
  53395=>"011010000",
  53396=>"001101000",
  53397=>"110011011",
  53398=>"110010000",
  53399=>"110111111",
  53400=>"010000011",
  53401=>"001001111",
  53402=>"101111010",
  53403=>"110110111",
  53404=>"000100111",
  53405=>"000001101",
  53406=>"001100101",
  53407=>"111100101",
  53408=>"010000100",
  53409=>"110101001",
  53410=>"001011101",
  53411=>"101101111",
  53412=>"001111010",
  53413=>"110100100",
  53414=>"101101010",
  53415=>"011010011",
  53416=>"110010110",
  53417=>"001101010",
  53418=>"001110000",
  53419=>"101001000",
  53420=>"011100110",
  53421=>"000000000",
  53422=>"110000101",
  53423=>"100110000",
  53424=>"111110101",
  53425=>"011111010",
  53426=>"110101100",
  53427=>"110101111",
  53428=>"110001011",
  53429=>"000010101",
  53430=>"100111001",
  53431=>"001110000",
  53432=>"100000010",
  53433=>"001001000",
  53434=>"001101001",
  53435=>"101000000",
  53436=>"000111000",
  53437=>"011000011",
  53438=>"000001100",
  53439=>"110000100",
  53440=>"111111100",
  53441=>"000011011",
  53442=>"010001100",
  53443=>"110101001",
  53444=>"111000001",
  53445=>"001100011",
  53446=>"111101010",
  53447=>"000110011",
  53448=>"100100001",
  53449=>"000010010",
  53450=>"100000011",
  53451=>"111001111",
  53452=>"111001111",
  53453=>"010111111",
  53454=>"100110101",
  53455=>"010000010",
  53456=>"010011100",
  53457=>"010011011",
  53458=>"101010101",
  53459=>"101010010",
  53460=>"010110011",
  53461=>"001111000",
  53462=>"010011100",
  53463=>"010101101",
  53464=>"111111001",
  53465=>"001001101",
  53466=>"110000011",
  53467=>"001100000",
  53468=>"111011000",
  53469=>"001011011",
  53470=>"001001111",
  53471=>"101110010",
  53472=>"110001000",
  53473=>"111101010",
  53474=>"100010101",
  53475=>"010010110",
  53476=>"001110111",
  53477=>"010011111",
  53478=>"011011111",
  53479=>"111011111",
  53480=>"000110101",
  53481=>"001100110",
  53482=>"000000000",
  53483=>"001100011",
  53484=>"100010000",
  53485=>"001100110",
  53486=>"011011010",
  53487=>"001100001",
  53488=>"011101010",
  53489=>"011110000",
  53490=>"000011001",
  53491=>"010000110",
  53492=>"001110000",
  53493=>"000111010",
  53494=>"111100010",
  53495=>"100010101",
  53496=>"011010001",
  53497=>"111111101",
  53498=>"110001000",
  53499=>"000001001",
  53500=>"010001100",
  53501=>"000100000",
  53502=>"111100111",
  53503=>"010001001",
  53504=>"110011011",
  53505=>"111010001",
  53506=>"000011011",
  53507=>"100111100",
  53508=>"111100111",
  53509=>"001110100",
  53510=>"101101100",
  53511=>"110101110",
  53512=>"011010010",
  53513=>"000100001",
  53514=>"001111010",
  53515=>"100001101",
  53516=>"000010011",
  53517=>"110100010",
  53518=>"011010010",
  53519=>"011010111",
  53520=>"101100110",
  53521=>"000011011",
  53522=>"101110110",
  53523=>"100101011",
  53524=>"101000011",
  53525=>"001111100",
  53526=>"011011101",
  53527=>"000001100",
  53528=>"110110011",
  53529=>"001001011",
  53530=>"111111111",
  53531=>"011000010",
  53532=>"101000011",
  53533=>"110001001",
  53534=>"100101010",
  53535=>"100000001",
  53536=>"000001110",
  53537=>"101000100",
  53538=>"100011111",
  53539=>"110101100",
  53540=>"110000001",
  53541=>"001110110",
  53542=>"001011001",
  53543=>"000001100",
  53544=>"001101111",
  53545=>"010010010",
  53546=>"101100110",
  53547=>"000101010",
  53548=>"010101011",
  53549=>"100011001",
  53550=>"000000000",
  53551=>"010001111",
  53552=>"000100010",
  53553=>"011101000",
  53554=>"101011100",
  53555=>"000010101",
  53556=>"011010011",
  53557=>"101010010",
  53558=>"011001001",
  53559=>"111000100",
  53560=>"000000011",
  53561=>"001100011",
  53562=>"100011010",
  53563=>"010101100",
  53564=>"100010000",
  53565=>"110000011",
  53566=>"010000111",
  53567=>"101010000",
  53568=>"111000010",
  53569=>"100011101",
  53570=>"000100000",
  53571=>"110100000",
  53572=>"110100100",
  53573=>"100011101",
  53574=>"010111000",
  53575=>"001111110",
  53576=>"011100011",
  53577=>"000010001",
  53578=>"010100100",
  53579=>"001000000",
  53580=>"000011000",
  53581=>"110100100",
  53582=>"010000111",
  53583=>"111101111",
  53584=>"111111111",
  53585=>"101111011",
  53586=>"100000010",
  53587=>"011111100",
  53588=>"000011110",
  53589=>"111010111",
  53590=>"010111111",
  53591=>"100010111",
  53592=>"110100101",
  53593=>"000101111",
  53594=>"110011111",
  53595=>"101100011",
  53596=>"111010000",
  53597=>"001110000",
  53598=>"011111101",
  53599=>"000100100",
  53600=>"011111001",
  53601=>"111011010",
  53602=>"001101001",
  53603=>"000001001",
  53604=>"101111110",
  53605=>"011110111",
  53606=>"110101111",
  53607=>"110011001",
  53608=>"101101111",
  53609=>"000100111",
  53610=>"000000000",
  53611=>"000010010",
  53612=>"110011110",
  53613=>"000010110",
  53614=>"000000111",
  53615=>"100111001",
  53616=>"000011110",
  53617=>"100101011",
  53618=>"101110011",
  53619=>"110110111",
  53620=>"011101101",
  53621=>"001010110",
  53622=>"011010100",
  53623=>"001000111",
  53624=>"011000000",
  53625=>"010001011",
  53626=>"110010111",
  53627=>"101011001",
  53628=>"100100110",
  53629=>"110111100",
  53630=>"011111011",
  53631=>"111001100",
  53632=>"000100011",
  53633=>"001101001",
  53634=>"011111010",
  53635=>"011101111",
  53636=>"111100111",
  53637=>"001000100",
  53638=>"010100010",
  53639=>"110110000",
  53640=>"000010010",
  53641=>"110100111",
  53642=>"010010011",
  53643=>"001100110",
  53644=>"010011101",
  53645=>"001000111",
  53646=>"100011000",
  53647=>"101011001",
  53648=>"000000110",
  53649=>"101100111",
  53650=>"010001111",
  53651=>"011101100",
  53652=>"111100010",
  53653=>"011001010",
  53654=>"001001001",
  53655=>"001010101",
  53656=>"101011010",
  53657=>"001000010",
  53658=>"001100111",
  53659=>"011010010",
  53660=>"001000010",
  53661=>"010110011",
  53662=>"010011100",
  53663=>"001001011",
  53664=>"011010000",
  53665=>"111010010",
  53666=>"010111011",
  53667=>"010101111",
  53668=>"111100100",
  53669=>"011101011",
  53670=>"100000010",
  53671=>"111100101",
  53672=>"100100110",
  53673=>"110011000",
  53674=>"101001110",
  53675=>"001000001",
  53676=>"000001110",
  53677=>"001111010",
  53678=>"110111011",
  53679=>"101010001",
  53680=>"100001001",
  53681=>"110000000",
  53682=>"101110001",
  53683=>"001011110",
  53684=>"111011111",
  53685=>"101011101",
  53686=>"011000111",
  53687=>"101010110",
  53688=>"111101111",
  53689=>"110010000",
  53690=>"000100110",
  53691=>"010111011",
  53692=>"000111001",
  53693=>"011100111",
  53694=>"010000111",
  53695=>"100001101",
  53696=>"000001001",
  53697=>"101101011",
  53698=>"101111100",
  53699=>"110101100",
  53700=>"001001000",
  53701=>"111101111",
  53702=>"111100000",
  53703=>"001000001",
  53704=>"010010111",
  53705=>"100111110",
  53706=>"001101010",
  53707=>"001111010",
  53708=>"010110100",
  53709=>"100100111",
  53710=>"000101000",
  53711=>"100010001",
  53712=>"100110111",
  53713=>"000010000",
  53714=>"011011011",
  53715=>"000000000",
  53716=>"111010111",
  53717=>"100101000",
  53718=>"010010000",
  53719=>"001011010",
  53720=>"011001000",
  53721=>"011110101",
  53722=>"100001110",
  53723=>"010001101",
  53724=>"111101011",
  53725=>"001000001",
  53726=>"100100001",
  53727=>"100111111",
  53728=>"111101000",
  53729=>"111101000",
  53730=>"000111111",
  53731=>"101000110",
  53732=>"101101110",
  53733=>"000110000",
  53734=>"111001010",
  53735=>"000100010",
  53736=>"110100111",
  53737=>"011001000",
  53738=>"101100000",
  53739=>"000111101",
  53740=>"001000111",
  53741=>"111111000",
  53742=>"101111001",
  53743=>"100101001",
  53744=>"000110111",
  53745=>"100101111",
  53746=>"101011110",
  53747=>"010100000",
  53748=>"110100000",
  53749=>"110110101",
  53750=>"110111011",
  53751=>"101011011",
  53752=>"110010001",
  53753=>"111111101",
  53754=>"100000100",
  53755=>"010001000",
  53756=>"011011101",
  53757=>"110000010",
  53758=>"101110111",
  53759=>"111001100",
  53760=>"010011001",
  53761=>"001111110",
  53762=>"011101100",
  53763=>"001001101",
  53764=>"101110000",
  53765=>"001101101",
  53766=>"110100010",
  53767=>"011101100",
  53768=>"011010100",
  53769=>"011001111",
  53770=>"101001110",
  53771=>"010110111",
  53772=>"110000100",
  53773=>"110100110",
  53774=>"000111111",
  53775=>"001100011",
  53776=>"001001110",
  53777=>"101100111",
  53778=>"110111011",
  53779=>"110011111",
  53780=>"100100111",
  53781=>"110010001",
  53782=>"010101000",
  53783=>"000111111",
  53784=>"001101010",
  53785=>"001010010",
  53786=>"011001100",
  53787=>"110110101",
  53788=>"000011011",
  53789=>"100000110",
  53790=>"011100001",
  53791=>"000111000",
  53792=>"011011111",
  53793=>"001111011",
  53794=>"010001011",
  53795=>"110101000",
  53796=>"011010011",
  53797=>"110100101",
  53798=>"110110100",
  53799=>"100010000",
  53800=>"000001110",
  53801=>"000011010",
  53802=>"010110011",
  53803=>"101010000",
  53804=>"010000100",
  53805=>"110001111",
  53806=>"000001000",
  53807=>"001100110",
  53808=>"011100101",
  53809=>"110001111",
  53810=>"011100001",
  53811=>"101000000",
  53812=>"101010000",
  53813=>"010101110",
  53814=>"000100101",
  53815=>"110010110",
  53816=>"000110111",
  53817=>"100001001",
  53818=>"110111100",
  53819=>"011100111",
  53820=>"000101100",
  53821=>"010010000",
  53822=>"100010000",
  53823=>"001000111",
  53824=>"010001100",
  53825=>"111000011",
  53826=>"011000000",
  53827=>"001010011",
  53828=>"000000000",
  53829=>"011100100",
  53830=>"101001100",
  53831=>"010111101",
  53832=>"001000000",
  53833=>"110011101",
  53834=>"110010111",
  53835=>"001110000",
  53836=>"011101101",
  53837=>"101010100",
  53838=>"010101010",
  53839=>"101001001",
  53840=>"111001111",
  53841=>"011101010",
  53842=>"101000001",
  53843=>"101000010",
  53844=>"010101100",
  53845=>"001010001",
  53846=>"000001111",
  53847=>"001100110",
  53848=>"000100100",
  53849=>"100010000",
  53850=>"110100000",
  53851=>"000000110",
  53852=>"001111101",
  53853=>"100001110",
  53854=>"000111100",
  53855=>"001100011",
  53856=>"011110100",
  53857=>"010001110",
  53858=>"101101100",
  53859=>"001011010",
  53860=>"100001011",
  53861=>"101110101",
  53862=>"101110100",
  53863=>"001000100",
  53864=>"010010010",
  53865=>"111011010",
  53866=>"111000011",
  53867=>"001110100",
  53868=>"000110001",
  53869=>"111000110",
  53870=>"111000010",
  53871=>"110000000",
  53872=>"011000110",
  53873=>"001001011",
  53874=>"100110010",
  53875=>"101100001",
  53876=>"000101110",
  53877=>"000010100",
  53878=>"100010011",
  53879=>"000010111",
  53880=>"111101100",
  53881=>"010011000",
  53882=>"000000010",
  53883=>"000001101",
  53884=>"011111001",
  53885=>"101011100",
  53886=>"100010010",
  53887=>"111101110",
  53888=>"001011101",
  53889=>"111010111",
  53890=>"101001110",
  53891=>"000010010",
  53892=>"010101110",
  53893=>"100101001",
  53894=>"110011110",
  53895=>"110010111",
  53896=>"111000101",
  53897=>"011001011",
  53898=>"100001101",
  53899=>"110001101",
  53900=>"011000001",
  53901=>"000001011",
  53902=>"000101101",
  53903=>"000011001",
  53904=>"111100001",
  53905=>"110111111",
  53906=>"101111111",
  53907=>"001001111",
  53908=>"000111011",
  53909=>"100001111",
  53910=>"111001011",
  53911=>"101011011",
  53912=>"110111001",
  53913=>"100110101",
  53914=>"100010001",
  53915=>"101100100",
  53916=>"100101010",
  53917=>"010001011",
  53918=>"010010101",
  53919=>"000000110",
  53920=>"010101011",
  53921=>"011001001",
  53922=>"100111101",
  53923=>"101001011",
  53924=>"001000100",
  53925=>"010101101",
  53926=>"010010101",
  53927=>"001010010",
  53928=>"111101011",
  53929=>"010100001",
  53930=>"110100001",
  53931=>"111100000",
  53932=>"100110100",
  53933=>"111100001",
  53934=>"010001100",
  53935=>"001100011",
  53936=>"011110111",
  53937=>"010011010",
  53938=>"011001001",
  53939=>"001011101",
  53940=>"011101000",
  53941=>"100000011",
  53942=>"011001101",
  53943=>"101001101",
  53944=>"001000110",
  53945=>"110010000",
  53946=>"001011010",
  53947=>"011101100",
  53948=>"011111101",
  53949=>"001001011",
  53950=>"001001101",
  53951=>"100101101",
  53952=>"111011001",
  53953=>"101011111",
  53954=>"001100100",
  53955=>"100100000",
  53956=>"100100010",
  53957=>"100111110",
  53958=>"110101011",
  53959=>"110011101",
  53960=>"111000011",
  53961=>"000011110",
  53962=>"101001100",
  53963=>"011010111",
  53964=>"101111101",
  53965=>"111010100",
  53966=>"010100101",
  53967=>"101001010",
  53968=>"110100010",
  53969=>"101101101",
  53970=>"010000010",
  53971=>"011111111",
  53972=>"100010011",
  53973=>"101110101",
  53974=>"001010000",
  53975=>"111000010",
  53976=>"101110010",
  53977=>"110000111",
  53978=>"010011000",
  53979=>"010010000",
  53980=>"001100111",
  53981=>"100000010",
  53982=>"110001010",
  53983=>"110111110",
  53984=>"111011100",
  53985=>"100110110",
  53986=>"101011111",
  53987=>"111111000",
  53988=>"001101100",
  53989=>"100000001",
  53990=>"100010010",
  53991=>"000111001",
  53992=>"000100100",
  53993=>"011001101",
  53994=>"011011001",
  53995=>"010010010",
  53996=>"001110000",
  53997=>"011110000",
  53998=>"011111110",
  53999=>"011000101",
  54000=>"001001101",
  54001=>"011011000",
  54002=>"100100011",
  54003=>"011010000",
  54004=>"011100101",
  54005=>"110101010",
  54006=>"001111001",
  54007=>"011010111",
  54008=>"010111000",
  54009=>"001000000",
  54010=>"110011111",
  54011=>"010110011",
  54012=>"111010101",
  54013=>"001000000",
  54014=>"000101001",
  54015=>"010100000",
  54016=>"111011111",
  54017=>"000011000",
  54018=>"010011110",
  54019=>"101010110",
  54020=>"010010001",
  54021=>"100110011",
  54022=>"001101101",
  54023=>"011010001",
  54024=>"101100000",
  54025=>"010000110",
  54026=>"111110010",
  54027=>"000011010",
  54028=>"000100100",
  54029=>"010111111",
  54030=>"010000110",
  54031=>"011000100",
  54032=>"111000011",
  54033=>"010000000",
  54034=>"101111111",
  54035=>"111111111",
  54036=>"101000101",
  54037=>"100010001",
  54038=>"101100101",
  54039=>"110100010",
  54040=>"101100001",
  54041=>"011010100",
  54042=>"000010110",
  54043=>"011100100",
  54044=>"110001100",
  54045=>"111010101",
  54046=>"000000110",
  54047=>"011000100",
  54048=>"100000010",
  54049=>"000010110",
  54050=>"110111000",
  54051=>"001001100",
  54052=>"011011011",
  54053=>"001000110",
  54054=>"111011100",
  54055=>"101000101",
  54056=>"111110010",
  54057=>"000111001",
  54058=>"000101001",
  54059=>"000100111",
  54060=>"111100011",
  54061=>"000111001",
  54062=>"100100100",
  54063=>"011100101",
  54064=>"101111011",
  54065=>"110110101",
  54066=>"000110001",
  54067=>"001000110",
  54068=>"011011000",
  54069=>"100111100",
  54070=>"111100000",
  54071=>"111001010",
  54072=>"111011000",
  54073=>"001001011",
  54074=>"001001000",
  54075=>"001001010",
  54076=>"001000011",
  54077=>"100101000",
  54078=>"001000000",
  54079=>"000101010",
  54080=>"110010001",
  54081=>"011000111",
  54082=>"011111100",
  54083=>"011011110",
  54084=>"111100111",
  54085=>"100100010",
  54086=>"011011010",
  54087=>"101001111",
  54088=>"000001110",
  54089=>"111101100",
  54090=>"010010100",
  54091=>"010001001",
  54092=>"010000000",
  54093=>"110011000",
  54094=>"101011001",
  54095=>"010101010",
  54096=>"100111001",
  54097=>"010110110",
  54098=>"001001001",
  54099=>"000011011",
  54100=>"011011000",
  54101=>"110000101",
  54102=>"011010111",
  54103=>"000010011",
  54104=>"110010010",
  54105=>"111010000",
  54106=>"000110001",
  54107=>"101010000",
  54108=>"111001110",
  54109=>"010111111",
  54110=>"001011111",
  54111=>"000011101",
  54112=>"010001011",
  54113=>"110010001",
  54114=>"011011001",
  54115=>"101101010",
  54116=>"011111000",
  54117=>"110010000",
  54118=>"100100111",
  54119=>"001101010",
  54120=>"111001111",
  54121=>"110011111",
  54122=>"001011100",
  54123=>"101001111",
  54124=>"000100000",
  54125=>"111101101",
  54126=>"011010010",
  54127=>"011111010",
  54128=>"000000100",
  54129=>"111001010",
  54130=>"001010011",
  54131=>"001010010",
  54132=>"100000110",
  54133=>"010011100",
  54134=>"101110010",
  54135=>"000101000",
  54136=>"100000101",
  54137=>"000001000",
  54138=>"000100111",
  54139=>"100000000",
  54140=>"001001000",
  54141=>"010001001",
  54142=>"101010001",
  54143=>"110010110",
  54144=>"111011001",
  54145=>"010100110",
  54146=>"100011000",
  54147=>"000001100",
  54148=>"110111100",
  54149=>"111100010",
  54150=>"100110010",
  54151=>"110000010",
  54152=>"011111010",
  54153=>"000000001",
  54154=>"101111111",
  54155=>"101001011",
  54156=>"101001010",
  54157=>"010010010",
  54158=>"100111010",
  54159=>"100100000",
  54160=>"000011100",
  54161=>"110010001",
  54162=>"000011010",
  54163=>"111000010",
  54164=>"011101001",
  54165=>"110010011",
  54166=>"000010111",
  54167=>"110010100",
  54168=>"001100000",
  54169=>"000001110",
  54170=>"101000010",
  54171=>"111001011",
  54172=>"100001010",
  54173=>"000001101",
  54174=>"010100000",
  54175=>"010100111",
  54176=>"001101001",
  54177=>"100100000",
  54178=>"011100111",
  54179=>"100100001",
  54180=>"001011000",
  54181=>"110111100",
  54182=>"001100101",
  54183=>"000111011",
  54184=>"100001011",
  54185=>"011000001",
  54186=>"101100111",
  54187=>"101000100",
  54188=>"000011000",
  54189=>"101001010",
  54190=>"110110000",
  54191=>"010000010",
  54192=>"000110101",
  54193=>"111110111",
  54194=>"011101110",
  54195=>"100100000",
  54196=>"010110010",
  54197=>"100111110",
  54198=>"011011000",
  54199=>"110111011",
  54200=>"010101110",
  54201=>"101101010",
  54202=>"110111001",
  54203=>"110001010",
  54204=>"011100000",
  54205=>"111001100",
  54206=>"101000000",
  54207=>"010001000",
  54208=>"010001010",
  54209=>"011100111",
  54210=>"011101011",
  54211=>"010000111",
  54212=>"100010000",
  54213=>"011101110",
  54214=>"111101001",
  54215=>"000100001",
  54216=>"000110110",
  54217=>"110100000",
  54218=>"101100110",
  54219=>"101110110",
  54220=>"000011100",
  54221=>"110000100",
  54222=>"100010100",
  54223=>"001001011",
  54224=>"001001101",
  54225=>"001100000",
  54226=>"001111011",
  54227=>"010010001",
  54228=>"010100000",
  54229=>"001011000",
  54230=>"100010000",
  54231=>"100000101",
  54232=>"111000100",
  54233=>"001110101",
  54234=>"010101011",
  54235=>"111010011",
  54236=>"001010101",
  54237=>"010001010",
  54238=>"000011010",
  54239=>"000000000",
  54240=>"001101010",
  54241=>"011001100",
  54242=>"000111101",
  54243=>"001101100",
  54244=>"001010000",
  54245=>"000111000",
  54246=>"000011011",
  54247=>"001010101",
  54248=>"100001100",
  54249=>"010111010",
  54250=>"101000111",
  54251=>"100111101",
  54252=>"010110101",
  54253=>"000101010",
  54254=>"001001111",
  54255=>"000011111",
  54256=>"010001111",
  54257=>"111000000",
  54258=>"000001100",
  54259=>"010101101",
  54260=>"000000010",
  54261=>"000100111",
  54262=>"111000010",
  54263=>"011100001",
  54264=>"000011001",
  54265=>"010100010",
  54266=>"100001011",
  54267=>"101011100",
  54268=>"011000011",
  54269=>"100011011",
  54270=>"011001111",
  54271=>"001000111",
  54272=>"000000100",
  54273=>"110010001",
  54274=>"010100001",
  54275=>"110111101",
  54276=>"011110100",
  54277=>"010111100",
  54278=>"000100011",
  54279=>"110011000",
  54280=>"001101100",
  54281=>"100001100",
  54282=>"100101111",
  54283=>"110011100",
  54284=>"100000101",
  54285=>"110111100",
  54286=>"111101111",
  54287=>"000001111",
  54288=>"000010001",
  54289=>"001010110",
  54290=>"100001110",
  54291=>"001001100",
  54292=>"110010010",
  54293=>"011011111",
  54294=>"000110001",
  54295=>"100001010",
  54296=>"100010100",
  54297=>"010010100",
  54298=>"010001111",
  54299=>"001110100",
  54300=>"110100101",
  54301=>"000011000",
  54302=>"010110001",
  54303=>"101001111",
  54304=>"011011101",
  54305=>"101011010",
  54306=>"010011010",
  54307=>"101111000",
  54308=>"011011010",
  54309=>"111101000",
  54310=>"111101101",
  54311=>"001111011",
  54312=>"110010111",
  54313=>"111010010",
  54314=>"000010111",
  54315=>"000000000",
  54316=>"001111111",
  54317=>"111110111",
  54318=>"011001010",
  54319=>"111101101",
  54320=>"110001101",
  54321=>"010110101",
  54322=>"000101000",
  54323=>"101110101",
  54324=>"100000000",
  54325=>"001100111",
  54326=>"101000111",
  54327=>"111001010",
  54328=>"000010001",
  54329=>"011010010",
  54330=>"011001000",
  54331=>"011100010",
  54332=>"001100000",
  54333=>"100101010",
  54334=>"011010100",
  54335=>"000001110",
  54336=>"000101100",
  54337=>"100101000",
  54338=>"001000100",
  54339=>"100111001",
  54340=>"101011110",
  54341=>"010001101",
  54342=>"100000010",
  54343=>"100010000",
  54344=>"110010100",
  54345=>"001001000",
  54346=>"100010101",
  54347=>"010110011",
  54348=>"001010110",
  54349=>"100100100",
  54350=>"101111010",
  54351=>"010111110",
  54352=>"111110000",
  54353=>"101101110",
  54354=>"001000011",
  54355=>"111100101",
  54356=>"101111110",
  54357=>"100100110",
  54358=>"100111000",
  54359=>"000011111",
  54360=>"101111110",
  54361=>"010000101",
  54362=>"000111011",
  54363=>"010101001",
  54364=>"001110110",
  54365=>"100111001",
  54366=>"110011100",
  54367=>"011000011",
  54368=>"010000101",
  54369=>"100001100",
  54370=>"101110111",
  54371=>"111000001",
  54372=>"111100000",
  54373=>"110100000",
  54374=>"110011110",
  54375=>"101000000",
  54376=>"001001011",
  54377=>"000010011",
  54378=>"001000111",
  54379=>"111010100",
  54380=>"011010001",
  54381=>"101010010",
  54382=>"001110010",
  54383=>"011101000",
  54384=>"101001011",
  54385=>"000011001",
  54386=>"100011110",
  54387=>"101110000",
  54388=>"000110101",
  54389=>"110011010",
  54390=>"011011011",
  54391=>"100101001",
  54392=>"101011111",
  54393=>"000010110",
  54394=>"101011100",
  54395=>"110000010",
  54396=>"101100111",
  54397=>"101011100",
  54398=>"000000000",
  54399=>"010000001",
  54400=>"001000001",
  54401=>"000110101",
  54402=>"000011101",
  54403=>"000110111",
  54404=>"100110010",
  54405=>"011101101",
  54406=>"011001111",
  54407=>"011011001",
  54408=>"111111001",
  54409=>"001111011",
  54410=>"011110010",
  54411=>"001010000",
  54412=>"111011100",
  54413=>"100111011",
  54414=>"111000100",
  54415=>"111000000",
  54416=>"101000011",
  54417=>"100010111",
  54418=>"000001011",
  54419=>"010111110",
  54420=>"110100101",
  54421=>"110101110",
  54422=>"011100010",
  54423=>"001100100",
  54424=>"000100001",
  54425=>"110100000",
  54426=>"000000100",
  54427=>"001101001",
  54428=>"100110111",
  54429=>"001001000",
  54430=>"100010001",
  54431=>"111100011",
  54432=>"111111001",
  54433=>"110100011",
  54434=>"110111111",
  54435=>"001010110",
  54436=>"111110101",
  54437=>"000011000",
  54438=>"110100010",
  54439=>"101100011",
  54440=>"001100010",
  54441=>"010000101",
  54442=>"000011011",
  54443=>"011000101",
  54444=>"100100010",
  54445=>"111011011",
  54446=>"100110110",
  54447=>"100101001",
  54448=>"111100100",
  54449=>"100001100",
  54450=>"111110001",
  54451=>"101000001",
  54452=>"111110011",
  54453=>"100111111",
  54454=>"001100111",
  54455=>"001011111",
  54456=>"011101111",
  54457=>"101011011",
  54458=>"100001110",
  54459=>"011000101",
  54460=>"100000001",
  54461=>"111111111",
  54462=>"000111101",
  54463=>"011110100",
  54464=>"001110001",
  54465=>"011000000",
  54466=>"110110111",
  54467=>"100100000",
  54468=>"110110011",
  54469=>"001100100",
  54470=>"000110011",
  54471=>"000000000",
  54472=>"100000011",
  54473=>"010010110",
  54474=>"010001010",
  54475=>"100001011",
  54476=>"011001111",
  54477=>"011111101",
  54478=>"111101100",
  54479=>"111101101",
  54480=>"001100010",
  54481=>"110001010",
  54482=>"100000001",
  54483=>"101111100",
  54484=>"010111010",
  54485=>"000001010",
  54486=>"000111010",
  54487=>"011111111",
  54488=>"111110001",
  54489=>"101111110",
  54490=>"100000011",
  54491=>"100110111",
  54492=>"011010101",
  54493=>"000010101",
  54494=>"111101111",
  54495=>"011011010",
  54496=>"011111001",
  54497=>"111011111",
  54498=>"110100000",
  54499=>"001110101",
  54500=>"101101111",
  54501=>"001001001",
  54502=>"010000010",
  54503=>"101101010",
  54504=>"010011100",
  54505=>"001111011",
  54506=>"110111111",
  54507=>"101101001",
  54508=>"101110111",
  54509=>"001000001",
  54510=>"001001000",
  54511=>"011100001",
  54512=>"010001011",
  54513=>"111111111",
  54514=>"100001000",
  54515=>"010100010",
  54516=>"011001100",
  54517=>"000111110",
  54518=>"000000100",
  54519=>"101000011",
  54520=>"100010011",
  54521=>"100010101",
  54522=>"101001111",
  54523=>"011000111",
  54524=>"110111111",
  54525=>"111100101",
  54526=>"000001000",
  54527=>"011101000",
  54528=>"000111001",
  54529=>"000111100",
  54530=>"100101101",
  54531=>"111110001",
  54532=>"010011011",
  54533=>"000001111",
  54534=>"100001100",
  54535=>"111111111",
  54536=>"000000100",
  54537=>"001010100",
  54538=>"110111100",
  54539=>"100010011",
  54540=>"010001110",
  54541=>"111110110",
  54542=>"011001001",
  54543=>"111000100",
  54544=>"101100010",
  54545=>"101111111",
  54546=>"001011111",
  54547=>"010110011",
  54548=>"010111000",
  54549=>"000111111",
  54550=>"111010010",
  54551=>"000010111",
  54552=>"111001100",
  54553=>"110100000",
  54554=>"111001000",
  54555=>"010010001",
  54556=>"101010001",
  54557=>"010110010",
  54558=>"001010011",
  54559=>"011011110",
  54560=>"000011111",
  54561=>"110010100",
  54562=>"011001011",
  54563=>"000111111",
  54564=>"110100101",
  54565=>"110111001",
  54566=>"100001101",
  54567=>"101100110",
  54568=>"111100111",
  54569=>"001000111",
  54570=>"101010101",
  54571=>"010000010",
  54572=>"000001011",
  54573=>"000000010",
  54574=>"010110000",
  54575=>"100111000",
  54576=>"000011010",
  54577=>"101000000",
  54578=>"110101010",
  54579=>"000111101",
  54580=>"000101110",
  54581=>"001010011",
  54582=>"111101000",
  54583=>"101010111",
  54584=>"000001000",
  54585=>"111011000",
  54586=>"000000000",
  54587=>"001010111",
  54588=>"110000001",
  54589=>"110010001",
  54590=>"101100110",
  54591=>"100000110",
  54592=>"000101101",
  54593=>"001101110",
  54594=>"011000110",
  54595=>"001000100",
  54596=>"101111001",
  54597=>"001000001",
  54598=>"010001000",
  54599=>"111101011",
  54600=>"101110111",
  54601=>"011111001",
  54602=>"011011011",
  54603=>"011110000",
  54604=>"100010101",
  54605=>"010011001",
  54606=>"111110101",
  54607=>"100011111",
  54608=>"011011100",
  54609=>"000101001",
  54610=>"010010111",
  54611=>"101001011",
  54612=>"101010111",
  54613=>"100010001",
  54614=>"001111001",
  54615=>"110101000",
  54616=>"010000101",
  54617=>"011000010",
  54618=>"111110101",
  54619=>"111001010",
  54620=>"011101000",
  54621=>"111111001",
  54622=>"001010011",
  54623=>"111000011",
  54624=>"001001100",
  54625=>"110000100",
  54626=>"101001000",
  54627=>"010111100",
  54628=>"001010110",
  54629=>"010011000",
  54630=>"101111110",
  54631=>"111111101",
  54632=>"101001100",
  54633=>"101100101",
  54634=>"010001001",
  54635=>"010000101",
  54636=>"101100100",
  54637=>"111000100",
  54638=>"110000000",
  54639=>"101010000",
  54640=>"000101001",
  54641=>"110100010",
  54642=>"011111110",
  54643=>"111101010",
  54644=>"111110000",
  54645=>"011011100",
  54646=>"011001101",
  54647=>"101101100",
  54648=>"101000100",
  54649=>"110111000",
  54650=>"010110011",
  54651=>"110011010",
  54652=>"110110111",
  54653=>"111111111",
  54654=>"110011101",
  54655=>"010101111",
  54656=>"111111111",
  54657=>"101001010",
  54658=>"000101001",
  54659=>"011111111",
  54660=>"111100110",
  54661=>"001011111",
  54662=>"011010010",
  54663=>"000101010",
  54664=>"011110011",
  54665=>"110110110",
  54666=>"111010000",
  54667=>"111111111",
  54668=>"010001011",
  54669=>"000111111",
  54670=>"110000001",
  54671=>"110101001",
  54672=>"111101111",
  54673=>"100100001",
  54674=>"110101011",
  54675=>"010111101",
  54676=>"100001111",
  54677=>"000011001",
  54678=>"111000110",
  54679=>"010001101",
  54680=>"011001001",
  54681=>"010001111",
  54682=>"100111011",
  54683=>"010100110",
  54684=>"000001001",
  54685=>"010011011",
  54686=>"101100101",
  54687=>"111101000",
  54688=>"110100010",
  54689=>"000010101",
  54690=>"000011111",
  54691=>"010010100",
  54692=>"010100101",
  54693=>"010000001",
  54694=>"001010110",
  54695=>"010010100",
  54696=>"100110100",
  54697=>"111101110",
  54698=>"001000010",
  54699=>"111010011",
  54700=>"000110001",
  54701=>"001001000",
  54702=>"110011110",
  54703=>"100100000",
  54704=>"011111010",
  54705=>"101111110",
  54706=>"000100100",
  54707=>"001010110",
  54708=>"100000101",
  54709=>"010001000",
  54710=>"011100110",
  54711=>"001000001",
  54712=>"010000101",
  54713=>"111101100",
  54714=>"101000000",
  54715=>"001111001",
  54716=>"100111110",
  54717=>"000100000",
  54718=>"000010100",
  54719=>"010100011",
  54720=>"101101010",
  54721=>"111111011",
  54722=>"001010110",
  54723=>"111111110",
  54724=>"010000101",
  54725=>"101010110",
  54726=>"111011111",
  54727=>"110010010",
  54728=>"010001010",
  54729=>"000101100",
  54730=>"100000101",
  54731=>"101010001",
  54732=>"101010000",
  54733=>"101100010",
  54734=>"111100101",
  54735=>"110110110",
  54736=>"111001001",
  54737=>"000101000",
  54738=>"110010001",
  54739=>"010000011",
  54740=>"011010100",
  54741=>"011010001",
  54742=>"000111101",
  54743=>"000111111",
  54744=>"000111001",
  54745=>"101011000",
  54746=>"011011010",
  54747=>"000010000",
  54748=>"000111110",
  54749=>"101000110",
  54750=>"001011010",
  54751=>"000011111",
  54752=>"101111011",
  54753=>"111001001",
  54754=>"101110010",
  54755=>"101000101",
  54756=>"111010010",
  54757=>"011101000",
  54758=>"100001101",
  54759=>"101111101",
  54760=>"100000001",
  54761=>"110001001",
  54762=>"100100110",
  54763=>"000101011",
  54764=>"010001110",
  54765=>"010011011",
  54766=>"001010111",
  54767=>"010011110",
  54768=>"011011111",
  54769=>"101111011",
  54770=>"000110101",
  54771=>"000001011",
  54772=>"111001011",
  54773=>"011110010",
  54774=>"100011011",
  54775=>"001101010",
  54776=>"111101001",
  54777=>"100110111",
  54778=>"001001011",
  54779=>"001000011",
  54780=>"101000101",
  54781=>"101101110",
  54782=>"010010110",
  54783=>"000111001",
  54784=>"110010011",
  54785=>"110001001",
  54786=>"001101000",
  54787=>"110110101",
  54788=>"100000101",
  54789=>"101011110",
  54790=>"111000110",
  54791=>"110100110",
  54792=>"100011011",
  54793=>"011010110",
  54794=>"110111111",
  54795=>"000001010",
  54796=>"011010000",
  54797=>"100011010",
  54798=>"001100000",
  54799=>"011101011",
  54800=>"101111010",
  54801=>"000000001",
  54802=>"000010001",
  54803=>"111011101",
  54804=>"101011010",
  54805=>"101010111",
  54806=>"010111111",
  54807=>"010010110",
  54808=>"100010100",
  54809=>"000001010",
  54810=>"100001001",
  54811=>"100000000",
  54812=>"101101100",
  54813=>"101001111",
  54814=>"111110010",
  54815=>"100000111",
  54816=>"011010001",
  54817=>"011000011",
  54818=>"001110010",
  54819=>"100010001",
  54820=>"111011111",
  54821=>"001011001",
  54822=>"000010011",
  54823=>"010001000",
  54824=>"100000011",
  54825=>"101011011",
  54826=>"000011000",
  54827=>"000001110",
  54828=>"111010001",
  54829=>"001000100",
  54830=>"110011000",
  54831=>"010000101",
  54832=>"010111110",
  54833=>"000000101",
  54834=>"010110101",
  54835=>"011100000",
  54836=>"100001001",
  54837=>"010001011",
  54838=>"010010111",
  54839=>"110110000",
  54840=>"011000010",
  54841=>"000001000",
  54842=>"111000001",
  54843=>"110001101",
  54844=>"010010101",
  54845=>"110001100",
  54846=>"001001001",
  54847=>"000001001",
  54848=>"011110000",
  54849=>"100000000",
  54850=>"010001000",
  54851=>"010011011",
  54852=>"011110101",
  54853=>"010010100",
  54854=>"000010101",
  54855=>"101010011",
  54856=>"111111111",
  54857=>"011001110",
  54858=>"101101011",
  54859=>"111001000",
  54860=>"000001111",
  54861=>"000100001",
  54862=>"000110111",
  54863=>"111101110",
  54864=>"111010010",
  54865=>"011101111",
  54866=>"110000101",
  54867=>"100011101",
  54868=>"000100001",
  54869=>"011110000",
  54870=>"100111001",
  54871=>"011100011",
  54872=>"111001111",
  54873=>"101101011",
  54874=>"100110000",
  54875=>"110110111",
  54876=>"000001011",
  54877=>"000101100",
  54878=>"010110011",
  54879=>"000110000",
  54880=>"101010000",
  54881=>"000101001",
  54882=>"001110011",
  54883=>"010101000",
  54884=>"000000101",
  54885=>"111010110",
  54886=>"011101000",
  54887=>"110010101",
  54888=>"010001000",
  54889=>"100100000",
  54890=>"101100101",
  54891=>"011010111",
  54892=>"011100011",
  54893=>"011111011",
  54894=>"011011101",
  54895=>"000110111",
  54896=>"010111100",
  54897=>"110011101",
  54898=>"111110101",
  54899=>"100001000",
  54900=>"011110100",
  54901=>"010110111",
  54902=>"111101100",
  54903=>"110101101",
  54904=>"001001000",
  54905=>"111011101",
  54906=>"010000100",
  54907=>"101101000",
  54908=>"111110001",
  54909=>"110001010",
  54910=>"111010100",
  54911=>"111111000",
  54912=>"111000110",
  54913=>"100000101",
  54914=>"101010000",
  54915=>"010000000",
  54916=>"111001111",
  54917=>"101101111",
  54918=>"100100101",
  54919=>"111101001",
  54920=>"110010101",
  54921=>"001100110",
  54922=>"101010000",
  54923=>"101101110",
  54924=>"011010000",
  54925=>"011010100",
  54926=>"010001001",
  54927=>"001111011",
  54928=>"110110101",
  54929=>"000001010",
  54930=>"011011101",
  54931=>"110000110",
  54932=>"111111111",
  54933=>"100100000",
  54934=>"000010100",
  54935=>"000111001",
  54936=>"000110011",
  54937=>"101110001",
  54938=>"010100111",
  54939=>"111100000",
  54940=>"001000011",
  54941=>"011001101",
  54942=>"110000011",
  54943=>"110101111",
  54944=>"001000011",
  54945=>"000101111",
  54946=>"111000110",
  54947=>"100110001",
  54948=>"001111100",
  54949=>"111011011",
  54950=>"111101000",
  54951=>"101000101",
  54952=>"111001110",
  54953=>"110010111",
  54954=>"111001000",
  54955=>"000100100",
  54956=>"000110010",
  54957=>"011100110",
  54958=>"011000110",
  54959=>"111111010",
  54960=>"111110010",
  54961=>"110110110",
  54962=>"100001111",
  54963=>"100111101",
  54964=>"011100001",
  54965=>"110101100",
  54966=>"001110111",
  54967=>"111110110",
  54968=>"100001100",
  54969=>"011001011",
  54970=>"111111001",
  54971=>"010110111",
  54972=>"111001111",
  54973=>"001010001",
  54974=>"000000101",
  54975=>"010110110",
  54976=>"101100011",
  54977=>"010011110",
  54978=>"111010110",
  54979=>"011010000",
  54980=>"101000100",
  54981=>"100111001",
  54982=>"101100111",
  54983=>"110001111",
  54984=>"000001010",
  54985=>"111000111",
  54986=>"000001011",
  54987=>"111101011",
  54988=>"001010100",
  54989=>"010111000",
  54990=>"001000111",
  54991=>"000011111",
  54992=>"111011011",
  54993=>"111100101",
  54994=>"110000100",
  54995=>"001001100",
  54996=>"111011000",
  54997=>"000100111",
  54998=>"000011010",
  54999=>"110001010",
  55000=>"110111001",
  55001=>"101110001",
  55002=>"011111100",
  55003=>"110101001",
  55004=>"111111101",
  55005=>"010001010",
  55006=>"001000011",
  55007=>"010100011",
  55008=>"011101110",
  55009=>"101100110",
  55010=>"111011011",
  55011=>"001001110",
  55012=>"111111001",
  55013=>"010100101",
  55014=>"001001100",
  55015=>"001011010",
  55016=>"010000010",
  55017=>"011011010",
  55018=>"011000010",
  55019=>"110110010",
  55020=>"000000101",
  55021=>"101011111",
  55022=>"010010100",
  55023=>"010110110",
  55024=>"100011010",
  55025=>"000000111",
  55026=>"000011101",
  55027=>"011001111",
  55028=>"010101010",
  55029=>"010111110",
  55030=>"110110100",
  55031=>"111000001",
  55032=>"001001001",
  55033=>"100110011",
  55034=>"000111100",
  55035=>"000010101",
  55036=>"110010000",
  55037=>"010001001",
  55038=>"001101100",
  55039=>"111100111",
  55040=>"011001110",
  55041=>"001011000",
  55042=>"111000110",
  55043=>"001000010",
  55044=>"011010100",
  55045=>"101000010",
  55046=>"011110101",
  55047=>"011010000",
  55048=>"100110000",
  55049=>"000111111",
  55050=>"011001110",
  55051=>"101111010",
  55052=>"010001111",
  55053=>"100010011",
  55054=>"100000001",
  55055=>"101010100",
  55056=>"110000011",
  55057=>"010111100",
  55058=>"000011110",
  55059=>"100010000",
  55060=>"000010111",
  55061=>"110110010",
  55062=>"100111010",
  55063=>"000100101",
  55064=>"011100011",
  55065=>"110010000",
  55066=>"000000111",
  55067=>"110110000",
  55068=>"010010110",
  55069=>"001100010",
  55070=>"100100111",
  55071=>"011101001",
  55072=>"111111011",
  55073=>"010101111",
  55074=>"010011010",
  55075=>"110100000",
  55076=>"111010010",
  55077=>"100010011",
  55078=>"001101110",
  55079=>"110111101",
  55080=>"100001100",
  55081=>"110110000",
  55082=>"111111011",
  55083=>"101010100",
  55084=>"101010000",
  55085=>"000110110",
  55086=>"011111001",
  55087=>"110100010",
  55088=>"001001011",
  55089=>"001110010",
  55090=>"101010101",
  55091=>"100101101",
  55092=>"101110110",
  55093=>"101101010",
  55094=>"100010111",
  55095=>"100000010",
  55096=>"011001000",
  55097=>"110100000",
  55098=>"000011001",
  55099=>"100110111",
  55100=>"111100100",
  55101=>"011101111",
  55102=>"111101000",
  55103=>"110100101",
  55104=>"110000001",
  55105=>"110011110",
  55106=>"010110110",
  55107=>"111100011",
  55108=>"011011001",
  55109=>"110101000",
  55110=>"000101010",
  55111=>"100011111",
  55112=>"101000000",
  55113=>"011001010",
  55114=>"001111110",
  55115=>"011001111",
  55116=>"010111001",
  55117=>"101111101",
  55118=>"110001000",
  55119=>"111000010",
  55120=>"010010010",
  55121=>"011111111",
  55122=>"000110010",
  55123=>"000000000",
  55124=>"000101110",
  55125=>"010000010",
  55126=>"110000110",
  55127=>"000101001",
  55128=>"010000100",
  55129=>"010011011",
  55130=>"111111000",
  55131=>"000000000",
  55132=>"001100101",
  55133=>"001011110",
  55134=>"110100000",
  55135=>"000001101",
  55136=>"001000100",
  55137=>"110100101",
  55138=>"101000111",
  55139=>"011101101",
  55140=>"001010110",
  55141=>"100000001",
  55142=>"011001001",
  55143=>"101010001",
  55144=>"010000111",
  55145=>"000010110",
  55146=>"000001011",
  55147=>"011001100",
  55148=>"000100100",
  55149=>"100011100",
  55150=>"000011010",
  55151=>"100000001",
  55152=>"101011001",
  55153=>"111001101",
  55154=>"010001101",
  55155=>"011100100",
  55156=>"000000100",
  55157=>"111000000",
  55158=>"001000001",
  55159=>"011001001",
  55160=>"001111001",
  55161=>"001110010",
  55162=>"101101101",
  55163=>"100110010",
  55164=>"111100110",
  55165=>"000100110",
  55166=>"100111010",
  55167=>"000101011",
  55168=>"010101100",
  55169=>"111111001",
  55170=>"010101110",
  55171=>"101011001",
  55172=>"010011010",
  55173=>"100101011",
  55174=>"010011100",
  55175=>"001011110",
  55176=>"010010011",
  55177=>"111100011",
  55178=>"111010101",
  55179=>"000100001",
  55180=>"010110101",
  55181=>"001110101",
  55182=>"101000000",
  55183=>"101010111",
  55184=>"010110010",
  55185=>"100100111",
  55186=>"000100111",
  55187=>"111111101",
  55188=>"000011000",
  55189=>"110010001",
  55190=>"111011011",
  55191=>"010100001",
  55192=>"011000111",
  55193=>"010010000",
  55194=>"110010000",
  55195=>"001010010",
  55196=>"001011001",
  55197=>"101010000",
  55198=>"000011110",
  55199=>"000010010",
  55200=>"000100100",
  55201=>"001011101",
  55202=>"010111100",
  55203=>"111110010",
  55204=>"101111010",
  55205=>"101000100",
  55206=>"011111110",
  55207=>"000001000",
  55208=>"001101010",
  55209=>"110000111",
  55210=>"001101001",
  55211=>"111001110",
  55212=>"000110110",
  55213=>"010100100",
  55214=>"011000111",
  55215=>"100011000",
  55216=>"100011111",
  55217=>"110001000",
  55218=>"101001101",
  55219=>"100000000",
  55220=>"001011011",
  55221=>"100111011",
  55222=>"001000000",
  55223=>"111110010",
  55224=>"010000101",
  55225=>"111001000",
  55226=>"110110111",
  55227=>"100010111",
  55228=>"101100010",
  55229=>"110110011",
  55230=>"010110100",
  55231=>"111010101",
  55232=>"001110000",
  55233=>"111011110",
  55234=>"101110000",
  55235=>"011110111",
  55236=>"111111010",
  55237=>"110000111",
  55238=>"001101101",
  55239=>"000011010",
  55240=>"110011011",
  55241=>"001011000",
  55242=>"000110011",
  55243=>"000000001",
  55244=>"011001100",
  55245=>"100111001",
  55246=>"011001100",
  55247=>"000000111",
  55248=>"011001101",
  55249=>"100010000",
  55250=>"111011110",
  55251=>"101000001",
  55252=>"111111000",
  55253=>"101101001",
  55254=>"010010001",
  55255=>"011011011",
  55256=>"011001100",
  55257=>"110000111",
  55258=>"010111111",
  55259=>"110000011",
  55260=>"101011001",
  55261=>"101001100",
  55262=>"001010001",
  55263=>"001001001",
  55264=>"111100011",
  55265=>"011001001",
  55266=>"110101001",
  55267=>"101100110",
  55268=>"101001000",
  55269=>"100100100",
  55270=>"001101111",
  55271=>"101011100",
  55272=>"100101000",
  55273=>"111001101",
  55274=>"010011011",
  55275=>"111010100",
  55276=>"010110111",
  55277=>"001011100",
  55278=>"100101101",
  55279=>"101101000",
  55280=>"001101010",
  55281=>"000001111",
  55282=>"100001101",
  55283=>"111100011",
  55284=>"000111001",
  55285=>"011101000",
  55286=>"101101111",
  55287=>"011110001",
  55288=>"010011110",
  55289=>"011100100",
  55290=>"000001100",
  55291=>"111010010",
  55292=>"101110001",
  55293=>"000010010",
  55294=>"010001110",
  55295=>"000000110",
  55296=>"001110001",
  55297=>"001010010",
  55298=>"110011111",
  55299=>"000011100",
  55300=>"000011100",
  55301=>"100001010",
  55302=>"100100111",
  55303=>"010011010",
  55304=>"010101111",
  55305=>"001101110",
  55306=>"001110000",
  55307=>"111110001",
  55308=>"110100010",
  55309=>"011011010",
  55310=>"011100000",
  55311=>"001101010",
  55312=>"010111100",
  55313=>"001011011",
  55314=>"100000101",
  55315=>"100110010",
  55316=>"100000111",
  55317=>"011011010",
  55318=>"111011111",
  55319=>"000001000",
  55320=>"101111101",
  55321=>"000110000",
  55322=>"000001011",
  55323=>"000001100",
  55324=>"110001101",
  55325=>"001010010",
  55326=>"101100000",
  55327=>"110100010",
  55328=>"001111011",
  55329=>"001111110",
  55330=>"011000101",
  55331=>"100000110",
  55332=>"001011111",
  55333=>"101000111",
  55334=>"001101001",
  55335=>"011101000",
  55336=>"001010010",
  55337=>"110010010",
  55338=>"111100010",
  55339=>"001111111",
  55340=>"010100110",
  55341=>"010001100",
  55342=>"010010101",
  55343=>"011001110",
  55344=>"111011000",
  55345=>"101100110",
  55346=>"001010101",
  55347=>"110010011",
  55348=>"100110001",
  55349=>"100000100",
  55350=>"000110101",
  55351=>"001111111",
  55352=>"001101011",
  55353=>"100110000",
  55354=>"000100100",
  55355=>"100000101",
  55356=>"100101110",
  55357=>"101001000",
  55358=>"010100101",
  55359=>"000001111",
  55360=>"001101001",
  55361=>"010100111",
  55362=>"001110110",
  55363=>"000010111",
  55364=>"000011001",
  55365=>"001111101",
  55366=>"000011111",
  55367=>"000001010",
  55368=>"011001100",
  55369=>"101101111",
  55370=>"100001010",
  55371=>"110000111",
  55372=>"101001111",
  55373=>"111001111",
  55374=>"011011110",
  55375=>"010111011",
  55376=>"011011111",
  55377=>"110011011",
  55378=>"111010110",
  55379=>"000001110",
  55380=>"110111010",
  55381=>"000100000",
  55382=>"001101111",
  55383=>"100100001",
  55384=>"101001111",
  55385=>"100011111",
  55386=>"101001100",
  55387=>"100000001",
  55388=>"100101101",
  55389=>"100111001",
  55390=>"111010110",
  55391=>"111111011",
  55392=>"101101111",
  55393=>"110011010",
  55394=>"100100110",
  55395=>"001010000",
  55396=>"000100111",
  55397=>"101000010",
  55398=>"100110000",
  55399=>"000011100",
  55400=>"000010100",
  55401=>"111000010",
  55402=>"100100011",
  55403=>"111010000",
  55404=>"110011001",
  55405=>"111101100",
  55406=>"011110110",
  55407=>"110010010",
  55408=>"000111010",
  55409=>"001011011",
  55410=>"010100001",
  55411=>"010011111",
  55412=>"000111001",
  55413=>"100001000",
  55414=>"101000110",
  55415=>"001010001",
  55416=>"001011000",
  55417=>"001101010",
  55418=>"100010110",
  55419=>"000010110",
  55420=>"100001101",
  55421=>"110001000",
  55422=>"101100101",
  55423=>"001101000",
  55424=>"011000000",
  55425=>"111000001",
  55426=>"101010101",
  55427=>"010111010",
  55428=>"001000001",
  55429=>"110000101",
  55430=>"000001001",
  55431=>"011111100",
  55432=>"011001011",
  55433=>"100010111",
  55434=>"001010000",
  55435=>"001000001",
  55436=>"100111100",
  55437=>"000101110",
  55438=>"001000100",
  55439=>"111110101",
  55440=>"001000111",
  55441=>"010110111",
  55442=>"100101110",
  55443=>"001001100",
  55444=>"110001100",
  55445=>"110010110",
  55446=>"001010001",
  55447=>"011011011",
  55448=>"110001011",
  55449=>"100100101",
  55450=>"110111001",
  55451=>"100100011",
  55452=>"100111110",
  55453=>"110110110",
  55454=>"100101010",
  55455=>"010010101",
  55456=>"101100111",
  55457=>"111101001",
  55458=>"011001001",
  55459=>"100111011",
  55460=>"101010111",
  55461=>"001000011",
  55462=>"101110111",
  55463=>"000000110",
  55464=>"100010010",
  55465=>"110010000",
  55466=>"101011100",
  55467=>"010010001",
  55468=>"111011010",
  55469=>"101111101",
  55470=>"101000010",
  55471=>"110111010",
  55472=>"110111010",
  55473=>"101001101",
  55474=>"110110001",
  55475=>"001010110",
  55476=>"100000000",
  55477=>"101111011",
  55478=>"001000101",
  55479=>"010010000",
  55480=>"001001011",
  55481=>"010000001",
  55482=>"001011111",
  55483=>"111011101",
  55484=>"000110000",
  55485=>"101010010",
  55486=>"011110010",
  55487=>"100001000",
  55488=>"111111101",
  55489=>"100110010",
  55490=>"110100111",
  55491=>"010000011",
  55492=>"001110011",
  55493=>"000110111",
  55494=>"101101111",
  55495=>"010101111",
  55496=>"101101010",
  55497=>"001000100",
  55498=>"111010111",
  55499=>"001001001",
  55500=>"001010000",
  55501=>"001110011",
  55502=>"100011011",
  55503=>"001100011",
  55504=>"011100011",
  55505=>"100011100",
  55506=>"100101011",
  55507=>"110100110",
  55508=>"100010100",
  55509=>"010001111",
  55510=>"001000100",
  55511=>"000110000",
  55512=>"110111000",
  55513=>"110110010",
  55514=>"110010010",
  55515=>"110101010",
  55516=>"100000010",
  55517=>"100011110",
  55518=>"110111010",
  55519=>"100010110",
  55520=>"100100100",
  55521=>"100110111",
  55522=>"110111110",
  55523=>"100000010",
  55524=>"011101000",
  55525=>"010010111",
  55526=>"000101111",
  55527=>"011011111",
  55528=>"001001010",
  55529=>"101110000",
  55530=>"001011011",
  55531=>"111001000",
  55532=>"111000011",
  55533=>"000100110",
  55534=>"111001111",
  55535=>"001001001",
  55536=>"001110010",
  55537=>"111100111",
  55538=>"010011101",
  55539=>"111110010",
  55540=>"010110111",
  55541=>"010111111",
  55542=>"011100100",
  55543=>"001111011",
  55544=>"100000100",
  55545=>"001111110",
  55546=>"000111110",
  55547=>"100010111",
  55548=>"110111111",
  55549=>"110101010",
  55550=>"110010000",
  55551=>"100111111",
  55552=>"110101000",
  55553=>"111010100",
  55554=>"100100110",
  55555=>"010101000",
  55556=>"001011100",
  55557=>"000001100",
  55558=>"011001101",
  55559=>"100000100",
  55560=>"100111011",
  55561=>"111111000",
  55562=>"010111011",
  55563=>"000101110",
  55564=>"110011000",
  55565=>"001000001",
  55566=>"100110100",
  55567=>"001010110",
  55568=>"011101101",
  55569=>"111110001",
  55570=>"110101010",
  55571=>"101001100",
  55572=>"010110111",
  55573=>"001111001",
  55574=>"110011010",
  55575=>"101001100",
  55576=>"100001000",
  55577=>"001110011",
  55578=>"011011010",
  55579=>"100010101",
  55580=>"110011010",
  55581=>"000000011",
  55582=>"111000001",
  55583=>"110011000",
  55584=>"000000110",
  55585=>"111110011",
  55586=>"000011111",
  55587=>"101101010",
  55588=>"000000011",
  55589=>"101001010",
  55590=>"000100101",
  55591=>"001100110",
  55592=>"110100011",
  55593=>"101010000",
  55594=>"100100100",
  55595=>"010011000",
  55596=>"110000111",
  55597=>"010010101",
  55598=>"101001111",
  55599=>"000011000",
  55600=>"101000100",
  55601=>"000100111",
  55602=>"000001011",
  55603=>"001011110",
  55604=>"001001100",
  55605=>"100101100",
  55606=>"001000110",
  55607=>"110101001",
  55608=>"001101011",
  55609=>"111000001",
  55610=>"001010111",
  55611=>"010001001",
  55612=>"100101100",
  55613=>"101101011",
  55614=>"110110100",
  55615=>"111111101",
  55616=>"110010101",
  55617=>"110001111",
  55618=>"100101010",
  55619=>"110101100",
  55620=>"001110001",
  55621=>"011011001",
  55622=>"000000110",
  55623=>"110010010",
  55624=>"101111000",
  55625=>"010111000",
  55626=>"001101010",
  55627=>"010100101",
  55628=>"000011111",
  55629=>"100111111",
  55630=>"010100101",
  55631=>"010111111",
  55632=>"110100101",
  55633=>"101110010",
  55634=>"100010101",
  55635=>"111100111",
  55636=>"101100011",
  55637=>"001111101",
  55638=>"011101010",
  55639=>"001100110",
  55640=>"000101010",
  55641=>"011111111",
  55642=>"000101101",
  55643=>"111011011",
  55644=>"001010110",
  55645=>"000110100",
  55646=>"000010010",
  55647=>"111110101",
  55648=>"100110101",
  55649=>"000010110",
  55650=>"000010010",
  55651=>"000110111",
  55652=>"010010001",
  55653=>"101101101",
  55654=>"000111111",
  55655=>"000011011",
  55656=>"101111000",
  55657=>"000101010",
  55658=>"110000100",
  55659=>"111011000",
  55660=>"011011100",
  55661=>"111011010",
  55662=>"101101110",
  55663=>"010111100",
  55664=>"000010001",
  55665=>"111010000",
  55666=>"111101001",
  55667=>"111001101",
  55668=>"010111010",
  55669=>"011111011",
  55670=>"110011111",
  55671=>"110111010",
  55672=>"010001010",
  55673=>"111111110",
  55674=>"110010101",
  55675=>"000110001",
  55676=>"010110111",
  55677=>"000110101",
  55678=>"110101100",
  55679=>"101100111",
  55680=>"011110001",
  55681=>"010111100",
  55682=>"010110001",
  55683=>"001100111",
  55684=>"101000110",
  55685=>"110000101",
  55686=>"000110111",
  55687=>"100010000",
  55688=>"111100011",
  55689=>"011010010",
  55690=>"001111000",
  55691=>"111001111",
  55692=>"010011110",
  55693=>"000011010",
  55694=>"101110000",
  55695=>"001001100",
  55696=>"100011000",
  55697=>"000100010",
  55698=>"000100101",
  55699=>"010111110",
  55700=>"010100101",
  55701=>"010000011",
  55702=>"111111100",
  55703=>"000001100",
  55704=>"001110110",
  55705=>"010101100",
  55706=>"111111100",
  55707=>"101011101",
  55708=>"100001001",
  55709=>"000110110",
  55710=>"010101010",
  55711=>"011111111",
  55712=>"111011111",
  55713=>"100010101",
  55714=>"000110001",
  55715=>"011100110",
  55716=>"001000101",
  55717=>"111000101",
  55718=>"110000011",
  55719=>"000001000",
  55720=>"010010011",
  55721=>"110001001",
  55722=>"101100110",
  55723=>"111000101",
  55724=>"001110111",
  55725=>"100001011",
  55726=>"110010110",
  55727=>"001101101",
  55728=>"010100000",
  55729=>"110101001",
  55730=>"010100011",
  55731=>"010110110",
  55732=>"010111011",
  55733=>"110010000",
  55734=>"100001100",
  55735=>"010011111",
  55736=>"011010000",
  55737=>"010001010",
  55738=>"110011001",
  55739=>"001000000",
  55740=>"110111010",
  55741=>"111110000",
  55742=>"001100010",
  55743=>"101110010",
  55744=>"011001001",
  55745=>"111010001",
  55746=>"010100100",
  55747=>"101001010",
  55748=>"100111000",
  55749=>"111011101",
  55750=>"110000011",
  55751=>"110110000",
  55752=>"010101100",
  55753=>"010011010",
  55754=>"011100011",
  55755=>"000101010",
  55756=>"101110111",
  55757=>"110110010",
  55758=>"110110101",
  55759=>"101111010",
  55760=>"001010110",
  55761=>"100110000",
  55762=>"101001100",
  55763=>"111110101",
  55764=>"011101100",
  55765=>"101001100",
  55766=>"101111101",
  55767=>"101100011",
  55768=>"111010101",
  55769=>"101100101",
  55770=>"000010001",
  55771=>"111010010",
  55772=>"010000001",
  55773=>"010100101",
  55774=>"010101111",
  55775=>"110111100",
  55776=>"101100111",
  55777=>"110111111",
  55778=>"110011001",
  55779=>"101011101",
  55780=>"101111100",
  55781=>"100100101",
  55782=>"101001011",
  55783=>"100110110",
  55784=>"001110100",
  55785=>"011101110",
  55786=>"101101111",
  55787=>"000010100",
  55788=>"101011101",
  55789=>"111111101",
  55790=>"101100101",
  55791=>"000001100",
  55792=>"000110011",
  55793=>"001101001",
  55794=>"000001011",
  55795=>"000000001",
  55796=>"010011111",
  55797=>"100110011",
  55798=>"100000101",
  55799=>"111101001",
  55800=>"000110011",
  55801=>"011111001",
  55802=>"010010010",
  55803=>"110010010",
  55804=>"110100111",
  55805=>"010000111",
  55806=>"101101010",
  55807=>"100111001",
  55808=>"001111110",
  55809=>"100111111",
  55810=>"111001001",
  55811=>"000000001",
  55812=>"101000100",
  55813=>"000010101",
  55814=>"010010001",
  55815=>"100000111",
  55816=>"001011110",
  55817=>"000001011",
  55818=>"111100110",
  55819=>"001000000",
  55820=>"100110011",
  55821=>"011100100",
  55822=>"111000111",
  55823=>"010000101",
  55824=>"011010100",
  55825=>"000111011",
  55826=>"110010101",
  55827=>"100101100",
  55828=>"101001110",
  55829=>"000001100",
  55830=>"101100111",
  55831=>"111101110",
  55832=>"100001011",
  55833=>"000100100",
  55834=>"010101100",
  55835=>"101001001",
  55836=>"110001100",
  55837=>"000100001",
  55838=>"100011111",
  55839=>"100010001",
  55840=>"010001000",
  55841=>"100000110",
  55842=>"110010011",
  55843=>"101101100",
  55844=>"000000101",
  55845=>"101001010",
  55846=>"000010000",
  55847=>"110101001",
  55848=>"000010000",
  55849=>"000011010",
  55850=>"111111011",
  55851=>"110100100",
  55852=>"100001110",
  55853=>"001001111",
  55854=>"010011001",
  55855=>"010010111",
  55856=>"011110110",
  55857=>"011101101",
  55858=>"101111100",
  55859=>"101000111",
  55860=>"101101101",
  55861=>"100010010",
  55862=>"000110001",
  55863=>"011011000",
  55864=>"100000110",
  55865=>"001010100",
  55866=>"010101001",
  55867=>"000001111",
  55868=>"001001011",
  55869=>"001000101",
  55870=>"110000001",
  55871=>"000101110",
  55872=>"100011100",
  55873=>"101111101",
  55874=>"010010111",
  55875=>"101011111",
  55876=>"010010000",
  55877=>"110001001",
  55878=>"100101110",
  55879=>"101001010",
  55880=>"110100110",
  55881=>"101111010",
  55882=>"100010100",
  55883=>"110101110",
  55884=>"111011111",
  55885=>"101100001",
  55886=>"110111111",
  55887=>"111101010",
  55888=>"000111010",
  55889=>"101011111",
  55890=>"011110111",
  55891=>"100011110",
  55892=>"110101010",
  55893=>"011010111",
  55894=>"100101001",
  55895=>"000011100",
  55896=>"011111011",
  55897=>"011100000",
  55898=>"001101110",
  55899=>"101000001",
  55900=>"101110100",
  55901=>"100111110",
  55902=>"010101000",
  55903=>"001000001",
  55904=>"111100001",
  55905=>"111010000",
  55906=>"101010101",
  55907=>"101111011",
  55908=>"001000101",
  55909=>"111011100",
  55910=>"010110100",
  55911=>"000110100",
  55912=>"000101001",
  55913=>"001011000",
  55914=>"010001101",
  55915=>"111001001",
  55916=>"010111111",
  55917=>"001101011",
  55918=>"110000110",
  55919=>"100000001",
  55920=>"001001000",
  55921=>"110101011",
  55922=>"011011100",
  55923=>"110101110",
  55924=>"110011010",
  55925=>"110100011",
  55926=>"001001100",
  55927=>"011011000",
  55928=>"010101111",
  55929=>"100001001",
  55930=>"001001100",
  55931=>"011100110",
  55932=>"100100011",
  55933=>"100100101",
  55934=>"000100000",
  55935=>"011101101",
  55936=>"001011010",
  55937=>"100111101",
  55938=>"101001000",
  55939=>"110100000",
  55940=>"011010001",
  55941=>"101011000",
  55942=>"000010101",
  55943=>"111011110",
  55944=>"011110100",
  55945=>"110100000",
  55946=>"001011110",
  55947=>"110111011",
  55948=>"111101001",
  55949=>"100010110",
  55950=>"110000000",
  55951=>"010101101",
  55952=>"101100101",
  55953=>"000110011",
  55954=>"101100000",
  55955=>"110111111",
  55956=>"110000011",
  55957=>"001011110",
  55958=>"111000001",
  55959=>"111111101",
  55960=>"011101101",
  55961=>"100101000",
  55962=>"110100101",
  55963=>"100001011",
  55964=>"110100000",
  55965=>"010001100",
  55966=>"000010010",
  55967=>"110010000",
  55968=>"111100101",
  55969=>"111101011",
  55970=>"110000000",
  55971=>"111001111",
  55972=>"010100101",
  55973=>"110010111",
  55974=>"101010100",
  55975=>"010001110",
  55976=>"010101011",
  55977=>"110011110",
  55978=>"011000111",
  55979=>"100010011",
  55980=>"011110111",
  55981=>"111010100",
  55982=>"011100000",
  55983=>"111111010",
  55984=>"110101100",
  55985=>"111011111",
  55986=>"100010010",
  55987=>"011010000",
  55988=>"010110011",
  55989=>"111101011",
  55990=>"010010101",
  55991=>"011011101",
  55992=>"100100000",
  55993=>"001111110",
  55994=>"111100001",
  55995=>"001110011",
  55996=>"011100111",
  55997=>"010110001",
  55998=>"100000001",
  55999=>"111111011",
  56000=>"000010110",
  56001=>"001011000",
  56002=>"010001110",
  56003=>"000001011",
  56004=>"001000000",
  56005=>"110101011",
  56006=>"111001100",
  56007=>"111110001",
  56008=>"110101100",
  56009=>"001000011",
  56010=>"111001011",
  56011=>"010000011",
  56012=>"101110100",
  56013=>"000101101",
  56014=>"101011111",
  56015=>"110111011",
  56016=>"101001001",
  56017=>"010110110",
  56018=>"001001000",
  56019=>"010101100",
  56020=>"110111111",
  56021=>"001000001",
  56022=>"110001001",
  56023=>"010001010",
  56024=>"111110010",
  56025=>"101111100",
  56026=>"110010111",
  56027=>"001111110",
  56028=>"100100110",
  56029=>"110101010",
  56030=>"101110101",
  56031=>"111100001",
  56032=>"010100001",
  56033=>"111001000",
  56034=>"011000001",
  56035=>"101011110",
  56036=>"011010111",
  56037=>"111001100",
  56038=>"000101111",
  56039=>"100010110",
  56040=>"100110110",
  56041=>"010010110",
  56042=>"111000001",
  56043=>"001111001",
  56044=>"100000110",
  56045=>"100111110",
  56046=>"001011111",
  56047=>"010010110",
  56048=>"100111010",
  56049=>"000011110",
  56050=>"101001110",
  56051=>"101011111",
  56052=>"010001100",
  56053=>"001001000",
  56054=>"100110000",
  56055=>"011101111",
  56056=>"000110001",
  56057=>"000110110",
  56058=>"111101011",
  56059=>"110001111",
  56060=>"001001011",
  56061=>"100100010",
  56062=>"111011101",
  56063=>"010010101",
  56064=>"101110110",
  56065=>"100111101",
  56066=>"011010110",
  56067=>"001001111",
  56068=>"011001001",
  56069=>"001111011",
  56070=>"101011110",
  56071=>"111111001",
  56072=>"110001010",
  56073=>"001100001",
  56074=>"100111111",
  56075=>"001001111",
  56076=>"011001010",
  56077=>"000100110",
  56078=>"111000001",
  56079=>"011110001",
  56080=>"001001101",
  56081=>"001011101",
  56082=>"000101001",
  56083=>"110000101",
  56084=>"100000011",
  56085=>"101010001",
  56086=>"010001011",
  56087=>"100101101",
  56088=>"100101000",
  56089=>"011100001",
  56090=>"000001111",
  56091=>"011101010",
  56092=>"101001001",
  56093=>"111010110",
  56094=>"101110000",
  56095=>"000000111",
  56096=>"110001011",
  56097=>"000100111",
  56098=>"111010001",
  56099=>"101110010",
  56100=>"101010100",
  56101=>"111111111",
  56102=>"001101010",
  56103=>"010111100",
  56104=>"111011100",
  56105=>"010100010",
  56106=>"000110011",
  56107=>"111101100",
  56108=>"101011001",
  56109=>"101001011",
  56110=>"100010110",
  56111=>"100100100",
  56112=>"111101001",
  56113=>"011001101",
  56114=>"100010111",
  56115=>"011011111",
  56116=>"010000100",
  56117=>"101011111",
  56118=>"000100110",
  56119=>"001010111",
  56120=>"011101011",
  56121=>"010010110",
  56122=>"110101011",
  56123=>"110010011",
  56124=>"101110011",
  56125=>"001101011",
  56126=>"001110000",
  56127=>"000100011",
  56128=>"101000000",
  56129=>"101111001",
  56130=>"000110111",
  56131=>"110100111",
  56132=>"111110111",
  56133=>"000001010",
  56134=>"101101100",
  56135=>"111001001",
  56136=>"010100101",
  56137=>"010101000",
  56138=>"100100101",
  56139=>"001000010",
  56140=>"101011011",
  56141=>"101110010",
  56142=>"001110110",
  56143=>"001110010",
  56144=>"111111110",
  56145=>"001110011",
  56146=>"000001010",
  56147=>"000100111",
  56148=>"101011001",
  56149=>"001100111",
  56150=>"010101111",
  56151=>"101101010",
  56152=>"000110111",
  56153=>"100011101",
  56154=>"011011101",
  56155=>"110100110",
  56156=>"001101010",
  56157=>"001110110",
  56158=>"010100110",
  56159=>"011110010",
  56160=>"001100001",
  56161=>"101111001",
  56162=>"101110110",
  56163=>"010010001",
  56164=>"011011110",
  56165=>"111000010",
  56166=>"001110111",
  56167=>"111100011",
  56168=>"000000000",
  56169=>"100011110",
  56170=>"000100011",
  56171=>"100000111",
  56172=>"101110000",
  56173=>"101100100",
  56174=>"000100100",
  56175=>"100011000",
  56176=>"011101111",
  56177=>"110011011",
  56178=>"000000101",
  56179=>"000011010",
  56180=>"100101101",
  56181=>"111111101",
  56182=>"100100000",
  56183=>"000111011",
  56184=>"001100010",
  56185=>"000001010",
  56186=>"100000000",
  56187=>"101000010",
  56188=>"000101000",
  56189=>"110000000",
  56190=>"111101111",
  56191=>"000011011",
  56192=>"001000000",
  56193=>"011110001",
  56194=>"100101110",
  56195=>"011010100",
  56196=>"001110011",
  56197=>"100000101",
  56198=>"111000101",
  56199=>"000100000",
  56200=>"110110111",
  56201=>"010001001",
  56202=>"100111100",
  56203=>"000110100",
  56204=>"010111100",
  56205=>"111100110",
  56206=>"010111111",
  56207=>"110011000",
  56208=>"000011010",
  56209=>"001110000",
  56210=>"001100100",
  56211=>"010011101",
  56212=>"000011000",
  56213=>"111010000",
  56214=>"100100010",
  56215=>"100011101",
  56216=>"001100100",
  56217=>"110001111",
  56218=>"110011000",
  56219=>"010111110",
  56220=>"000001101",
  56221=>"011011110",
  56222=>"000010111",
  56223=>"100111001",
  56224=>"010101001",
  56225=>"011100111",
  56226=>"011000101",
  56227=>"101001100",
  56228=>"101000011",
  56229=>"010011100",
  56230=>"100101000",
  56231=>"010100001",
  56232=>"000000010",
  56233=>"010001100",
  56234=>"011000110",
  56235=>"011101001",
  56236=>"110110001",
  56237=>"111011101",
  56238=>"110101110",
  56239=>"101010110",
  56240=>"011010110",
  56241=>"001110011",
  56242=>"011001101",
  56243=>"001010010",
  56244=>"010000101",
  56245=>"000100011",
  56246=>"011111000",
  56247=>"000011101",
  56248=>"101000100",
  56249=>"101000000",
  56250=>"110011001",
  56251=>"011110101",
  56252=>"111010101",
  56253=>"000000100",
  56254=>"000110001",
  56255=>"100111111",
  56256=>"110100100",
  56257=>"001010001",
  56258=>"110000010",
  56259=>"100101101",
  56260=>"000000011",
  56261=>"010000011",
  56262=>"111010011",
  56263=>"011110001",
  56264=>"001011010",
  56265=>"100100010",
  56266=>"101000001",
  56267=>"001110101",
  56268=>"011110111",
  56269=>"111101101",
  56270=>"100111010",
  56271=>"101010000",
  56272=>"100100001",
  56273=>"011110001",
  56274=>"111100111",
  56275=>"110100011",
  56276=>"101100000",
  56277=>"100111000",
  56278=>"001010011",
  56279=>"101011111",
  56280=>"110100100",
  56281=>"000011001",
  56282=>"010000010",
  56283=>"111100111",
  56284=>"000011101",
  56285=>"110111000",
  56286=>"101010011",
  56287=>"010100000",
  56288=>"100010000",
  56289=>"010010100",
  56290=>"001001001",
  56291=>"010000101",
  56292=>"010000100",
  56293=>"100010011",
  56294=>"111000011",
  56295=>"100000010",
  56296=>"100100100",
  56297=>"001110111",
  56298=>"010001010",
  56299=>"001101111",
  56300=>"010110000",
  56301=>"101111111",
  56302=>"111100010",
  56303=>"011000110",
  56304=>"101101110",
  56305=>"010000101",
  56306=>"111110101",
  56307=>"111111010",
  56308=>"000001000",
  56309=>"101110010",
  56310=>"101001101",
  56311=>"111111111",
  56312=>"100000010",
  56313=>"110110111",
  56314=>"001010110",
  56315=>"011010000",
  56316=>"100010111",
  56317=>"000001111",
  56318=>"000000011",
  56319=>"001100001",
  56320=>"000001000",
  56321=>"010110001",
  56322=>"110001001",
  56323=>"000011110",
  56324=>"101000010",
  56325=>"000011110",
  56326=>"000000011",
  56327=>"001101111",
  56328=>"101011000",
  56329=>"000110101",
  56330=>"110101100",
  56331=>"011111010",
  56332=>"101110110",
  56333=>"101001111",
  56334=>"000000001",
  56335=>"011000010",
  56336=>"111000110",
  56337=>"000100001",
  56338=>"000000010",
  56339=>"000110101",
  56340=>"100011010",
  56341=>"110101100",
  56342=>"000010010",
  56343=>"101000100",
  56344=>"011111000",
  56345=>"000101000",
  56346=>"111000111",
  56347=>"110101111",
  56348=>"101110000",
  56349=>"001101100",
  56350=>"010111001",
  56351=>"001010011",
  56352=>"011000100",
  56353=>"000110111",
  56354=>"111111001",
  56355=>"010001100",
  56356=>"000001011",
  56357=>"111000110",
  56358=>"101111011",
  56359=>"010001011",
  56360=>"011011110",
  56361=>"100101000",
  56362=>"110110010",
  56363=>"001010110",
  56364=>"010001010",
  56365=>"111010001",
  56366=>"000111010",
  56367=>"111000111",
  56368=>"100110101",
  56369=>"110100011",
  56370=>"101000100",
  56371=>"000110110",
  56372=>"000110000",
  56373=>"001001110",
  56374=>"000011000",
  56375=>"101111100",
  56376=>"001111011",
  56377=>"001001011",
  56378=>"001100011",
  56379=>"000011111",
  56380=>"111011100",
  56381=>"111010100",
  56382=>"100000000",
  56383=>"001001110",
  56384=>"111011110",
  56385=>"001001111",
  56386=>"001101011",
  56387=>"101000001",
  56388=>"001101011",
  56389=>"000110101",
  56390=>"111111010",
  56391=>"011101110",
  56392=>"000001101",
  56393=>"010010000",
  56394=>"100100000",
  56395=>"010111110",
  56396=>"111111110",
  56397=>"000110111",
  56398=>"001000111",
  56399=>"011110000",
  56400=>"100110000",
  56401=>"000110110",
  56402=>"110110100",
  56403=>"011101100",
  56404=>"001000010",
  56405=>"100001101",
  56406=>"100111000",
  56407=>"101101101",
  56408=>"010100101",
  56409=>"100010111",
  56410=>"001111111",
  56411=>"010010001",
  56412=>"100110000",
  56413=>"100100001",
  56414=>"000011011",
  56415=>"111100010",
  56416=>"000110001",
  56417=>"111101010",
  56418=>"101100101",
  56419=>"101110011",
  56420=>"101100001",
  56421=>"100101010",
  56422=>"100010110",
  56423=>"001110010",
  56424=>"100011111",
  56425=>"101111111",
  56426=>"110111101",
  56427=>"110000010",
  56428=>"110100000",
  56429=>"111010011",
  56430=>"101000100",
  56431=>"110111010",
  56432=>"000111010",
  56433=>"100001110",
  56434=>"101000000",
  56435=>"000101101",
  56436=>"110001000",
  56437=>"001101100",
  56438=>"110001101",
  56439=>"001101001",
  56440=>"000001111",
  56441=>"110011010",
  56442=>"010100101",
  56443=>"000000000",
  56444=>"001001000",
  56445=>"110110010",
  56446=>"110100001",
  56447=>"000100110",
  56448=>"011010111",
  56449=>"101100010",
  56450=>"001001100",
  56451=>"010111011",
  56452=>"001011101",
  56453=>"001111001",
  56454=>"001001100",
  56455=>"101010111",
  56456=>"011011101",
  56457=>"110010100",
  56458=>"100111100",
  56459=>"111110000",
  56460=>"000001011",
  56461=>"010000100",
  56462=>"111101111",
  56463=>"111000011",
  56464=>"000100010",
  56465=>"111111001",
  56466=>"101101101",
  56467=>"010011111",
  56468=>"000111101",
  56469=>"001001110",
  56470=>"111010110",
  56471=>"010010111",
  56472=>"111010101",
  56473=>"101001111",
  56474=>"111110000",
  56475=>"000101101",
  56476=>"101000111",
  56477=>"100101101",
  56478=>"100000010",
  56479=>"001100111",
  56480=>"110110000",
  56481=>"110000010",
  56482=>"101000110",
  56483=>"010111100",
  56484=>"100011000",
  56485=>"101011101",
  56486=>"101000010",
  56487=>"000100101",
  56488=>"011011011",
  56489=>"110000000",
  56490=>"111110001",
  56491=>"011101000",
  56492=>"010000011",
  56493=>"000001101",
  56494=>"101111110",
  56495=>"001110011",
  56496=>"001011000",
  56497=>"110010000",
  56498=>"101011000",
  56499=>"000000011",
  56500=>"000100010",
  56501=>"011111010",
  56502=>"011000001",
  56503=>"110110100",
  56504=>"000010011",
  56505=>"100100110",
  56506=>"101010100",
  56507=>"101101111",
  56508=>"100111101",
  56509=>"011111000",
  56510=>"111010111",
  56511=>"000100010",
  56512=>"110110001",
  56513=>"011111111",
  56514=>"100011000",
  56515=>"010000100",
  56516=>"111010011",
  56517=>"001111110",
  56518=>"001111111",
  56519=>"100111111",
  56520=>"110110001",
  56521=>"011010000",
  56522=>"000000000",
  56523=>"000101100",
  56524=>"001101110",
  56525=>"110001100",
  56526=>"011011110",
  56527=>"110011111",
  56528=>"000010000",
  56529=>"011010000",
  56530=>"000111111",
  56531=>"110100010",
  56532=>"011000010",
  56533=>"011111101",
  56534=>"110001001",
  56535=>"111010000",
  56536=>"000100000",
  56537=>"000111011",
  56538=>"101101011",
  56539=>"101011010",
  56540=>"011001100",
  56541=>"000110010",
  56542=>"011100001",
  56543=>"011100001",
  56544=>"111001101",
  56545=>"100110011",
  56546=>"110100000",
  56547=>"111010001",
  56548=>"101010111",
  56549=>"110110110",
  56550=>"111001110",
  56551=>"111101010",
  56552=>"100101111",
  56553=>"110111011",
  56554=>"000101010",
  56555=>"001110111",
  56556=>"110011001",
  56557=>"110100001",
  56558=>"111111101",
  56559=>"110000100",
  56560=>"000001000",
  56561=>"100001101",
  56562=>"110111111",
  56563=>"101110011",
  56564=>"001011001",
  56565=>"000010000",
  56566=>"001101101",
  56567=>"000101111",
  56568=>"000010000",
  56569=>"011111011",
  56570=>"111110011",
  56571=>"001111101",
  56572=>"011011110",
  56573=>"010011011",
  56574=>"000001100",
  56575=>"001000111",
  56576=>"001001010",
  56577=>"010101001",
  56578=>"110001001",
  56579=>"000000111",
  56580=>"101101111",
  56581=>"000000010",
  56582=>"111100010",
  56583=>"100010000",
  56584=>"100100111",
  56585=>"001110000",
  56586=>"110000011",
  56587=>"011111000",
  56588=>"100000000",
  56589=>"011000001",
  56590=>"100010001",
  56591=>"000110011",
  56592=>"000001000",
  56593=>"111001011",
  56594=>"111000000",
  56595=>"101110000",
  56596=>"100010100",
  56597=>"001001010",
  56598=>"111110111",
  56599=>"100100100",
  56600=>"110111010",
  56601=>"010001010",
  56602=>"000001000",
  56603=>"010100111",
  56604=>"100010000",
  56605=>"111011110",
  56606=>"100111001",
  56607=>"100101000",
  56608=>"011100001",
  56609=>"011001011",
  56610=>"110110000",
  56611=>"001111001",
  56612=>"011111110",
  56613=>"111011001",
  56614=>"000001100",
  56615=>"100011010",
  56616=>"001010011",
  56617=>"000111010",
  56618=>"100001000",
  56619=>"010010011",
  56620=>"011011001",
  56621=>"110011111",
  56622=>"001101010",
  56623=>"011001000",
  56624=>"101101001",
  56625=>"110001000",
  56626=>"001011011",
  56627=>"110011001",
  56628=>"010001010",
  56629=>"100011011",
  56630=>"101111100",
  56631=>"101011001",
  56632=>"001111111",
  56633=>"111000110",
  56634=>"110111111",
  56635=>"101001000",
  56636=>"000111011",
  56637=>"101101011",
  56638=>"111101100",
  56639=>"111001101",
  56640=>"010101011",
  56641=>"001111100",
  56642=>"000100000",
  56643=>"010110000",
  56644=>"101110001",
  56645=>"001011110",
  56646=>"111100000",
  56647=>"111000011",
  56648=>"101100110",
  56649=>"101000101",
  56650=>"011010000",
  56651=>"011100011",
  56652=>"111110010",
  56653=>"111001011",
  56654=>"011111111",
  56655=>"101010000",
  56656=>"001100110",
  56657=>"010100100",
  56658=>"010010011",
  56659=>"000010011",
  56660=>"101100010",
  56661=>"000001000",
  56662=>"111100100",
  56663=>"001000010",
  56664=>"110100101",
  56665=>"101101111",
  56666=>"011000001",
  56667=>"100100011",
  56668=>"011111101",
  56669=>"010110101",
  56670=>"011000100",
  56671=>"100101000",
  56672=>"111101001",
  56673=>"110001000",
  56674=>"010010010",
  56675=>"001001011",
  56676=>"101111111",
  56677=>"100100101",
  56678=>"100111011",
  56679=>"100100010",
  56680=>"111000100",
  56681=>"100110000",
  56682=>"110011101",
  56683=>"100100100",
  56684=>"100000110",
  56685=>"111000101",
  56686=>"000011110",
  56687=>"110101110",
  56688=>"001001111",
  56689=>"010100000",
  56690=>"100001010",
  56691=>"111011100",
  56692=>"111101100",
  56693=>"001100001",
  56694=>"110100010",
  56695=>"010000110",
  56696=>"010000001",
  56697=>"001001011",
  56698=>"001111101",
  56699=>"001011100",
  56700=>"100111011",
  56701=>"100111110",
  56702=>"111001011",
  56703=>"101100111",
  56704=>"101011111",
  56705=>"010111010",
  56706=>"011110100",
  56707=>"100110010",
  56708=>"101010110",
  56709=>"111011110",
  56710=>"111010011",
  56711=>"111110111",
  56712=>"001000000",
  56713=>"000101111",
  56714=>"111000001",
  56715=>"001000110",
  56716=>"001000010",
  56717=>"000110000",
  56718=>"111101110",
  56719=>"111011001",
  56720=>"011010111",
  56721=>"100001110",
  56722=>"001101011",
  56723=>"001000100",
  56724=>"100110000",
  56725=>"010001011",
  56726=>"100010111",
  56727=>"001000011",
  56728=>"101001100",
  56729=>"101100001",
  56730=>"011110110",
  56731=>"100110100",
  56732=>"111110110",
  56733=>"101001001",
  56734=>"100100101",
  56735=>"010110100",
  56736=>"011100111",
  56737=>"001101001",
  56738=>"000000001",
  56739=>"110011100",
  56740=>"000010101",
  56741=>"101011110",
  56742=>"011000011",
  56743=>"110010111",
  56744=>"001100101",
  56745=>"100100001",
  56746=>"101101100",
  56747=>"010111101",
  56748=>"111110010",
  56749=>"001011111",
  56750=>"000011000",
  56751=>"001101111",
  56752=>"111001101",
  56753=>"001000111",
  56754=>"111111111",
  56755=>"011101111",
  56756=>"000010111",
  56757=>"101000101",
  56758=>"001110011",
  56759=>"001010011",
  56760=>"110001011",
  56761=>"000101111",
  56762=>"110110010",
  56763=>"100011100",
  56764=>"001011000",
  56765=>"111010011",
  56766=>"100011100",
  56767=>"111101100",
  56768=>"001001001",
  56769=>"010100000",
  56770=>"100000110",
  56771=>"010011001",
  56772=>"100001000",
  56773=>"001100100",
  56774=>"110000110",
  56775=>"110100101",
  56776=>"011100001",
  56777=>"101100000",
  56778=>"000010000",
  56779=>"110001011",
  56780=>"010100000",
  56781=>"001100011",
  56782=>"000111100",
  56783=>"101011100",
  56784=>"000011010",
  56785=>"010011010",
  56786=>"010101011",
  56787=>"111111100",
  56788=>"110101011",
  56789=>"001110001",
  56790=>"000111100",
  56791=>"000110010",
  56792=>"000110110",
  56793=>"101000000",
  56794=>"001100100",
  56795=>"100100000",
  56796=>"001011101",
  56797=>"100100001",
  56798=>"011010101",
  56799=>"111110101",
  56800=>"110000011",
  56801=>"011111111",
  56802=>"110001001",
  56803=>"000110100",
  56804=>"001011010",
  56805=>"000001010",
  56806=>"001111101",
  56807=>"101010001",
  56808=>"110011001",
  56809=>"001101001",
  56810=>"000100001",
  56811=>"100101001",
  56812=>"111111100",
  56813=>"000100100",
  56814=>"011010010",
  56815=>"100000101",
  56816=>"101110101",
  56817=>"001101001",
  56818=>"000101011",
  56819=>"110101010",
  56820=>"111000110",
  56821=>"001001111",
  56822=>"001010010",
  56823=>"110000010",
  56824=>"000110100",
  56825=>"000011101",
  56826=>"100011010",
  56827=>"001110111",
  56828=>"010111111",
  56829=>"001001001",
  56830=>"010001110",
  56831=>"000101111",
  56832=>"000011000",
  56833=>"000100010",
  56834=>"111100101",
  56835=>"100101011",
  56836=>"101100011",
  56837=>"001000001",
  56838=>"100111111",
  56839=>"111111111",
  56840=>"100001000",
  56841=>"000001110",
  56842=>"111011100",
  56843=>"011110010",
  56844=>"010100111",
  56845=>"010100010",
  56846=>"110100100",
  56847=>"010110011",
  56848=>"100110010",
  56849=>"101111010",
  56850=>"100110111",
  56851=>"110011101",
  56852=>"000001011",
  56853=>"110011000",
  56854=>"101010101",
  56855=>"110001101",
  56856=>"000100001",
  56857=>"110100110",
  56858=>"000000001",
  56859=>"110001100",
  56860=>"000000011",
  56861=>"010110010",
  56862=>"000110100",
  56863=>"100101001",
  56864=>"011100000",
  56865=>"000100111",
  56866=>"011000100",
  56867=>"001001110",
  56868=>"010101111",
  56869=>"011011010",
  56870=>"111011110",
  56871=>"111111011",
  56872=>"000111000",
  56873=>"010101000",
  56874=>"100010011",
  56875=>"111000011",
  56876=>"000111101",
  56877=>"100000000",
  56878=>"111001001",
  56879=>"011010010",
  56880=>"010001011",
  56881=>"110101110",
  56882=>"011000010",
  56883=>"001100101",
  56884=>"001011111",
  56885=>"100110011",
  56886=>"000010000",
  56887=>"001100110",
  56888=>"001001010",
  56889=>"001100110",
  56890=>"001111011",
  56891=>"100111010",
  56892=>"000110101",
  56893=>"101001110",
  56894=>"101100011",
  56895=>"000000101",
  56896=>"010010111",
  56897=>"111001000",
  56898=>"000011101",
  56899=>"010011011",
  56900=>"110101011",
  56901=>"110100000",
  56902=>"010101101",
  56903=>"111110110",
  56904=>"101011010",
  56905=>"011100010",
  56906=>"111010111",
  56907=>"011011010",
  56908=>"000011000",
  56909=>"100101111",
  56910=>"010001011",
  56911=>"111101100",
  56912=>"110010001",
  56913=>"001101001",
  56914=>"000110110",
  56915=>"011010010",
  56916=>"001101100",
  56917=>"100111000",
  56918=>"000011010",
  56919=>"100000101",
  56920=>"110111001",
  56921=>"100011011",
  56922=>"111011110",
  56923=>"110101101",
  56924=>"001001100",
  56925=>"000100111",
  56926=>"001001101",
  56927=>"110010011",
  56928=>"000011010",
  56929=>"000010101",
  56930=>"010011011",
  56931=>"101011110",
  56932=>"011100001",
  56933=>"101001001",
  56934=>"011101000",
  56935=>"100100110",
  56936=>"100111100",
  56937=>"110011111",
  56938=>"111101101",
  56939=>"000110010",
  56940=>"001110100",
  56941=>"111100000",
  56942=>"100000110",
  56943=>"000100000",
  56944=>"100110001",
  56945=>"011100010",
  56946=>"111001000",
  56947=>"010000100",
  56948=>"111110111",
  56949=>"100001101",
  56950=>"001000111",
  56951=>"001001100",
  56952=>"111100010",
  56953=>"100000001",
  56954=>"110011011",
  56955=>"110000101",
  56956=>"000111100",
  56957=>"110110000",
  56958=>"011110011",
  56959=>"011100100",
  56960=>"010110011",
  56961=>"111111010",
  56962=>"110110000",
  56963=>"001111010",
  56964=>"010000010",
  56965=>"101100010",
  56966=>"001110010",
  56967=>"101000000",
  56968=>"010100000",
  56969=>"111000111",
  56970=>"001011100",
  56971=>"111000111",
  56972=>"100011111",
  56973=>"011111001",
  56974=>"111011100",
  56975=>"011110110",
  56976=>"110011011",
  56977=>"011111100",
  56978=>"001101000",
  56979=>"010001001",
  56980=>"100011000",
  56981=>"001011000",
  56982=>"000100111",
  56983=>"100011001",
  56984=>"000100010",
  56985=>"010001101",
  56986=>"100000110",
  56987=>"110001010",
  56988=>"100101111",
  56989=>"101010100",
  56990=>"000111100",
  56991=>"111100101",
  56992=>"100110100",
  56993=>"111001000",
  56994=>"000001110",
  56995=>"110000011",
  56996=>"000010100",
  56997=>"111101011",
  56998=>"101010101",
  56999=>"101011001",
  57000=>"100001001",
  57001=>"001000000",
  57002=>"110001111",
  57003=>"100001110",
  57004=>"111010010",
  57005=>"011001011",
  57006=>"010000110",
  57007=>"101011101",
  57008=>"011011000",
  57009=>"111110110",
  57010=>"010011010",
  57011=>"111010000",
  57012=>"100101010",
  57013=>"110110101",
  57014=>"100111110",
  57015=>"111110101",
  57016=>"101010010",
  57017=>"010000101",
  57018=>"011001100",
  57019=>"100101001",
  57020=>"001110100",
  57021=>"011100101",
  57022=>"101101101",
  57023=>"111100011",
  57024=>"001000101",
  57025=>"010010000",
  57026=>"100011101",
  57027=>"111111110",
  57028=>"010000000",
  57029=>"010100110",
  57030=>"111111000",
  57031=>"000010110",
  57032=>"011100100",
  57033=>"110101100",
  57034=>"000000100",
  57035=>"001000101",
  57036=>"101011010",
  57037=>"010110100",
  57038=>"000111111",
  57039=>"011111111",
  57040=>"100101101",
  57041=>"101011100",
  57042=>"110010111",
  57043=>"100001101",
  57044=>"100000100",
  57045=>"110010111",
  57046=>"111010101",
  57047=>"000011001",
  57048=>"001011111",
  57049=>"000000011",
  57050=>"001010001",
  57051=>"000000001",
  57052=>"001010101",
  57053=>"100101101",
  57054=>"100110000",
  57055=>"100001000",
  57056=>"001101111",
  57057=>"000000000",
  57058=>"111110100",
  57059=>"101111111",
  57060=>"110111010",
  57061=>"101000100",
  57062=>"100010111",
  57063=>"111011111",
  57064=>"010111010",
  57065=>"010110010",
  57066=>"001001111",
  57067=>"000010001",
  57068=>"001001111",
  57069=>"110101001",
  57070=>"100010011",
  57071=>"000001001",
  57072=>"011110101",
  57073=>"110011110",
  57074=>"100111100",
  57075=>"001000000",
  57076=>"101100100",
  57077=>"011010000",
  57078=>"111000100",
  57079=>"111101111",
  57080=>"000000011",
  57081=>"101101000",
  57082=>"101111011",
  57083=>"001010011",
  57084=>"001011001",
  57085=>"100010010",
  57086=>"111100101",
  57087=>"000111000",
  57088=>"000000001",
  57089=>"001000000",
  57090=>"101000101",
  57091=>"011100000",
  57092=>"000010001",
  57093=>"110000100",
  57094=>"111101111",
  57095=>"100110010",
  57096=>"001010010",
  57097=>"011110001",
  57098=>"000011010",
  57099=>"101111011",
  57100=>"111000011",
  57101=>"010110000",
  57102=>"100100101",
  57103=>"001111001",
  57104=>"111010100",
  57105=>"110000011",
  57106=>"000010000",
  57107=>"111110001",
  57108=>"110011110",
  57109=>"001000011",
  57110=>"100000111",
  57111=>"101000100",
  57112=>"101101100",
  57113=>"100110010",
  57114=>"010101111",
  57115=>"101111101",
  57116=>"001110001",
  57117=>"001110110",
  57118=>"100000010",
  57119=>"111001001",
  57120=>"000011011",
  57121=>"000010010",
  57122=>"111110101",
  57123=>"111010001",
  57124=>"011001001",
  57125=>"001101000",
  57126=>"000100101",
  57127=>"110101000",
  57128=>"111110111",
  57129=>"111010110",
  57130=>"111100100",
  57131=>"101100010",
  57132=>"101110000",
  57133=>"111100101",
  57134=>"101010110",
  57135=>"000000011",
  57136=>"000010011",
  57137=>"001101001",
  57138=>"011111000",
  57139=>"001100011",
  57140=>"011100000",
  57141=>"110010010",
  57142=>"110101110",
  57143=>"100111111",
  57144=>"101010001",
  57145=>"001010111",
  57146=>"011110011",
  57147=>"101001101",
  57148=>"010110000",
  57149=>"110101100",
  57150=>"110001011",
  57151=>"001100100",
  57152=>"010001000",
  57153=>"001001000",
  57154=>"001100001",
  57155=>"111111001",
  57156=>"001100110",
  57157=>"110100001",
  57158=>"011111111",
  57159=>"111000011",
  57160=>"011000111",
  57161=>"111011011",
  57162=>"100000010",
  57163=>"000100010",
  57164=>"011000001",
  57165=>"011110001",
  57166=>"101011011",
  57167=>"001111111",
  57168=>"101100011",
  57169=>"001101100",
  57170=>"101100101",
  57171=>"011110100",
  57172=>"100100101",
  57173=>"001000001",
  57174=>"010000011",
  57175=>"001000010",
  57176=>"111010011",
  57177=>"011001101",
  57178=>"100100111",
  57179=>"000010110",
  57180=>"010000010",
  57181=>"111110101",
  57182=>"001111100",
  57183=>"101001010",
  57184=>"000101010",
  57185=>"000001001",
  57186=>"011010001",
  57187=>"111101111",
  57188=>"110000101",
  57189=>"111110101",
  57190=>"000100010",
  57191=>"111101011",
  57192=>"000010111",
  57193=>"001100011",
  57194=>"001000011",
  57195=>"110001100",
  57196=>"101100101",
  57197=>"001011101",
  57198=>"001110011",
  57199=>"011000001",
  57200=>"001100010",
  57201=>"111011111",
  57202=>"100001000",
  57203=>"111011111",
  57204=>"011101111",
  57205=>"111111111",
  57206=>"100111111",
  57207=>"110010111",
  57208=>"000011110",
  57209=>"010011011",
  57210=>"010101011",
  57211=>"001101001",
  57212=>"101000100",
  57213=>"010100101",
  57214=>"111100010",
  57215=>"000110001",
  57216=>"011100110",
  57217=>"011010001",
  57218=>"111101011",
  57219=>"001111101",
  57220=>"001000010",
  57221=>"101111010",
  57222=>"010100101",
  57223=>"010110100",
  57224=>"001011011",
  57225=>"010010010",
  57226=>"110101011",
  57227=>"111011100",
  57228=>"001101000",
  57229=>"011010000",
  57230=>"110001101",
  57231=>"101000110",
  57232=>"111111001",
  57233=>"011101000",
  57234=>"100110010",
  57235=>"110001001",
  57236=>"000001001",
  57237=>"000000111",
  57238=>"111110101",
  57239=>"101101001",
  57240=>"101101111",
  57241=>"101111111",
  57242=>"111110000",
  57243=>"011110100",
  57244=>"101101111",
  57245=>"001010101",
  57246=>"000010100",
  57247=>"101011110",
  57248=>"100001111",
  57249=>"111011100",
  57250=>"011001111",
  57251=>"001101010",
  57252=>"110111100",
  57253=>"100010001",
  57254=>"111101001",
  57255=>"000101101",
  57256=>"000000001",
  57257=>"101101101",
  57258=>"111101111",
  57259=>"111110110",
  57260=>"110101101",
  57261=>"011011001",
  57262=>"101111010",
  57263=>"100100001",
  57264=>"001110100",
  57265=>"000110110",
  57266=>"111000000",
  57267=>"011010011",
  57268=>"110110000",
  57269=>"011001011",
  57270=>"010001011",
  57271=>"101000101",
  57272=>"000001010",
  57273=>"010001110",
  57274=>"110110010",
  57275=>"000100011",
  57276=>"111001101",
  57277=>"000110000",
  57278=>"111011111",
  57279=>"010010101",
  57280=>"010000100",
  57281=>"111010100",
  57282=>"010111011",
  57283=>"111001000",
  57284=>"110101001",
  57285=>"001101101",
  57286=>"110001100",
  57287=>"110100110",
  57288=>"111101000",
  57289=>"110001001",
  57290=>"001011100",
  57291=>"001101110",
  57292=>"001101100",
  57293=>"100100100",
  57294=>"001100111",
  57295=>"000111101",
  57296=>"111010110",
  57297=>"011101110",
  57298=>"100010000",
  57299=>"100011001",
  57300=>"000000000",
  57301=>"010000110",
  57302=>"000000010",
  57303=>"001110011",
  57304=>"010101010",
  57305=>"111111101",
  57306=>"011011001",
  57307=>"101110110",
  57308=>"010100101",
  57309=>"001100010",
  57310=>"110101001",
  57311=>"011101000",
  57312=>"000010101",
  57313=>"000000101",
  57314=>"111011011",
  57315=>"110100001",
  57316=>"000000111",
  57317=>"011110100",
  57318=>"101011011",
  57319=>"100111000",
  57320=>"100101101",
  57321=>"000000001",
  57322=>"110100100",
  57323=>"100101101",
  57324=>"010110000",
  57325=>"101011100",
  57326=>"000011011",
  57327=>"101101001",
  57328=>"001101001",
  57329=>"100101001",
  57330=>"100100001",
  57331=>"001010111",
  57332=>"101010110",
  57333=>"101010010",
  57334=>"000011011",
  57335=>"111001000",
  57336=>"000010101",
  57337=>"101111000",
  57338=>"101111110",
  57339=>"010011101",
  57340=>"111110011",
  57341=>"111110001",
  57342=>"001011100",
  57343=>"111011000",
  57344=>"000000011",
  57345=>"100111001",
  57346=>"101011010",
  57347=>"101011100",
  57348=>"111100100",
  57349=>"110011010",
  57350=>"111000011",
  57351=>"110011100",
  57352=>"000010101",
  57353=>"100000011",
  57354=>"010010000",
  57355=>"011011101",
  57356=>"011111000",
  57357=>"001110110",
  57358=>"001100000",
  57359=>"111010100",
  57360=>"111011010",
  57361=>"110110110",
  57362=>"011000010",
  57363=>"110000000",
  57364=>"001100110",
  57365=>"001001010",
  57366=>"011110110",
  57367=>"011000010",
  57368=>"010111101",
  57369=>"000101010",
  57370=>"011110101",
  57371=>"000011111",
  57372=>"111101110",
  57373=>"011000100",
  57374=>"010111000",
  57375=>"010111001",
  57376=>"100100111",
  57377=>"001100100",
  57378=>"110111101",
  57379=>"001000111",
  57380=>"101001110",
  57381=>"011000101",
  57382=>"010101110",
  57383=>"111011111",
  57384=>"111001101",
  57385=>"111000111",
  57386=>"010000011",
  57387=>"111100001",
  57388=>"101011101",
  57389=>"011000010",
  57390=>"111000000",
  57391=>"101001011",
  57392=>"111111001",
  57393=>"110101110",
  57394=>"110001101",
  57395=>"111001111",
  57396=>"001000001",
  57397=>"010000111",
  57398=>"111010111",
  57399=>"110101000",
  57400=>"010110000",
  57401=>"100111000",
  57402=>"000010100",
  57403=>"110111111",
  57404=>"100010110",
  57405=>"010111000",
  57406=>"101111001",
  57407=>"000011001",
  57408=>"100001101",
  57409=>"011101100",
  57410=>"111001101",
  57411=>"110010110",
  57412=>"111000011",
  57413=>"010100010",
  57414=>"011000000",
  57415=>"100111011",
  57416=>"101001110",
  57417=>"101010110",
  57418=>"000100101",
  57419=>"011001011",
  57420=>"111110110",
  57421=>"111100110",
  57422=>"100101011",
  57423=>"111111100",
  57424=>"110111100",
  57425=>"111101101",
  57426=>"101000011",
  57427=>"101101000",
  57428=>"111101100",
  57429=>"000010101",
  57430=>"001111111",
  57431=>"110011110",
  57432=>"000111110",
  57433=>"010010100",
  57434=>"010001001",
  57435=>"001011100",
  57436=>"011000101",
  57437=>"010001010",
  57438=>"010111000",
  57439=>"010100111",
  57440=>"100000010",
  57441=>"011001101",
  57442=>"001011001",
  57443=>"100010011",
  57444=>"010110101",
  57445=>"001110011",
  57446=>"100100010",
  57447=>"101111011",
  57448=>"101010000",
  57449=>"011010101",
  57450=>"101011001",
  57451=>"011001011",
  57452=>"111000000",
  57453=>"111011101",
  57454=>"101010111",
  57455=>"110000011",
  57456=>"101001111",
  57457=>"111000110",
  57458=>"111101111",
  57459=>"001110010",
  57460=>"110001001",
  57461=>"100111100",
  57462=>"011100111",
  57463=>"110000010",
  57464=>"111101101",
  57465=>"111111100",
  57466=>"100111101",
  57467=>"101000111",
  57468=>"111100001",
  57469=>"101101010",
  57470=>"000001010",
  57471=>"110001000",
  57472=>"110101011",
  57473=>"000100111",
  57474=>"000000110",
  57475=>"000100011",
  57476=>"110011000",
  57477=>"111110011",
  57478=>"100111010",
  57479=>"011101010",
  57480=>"111111100",
  57481=>"100011000",
  57482=>"010011010",
  57483=>"010001100",
  57484=>"110101000",
  57485=>"010111101",
  57486=>"100100111",
  57487=>"111100001",
  57488=>"101001001",
  57489=>"111100110",
  57490=>"100011010",
  57491=>"010011010",
  57492=>"110010000",
  57493=>"100101011",
  57494=>"111100111",
  57495=>"010001111",
  57496=>"101010010",
  57497=>"011111000",
  57498=>"000000000",
  57499=>"001111110",
  57500=>"100101100",
  57501=>"000001101",
  57502=>"100110001",
  57503=>"111011011",
  57504=>"000011101",
  57505=>"001000011",
  57506=>"110100001",
  57507=>"000011000",
  57508=>"101101111",
  57509=>"010111000",
  57510=>"010010110",
  57511=>"000110111",
  57512=>"010110101",
  57513=>"110111111",
  57514=>"111011111",
  57515=>"000101010",
  57516=>"010000011",
  57517=>"001110000",
  57518=>"111011011",
  57519=>"110000100",
  57520=>"111011000",
  57521=>"000000000",
  57522=>"011111111",
  57523=>"100011100",
  57524=>"000100010",
  57525=>"000001001",
  57526=>"010111101",
  57527=>"110101001",
  57528=>"100011000",
  57529=>"010000010",
  57530=>"010000001",
  57531=>"011100100",
  57532=>"111101101",
  57533=>"111100101",
  57534=>"011101101",
  57535=>"010011000",
  57536=>"100110001",
  57537=>"100100110",
  57538=>"010111101",
  57539=>"100101011",
  57540=>"001000010",
  57541=>"110111011",
  57542=>"000101001",
  57543=>"011000100",
  57544=>"000011111",
  57545=>"110001110",
  57546=>"010000011",
  57547=>"111111000",
  57548=>"000111001",
  57549=>"111001110",
  57550=>"010111010",
  57551=>"101001011",
  57552=>"011011010",
  57553=>"110010011",
  57554=>"100010000",
  57555=>"101111110",
  57556=>"010110111",
  57557=>"011111001",
  57558=>"101100001",
  57559=>"110000111",
  57560=>"001011110",
  57561=>"101000111",
  57562=>"000100000",
  57563=>"101100010",
  57564=>"001110010",
  57565=>"011011110",
  57566=>"100011000",
  57567=>"111110111",
  57568=>"011000110",
  57569=>"001111000",
  57570=>"101001111",
  57571=>"100110001",
  57572=>"100110000",
  57573=>"100001100",
  57574=>"000000010",
  57575=>"101111100",
  57576=>"001101001",
  57577=>"111111100",
  57578=>"011110001",
  57579=>"000100000",
  57580=>"101110110",
  57581=>"111100010",
  57582=>"000000011",
  57583=>"101010001",
  57584=>"101111101",
  57585=>"110100001",
  57586=>"111001011",
  57587=>"000010011",
  57588=>"101110111",
  57589=>"001011100",
  57590=>"011110110",
  57591=>"111001011",
  57592=>"111011011",
  57593=>"111110110",
  57594=>"100111100",
  57595=>"000001001",
  57596=>"101010111",
  57597=>"001001110",
  57598=>"110001001",
  57599=>"110101011",
  57600=>"000011111",
  57601=>"101000100",
  57602=>"001000111",
  57603=>"000010010",
  57604=>"011110011",
  57605=>"110011101",
  57606=>"001100101",
  57607=>"111110011",
  57608=>"101100101",
  57609=>"000010011",
  57610=>"000010000",
  57611=>"110110001",
  57612=>"101110111",
  57613=>"010001000",
  57614=>"111010010",
  57615=>"101010000",
  57616=>"000010010",
  57617=>"101011110",
  57618=>"001111111",
  57619=>"000010011",
  57620=>"001101000",
  57621=>"100010000",
  57622=>"100110111",
  57623=>"011001101",
  57624=>"010111010",
  57625=>"011011100",
  57626=>"100100010",
  57627=>"001010001",
  57628=>"001011010",
  57629=>"101000011",
  57630=>"000101000",
  57631=>"111010000",
  57632=>"100001001",
  57633=>"001011101",
  57634=>"011101011",
  57635=>"001000100",
  57636=>"111000101",
  57637=>"011110111",
  57638=>"110000010",
  57639=>"111000110",
  57640=>"100010010",
  57641=>"101001010",
  57642=>"111011110",
  57643=>"011110000",
  57644=>"111110010",
  57645=>"011000000",
  57646=>"011010011",
  57647=>"010110001",
  57648=>"000010001",
  57649=>"100101110",
  57650=>"111101011",
  57651=>"101000110",
  57652=>"110111001",
  57653=>"101010011",
  57654=>"001111100",
  57655=>"101001001",
  57656=>"101011011",
  57657=>"111010011",
  57658=>"101001100",
  57659=>"100001111",
  57660=>"111000000",
  57661=>"001000000",
  57662=>"000001110",
  57663=>"001101011",
  57664=>"001001000",
  57665=>"010010101",
  57666=>"110111110",
  57667=>"110000000",
  57668=>"010011111",
  57669=>"001101000",
  57670=>"011010001",
  57671=>"100011111",
  57672=>"111011011",
  57673=>"011101000",
  57674=>"011110011",
  57675=>"001010011",
  57676=>"110010101",
  57677=>"100111101",
  57678=>"010111100",
  57679=>"100100011",
  57680=>"110101101",
  57681=>"110010011",
  57682=>"000110001",
  57683=>"101110011",
  57684=>"111101001",
  57685=>"001010011",
  57686=>"010110011",
  57687=>"101010000",
  57688=>"001001110",
  57689=>"011011000",
  57690=>"011011101",
  57691=>"000011010",
  57692=>"010110111",
  57693=>"011100010",
  57694=>"000110011",
  57695=>"001000101",
  57696=>"111110011",
  57697=>"110111010",
  57698=>"010010000",
  57699=>"101000100",
  57700=>"001111111",
  57701=>"010000000",
  57702=>"111001111",
  57703=>"010001010",
  57704=>"011101011",
  57705=>"000010100",
  57706=>"110100010",
  57707=>"100001100",
  57708=>"001001001",
  57709=>"101011011",
  57710=>"010010111",
  57711=>"111100000",
  57712=>"000100000",
  57713=>"011111001",
  57714=>"001010111",
  57715=>"100011101",
  57716=>"110011101",
  57717=>"011000100",
  57718=>"101000101",
  57719=>"010110110",
  57720=>"101100100",
  57721=>"000000000",
  57722=>"011110010",
  57723=>"111100000",
  57724=>"001000010",
  57725=>"011100010",
  57726=>"100110111",
  57727=>"111110000",
  57728=>"100010100",
  57729=>"110111010",
  57730=>"001010111",
  57731=>"000101111",
  57732=>"010110110",
  57733=>"010100000",
  57734=>"000101110",
  57735=>"111000100",
  57736=>"001001100",
  57737=>"011001110",
  57738=>"101011001",
  57739=>"000101110",
  57740=>"110111011",
  57741=>"000011001",
  57742=>"111110011",
  57743=>"101110011",
  57744=>"101100000",
  57745=>"000111111",
  57746=>"000110010",
  57747=>"110000000",
  57748=>"010101011",
  57749=>"110010010",
  57750=>"110001010",
  57751=>"101110110",
  57752=>"100000110",
  57753=>"011001110",
  57754=>"000110011",
  57755=>"110101001",
  57756=>"101110010",
  57757=>"001010000",
  57758=>"010101101",
  57759=>"011000110",
  57760=>"010010001",
  57761=>"010110111",
  57762=>"000010110",
  57763=>"011110111",
  57764=>"000011101",
  57765=>"100100101",
  57766=>"011010000",
  57767=>"000100011",
  57768=>"000001011",
  57769=>"010011111",
  57770=>"010010011",
  57771=>"100101011",
  57772=>"110010101",
  57773=>"111000000",
  57774=>"100110011",
  57775=>"110000010",
  57776=>"010011000",
  57777=>"011001101",
  57778=>"010100011",
  57779=>"001000110",
  57780=>"110111001",
  57781=>"111110011",
  57782=>"000010101",
  57783=>"011001010",
  57784=>"000100110",
  57785=>"011100001",
  57786=>"000110101",
  57787=>"011011110",
  57788=>"001111110",
  57789=>"000111101",
  57790=>"001000010",
  57791=>"011010001",
  57792=>"011010111",
  57793=>"100000001",
  57794=>"101111001",
  57795=>"101000001",
  57796=>"000001100",
  57797=>"110101101",
  57798=>"011100111",
  57799=>"010001111",
  57800=>"101001100",
  57801=>"010011110",
  57802=>"111001100",
  57803=>"011111111",
  57804=>"011101111",
  57805=>"111101110",
  57806=>"011111110",
  57807=>"100011000",
  57808=>"111101001",
  57809=>"011101111",
  57810=>"111010000",
  57811=>"000100010",
  57812=>"000010100",
  57813=>"000111110",
  57814=>"010001010",
  57815=>"101110011",
  57816=>"111100101",
  57817=>"110000101",
  57818=>"010111111",
  57819=>"010001010",
  57820=>"110010100",
  57821=>"101001110",
  57822=>"101011111",
  57823=>"111100110",
  57824=>"111001110",
  57825=>"000100100",
  57826=>"011001000",
  57827=>"010111110",
  57828=>"111000000",
  57829=>"101011000",
  57830=>"100010001",
  57831=>"101110011",
  57832=>"101010000",
  57833=>"100010011",
  57834=>"001010111",
  57835=>"001001111",
  57836=>"011010110",
  57837=>"000100000",
  57838=>"001110011",
  57839=>"010100110",
  57840=>"111111010",
  57841=>"011000010",
  57842=>"010001010",
  57843=>"111110111",
  57844=>"010100000",
  57845=>"001111101",
  57846=>"111101101",
  57847=>"110000100",
  57848=>"010001011",
  57849=>"011000101",
  57850=>"010110000",
  57851=>"001000110",
  57852=>"111000101",
  57853=>"111001100",
  57854=>"000001111",
  57855=>"101000111",
  57856=>"010100001",
  57857=>"000010111",
  57858=>"111101101",
  57859=>"010110011",
  57860=>"100000010",
  57861=>"110101011",
  57862=>"000101011",
  57863=>"010101100",
  57864=>"000001110",
  57865=>"000001000",
  57866=>"111101000",
  57867=>"010100110",
  57868=>"101101111",
  57869=>"011010100",
  57870=>"110101111",
  57871=>"010110111",
  57872=>"010110010",
  57873=>"111011111",
  57874=>"110000111",
  57875=>"000010110",
  57876=>"000000001",
  57877=>"010010001",
  57878=>"101100010",
  57879=>"111110001",
  57880=>"111011101",
  57881=>"011010101",
  57882=>"110011011",
  57883=>"001111101",
  57884=>"111001000",
  57885=>"000101001",
  57886=>"100111011",
  57887=>"001010101",
  57888=>"101100000",
  57889=>"010011000",
  57890=>"001110111",
  57891=>"100000000",
  57892=>"111110111",
  57893=>"000001010",
  57894=>"001000011",
  57895=>"111110010",
  57896=>"101110110",
  57897=>"010001000",
  57898=>"011000100",
  57899=>"001000010",
  57900=>"001001110",
  57901=>"011000001",
  57902=>"101100100",
  57903=>"001000010",
  57904=>"000011100",
  57905=>"000111111",
  57906=>"110101110",
  57907=>"101000011",
  57908=>"110110000",
  57909=>"110111101",
  57910=>"101101100",
  57911=>"111100111",
  57912=>"010000001",
  57913=>"000011101",
  57914=>"001001001",
  57915=>"110000101",
  57916=>"010101100",
  57917=>"010100100",
  57918=>"011001111",
  57919=>"010011101",
  57920=>"000101000",
  57921=>"011100000",
  57922=>"110001000",
  57923=>"001011000",
  57924=>"100100011",
  57925=>"111000011",
  57926=>"100001100",
  57927=>"111011111",
  57928=>"111010111",
  57929=>"001100101",
  57930=>"101001101",
  57931=>"010000110",
  57932=>"011000110",
  57933=>"110001111",
  57934=>"101111010",
  57935=>"111100101",
  57936=>"100100010",
  57937=>"011111110",
  57938=>"110110101",
  57939=>"001110010",
  57940=>"000101001",
  57941=>"000110101",
  57942=>"011110111",
  57943=>"111001010",
  57944=>"000100011",
  57945=>"110001011",
  57946=>"010000110",
  57947=>"111111010",
  57948=>"010000000",
  57949=>"000101001",
  57950=>"000011011",
  57951=>"010101100",
  57952=>"110010011",
  57953=>"011100011",
  57954=>"010110100",
  57955=>"110110011",
  57956=>"000000001",
  57957=>"000111001",
  57958=>"100100011",
  57959=>"011100111",
  57960=>"100010110",
  57961=>"101110111",
  57962=>"100110111",
  57963=>"000101111",
  57964=>"000101111",
  57965=>"100000000",
  57966=>"111011010",
  57967=>"001010110",
  57968=>"001000010",
  57969=>"000110110",
  57970=>"101110010",
  57971=>"001010011",
  57972=>"110101100",
  57973=>"010001101",
  57974=>"001010011",
  57975=>"111000010",
  57976=>"111010011",
  57977=>"011010001",
  57978=>"000011101",
  57979=>"100000001",
  57980=>"111010000",
  57981=>"000001011",
  57982=>"001001111",
  57983=>"110100000",
  57984=>"010011010",
  57985=>"101110101",
  57986=>"010010001",
  57987=>"110101010",
  57988=>"010111111",
  57989=>"001111001",
  57990=>"110001010",
  57991=>"101111010",
  57992=>"101000100",
  57993=>"000101101",
  57994=>"101111111",
  57995=>"011010101",
  57996=>"011000000",
  57997=>"000110110",
  57998=>"001101110",
  57999=>"000110111",
  58000=>"111001011",
  58001=>"100001100",
  58002=>"111110000",
  58003=>"000110010",
  58004=>"000001001",
  58005=>"101111110",
  58006=>"110010010",
  58007=>"101110111",
  58008=>"000011010",
  58009=>"000011001",
  58010=>"010000001",
  58011=>"110110110",
  58012=>"111110110",
  58013=>"100011100",
  58014=>"110010101",
  58015=>"001111010",
  58016=>"000010100",
  58017=>"111100010",
  58018=>"100111010",
  58019=>"101011011",
  58020=>"111111111",
  58021=>"110101110",
  58022=>"000010001",
  58023=>"001111110",
  58024=>"001110010",
  58025=>"000011001",
  58026=>"101101101",
  58027=>"011001101",
  58028=>"101000001",
  58029=>"101100010",
  58030=>"000110101",
  58031=>"110011100",
  58032=>"100100011",
  58033=>"110001100",
  58034=>"010100100",
  58035=>"101110010",
  58036=>"000010010",
  58037=>"001100000",
  58038=>"101111011",
  58039=>"010100111",
  58040=>"010001100",
  58041=>"010001000",
  58042=>"101010111",
  58043=>"010110101",
  58044=>"101100011",
  58045=>"110101111",
  58046=>"101101010",
  58047=>"010100001",
  58048=>"100111000",
  58049=>"111010010",
  58050=>"011010111",
  58051=>"001111000",
  58052=>"101100111",
  58053=>"100111111",
  58054=>"011101100",
  58055=>"001111010",
  58056=>"011110001",
  58057=>"101101001",
  58058=>"111000100",
  58059=>"000101000",
  58060=>"101001010",
  58061=>"000000001",
  58062=>"011100111",
  58063=>"101100110",
  58064=>"000000011",
  58065=>"100010000",
  58066=>"110001001",
  58067=>"110111000",
  58068=>"111000111",
  58069=>"101000011",
  58070=>"001110010",
  58071=>"100001100",
  58072=>"101010001",
  58073=>"100111000",
  58074=>"101100100",
  58075=>"001000111",
  58076=>"010111001",
  58077=>"110111101",
  58078=>"101010010",
  58079=>"001001011",
  58080=>"011010110",
  58081=>"001101101",
  58082=>"100000011",
  58083=>"010100111",
  58084=>"000001101",
  58085=>"100001000",
  58086=>"111011001",
  58087=>"101100111",
  58088=>"000100000",
  58089=>"111111111",
  58090=>"000110101",
  58091=>"110010000",
  58092=>"111011110",
  58093=>"001000001",
  58094=>"110111100",
  58095=>"010101001",
  58096=>"000100101",
  58097=>"100000111",
  58098=>"111110101",
  58099=>"111011011",
  58100=>"100111001",
  58101=>"001010101",
  58102=>"000100101",
  58103=>"110001111",
  58104=>"100110111",
  58105=>"000111011",
  58106=>"100011100",
  58107=>"011010001",
  58108=>"000101001",
  58109=>"101010000",
  58110=>"000110111",
  58111=>"000000000",
  58112=>"100001000",
  58113=>"001000110",
  58114=>"110100100",
  58115=>"011001110",
  58116=>"111001101",
  58117=>"011010100",
  58118=>"101101110",
  58119=>"100110010",
  58120=>"111100110",
  58121=>"001111111",
  58122=>"000011101",
  58123=>"111010011",
  58124=>"000000101",
  58125=>"100011001",
  58126=>"100010011",
  58127=>"000011110",
  58128=>"110101001",
  58129=>"011010010",
  58130=>"000011100",
  58131=>"110111011",
  58132=>"110101100",
  58133=>"110100101",
  58134=>"001000000",
  58135=>"001000001",
  58136=>"010000010",
  58137=>"111100111",
  58138=>"000111010",
  58139=>"100001111",
  58140=>"101101111",
  58141=>"010011000",
  58142=>"101100011",
  58143=>"111110100",
  58144=>"110001111",
  58145=>"010010010",
  58146=>"111011001",
  58147=>"011101100",
  58148=>"111101001",
  58149=>"111101010",
  58150=>"110001010",
  58151=>"111010111",
  58152=>"111000111",
  58153=>"101101101",
  58154=>"110111011",
  58155=>"010100100",
  58156=>"000011100",
  58157=>"000101110",
  58158=>"100010111",
  58159=>"011111100",
  58160=>"010101011",
  58161=>"110011101",
  58162=>"101110010",
  58163=>"010000100",
  58164=>"101101000",
  58165=>"101110000",
  58166=>"000010110",
  58167=>"111101101",
  58168=>"010100000",
  58169=>"101110000",
  58170=>"010101000",
  58171=>"011001010",
  58172=>"000000000",
  58173=>"111111010",
  58174=>"001001001",
  58175=>"010011101",
  58176=>"111010100",
  58177=>"010000010",
  58178=>"011111011",
  58179=>"001110000",
  58180=>"110010011",
  58181=>"111001100",
  58182=>"110011101",
  58183=>"011010111",
  58184=>"011100011",
  58185=>"000111011",
  58186=>"110010101",
  58187=>"010110011",
  58188=>"100001000",
  58189=>"000110101",
  58190=>"101101011",
  58191=>"100010001",
  58192=>"010111101",
  58193=>"111111111",
  58194=>"001101001",
  58195=>"101100111",
  58196=>"011111001",
  58197=>"011101010",
  58198=>"001011010",
  58199=>"001011001",
  58200=>"110111011",
  58201=>"111101001",
  58202=>"010101100",
  58203=>"000100011",
  58204=>"110100101",
  58205=>"110001011",
  58206=>"000001101",
  58207=>"100100000",
  58208=>"011100111",
  58209=>"100101101",
  58210=>"001000001",
  58211=>"101011111",
  58212=>"001101011",
  58213=>"110001001",
  58214=>"010100101",
  58215=>"000101000",
  58216=>"111001101",
  58217=>"011000001",
  58218=>"011011110",
  58219=>"100101011",
  58220=>"100001010",
  58221=>"010101101",
  58222=>"100111010",
  58223=>"111110100",
  58224=>"111101101",
  58225=>"110001101",
  58226=>"001101111",
  58227=>"010100101",
  58228=>"011001010",
  58229=>"001011000",
  58230=>"010111010",
  58231=>"100111110",
  58232=>"100101010",
  58233=>"001011000",
  58234=>"111001001",
  58235=>"010101100",
  58236=>"001100111",
  58237=>"100001100",
  58238=>"100011100",
  58239=>"000101100",
  58240=>"100010010",
  58241=>"010001010",
  58242=>"011001111",
  58243=>"001100000",
  58244=>"011111010",
  58245=>"101001101",
  58246=>"101011111",
  58247=>"110100101",
  58248=>"001101101",
  58249=>"000100100",
  58250=>"010001110",
  58251=>"111101110",
  58252=>"010111011",
  58253=>"101011010",
  58254=>"001100011",
  58255=>"000001100",
  58256=>"010011111",
  58257=>"010001010",
  58258=>"000101001",
  58259=>"010111011",
  58260=>"110000000",
  58261=>"000110110",
  58262=>"001000011",
  58263=>"011100001",
  58264=>"010101011",
  58265=>"111010110",
  58266=>"100101100",
  58267=>"001011011",
  58268=>"011010110",
  58269=>"011111110",
  58270=>"000001000",
  58271=>"011011100",
  58272=>"000000011",
  58273=>"000010001",
  58274=>"000110010",
  58275=>"000100011",
  58276=>"001000111",
  58277=>"011100010",
  58278=>"011001101",
  58279=>"000010011",
  58280=>"000101100",
  58281=>"011011101",
  58282=>"110000110",
  58283=>"110011010",
  58284=>"001000010",
  58285=>"100100111",
  58286=>"010011111",
  58287=>"110000111",
  58288=>"111011001",
  58289=>"111001011",
  58290=>"010110110",
  58291=>"010010110",
  58292=>"000010110",
  58293=>"001010100",
  58294=>"010101101",
  58295=>"000011010",
  58296=>"110001101",
  58297=>"000100110",
  58298=>"110011100",
  58299=>"010001110",
  58300=>"001011001",
  58301=>"010100001",
  58302=>"100001010",
  58303=>"000011100",
  58304=>"000000110",
  58305=>"101111101",
  58306=>"111000110",
  58307=>"010010101",
  58308=>"010010100",
  58309=>"101110001",
  58310=>"010010100",
  58311=>"010001100",
  58312=>"001011111",
  58313=>"010011101",
  58314=>"010101110",
  58315=>"011100100",
  58316=>"111001000",
  58317=>"010000010",
  58318=>"101000101",
  58319=>"111011100",
  58320=>"000010011",
  58321=>"011000010",
  58322=>"010111111",
  58323=>"001110101",
  58324=>"011100010",
  58325=>"001001100",
  58326=>"111000010",
  58327=>"111110000",
  58328=>"100010001",
  58329=>"101101111",
  58330=>"001010001",
  58331=>"000001100",
  58332=>"101110110",
  58333=>"011001111",
  58334=>"101101111",
  58335=>"111100110",
  58336=>"101001011",
  58337=>"011111000",
  58338=>"011100110",
  58339=>"001010011",
  58340=>"111100101",
  58341=>"111111110",
  58342=>"110111101",
  58343=>"100100000",
  58344=>"011100101",
  58345=>"111000100",
  58346=>"010000111",
  58347=>"110000111",
  58348=>"111010010",
  58349=>"010010101",
  58350=>"100100010",
  58351=>"000110101",
  58352=>"000110000",
  58353=>"011111001",
  58354=>"111101011",
  58355=>"000010010",
  58356=>"000100001",
  58357=>"001100111",
  58358=>"001111110",
  58359=>"001011100",
  58360=>"100010010",
  58361=>"100100000",
  58362=>"111000010",
  58363=>"001000110",
  58364=>"001000000",
  58365=>"111111111",
  58366=>"110011101",
  58367=>"001000001",
  58368=>"011100101",
  58369=>"010110011",
  58370=>"110100010",
  58371=>"111000111",
  58372=>"011011010",
  58373=>"110111100",
  58374=>"111011111",
  58375=>"011100101",
  58376=>"010100001",
  58377=>"110100011",
  58378=>"000110010",
  58379=>"101111101",
  58380=>"100000111",
  58381=>"111110001",
  58382=>"110001110",
  58383=>"001000100",
  58384=>"100010010",
  58385=>"000010101",
  58386=>"100111011",
  58387=>"000110110",
  58388=>"011101100",
  58389=>"001101100",
  58390=>"010110110",
  58391=>"011001111",
  58392=>"111010100",
  58393=>"101010010",
  58394=>"001101111",
  58395=>"001100100",
  58396=>"101001101",
  58397=>"111011111",
  58398=>"000001100",
  58399=>"010111011",
  58400=>"100000000",
  58401=>"101110011",
  58402=>"010000011",
  58403=>"010110101",
  58404=>"001101010",
  58405=>"110110010",
  58406=>"001011001",
  58407=>"101010000",
  58408=>"010011101",
  58409=>"101010010",
  58410=>"111000011",
  58411=>"011111100",
  58412=>"101010001",
  58413=>"000101110",
  58414=>"101111110",
  58415=>"000011001",
  58416=>"001101011",
  58417=>"010101011",
  58418=>"110011000",
  58419=>"000100001",
  58420=>"111111000",
  58421=>"010111010",
  58422=>"000100110",
  58423=>"111010111",
  58424=>"101110101",
  58425=>"000010001",
  58426=>"101111010",
  58427=>"000010100",
  58428=>"110000101",
  58429=>"000011110",
  58430=>"011011000",
  58431=>"001010101",
  58432=>"010000001",
  58433=>"110111101",
  58434=>"110010100",
  58435=>"000100110",
  58436=>"101111111",
  58437=>"111000100",
  58438=>"111001010",
  58439=>"001101111",
  58440=>"111010001",
  58441=>"101101101",
  58442=>"101110110",
  58443=>"110101110",
  58444=>"010101101",
  58445=>"100110000",
  58446=>"100111000",
  58447=>"101101010",
  58448=>"100101110",
  58449=>"000000100",
  58450=>"111110100",
  58451=>"000001111",
  58452=>"001001110",
  58453=>"011101100",
  58454=>"110011001",
  58455=>"101100010",
  58456=>"111000100",
  58457=>"010010111",
  58458=>"000010101",
  58459=>"100000100",
  58460=>"100010000",
  58461=>"000000111",
  58462=>"000101110",
  58463=>"010111010",
  58464=>"101011000",
  58465=>"001000101",
  58466=>"001010000",
  58467=>"001100011",
  58468=>"010000001",
  58469=>"100111111",
  58470=>"011000001",
  58471=>"000111111",
  58472=>"000010100",
  58473=>"111001001",
  58474=>"101000101",
  58475=>"001001110",
  58476=>"111101111",
  58477=>"000010101",
  58478=>"010100001",
  58479=>"001100110",
  58480=>"111000001",
  58481=>"000100001",
  58482=>"110000010",
  58483=>"110011100",
  58484=>"110110011",
  58485=>"011100110",
  58486=>"110011000",
  58487=>"011011010",
  58488=>"111011101",
  58489=>"000010100",
  58490=>"000100110",
  58491=>"011000000",
  58492=>"001101101",
  58493=>"011000100",
  58494=>"010001010",
  58495=>"100100101",
  58496=>"011010101",
  58497=>"010100110",
  58498=>"111100100",
  58499=>"010001100",
  58500=>"001000011",
  58501=>"000111110",
  58502=>"010110101",
  58503=>"010000101",
  58504=>"010100000",
  58505=>"110001101",
  58506=>"011001011",
  58507=>"111010111",
  58508=>"011011001",
  58509=>"101001110",
  58510=>"110011100",
  58511=>"000110110",
  58512=>"000110111",
  58513=>"011101111",
  58514=>"000110011",
  58515=>"101101011",
  58516=>"100011001",
  58517=>"000011000",
  58518=>"000011011",
  58519=>"011100101",
  58520=>"000101101",
  58521=>"001000110",
  58522=>"111011010",
  58523=>"000000000",
  58524=>"000001001",
  58525=>"000010000",
  58526=>"001001000",
  58527=>"011101111",
  58528=>"111010101",
  58529=>"111110001",
  58530=>"101000101",
  58531=>"110000110",
  58532=>"101111000",
  58533=>"110010010",
  58534=>"010011100",
  58535=>"111000011",
  58536=>"000111110",
  58537=>"011001010",
  58538=>"011011010",
  58539=>"101001110",
  58540=>"000010010",
  58541=>"100000011",
  58542=>"101110111",
  58543=>"100011110",
  58544=>"000110000",
  58545=>"000010011",
  58546=>"001111000",
  58547=>"010100100",
  58548=>"001111111",
  58549=>"000001101",
  58550=>"001100000",
  58551=>"000101110",
  58552=>"111000111",
  58553=>"101010010",
  58554=>"111001100",
  58555=>"000111010",
  58556=>"111001010",
  58557=>"010001100",
  58558=>"101101000",
  58559=>"111101010",
  58560=>"001101110",
  58561=>"001100101",
  58562=>"001000000",
  58563=>"111111110",
  58564=>"110101110",
  58565=>"100011011",
  58566=>"111010110",
  58567=>"101010110",
  58568=>"010011100",
  58569=>"111001101",
  58570=>"000000010",
  58571=>"100110101",
  58572=>"110001001",
  58573=>"100111101",
  58574=>"100011111",
  58575=>"000010001",
  58576=>"010010100",
  58577=>"010001111",
  58578=>"001000100",
  58579=>"111000110",
  58580=>"111000001",
  58581=>"010000100",
  58582=>"100100011",
  58583=>"101001101",
  58584=>"101011010",
  58585=>"101101011",
  58586=>"000000000",
  58587=>"000001001",
  58588=>"100111010",
  58589=>"011010000",
  58590=>"110011010",
  58591=>"011111011",
  58592=>"000011011",
  58593=>"011000100",
  58594=>"110101100",
  58595=>"010110001",
  58596=>"010111100",
  58597=>"001000001",
  58598=>"011000000",
  58599=>"000000011",
  58600=>"000101011",
  58601=>"101010100",
  58602=>"011001010",
  58603=>"001100001",
  58604=>"100111000",
  58605=>"111101000",
  58606=>"011011010",
  58607=>"110011101",
  58608=>"111111111",
  58609=>"000001010",
  58610=>"101100010",
  58611=>"010101010",
  58612=>"010110111",
  58613=>"001111111",
  58614=>"001100100",
  58615=>"010111001",
  58616=>"000011001",
  58617=>"100101111",
  58618=>"011001100",
  58619=>"000010111",
  58620=>"111011111",
  58621=>"010100110",
  58622=>"001111011",
  58623=>"010100100",
  58624=>"010110110",
  58625=>"111000111",
  58626=>"111011101",
  58627=>"001001000",
  58628=>"110111111",
  58629=>"010000111",
  58630=>"001000011",
  58631=>"111000001",
  58632=>"100111010",
  58633=>"001000001",
  58634=>"001111000",
  58635=>"101000011",
  58636=>"010001011",
  58637=>"111010000",
  58638=>"100010110",
  58639=>"100010101",
  58640=>"011100100",
  58641=>"100001101",
  58642=>"010110101",
  58643=>"010110101",
  58644=>"001110100",
  58645=>"110110010",
  58646=>"000010001",
  58647=>"101111110",
  58648=>"111110000",
  58649=>"001011110",
  58650=>"001010110",
  58651=>"000011100",
  58652=>"011111111",
  58653=>"010000000",
  58654=>"101101110",
  58655=>"100101011",
  58656=>"000110100",
  58657=>"011000000",
  58658=>"000111111",
  58659=>"101000010",
  58660=>"111000111",
  58661=>"101000101",
  58662=>"000011110",
  58663=>"000001101",
  58664=>"001101110",
  58665=>"101111001",
  58666=>"000001010",
  58667=>"000001100",
  58668=>"001110011",
  58669=>"111001100",
  58670=>"101101010",
  58671=>"111101110",
  58672=>"001001010",
  58673=>"000101001",
  58674=>"000001101",
  58675=>"000111101",
  58676=>"110011100",
  58677=>"000011110",
  58678=>"011010100",
  58679=>"111010101",
  58680=>"000100000",
  58681=>"101000010",
  58682=>"110001101",
  58683=>"101011111",
  58684=>"001001000",
  58685=>"110011011",
  58686=>"001001111",
  58687=>"111001111",
  58688=>"011001000",
  58689=>"011101111",
  58690=>"000110011",
  58691=>"000101010",
  58692=>"000000000",
  58693=>"101110111",
  58694=>"100000110",
  58695=>"100110101",
  58696=>"101000111",
  58697=>"010101011",
  58698=>"111100101",
  58699=>"011100000",
  58700=>"011001111",
  58701=>"111000111",
  58702=>"101100010",
  58703=>"000110100",
  58704=>"000011111",
  58705=>"011111000",
  58706=>"001010101",
  58707=>"111101000",
  58708=>"000000100",
  58709=>"100111101",
  58710=>"111000001",
  58711=>"001001100",
  58712=>"110111010",
  58713=>"100000011",
  58714=>"100011001",
  58715=>"011011111",
  58716=>"110110001",
  58717=>"010001011",
  58718=>"001101100",
  58719=>"100001001",
  58720=>"110001110",
  58721=>"100100100",
  58722=>"000010101",
  58723=>"000000111",
  58724=>"010110111",
  58725=>"101001111",
  58726=>"101110111",
  58727=>"010100111",
  58728=>"010100001",
  58729=>"001011011",
  58730=>"101001101",
  58731=>"001001101",
  58732=>"010101010",
  58733=>"001110101",
  58734=>"011001001",
  58735=>"111111010",
  58736=>"001001010",
  58737=>"011101010",
  58738=>"000010110",
  58739=>"110100010",
  58740=>"000111110",
  58741=>"000100100",
  58742=>"001010111",
  58743=>"010101110",
  58744=>"101011000",
  58745=>"000101010",
  58746=>"100111000",
  58747=>"100000001",
  58748=>"011101110",
  58749=>"001101010",
  58750=>"111011010",
  58751=>"000000010",
  58752=>"000001001",
  58753=>"000000000",
  58754=>"000010101",
  58755=>"100000110",
  58756=>"000000110",
  58757=>"010001001",
  58758=>"111010101",
  58759=>"100100111",
  58760=>"000000100",
  58761=>"111011010",
  58762=>"011111101",
  58763=>"000110111",
  58764=>"101011000",
  58765=>"000011100",
  58766=>"110011010",
  58767=>"000100100",
  58768=>"111101100",
  58769=>"001000010",
  58770=>"001001110",
  58771=>"001111011",
  58772=>"001111011",
  58773=>"011111101",
  58774=>"010110000",
  58775=>"101000000",
  58776=>"001110110",
  58777=>"101001001",
  58778=>"111100111",
  58779=>"001000101",
  58780=>"010000001",
  58781=>"010101100",
  58782=>"100100011",
  58783=>"100100001",
  58784=>"110111110",
  58785=>"000000111",
  58786=>"001100110",
  58787=>"101111101",
  58788=>"100101000",
  58789=>"011110100",
  58790=>"100001111",
  58791=>"111111000",
  58792=>"111110110",
  58793=>"011101010",
  58794=>"001100011",
  58795=>"000101001",
  58796=>"010001000",
  58797=>"101010101",
  58798=>"110101101",
  58799=>"101011000",
  58800=>"010110010",
  58801=>"000000011",
  58802=>"111000010",
  58803=>"001000001",
  58804=>"110011111",
  58805=>"001100111",
  58806=>"010001000",
  58807=>"100100110",
  58808=>"101100000",
  58809=>"100101110",
  58810=>"010000111",
  58811=>"010111000",
  58812=>"101001011",
  58813=>"010010001",
  58814=>"011110000",
  58815=>"101011101",
  58816=>"001101111",
  58817=>"100001010",
  58818=>"001101001",
  58819=>"011110010",
  58820=>"000000010",
  58821=>"110001011",
  58822=>"011011110",
  58823=>"110001001",
  58824=>"110100010",
  58825=>"001001001",
  58826=>"001100011",
  58827=>"101110111",
  58828=>"100011101",
  58829=>"100100001",
  58830=>"000010001",
  58831=>"100000100",
  58832=>"100111110",
  58833=>"010010100",
  58834=>"011101010",
  58835=>"100010000",
  58836=>"101011010",
  58837=>"101001100",
  58838=>"101101001",
  58839=>"000100001",
  58840=>"010010110",
  58841=>"111101101",
  58842=>"101010001",
  58843=>"001111100",
  58844=>"001110011",
  58845=>"101111110",
  58846=>"100000000",
  58847=>"000100110",
  58848=>"101110011",
  58849=>"011110110",
  58850=>"001011000",
  58851=>"110110100",
  58852=>"111110101",
  58853=>"001000110",
  58854=>"100111000",
  58855=>"011010001",
  58856=>"110110111",
  58857=>"100000001",
  58858=>"000110011",
  58859=>"010000001",
  58860=>"010011010",
  58861=>"010010101",
  58862=>"100110001",
  58863=>"101010100",
  58864=>"111111001",
  58865=>"111110010",
  58866=>"010011111",
  58867=>"010011011",
  58868=>"110010111",
  58869=>"000010000",
  58870=>"111101011",
  58871=>"010111011",
  58872=>"010111001",
  58873=>"011011101",
  58874=>"101000001",
  58875=>"000101001",
  58876=>"111011100",
  58877=>"000010110",
  58878=>"000111001",
  58879=>"000100100",
  58880=>"100110011",
  58881=>"011000011",
  58882=>"100101101",
  58883=>"000010001",
  58884=>"111110111",
  58885=>"100011110",
  58886=>"010111100",
  58887=>"010100010",
  58888=>"000100010",
  58889=>"001000100",
  58890=>"000011100",
  58891=>"011110111",
  58892=>"110111111",
  58893=>"000010111",
  58894=>"011001011",
  58895=>"100101101",
  58896=>"011110001",
  58897=>"011001010",
  58898=>"111100110",
  58899=>"110010010",
  58900=>"010000001",
  58901=>"001000011",
  58902=>"011100110",
  58903=>"010101110",
  58904=>"000000111",
  58905=>"010100111",
  58906=>"000001111",
  58907=>"110101101",
  58908=>"101100000",
  58909=>"001101001",
  58910=>"001001001",
  58911=>"010010101",
  58912=>"100010010",
  58913=>"111111010",
  58914=>"001101110",
  58915=>"000101010",
  58916=>"000111001",
  58917=>"011101110",
  58918=>"010000101",
  58919=>"000000010",
  58920=>"010100000",
  58921=>"011111101",
  58922=>"101001111",
  58923=>"100100001",
  58924=>"110010100",
  58925=>"010111000",
  58926=>"100100001",
  58927=>"111010011",
  58928=>"000000001",
  58929=>"011001010",
  58930=>"001110001",
  58931=>"000001000",
  58932=>"110011000",
  58933=>"110110011",
  58934=>"110100001",
  58935=>"011111011",
  58936=>"001010010",
  58937=>"001001000",
  58938=>"100010001",
  58939=>"000100010",
  58940=>"110101100",
  58941=>"010011110",
  58942=>"001110001",
  58943=>"100001111",
  58944=>"000000111",
  58945=>"001010101",
  58946=>"010110100",
  58947=>"110100011",
  58948=>"000000101",
  58949=>"000101111",
  58950=>"001100001",
  58951=>"000011111",
  58952=>"110110010",
  58953=>"100010011",
  58954=>"100110100",
  58955=>"110111101",
  58956=>"010111110",
  58957=>"101110110",
  58958=>"111100100",
  58959=>"110011100",
  58960=>"101001111",
  58961=>"010101000",
  58962=>"110110001",
  58963=>"110000110",
  58964=>"110110010",
  58965=>"000000000",
  58966=>"000001110",
  58967=>"000011111",
  58968=>"111010101",
  58969=>"111100011",
  58970=>"101000111",
  58971=>"110000101",
  58972=>"101000011",
  58973=>"000000001",
  58974=>"001111100",
  58975=>"010110100",
  58976=>"110000011",
  58977=>"011000001",
  58978=>"101111011",
  58979=>"001110101",
  58980=>"000011000",
  58981=>"111000001",
  58982=>"110011001",
  58983=>"101010101",
  58984=>"100110101",
  58985=>"100111001",
  58986=>"010101110",
  58987=>"100011001",
  58988=>"101110110",
  58989=>"110111110",
  58990=>"100111010",
  58991=>"011101111",
  58992=>"010111101",
  58993=>"100011011",
  58994=>"100101110",
  58995=>"010101111",
  58996=>"111110010",
  58997=>"101011100",
  58998=>"011010110",
  58999=>"110001010",
  59000=>"010010000",
  59001=>"001011001",
  59002=>"110000011",
  59003=>"011101010",
  59004=>"101101110",
  59005=>"011100101",
  59006=>"000000100",
  59007=>"011101111",
  59008=>"101100011",
  59009=>"111110010",
  59010=>"010011100",
  59011=>"000101101",
  59012=>"001010111",
  59013=>"011110110",
  59014=>"110100101",
  59015=>"000101101",
  59016=>"101111110",
  59017=>"110100000",
  59018=>"001001110",
  59019=>"101111110",
  59020=>"000101101",
  59021=>"001011010",
  59022=>"111001011",
  59023=>"010001111",
  59024=>"111011110",
  59025=>"110011011",
  59026=>"101101011",
  59027=>"111111010",
  59028=>"001101100",
  59029=>"100000011",
  59030=>"101010011",
  59031=>"110001010",
  59032=>"110001010",
  59033=>"110110110",
  59034=>"011011010",
  59035=>"010111110",
  59036=>"011010010",
  59037=>"111110110",
  59038=>"101111110",
  59039=>"011100010",
  59040=>"100011110",
  59041=>"000010001",
  59042=>"111110100",
  59043=>"111001011",
  59044=>"010011100",
  59045=>"111010111",
  59046=>"001000001",
  59047=>"010011001",
  59048=>"110010011",
  59049=>"110100111",
  59050=>"010101001",
  59051=>"010001000",
  59052=>"110010001",
  59053=>"100000011",
  59054=>"001100101",
  59055=>"110000000",
  59056=>"010011111",
  59057=>"101001100",
  59058=>"000000101",
  59059=>"110101000",
  59060=>"111111010",
  59061=>"010010101",
  59062=>"110000000",
  59063=>"001101000",
  59064=>"101100000",
  59065=>"000011010",
  59066=>"101001010",
  59067=>"100111111",
  59068=>"010010110",
  59069=>"001001100",
  59070=>"000000100",
  59071=>"000100010",
  59072=>"100101110",
  59073=>"111100011",
  59074=>"000100100",
  59075=>"111111100",
  59076=>"100111010",
  59077=>"011000011",
  59078=>"110000111",
  59079=>"100110000",
  59080=>"000001001",
  59081=>"111110111",
  59082=>"001000000",
  59083=>"001000101",
  59084=>"001011100",
  59085=>"100101011",
  59086=>"111100000",
  59087=>"110011011",
  59088=>"110110001",
  59089=>"000000010",
  59090=>"001000100",
  59091=>"000001110",
  59092=>"001100000",
  59093=>"000110010",
  59094=>"011110001",
  59095=>"010100111",
  59096=>"110000111",
  59097=>"111001100",
  59098=>"011010110",
  59099=>"100100100",
  59100=>"001101110",
  59101=>"010100010",
  59102=>"001101010",
  59103=>"000100100",
  59104=>"000111000",
  59105=>"000010011",
  59106=>"000111100",
  59107=>"010001010",
  59108=>"011000101",
  59109=>"111011100",
  59110=>"000101011",
  59111=>"101001111",
  59112=>"110101110",
  59113=>"101111000",
  59114=>"101110001",
  59115=>"111110101",
  59116=>"111101000",
  59117=>"101101111",
  59118=>"111101100",
  59119=>"010000011",
  59120=>"001100100",
  59121=>"110011100",
  59122=>"000010111",
  59123=>"001101111",
  59124=>"011101111",
  59125=>"101110101",
  59126=>"000101001",
  59127=>"100001011",
  59128=>"110011011",
  59129=>"101010100",
  59130=>"000101110",
  59131=>"010010001",
  59132=>"110110001",
  59133=>"010100011",
  59134=>"110010010",
  59135=>"000111001",
  59136=>"010011110",
  59137=>"001110110",
  59138=>"010000100",
  59139=>"000010111",
  59140=>"110110001",
  59141=>"100101100",
  59142=>"100010001",
  59143=>"111100111",
  59144=>"110000100",
  59145=>"101100101",
  59146=>"011101011",
  59147=>"010010100",
  59148=>"110000000",
  59149=>"011101111",
  59150=>"100110111",
  59151=>"101111111",
  59152=>"000100000",
  59153=>"101010100",
  59154=>"101111001",
  59155=>"111101011",
  59156=>"000000010",
  59157=>"010011100",
  59158=>"111011101",
  59159=>"101111110",
  59160=>"000100011",
  59161=>"111000110",
  59162=>"111000111",
  59163=>"101101100",
  59164=>"101101111",
  59165=>"001010110",
  59166=>"100000001",
  59167=>"111011100",
  59168=>"000001110",
  59169=>"110011100",
  59170=>"010111010",
  59171=>"011010101",
  59172=>"111011110",
  59173=>"011010000",
  59174=>"011010100",
  59175=>"010011111",
  59176=>"000100011",
  59177=>"010001000",
  59178=>"100000011",
  59179=>"011100010",
  59180=>"101011001",
  59181=>"111010111",
  59182=>"100101101",
  59183=>"110001000",
  59184=>"001001010",
  59185=>"100110111",
  59186=>"101111001",
  59187=>"000101100",
  59188=>"011000000",
  59189=>"111011101",
  59190=>"001100101",
  59191=>"110101111",
  59192=>"110100000",
  59193=>"000001010",
  59194=>"000000011",
  59195=>"001101000",
  59196=>"111001101",
  59197=>"110001011",
  59198=>"000100100",
  59199=>"010100000",
  59200=>"101100101",
  59201=>"010100011",
  59202=>"110101010",
  59203=>"010111101",
  59204=>"000101001",
  59205=>"011000011",
  59206=>"000010101",
  59207=>"000000101",
  59208=>"001011001",
  59209=>"111000001",
  59210=>"100110111",
  59211=>"010111101",
  59212=>"000011010",
  59213=>"010101010",
  59214=>"100111011",
  59215=>"111000010",
  59216=>"010111011",
  59217=>"100100011",
  59218=>"101110111",
  59219=>"100010010",
  59220=>"111101001",
  59221=>"001001111",
  59222=>"000000100",
  59223=>"011110101",
  59224=>"100110111",
  59225=>"111001110",
  59226=>"001101000",
  59227=>"101111110",
  59228=>"101011000",
  59229=>"001000001",
  59230=>"011100111",
  59231=>"001100100",
  59232=>"000000011",
  59233=>"000100001",
  59234=>"001010010",
  59235=>"001011110",
  59236=>"010000010",
  59237=>"100110000",
  59238=>"100010110",
  59239=>"110110010",
  59240=>"101110100",
  59241=>"010111111",
  59242=>"000000001",
  59243=>"000010010",
  59244=>"111111010",
  59245=>"101010101",
  59246=>"101011001",
  59247=>"010101101",
  59248=>"101110101",
  59249=>"001110110",
  59250=>"011101001",
  59251=>"010000100",
  59252=>"100100000",
  59253=>"101111111",
  59254=>"000110111",
  59255=>"000000011",
  59256=>"000010001",
  59257=>"100101001",
  59258=>"101100100",
  59259=>"111011101",
  59260=>"010110000",
  59261=>"101100000",
  59262=>"011011011",
  59263=>"010100101",
  59264=>"000111111",
  59265=>"010000111",
  59266=>"011010011",
  59267=>"000011111",
  59268=>"000001100",
  59269=>"111100000",
  59270=>"110001100",
  59271=>"111000010",
  59272=>"000010000",
  59273=>"111001001",
  59274=>"001001000",
  59275=>"010001010",
  59276=>"011111111",
  59277=>"000101111",
  59278=>"010111000",
  59279=>"111001110",
  59280=>"000010101",
  59281=>"000110000",
  59282=>"000000000",
  59283=>"111000011",
  59284=>"110001100",
  59285=>"001000100",
  59286=>"100000111",
  59287=>"011011000",
  59288=>"100000111",
  59289=>"110011010",
  59290=>"001111110",
  59291=>"100100011",
  59292=>"100001100",
  59293=>"110101101",
  59294=>"110111001",
  59295=>"010001110",
  59296=>"101000001",
  59297=>"111001100",
  59298=>"011101001",
  59299=>"110101011",
  59300=>"001000000",
  59301=>"010111111",
  59302=>"010111000",
  59303=>"110111001",
  59304=>"011011000",
  59305=>"010011010",
  59306=>"011111110",
  59307=>"110011100",
  59308=>"000100111",
  59309=>"110000110",
  59310=>"001111100",
  59311=>"100101001",
  59312=>"000010100",
  59313=>"111010110",
  59314=>"010100001",
  59315=>"011100000",
  59316=>"100100100",
  59317=>"000000000",
  59318=>"111111101",
  59319=>"110000001",
  59320=>"111100101",
  59321=>"001111110",
  59322=>"001000000",
  59323=>"110010010",
  59324=>"000111101",
  59325=>"010100001",
  59326=>"110100000",
  59327=>"001110011",
  59328=>"000110011",
  59329=>"000011010",
  59330=>"111100100",
  59331=>"100111110",
  59332=>"010000100",
  59333=>"111101110",
  59334=>"100011111",
  59335=>"011110110",
  59336=>"011001010",
  59337=>"101010110",
  59338=>"111111000",
  59339=>"000100101",
  59340=>"011110111",
  59341=>"101100101",
  59342=>"100010011",
  59343=>"110001110",
  59344=>"000110001",
  59345=>"011010010",
  59346=>"100011111",
  59347=>"110100111",
  59348=>"000110110",
  59349=>"000000111",
  59350=>"011101011",
  59351=>"111001110",
  59352=>"111010000",
  59353=>"010110110",
  59354=>"010010100",
  59355=>"110111111",
  59356=>"111101100",
  59357=>"011100001",
  59358=>"000110101",
  59359=>"001001011",
  59360=>"111101111",
  59361=>"010000111",
  59362=>"111000001",
  59363=>"111101001",
  59364=>"001101111",
  59365=>"010101111",
  59366=>"110110101",
  59367=>"011011001",
  59368=>"100100001",
  59369=>"110111010",
  59370=>"000011001",
  59371=>"100101111",
  59372=>"010110110",
  59373=>"101101000",
  59374=>"011100110",
  59375=>"011001111",
  59376=>"111101010",
  59377=>"000101100",
  59378=>"100100110",
  59379=>"101110000",
  59380=>"010001101",
  59381=>"010010110",
  59382=>"111111101",
  59383=>"000110010",
  59384=>"110110111",
  59385=>"110010010",
  59386=>"001110011",
  59387=>"001010110",
  59388=>"000001010",
  59389=>"011110110",
  59390=>"110110101",
  59391=>"011000100",
  59392=>"001101001",
  59393=>"110010010",
  59394=>"000000111",
  59395=>"111011001",
  59396=>"110011110",
  59397=>"011010010",
  59398=>"110101000",
  59399=>"101110001",
  59400=>"101000001",
  59401=>"001110100",
  59402=>"110111111",
  59403=>"010100010",
  59404=>"011011011",
  59405=>"000001001",
  59406=>"110001010",
  59407=>"101111101",
  59408=>"100000000",
  59409=>"001010000",
  59410=>"000001000",
  59411=>"111001010",
  59412=>"000100000",
  59413=>"110011101",
  59414=>"101001100",
  59415=>"111001100",
  59416=>"011110110",
  59417=>"010001000",
  59418=>"010011110",
  59419=>"000011000",
  59420=>"000111010",
  59421=>"101100101",
  59422=>"001110110",
  59423=>"111001010",
  59424=>"010010101",
  59425=>"010100011",
  59426=>"110001111",
  59427=>"101101100",
  59428=>"001111001",
  59429=>"101010101",
  59430=>"111001000",
  59431=>"010001000",
  59432=>"101111001",
  59433=>"001011000",
  59434=>"100010110",
  59435=>"100101101",
  59436=>"101100001",
  59437=>"111110011",
  59438=>"001011110",
  59439=>"110001101",
  59440=>"010100111",
  59441=>"011101111",
  59442=>"000111000",
  59443=>"100000110",
  59444=>"010110110",
  59445=>"111010110",
  59446=>"000100010",
  59447=>"010110110",
  59448=>"101000010",
  59449=>"001110011",
  59450=>"110010110",
  59451=>"100111111",
  59452=>"111100101",
  59453=>"100111001",
  59454=>"100100010",
  59455=>"110000010",
  59456=>"011111001",
  59457=>"001000100",
  59458=>"100000010",
  59459=>"010101010",
  59460=>"001100000",
  59461=>"111111110",
  59462=>"000101101",
  59463=>"111000101",
  59464=>"011101000",
  59465=>"100010000",
  59466=>"101110111",
  59467=>"111010100",
  59468=>"001001000",
  59469=>"101101100",
  59470=>"110110010",
  59471=>"010101011",
  59472=>"000111011",
  59473=>"101101011",
  59474=>"011000000",
  59475=>"011001111",
  59476=>"111101000",
  59477=>"001101000",
  59478=>"110100110",
  59479=>"101111011",
  59480=>"110110100",
  59481=>"011001000",
  59482=>"001011001",
  59483=>"100101101",
  59484=>"110000000",
  59485=>"100100010",
  59486=>"001111000",
  59487=>"000100001",
  59488=>"001101110",
  59489=>"001000101",
  59490=>"000111101",
  59491=>"000101011",
  59492=>"110111101",
  59493=>"110101000",
  59494=>"100100111",
  59495=>"010100101",
  59496=>"001001110",
  59497=>"010011101",
  59498=>"011100011",
  59499=>"010000110",
  59500=>"100100001",
  59501=>"100110100",
  59502=>"011001101",
  59503=>"100111111",
  59504=>"110111110",
  59505=>"001001101",
  59506=>"010110010",
  59507=>"111111001",
  59508=>"100011110",
  59509=>"000010001",
  59510=>"111110100",
  59511=>"101100001",
  59512=>"101010110",
  59513=>"101100101",
  59514=>"010011001",
  59515=>"000111000",
  59516=>"110110101",
  59517=>"101101100",
  59518=>"111011101",
  59519=>"011110111",
  59520=>"100000011",
  59521=>"010100011",
  59522=>"010110111",
  59523=>"110111011",
  59524=>"101011100",
  59525=>"100111100",
  59526=>"110111110",
  59527=>"110000010",
  59528=>"000101010",
  59529=>"100000110",
  59530=>"111001001",
  59531=>"111101001",
  59532=>"100001110",
  59533=>"000011000",
  59534=>"101100000",
  59535=>"001001101",
  59536=>"010111111",
  59537=>"101010100",
  59538=>"011111011",
  59539=>"101110000",
  59540=>"000000001",
  59541=>"100001111",
  59542=>"000001000",
  59543=>"101110010",
  59544=>"001011101",
  59545=>"110000101",
  59546=>"001110111",
  59547=>"011101001",
  59548=>"101111001",
  59549=>"101110111",
  59550=>"101111001",
  59551=>"000110100",
  59552=>"000110111",
  59553=>"111111111",
  59554=>"101000101",
  59555=>"110101000",
  59556=>"111101001",
  59557=>"010110001",
  59558=>"111111101",
  59559=>"011001000",
  59560=>"100010101",
  59561=>"111001001",
  59562=>"110101010",
  59563=>"010011100",
  59564=>"101000011",
  59565=>"011001001",
  59566=>"111111010",
  59567=>"010101000",
  59568=>"011110101",
  59569=>"011100000",
  59570=>"100011101",
  59571=>"000001011",
  59572=>"010001001",
  59573=>"110110001",
  59574=>"100000001",
  59575=>"000100110",
  59576=>"000101100",
  59577=>"000010010",
  59578=>"010010111",
  59579=>"110001110",
  59580=>"100010000",
  59581=>"111101000",
  59582=>"000001010",
  59583=>"000001000",
  59584=>"111110111",
  59585=>"010100000",
  59586=>"010011001",
  59587=>"110000100",
  59588=>"001111001",
  59589=>"010111011",
  59590=>"101111010",
  59591=>"111111111",
  59592=>"011001000",
  59593=>"000100100",
  59594=>"000011011",
  59595=>"000100100",
  59596=>"011110110",
  59597=>"000011111",
  59598=>"100011100",
  59599=>"001100100",
  59600=>"100011110",
  59601=>"100010101",
  59602=>"101001010",
  59603=>"000101100",
  59604=>"000110100",
  59605=>"111101111",
  59606=>"011000000",
  59607=>"011100100",
  59608=>"010111001",
  59609=>"010010000",
  59610=>"010100111",
  59611=>"001010010",
  59612=>"111111100",
  59613=>"111001101",
  59614=>"101100000",
  59615=>"111101101",
  59616=>"001100111",
  59617=>"011000101",
  59618=>"000000110",
  59619=>"001100110",
  59620=>"011111100",
  59621=>"000000100",
  59622=>"101010010",
  59623=>"000011011",
  59624=>"101111110",
  59625=>"011111011",
  59626=>"110111100",
  59627=>"101100111",
  59628=>"111110011",
  59629=>"000010010",
  59630=>"011110110",
  59631=>"100001011",
  59632=>"000001111",
  59633=>"010101011",
  59634=>"000100110",
  59635=>"110100001",
  59636=>"100000000",
  59637=>"100001011",
  59638=>"000100110",
  59639=>"010010111",
  59640=>"010110100",
  59641=>"100111010",
  59642=>"100110011",
  59643=>"110100000",
  59644=>"101111011",
  59645=>"110000000",
  59646=>"011010101",
  59647=>"111101101",
  59648=>"000101100",
  59649=>"110111011",
  59650=>"100100000",
  59651=>"001111110",
  59652=>"110101011",
  59653=>"010101111",
  59654=>"001001100",
  59655=>"111111000",
  59656=>"010111000",
  59657=>"100111111",
  59658=>"011111110",
  59659=>"111010010",
  59660=>"010011100",
  59661=>"101001010",
  59662=>"001010000",
  59663=>"100101010",
  59664=>"101100111",
  59665=>"000101000",
  59666=>"010001100",
  59667=>"001110110",
  59668=>"110000110",
  59669=>"101001110",
  59670=>"000110111",
  59671=>"101011111",
  59672=>"110100110",
  59673=>"000001011",
  59674=>"111000011",
  59675=>"101110111",
  59676=>"011000111",
  59677=>"110110101",
  59678=>"000111110",
  59679=>"010001101",
  59680=>"010100011",
  59681=>"011011101",
  59682=>"000010110",
  59683=>"010110100",
  59684=>"110111001",
  59685=>"000111010",
  59686=>"000111001",
  59687=>"000100011",
  59688=>"010100011",
  59689=>"001111000",
  59690=>"111110110",
  59691=>"010110010",
  59692=>"010100100",
  59693=>"011111100",
  59694=>"010101111",
  59695=>"010000000",
  59696=>"111000111",
  59697=>"011011001",
  59698=>"001001110",
  59699=>"110011101",
  59700=>"111100110",
  59701=>"001001010",
  59702=>"000000000",
  59703=>"100100010",
  59704=>"001100011",
  59705=>"011011100",
  59706=>"010001111",
  59707=>"001000010",
  59708=>"001001001",
  59709=>"001001011",
  59710=>"111010001",
  59711=>"001111100",
  59712=>"111001010",
  59713=>"100111100",
  59714=>"100000111",
  59715=>"110111100",
  59716=>"000000001",
  59717=>"010111001",
  59718=>"101011010",
  59719=>"000001010",
  59720=>"000010010",
  59721=>"000111000",
  59722=>"010000111",
  59723=>"011000110",
  59724=>"001000011",
  59725=>"001101111",
  59726=>"000010101",
  59727=>"010010001",
  59728=>"110011000",
  59729=>"111000001",
  59730=>"111011001",
  59731=>"001110011",
  59732=>"010000110",
  59733=>"001010000",
  59734=>"100011010",
  59735=>"100100101",
  59736=>"101001111",
  59737=>"100011101",
  59738=>"111001111",
  59739=>"110000101",
  59740=>"111010111",
  59741=>"110111000",
  59742=>"011010001",
  59743=>"100111000",
  59744=>"101011010",
  59745=>"010010010",
  59746=>"100111110",
  59747=>"100010100",
  59748=>"001111011",
  59749=>"101111101",
  59750=>"100111000",
  59751=>"000101000",
  59752=>"000101010",
  59753=>"011101011",
  59754=>"100110001",
  59755=>"100001101",
  59756=>"111110111",
  59757=>"110100100",
  59758=>"101101110",
  59759=>"110101100",
  59760=>"101010011",
  59761=>"100000111",
  59762=>"010000100",
  59763=>"001100010",
  59764=>"111111101",
  59765=>"011100011",
  59766=>"101010001",
  59767=>"110111001",
  59768=>"001101101",
  59769=>"111010000",
  59770=>"111011000",
  59771=>"111011010",
  59772=>"110110101",
  59773=>"000001100",
  59774=>"000111100",
  59775=>"101101011",
  59776=>"000101001",
  59777=>"000110001",
  59778=>"110000101",
  59779=>"000110001",
  59780=>"011101011",
  59781=>"101010000",
  59782=>"110101100",
  59783=>"011110111",
  59784=>"100110100",
  59785=>"111110001",
  59786=>"100001000",
  59787=>"100011110",
  59788=>"000111000",
  59789=>"111000111",
  59790=>"010100001",
  59791=>"011101110",
  59792=>"101010000",
  59793=>"101110100",
  59794=>"101111010",
  59795=>"000000010",
  59796=>"000101100",
  59797=>"001001111",
  59798=>"100001011",
  59799=>"101100000",
  59800=>"011100000",
  59801=>"000101101",
  59802=>"001001010",
  59803=>"001100111",
  59804=>"111010010",
  59805=>"101110110",
  59806=>"110100111",
  59807=>"110110110",
  59808=>"100111110",
  59809=>"101100001",
  59810=>"011101010",
  59811=>"000010110",
  59812=>"101110110",
  59813=>"011101000",
  59814=>"000010000",
  59815=>"100111011",
  59816=>"000100000",
  59817=>"001001010",
  59818=>"100011101",
  59819=>"011000010",
  59820=>"100001101",
  59821=>"111011101",
  59822=>"011100100",
  59823=>"011111011",
  59824=>"110100110",
  59825=>"000011010",
  59826=>"110010101",
  59827=>"111001100",
  59828=>"111111001",
  59829=>"010001101",
  59830=>"100110011",
  59831=>"001000101",
  59832=>"111000111",
  59833=>"010010001",
  59834=>"101110110",
  59835=>"101110001",
  59836=>"111000101",
  59837=>"110101011",
  59838=>"001110100",
  59839=>"110111001",
  59840=>"110010101",
  59841=>"100111011",
  59842=>"110111101",
  59843=>"110000111",
  59844=>"100000001",
  59845=>"110000011",
  59846=>"001000000",
  59847=>"010010001",
  59848=>"101100001",
  59849=>"011100100",
  59850=>"101111111",
  59851=>"000010010",
  59852=>"111011101",
  59853=>"000001010",
  59854=>"010101001",
  59855=>"110001001",
  59856=>"100000110",
  59857=>"011100000",
  59858=>"101010010",
  59859=>"011111100",
  59860=>"011011001",
  59861=>"100000000",
  59862=>"000110101",
  59863=>"001100110",
  59864=>"101110100",
  59865=>"001010011",
  59866=>"000000001",
  59867=>"110000110",
  59868=>"010111011",
  59869=>"001000000",
  59870=>"111000101",
  59871=>"011000111",
  59872=>"111000011",
  59873=>"101011101",
  59874=>"110010100",
  59875=>"011101000",
  59876=>"101011111",
  59877=>"100101111",
  59878=>"110110101",
  59879=>"101101111",
  59880=>"101000010",
  59881=>"011001101",
  59882=>"100011011",
  59883=>"111110000",
  59884=>"010111000",
  59885=>"110100110",
  59886=>"110111111",
  59887=>"101000100",
  59888=>"001100111",
  59889=>"111111101",
  59890=>"110000111",
  59891=>"001000000",
  59892=>"110110001",
  59893=>"000011010",
  59894=>"111011000",
  59895=>"110000011",
  59896=>"000000010",
  59897=>"010011111",
  59898=>"110011011",
  59899=>"111011010",
  59900=>"111101001",
  59901=>"100111100",
  59902=>"101011100",
  59903=>"111111101",
  59904=>"000000000",
  59905=>"010001011",
  59906=>"010101000",
  59907=>"010000010",
  59908=>"111010101",
  59909=>"000011000",
  59910=>"110001110",
  59911=>"101001111",
  59912=>"101110110",
  59913=>"101101101",
  59914=>"111011110",
  59915=>"001101110",
  59916=>"010011101",
  59917=>"001001100",
  59918=>"101110010",
  59919=>"000000111",
  59920=>"000111101",
  59921=>"010011000",
  59922=>"001010111",
  59923=>"110001111",
  59924=>"001101110",
  59925=>"011110000",
  59926=>"110001101",
  59927=>"111001000",
  59928=>"101000000",
  59929=>"010110110",
  59930=>"110101000",
  59931=>"010011111",
  59932=>"000101000",
  59933=>"110111100",
  59934=>"111101010",
  59935=>"100110101",
  59936=>"001011100",
  59937=>"101110110",
  59938=>"011000101",
  59939=>"100000001",
  59940=>"110100110",
  59941=>"101011000",
  59942=>"111001010",
  59943=>"100111110",
  59944=>"001000011",
  59945=>"111000111",
  59946=>"101010100",
  59947=>"111110000",
  59948=>"111011110",
  59949=>"011110000",
  59950=>"111000001",
  59951=>"011101110",
  59952=>"000100101",
  59953=>"101101100",
  59954=>"000100110",
  59955=>"001010011",
  59956=>"001011010",
  59957=>"000110001",
  59958=>"001000011",
  59959=>"000011110",
  59960=>"110111001",
  59961=>"010010001",
  59962=>"011011110",
  59963=>"011001101",
  59964=>"000111001",
  59965=>"100110111",
  59966=>"001000011",
  59967=>"000110110",
  59968=>"111000111",
  59969=>"100111010",
  59970=>"001000000",
  59971=>"011001110",
  59972=>"100110110",
  59973=>"011001000",
  59974=>"100110011",
  59975=>"010001010",
  59976=>"110001111",
  59977=>"100000000",
  59978=>"100000010",
  59979=>"100000000",
  59980=>"100000001",
  59981=>"111010011",
  59982=>"101000010",
  59983=>"111110101",
  59984=>"010100100",
  59985=>"000110011",
  59986=>"101000110",
  59987=>"010011010",
  59988=>"001011111",
  59989=>"000111010",
  59990=>"110111101",
  59991=>"100101011",
  59992=>"000100001",
  59993=>"100011011",
  59994=>"000101011",
  59995=>"000111010",
  59996=>"010010111",
  59997=>"110011101",
  59998=>"000111010",
  59999=>"101010001",
  60000=>"111011010",
  60001=>"100010101",
  60002=>"000000000",
  60003=>"000010101",
  60004=>"100111110",
  60005=>"101101010",
  60006=>"010101101",
  60007=>"001100100",
  60008=>"110100111",
  60009=>"110111010",
  60010=>"111111100",
  60011=>"100111111",
  60012=>"001110110",
  60013=>"111110111",
  60014=>"000110110",
  60015=>"111110000",
  60016=>"000101001",
  60017=>"010000010",
  60018=>"110001011",
  60019=>"001111101",
  60020=>"110101100",
  60021=>"000101000",
  60022=>"100010011",
  60023=>"110111101",
  60024=>"101011011",
  60025=>"010000100",
  60026=>"010100011",
  60027=>"101100001",
  60028=>"000110101",
  60029=>"011111011",
  60030=>"010110100",
  60031=>"011010010",
  60032=>"110110110",
  60033=>"110001011",
  60034=>"010111010",
  60035=>"110101011",
  60036=>"010110100",
  60037=>"001001010",
  60038=>"101111110",
  60039=>"000111000",
  60040=>"011001001",
  60041=>"101101011",
  60042=>"000011100",
  60043=>"011111011",
  60044=>"100111001",
  60045=>"000101110",
  60046=>"101010101",
  60047=>"001001000",
  60048=>"100111010",
  60049=>"101110011",
  60050=>"010111100",
  60051=>"000101010",
  60052=>"111100110",
  60053=>"110101101",
  60054=>"011111111",
  60055=>"001110011",
  60056=>"101111101",
  60057=>"001000100",
  60058=>"110011010",
  60059=>"011000100",
  60060=>"101011010",
  60061=>"110100011",
  60062=>"110000011",
  60063=>"010000100",
  60064=>"110101000",
  60065=>"011001110",
  60066=>"000011010",
  60067=>"111000100",
  60068=>"010111110",
  60069=>"011110110",
  60070=>"100101010",
  60071=>"010001000",
  60072=>"001010001",
  60073=>"101110100",
  60074=>"110001110",
  60075=>"101010100",
  60076=>"111100111",
  60077=>"110010111",
  60078=>"101110111",
  60079=>"101010010",
  60080=>"100100111",
  60081=>"000011000",
  60082=>"101010000",
  60083=>"001010000",
  60084=>"101000010",
  60085=>"111111101",
  60086=>"101010100",
  60087=>"100001110",
  60088=>"010001101",
  60089=>"001100100",
  60090=>"000011101",
  60091=>"010100101",
  60092=>"011100000",
  60093=>"110111100",
  60094=>"111000100",
  60095=>"101000000",
  60096=>"111101001",
  60097=>"111010111",
  60098=>"000000011",
  60099=>"001111101",
  60100=>"011111010",
  60101=>"110011000",
  60102=>"101110110",
  60103=>"001011100",
  60104=>"111011010",
  60105=>"000000010",
  60106=>"001010011",
  60107=>"110100110",
  60108=>"000001101",
  60109=>"011011100",
  60110=>"010100001",
  60111=>"001101011",
  60112=>"100101001",
  60113=>"000101110",
  60114=>"011111010",
  60115=>"011011000",
  60116=>"001100000",
  60117=>"000001101",
  60118=>"000110010",
  60119=>"010101010",
  60120=>"000000001",
  60121=>"100001010",
  60122=>"100100000",
  60123=>"011001110",
  60124=>"111101100",
  60125=>"111111100",
  60126=>"110101100",
  60127=>"110110010",
  60128=>"111011001",
  60129=>"100010111",
  60130=>"111100000",
  60131=>"000111001",
  60132=>"100110100",
  60133=>"111110000",
  60134=>"100111011",
  60135=>"100111001",
  60136=>"001001000",
  60137=>"101001101",
  60138=>"110010110",
  60139=>"000011100",
  60140=>"110001010",
  60141=>"101010111",
  60142=>"100110010",
  60143=>"011010011",
  60144=>"110000111",
  60145=>"100111111",
  60146=>"011010110",
  60147=>"000111100",
  60148=>"111011100",
  60149=>"000001011",
  60150=>"111111101",
  60151=>"111101010",
  60152=>"011101000",
  60153=>"000001110",
  60154=>"110000001",
  60155=>"110011101",
  60156=>"111001001",
  60157=>"001000111",
  60158=>"001111010",
  60159=>"110110110",
  60160=>"001100011",
  60161=>"110010010",
  60162=>"111111010",
  60163=>"001000000",
  60164=>"110000110",
  60165=>"101111111",
  60166=>"000100010",
  60167=>"101000101",
  60168=>"110000000",
  60169=>"110000111",
  60170=>"001101001",
  60171=>"000111000",
  60172=>"001100110",
  60173=>"000111011",
  60174=>"000010010",
  60175=>"010000110",
  60176=>"010111000",
  60177=>"111010111",
  60178=>"100101010",
  60179=>"110011011",
  60180=>"111001110",
  60181=>"101101100",
  60182=>"101011010",
  60183=>"100001000",
  60184=>"100000111",
  60185=>"100001111",
  60186=>"111010100",
  60187=>"000101101",
  60188=>"001110111",
  60189=>"111001000",
  60190=>"000011100",
  60191=>"011000111",
  60192=>"010001101",
  60193=>"011011101",
  60194=>"011101111",
  60195=>"111110111",
  60196=>"011010100",
  60197=>"010000001",
  60198=>"111111101",
  60199=>"111000000",
  60200=>"100101000",
  60201=>"000101011",
  60202=>"100100011",
  60203=>"110100101",
  60204=>"110111111",
  60205=>"111010101",
  60206=>"000000011",
  60207=>"110000000",
  60208=>"110100111",
  60209=>"010101011",
  60210=>"011000011",
  60211=>"101101100",
  60212=>"110111100",
  60213=>"101111110",
  60214=>"111110100",
  60215=>"101100111",
  60216=>"110101000",
  60217=>"011001001",
  60218=>"001001100",
  60219=>"111100100",
  60220=>"010111110",
  60221=>"110000011",
  60222=>"000001000",
  60223=>"111110101",
  60224=>"011101111",
  60225=>"010011000",
  60226=>"100110000",
  60227=>"101110011",
  60228=>"111000100",
  60229=>"010010001",
  60230=>"010000011",
  60231=>"011111111",
  60232=>"001000000",
  60233=>"111110101",
  60234=>"011001111",
  60235=>"001010110",
  60236=>"001110000",
  60237=>"101000011",
  60238=>"000011000",
  60239=>"011100001",
  60240=>"000001010",
  60241=>"111000110",
  60242=>"000110101",
  60243=>"111110000",
  60244=>"110101010",
  60245=>"110101000",
  60246=>"011111111",
  60247=>"011100101",
  60248=>"101000110",
  60249=>"000110101",
  60250=>"010100100",
  60251=>"110111001",
  60252=>"001101010",
  60253=>"000010111",
  60254=>"101001111",
  60255=>"111101010",
  60256=>"011100010",
  60257=>"001100000",
  60258=>"100010100",
  60259=>"010011000",
  60260=>"111110110",
  60261=>"010010101",
  60262=>"110111001",
  60263=>"000001001",
  60264=>"111001010",
  60265=>"001000010",
  60266=>"001100001",
  60267=>"011001101",
  60268=>"000011111",
  60269=>"001100101",
  60270=>"011110000",
  60271=>"011110001",
  60272=>"100000111",
  60273=>"010101010",
  60274=>"001110000",
  60275=>"100001000",
  60276=>"010010110",
  60277=>"001000011",
  60278=>"101110010",
  60279=>"000110110",
  60280=>"111110110",
  60281=>"110000000",
  60282=>"100111000",
  60283=>"110011001",
  60284=>"010010010",
  60285=>"101111010",
  60286=>"101001000",
  60287=>"110111000",
  60288=>"010101000",
  60289=>"000101100",
  60290=>"001100010",
  60291=>"000111100",
  60292=>"110001001",
  60293=>"011001001",
  60294=>"011111111",
  60295=>"001110011",
  60296=>"100100111",
  60297=>"011110110",
  60298=>"001110101",
  60299=>"011011000",
  60300=>"100010000",
  60301=>"110101101",
  60302=>"110101011",
  60303=>"101010111",
  60304=>"010111101",
  60305=>"111011011",
  60306=>"010110100",
  60307=>"100100111",
  60308=>"110000011",
  60309=>"010100010",
  60310=>"110001111",
  60311=>"111101001",
  60312=>"010100000",
  60313=>"100111011",
  60314=>"101101001",
  60315=>"100000100",
  60316=>"000111110",
  60317=>"011010001",
  60318=>"110000111",
  60319=>"111110001",
  60320=>"101100110",
  60321=>"011110100",
  60322=>"010101111",
  60323=>"101101100",
  60324=>"111011110",
  60325=>"110011000",
  60326=>"110010100",
  60327=>"110110010",
  60328=>"100000001",
  60329=>"000100001",
  60330=>"000111011",
  60331=>"011010000",
  60332=>"010001011",
  60333=>"100000000",
  60334=>"101111111",
  60335=>"101001011",
  60336=>"010100011",
  60337=>"001101111",
  60338=>"010111111",
  60339=>"000100001",
  60340=>"001010100",
  60341=>"110001101",
  60342=>"011100001",
  60343=>"000110110",
  60344=>"011110101",
  60345=>"101101010",
  60346=>"110000000",
  60347=>"110100100",
  60348=>"000111111",
  60349=>"100111111",
  60350=>"011000101",
  60351=>"001001101",
  60352=>"001111011",
  60353=>"110010001",
  60354=>"100100111",
  60355=>"100100010",
  60356=>"001010100",
  60357=>"010011000",
  60358=>"001000011",
  60359=>"000100110",
  60360=>"110101001",
  60361=>"011000000",
  60362=>"011100001",
  60363=>"111111000",
  60364=>"011110101",
  60365=>"100001100",
  60366=>"000110111",
  60367=>"010101111",
  60368=>"101101100",
  60369=>"000101011",
  60370=>"011110010",
  60371=>"100000010",
  60372=>"101011010",
  60373=>"010001100",
  60374=>"101000000",
  60375=>"101000000",
  60376=>"010001001",
  60377=>"110111111",
  60378=>"101111100",
  60379=>"000000100",
  60380=>"110000010",
  60381=>"000000100",
  60382=>"111101010",
  60383=>"111100110",
  60384=>"100011001",
  60385=>"111101000",
  60386=>"010101001",
  60387=>"000111011",
  60388=>"111100101",
  60389=>"000111111",
  60390=>"011100000",
  60391=>"101111111",
  60392=>"101100101",
  60393=>"011011110",
  60394=>"000010100",
  60395=>"000000111",
  60396=>"011011111",
  60397=>"110111000",
  60398=>"001001010",
  60399=>"011010010",
  60400=>"110111011",
  60401=>"110010011",
  60402=>"000001001",
  60403=>"101101010",
  60404=>"001101111",
  60405=>"011110010",
  60406=>"011110011",
  60407=>"010011011",
  60408=>"010010011",
  60409=>"001101000",
  60410=>"010111001",
  60411=>"000110000",
  60412=>"001111100",
  60413=>"110011011",
  60414=>"101000101",
  60415=>"000001101",
  60416=>"101110010",
  60417=>"010110101",
  60418=>"001000000",
  60419=>"000000010",
  60420=>"100100001",
  60421=>"100000001",
  60422=>"010110000",
  60423=>"110111001",
  60424=>"000000011",
  60425=>"110101101",
  60426=>"011101101",
  60427=>"001001011",
  60428=>"101100010",
  60429=>"011110100",
  60430=>"001100000",
  60431=>"000110000",
  60432=>"100011101",
  60433=>"011110110",
  60434=>"101001000",
  60435=>"111111110",
  60436=>"100011011",
  60437=>"001101101",
  60438=>"010110001",
  60439=>"010000000",
  60440=>"011000010",
  60441=>"011011000",
  60442=>"110110010",
  60443=>"001001011",
  60444=>"100001111",
  60445=>"011010101",
  60446=>"101011010",
  60447=>"111000100",
  60448=>"100010001",
  60449=>"001000111",
  60450=>"000000011",
  60451=>"110001011",
  60452=>"111000111",
  60453=>"000011100",
  60454=>"001110000",
  60455=>"000111110",
  60456=>"100010101",
  60457=>"000101001",
  60458=>"101001001",
  60459=>"010101010",
  60460=>"111011001",
  60461=>"110011110",
  60462=>"100111100",
  60463=>"101010111",
  60464=>"010010011",
  60465=>"010011001",
  60466=>"011011110",
  60467=>"111111100",
  60468=>"010111010",
  60469=>"101001100",
  60470=>"000011000",
  60471=>"101010000",
  60472=>"000100011",
  60473=>"000000011",
  60474=>"011110011",
  60475=>"101000011",
  60476=>"111111111",
  60477=>"101001111",
  60478=>"000110111",
  60479=>"001111100",
  60480=>"011010100",
  60481=>"101000111",
  60482=>"111101000",
  60483=>"011010001",
  60484=>"010100000",
  60485=>"101110001",
  60486=>"010111001",
  60487=>"011101010",
  60488=>"001011001",
  60489=>"100100111",
  60490=>"100101001",
  60491=>"000001011",
  60492=>"101010011",
  60493=>"011111101",
  60494=>"110100001",
  60495=>"011101110",
  60496=>"100011000",
  60497=>"100100100",
  60498=>"000110010",
  60499=>"101001011",
  60500=>"010010101",
  60501=>"101100000",
  60502=>"001100101",
  60503=>"000010010",
  60504=>"110001001",
  60505=>"110101101",
  60506=>"011100010",
  60507=>"000011100",
  60508=>"100110111",
  60509=>"001101100",
  60510=>"110110100",
  60511=>"000011101",
  60512=>"000100100",
  60513=>"110000011",
  60514=>"000010100",
  60515=>"101100001",
  60516=>"011101111",
  60517=>"111101100",
  60518=>"101101100",
  60519=>"000101100",
  60520=>"110101111",
  60521=>"101001110",
  60522=>"100101101",
  60523=>"100001111",
  60524=>"011001111",
  60525=>"101110000",
  60526=>"101111100",
  60527=>"010101010",
  60528=>"001101111",
  60529=>"010111111",
  60530=>"001101001",
  60531=>"011000100",
  60532=>"100101001",
  60533=>"110001001",
  60534=>"101100110",
  60535=>"001100110",
  60536=>"111000010",
  60537=>"011010111",
  60538=>"111110111",
  60539=>"100000101",
  60540=>"010100000",
  60541=>"110110110",
  60542=>"000100000",
  60543=>"111011111",
  60544=>"101011001",
  60545=>"111011010",
  60546=>"111100100",
  60547=>"011111110",
  60548=>"101010110",
  60549=>"111011100",
  60550=>"111001001",
  60551=>"010010010",
  60552=>"110111111",
  60553=>"011100000",
  60554=>"011111100",
  60555=>"110101101",
  60556=>"100010100",
  60557=>"011110100",
  60558=>"100110101",
  60559=>"100010101",
  60560=>"110101000",
  60561=>"110100001",
  60562=>"111100001",
  60563=>"110111111",
  60564=>"111011110",
  60565=>"100001011",
  60566=>"010001110",
  60567=>"011011010",
  60568=>"101110100",
  60569=>"111001010",
  60570=>"011011010",
  60571=>"110011111",
  60572=>"110001100",
  60573=>"111111011",
  60574=>"110010010",
  60575=>"011111111",
  60576=>"110001010",
  60577=>"000100001",
  60578=>"010010010",
  60579=>"100111111",
  60580=>"011010010",
  60581=>"111011101",
  60582=>"100010000",
  60583=>"000111010",
  60584=>"100000101",
  60585=>"101011001",
  60586=>"010110011",
  60587=>"111101111",
  60588=>"100010010",
  60589=>"000110010",
  60590=>"111110111",
  60591=>"100001111",
  60592=>"111111111",
  60593=>"010110100",
  60594=>"011111000",
  60595=>"111011111",
  60596=>"011101100",
  60597=>"010010101",
  60598=>"111001000",
  60599=>"111100011",
  60600=>"111010100",
  60601=>"101111100",
  60602=>"000110010",
  60603=>"100101101",
  60604=>"111011101",
  60605=>"111101011",
  60606=>"000001111",
  60607=>"001111000",
  60608=>"011011101",
  60609=>"101111100",
  60610=>"001111110",
  60611=>"000000001",
  60612=>"000001110",
  60613=>"111101111",
  60614=>"000010101",
  60615=>"010011101",
  60616=>"011010110",
  60617=>"111010000",
  60618=>"111010010",
  60619=>"000000010",
  60620=>"000001101",
  60621=>"000011000",
  60622=>"110000100",
  60623=>"101111100",
  60624=>"011010010",
  60625=>"000000000",
  60626=>"000101000",
  60627=>"011010110",
  60628=>"010110001",
  60629=>"011100110",
  60630=>"100010111",
  60631=>"010000010",
  60632=>"111000010",
  60633=>"000010101",
  60634=>"011110001",
  60635=>"011000110",
  60636=>"110000010",
  60637=>"011011010",
  60638=>"110011100",
  60639=>"110110100",
  60640=>"000111000",
  60641=>"000111000",
  60642=>"011011111",
  60643=>"000001001",
  60644=>"000111101",
  60645=>"111111100",
  60646=>"111111111",
  60647=>"101000111",
  60648=>"010100101",
  60649=>"010001000",
  60650=>"000010000",
  60651=>"010000101",
  60652=>"010010010",
  60653=>"001110100",
  60654=>"010000111",
  60655=>"011010100",
  60656=>"000100011",
  60657=>"110111000",
  60658=>"101101111",
  60659=>"001011110",
  60660=>"100111111",
  60661=>"111111000",
  60662=>"111010100",
  60663=>"101010000",
  60664=>"011101011",
  60665=>"001010000",
  60666=>"000100100",
  60667=>"111110000",
  60668=>"110110000",
  60669=>"000010000",
  60670=>"001111000",
  60671=>"111100111",
  60672=>"010100000",
  60673=>"101000101",
  60674=>"110101000",
  60675=>"000010001",
  60676=>"101011011",
  60677=>"010100001",
  60678=>"111010010",
  60679=>"101010101",
  60680=>"101111011",
  60681=>"010000010",
  60682=>"001100101",
  60683=>"001010000",
  60684=>"000011110",
  60685=>"010000011",
  60686=>"001010001",
  60687=>"000101101",
  60688=>"100100100",
  60689=>"000111111",
  60690=>"001000100",
  60691=>"111001000",
  60692=>"010101010",
  60693=>"111001010",
  60694=>"111111001",
  60695=>"001001100",
  60696=>"110001011",
  60697=>"010110111",
  60698=>"011111101",
  60699=>"111111011",
  60700=>"110001101",
  60701=>"110001101",
  60702=>"111111110",
  60703=>"010000010",
  60704=>"011011011",
  60705=>"011101111",
  60706=>"110000001",
  60707=>"111100101",
  60708=>"011001010",
  60709=>"011101001",
  60710=>"010111100",
  60711=>"011101111",
  60712=>"111010011",
  60713=>"011111110",
  60714=>"100000101",
  60715=>"000110001",
  60716=>"111010110",
  60717=>"001101001",
  60718=>"001101000",
  60719=>"010001101",
  60720=>"110101111",
  60721=>"010000001",
  60722=>"001010111",
  60723=>"000010101",
  60724=>"000000010",
  60725=>"100111010",
  60726=>"111101011",
  60727=>"011100101",
  60728=>"111010101",
  60729=>"111000101",
  60730=>"001111101",
  60731=>"100101000",
  60732=>"001110110",
  60733=>"101011001",
  60734=>"110110101",
  60735=>"110000100",
  60736=>"111001110",
  60737=>"111110110",
  60738=>"011000011",
  60739=>"101000111",
  60740=>"110100000",
  60741=>"100101010",
  60742=>"101000100",
  60743=>"101010101",
  60744=>"000010001",
  60745=>"100000001",
  60746=>"010110000",
  60747=>"111110101",
  60748=>"000101011",
  60749=>"111111100",
  60750=>"110010001",
  60751=>"000100101",
  60752=>"100111111",
  60753=>"001001000",
  60754=>"001010010",
  60755=>"100101111",
  60756=>"100010111",
  60757=>"011000011",
  60758=>"000001001",
  60759=>"100111100",
  60760=>"010100111",
  60761=>"110110001",
  60762=>"000000110",
  60763=>"111011001",
  60764=>"010111101",
  60765=>"100111110",
  60766=>"010101000",
  60767=>"000011000",
  60768=>"001100010",
  60769=>"110001011",
  60770=>"011100101",
  60771=>"100010100",
  60772=>"111101111",
  60773=>"010111101",
  60774=>"001100001",
  60775=>"100001110",
  60776=>"011101100",
  60777=>"011000100",
  60778=>"100111101",
  60779=>"011110110",
  60780=>"010100000",
  60781=>"000011011",
  60782=>"101110100",
  60783=>"010110111",
  60784=>"101011011",
  60785=>"000111000",
  60786=>"000000111",
  60787=>"101001010",
  60788=>"110010110",
  60789=>"011011100",
  60790=>"011010100",
  60791=>"101101011",
  60792=>"010011101",
  60793=>"110111011",
  60794=>"010110010",
  60795=>"010111101",
  60796=>"111001011",
  60797=>"001011000",
  60798=>"111010110",
  60799=>"000100111",
  60800=>"010001100",
  60801=>"010000011",
  60802=>"100001101",
  60803=>"110100011",
  60804=>"011110000",
  60805=>"010010111",
  60806=>"001001111",
  60807=>"010010000",
  60808=>"100011011",
  60809=>"101011101",
  60810=>"011001110",
  60811=>"101111011",
  60812=>"110111011",
  60813=>"111110100",
  60814=>"101101100",
  60815=>"111011101",
  60816=>"010111100",
  60817=>"010111111",
  60818=>"011000011",
  60819=>"100111010",
  60820=>"101010111",
  60821=>"000010001",
  60822=>"111101100",
  60823=>"011100001",
  60824=>"110101100",
  60825=>"011001111",
  60826=>"000111100",
  60827=>"110100010",
  60828=>"111011111",
  60829=>"011000100",
  60830=>"101110111",
  60831=>"010110110",
  60832=>"101101111",
  60833=>"001111011",
  60834=>"100010101",
  60835=>"011001010",
  60836=>"100000010",
  60837=>"001100110",
  60838=>"110110011",
  60839=>"001110000",
  60840=>"110011011",
  60841=>"100011111",
  60842=>"000111100",
  60843=>"111010011",
  60844=>"101101110",
  60845=>"100110001",
  60846=>"101001101",
  60847=>"111100010",
  60848=>"001100100",
  60849=>"101100100",
  60850=>"010011001",
  60851=>"100110010",
  60852=>"010111101",
  60853=>"111010010",
  60854=>"100001011",
  60855=>"000001100",
  60856=>"111000000",
  60857=>"111010100",
  60858=>"000000011",
  60859=>"010001010",
  60860=>"101101100",
  60861=>"011000101",
  60862=>"110111010",
  60863=>"100010100",
  60864=>"001100010",
  60865=>"100001110",
  60866=>"111111010",
  60867=>"111101110",
  60868=>"000101001",
  60869=>"111001111",
  60870=>"010101101",
  60871=>"101111011",
  60872=>"010010011",
  60873=>"110010010",
  60874=>"010010000",
  60875=>"000001010",
  60876=>"100011100",
  60877=>"111001010",
  60878=>"111101100",
  60879=>"100100010",
  60880=>"110100100",
  60881=>"110111101",
  60882=>"100000001",
  60883=>"110101000",
  60884=>"011101100",
  60885=>"101111110",
  60886=>"101001110",
  60887=>"100010010",
  60888=>"101001101",
  60889=>"101111101",
  60890=>"011001101",
  60891=>"110001001",
  60892=>"100010110",
  60893=>"100111000",
  60894=>"001100101",
  60895=>"111000111",
  60896=>"110110100",
  60897=>"101111111",
  60898=>"010101111",
  60899=>"100111110",
  60900=>"110001001",
  60901=>"000100100",
  60902=>"011111001",
  60903=>"010010010",
  60904=>"001101001",
  60905=>"000111001",
  60906=>"010011111",
  60907=>"101100101",
  60908=>"000000011",
  60909=>"000111110",
  60910=>"100111010",
  60911=>"000010010",
  60912=>"001010001",
  60913=>"001011100",
  60914=>"110100100",
  60915=>"000100001",
  60916=>"110110001",
  60917=>"101010000",
  60918=>"100111110",
  60919=>"001010010",
  60920=>"011001001",
  60921=>"100110010",
  60922=>"100100101",
  60923=>"100001101",
  60924=>"100110110",
  60925=>"000101100",
  60926=>"010010011",
  60927=>"011001010",
  60928=>"111101001",
  60929=>"000001000",
  60930=>"100111011",
  60931=>"111101101",
  60932=>"101101100",
  60933=>"000101000",
  60934=>"110010000",
  60935=>"001111110",
  60936=>"100110000",
  60937=>"000111101",
  60938=>"111010010",
  60939=>"101001100",
  60940=>"111000001",
  60941=>"110111000",
  60942=>"111100000",
  60943=>"001111100",
  60944=>"100100010",
  60945=>"100001100",
  60946=>"111011111",
  60947=>"111011111",
  60948=>"111000000",
  60949=>"000001101",
  60950=>"111100001",
  60951=>"010011110",
  60952=>"100111011",
  60953=>"111100010",
  60954=>"000100000",
  60955=>"100110111",
  60956=>"101110111",
  60957=>"011001111",
  60958=>"110010011",
  60959=>"001111011",
  60960=>"000010110",
  60961=>"010000011",
  60962=>"011001001",
  60963=>"111000100",
  60964=>"010001100",
  60965=>"111101001",
  60966=>"001000110",
  60967=>"110000110",
  60968=>"101100110",
  60969=>"101100001",
  60970=>"101011101",
  60971=>"100111101",
  60972=>"110010111",
  60973=>"000100100",
  60974=>"011111000",
  60975=>"101011101",
  60976=>"101111101",
  60977=>"010011010",
  60978=>"100110000",
  60979=>"010110001",
  60980=>"100001111",
  60981=>"001101100",
  60982=>"111001010",
  60983=>"101100111",
  60984=>"101111011",
  60985=>"100000000",
  60986=>"010110101",
  60987=>"100111010",
  60988=>"111111001",
  60989=>"000111100",
  60990=>"000001011",
  60991=>"110011001",
  60992=>"011001010",
  60993=>"111000100",
  60994=>"110011000",
  60995=>"010101000",
  60996=>"001000001",
  60997=>"001110111",
  60998=>"000010000",
  60999=>"001001011",
  61000=>"000000011",
  61001=>"101011011",
  61002=>"110100011",
  61003=>"010011011",
  61004=>"101011111",
  61005=>"001001000",
  61006=>"100010011",
  61007=>"001011110",
  61008=>"000111101",
  61009=>"000001100",
  61010=>"010101100",
  61011=>"011100110",
  61012=>"100110110",
  61013=>"011101001",
  61014=>"111011001",
  61015=>"111101001",
  61016=>"010100010",
  61017=>"000101111",
  61018=>"000011001",
  61019=>"010111101",
  61020=>"011010000",
  61021=>"010000000",
  61022=>"000000001",
  61023=>"100101110",
  61024=>"101111010",
  61025=>"001100001",
  61026=>"011010010",
  61027=>"001011000",
  61028=>"010000101",
  61029=>"110111100",
  61030=>"111010101",
  61031=>"111000111",
  61032=>"101000101",
  61033=>"111010000",
  61034=>"001001101",
  61035=>"110011001",
  61036=>"101011110",
  61037=>"101100010",
  61038=>"101111110",
  61039=>"010000010",
  61040=>"100010000",
  61041=>"110000000",
  61042=>"000000011",
  61043=>"110111111",
  61044=>"110000000",
  61045=>"000000100",
  61046=>"111000000",
  61047=>"110011100",
  61048=>"011011101",
  61049=>"111100001",
  61050=>"111101110",
  61051=>"111101000",
  61052=>"001111110",
  61053=>"000110111",
  61054=>"010000100",
  61055=>"111111101",
  61056=>"100001111",
  61057=>"111000001",
  61058=>"110111111",
  61059=>"010010111",
  61060=>"001100110",
  61061=>"010000010",
  61062=>"111010111",
  61063=>"000011011",
  61064=>"000101000",
  61065=>"011010110",
  61066=>"010101011",
  61067=>"010101010",
  61068=>"000010011",
  61069=>"100011000",
  61070=>"010110110",
  61071=>"100100011",
  61072=>"101111001",
  61073=>"011011000",
  61074=>"100111000",
  61075=>"001110010",
  61076=>"010111010",
  61077=>"000101101",
  61078=>"100101001",
  61079=>"110111101",
  61080=>"000101010",
  61081=>"111100101",
  61082=>"010101101",
  61083=>"110000111",
  61084=>"111011000",
  61085=>"100101100",
  61086=>"100000010",
  61087=>"100001101",
  61088=>"110100111",
  61089=>"111100000",
  61090=>"011100100",
  61091=>"100011110",
  61092=>"100011010",
  61093=>"010101000",
  61094=>"001111111",
  61095=>"111000001",
  61096=>"111101111",
  61097=>"100100010",
  61098=>"011110101",
  61099=>"111110011",
  61100=>"100111111",
  61101=>"111010100",
  61102=>"010111001",
  61103=>"100010110",
  61104=>"001101010",
  61105=>"101101101",
  61106=>"101101111",
  61107=>"001110101",
  61108=>"000110111",
  61109=>"111000010",
  61110=>"011010000",
  61111=>"111011001",
  61112=>"101010111",
  61113=>"111000010",
  61114=>"000110001",
  61115=>"000000100",
  61116=>"101000101",
  61117=>"001011000",
  61118=>"111110110",
  61119=>"011000010",
  61120=>"111110000",
  61121=>"111000110",
  61122=>"010111000",
  61123=>"100111101",
  61124=>"001111011",
  61125=>"010110000",
  61126=>"110000000",
  61127=>"001111100",
  61128=>"001001000",
  61129=>"101101101",
  61130=>"000101000",
  61131=>"100001000",
  61132=>"110011001",
  61133=>"101110001",
  61134=>"100100111",
  61135=>"011101110",
  61136=>"001000001",
  61137=>"001010010",
  61138=>"001110101",
  61139=>"001111110",
  61140=>"010100100",
  61141=>"100011111",
  61142=>"100111010",
  61143=>"110111110",
  61144=>"000100001",
  61145=>"000011001",
  61146=>"101001011",
  61147=>"010001101",
  61148=>"010001000",
  61149=>"111100000",
  61150=>"000000010",
  61151=>"000001010",
  61152=>"010011001",
  61153=>"100010111",
  61154=>"110101100",
  61155=>"000000101",
  61156=>"000001110",
  61157=>"001101111",
  61158=>"000010001",
  61159=>"000001111",
  61160=>"000100000",
  61161=>"010110110",
  61162=>"101111100",
  61163=>"110011111",
  61164=>"010011110",
  61165=>"000011110",
  61166=>"000101110",
  61167=>"111001111",
  61168=>"110100011",
  61169=>"010100011",
  61170=>"111111110",
  61171=>"000101100",
  61172=>"101110011",
  61173=>"011001100",
  61174=>"111101111",
  61175=>"001000110",
  61176=>"011101011",
  61177=>"010000110",
  61178=>"111010000",
  61179=>"010110011",
  61180=>"100100100",
  61181=>"110011101",
  61182=>"100000000",
  61183=>"101000110",
  61184=>"111010010",
  61185=>"110110111",
  61186=>"100111101",
  61187=>"111000110",
  61188=>"000011000",
  61189=>"011010110",
  61190=>"110101011",
  61191=>"111011011",
  61192=>"111101111",
  61193=>"000010010",
  61194=>"010111000",
  61195=>"000100101",
  61196=>"000001101",
  61197=>"111111111",
  61198=>"101000010",
  61199=>"111111011",
  61200=>"001100110",
  61201=>"010000100",
  61202=>"110011011",
  61203=>"111000110",
  61204=>"010111100",
  61205=>"110011111",
  61206=>"110011111",
  61207=>"110001011",
  61208=>"111111111",
  61209=>"000010001",
  61210=>"111000001",
  61211=>"011000101",
  61212=>"100001000",
  61213=>"111011101",
  61214=>"001100000",
  61215=>"001001000",
  61216=>"001111110",
  61217=>"110011100",
  61218=>"110000111",
  61219=>"001100111",
  61220=>"101111010",
  61221=>"000101000",
  61222=>"011101110",
  61223=>"000011000",
  61224=>"100100010",
  61225=>"111010111",
  61226=>"001101010",
  61227=>"001001010",
  61228=>"101001101",
  61229=>"101000000",
  61230=>"011001001",
  61231=>"111011110",
  61232=>"000000000",
  61233=>"111011101",
  61234=>"100100001",
  61235=>"001010111",
  61236=>"101010111",
  61237=>"010100110",
  61238=>"100100100",
  61239=>"010110111",
  61240=>"000001000",
  61241=>"001111011",
  61242=>"110101000",
  61243=>"001100011",
  61244=>"001101001",
  61245=>"000001000",
  61246=>"101001000",
  61247=>"010100101",
  61248=>"000001100",
  61249=>"111100001",
  61250=>"110110010",
  61251=>"101111110",
  61252=>"111000100",
  61253=>"111100100",
  61254=>"001000010",
  61255=>"000001101",
  61256=>"111011101",
  61257=>"001101000",
  61258=>"010110101",
  61259=>"001001000",
  61260=>"101111110",
  61261=>"100010001",
  61262=>"110000000",
  61263=>"001101010",
  61264=>"000110100",
  61265=>"100100111",
  61266=>"001011101",
  61267=>"011110101",
  61268=>"000011110",
  61269=>"011010011",
  61270=>"111100110",
  61271=>"110110010",
  61272=>"110101001",
  61273=>"110000110",
  61274=>"110111010",
  61275=>"110110100",
  61276=>"110000110",
  61277=>"100000101",
  61278=>"011111111",
  61279=>"001000100",
  61280=>"011010111",
  61281=>"100111001",
  61282=>"101110010",
  61283=>"011110000",
  61284=>"111100100",
  61285=>"100001110",
  61286=>"101011100",
  61287=>"001000001",
  61288=>"101110010",
  61289=>"000000011",
  61290=>"111010101",
  61291=>"111001000",
  61292=>"100111110",
  61293=>"101100001",
  61294=>"011000111",
  61295=>"001101101",
  61296=>"110111011",
  61297=>"111101100",
  61298=>"110000111",
  61299=>"110000101",
  61300=>"001100101",
  61301=>"011111000",
  61302=>"000011000",
  61303=>"000001101",
  61304=>"100110011",
  61305=>"010000100",
  61306=>"110101001",
  61307=>"110110000",
  61308=>"111101011",
  61309=>"001111011",
  61310=>"111011001",
  61311=>"111100101",
  61312=>"010100010",
  61313=>"010110110",
  61314=>"001101011",
  61315=>"111000010",
  61316=>"100001000",
  61317=>"000010010",
  61318=>"011011111",
  61319=>"001001001",
  61320=>"110110000",
  61321=>"000110111",
  61322=>"100000010",
  61323=>"111110110",
  61324=>"001110101",
  61325=>"101000111",
  61326=>"010000010",
  61327=>"100100111",
  61328=>"010011100",
  61329=>"101111011",
  61330=>"000111100",
  61331=>"010011010",
  61332=>"100101110",
  61333=>"100000101",
  61334=>"011101101",
  61335=>"110001100",
  61336=>"001100011",
  61337=>"011001001",
  61338=>"001110101",
  61339=>"101110101",
  61340=>"101010001",
  61341=>"011111101",
  61342=>"110010001",
  61343=>"100111000",
  61344=>"010111110",
  61345=>"110000101",
  61346=>"100110100",
  61347=>"001010111",
  61348=>"000010000",
  61349=>"111011000",
  61350=>"010011000",
  61351=>"110000010",
  61352=>"011101000",
  61353=>"011111101",
  61354=>"111011001",
  61355=>"101011001",
  61356=>"110101011",
  61357=>"111001010",
  61358=>"111001010",
  61359=>"000010000",
  61360=>"011110111",
  61361=>"010110100",
  61362=>"011011011",
  61363=>"010111111",
  61364=>"100110011",
  61365=>"101111100",
  61366=>"111110110",
  61367=>"110010110",
  61368=>"111011000",
  61369=>"110010000",
  61370=>"011111110",
  61371=>"000010111",
  61372=>"000010001",
  61373=>"000010110",
  61374=>"011110101",
  61375=>"101111101",
  61376=>"101001111",
  61377=>"010000000",
  61378=>"000100111",
  61379=>"000100101",
  61380=>"101001010",
  61381=>"001011101",
  61382=>"011100001",
  61383=>"110010001",
  61384=>"101001011",
  61385=>"000111111",
  61386=>"011101111",
  61387=>"101101101",
  61388=>"000001010",
  61389=>"111101001",
  61390=>"011011101",
  61391=>"111000001",
  61392=>"010111000",
  61393=>"100110011",
  61394=>"111010110",
  61395=>"010010001",
  61396=>"101111000",
  61397=>"010000100",
  61398=>"101000100",
  61399=>"010100111",
  61400=>"111101000",
  61401=>"010010011",
  61402=>"101101100",
  61403=>"001011101",
  61404=>"111111110",
  61405=>"001100100",
  61406=>"111110101",
  61407=>"010001001",
  61408=>"100000100",
  61409=>"001100110",
  61410=>"111110011",
  61411=>"110010110",
  61412=>"000110000",
  61413=>"111001101",
  61414=>"001001000",
  61415=>"001000010",
  61416=>"101100011",
  61417=>"100011111",
  61418=>"000000011",
  61419=>"111100001",
  61420=>"100100101",
  61421=>"001011100",
  61422=>"111101111",
  61423=>"100010000",
  61424=>"101111011",
  61425=>"101100010",
  61426=>"010011010",
  61427=>"000101010",
  61428=>"111110100",
  61429=>"110001000",
  61430=>"100011101",
  61431=>"010000001",
  61432=>"110110010",
  61433=>"100100100",
  61434=>"110000110",
  61435=>"100110111",
  61436=>"100101001",
  61437=>"100110110",
  61438=>"111111001",
  61439=>"001110110",
  61440=>"111001011",
  61441=>"000100100",
  61442=>"010111110",
  61443=>"100011110",
  61444=>"001011001",
  61445=>"010001101",
  61446=>"010110111",
  61447=>"000101100",
  61448=>"000000001",
  61449=>"000111001",
  61450=>"011000001",
  61451=>"100111111",
  61452=>"001011010",
  61453=>"110000011",
  61454=>"010011111",
  61455=>"000001100",
  61456=>"000101110",
  61457=>"100000111",
  61458=>"010101100",
  61459=>"000111000",
  61460=>"000000111",
  61461=>"101110000",
  61462=>"101010111",
  61463=>"010000100",
  61464=>"011110110",
  61465=>"111110011",
  61466=>"100010101",
  61467=>"101001000",
  61468=>"011001100",
  61469=>"100111001",
  61470=>"000000011",
  61471=>"101110100",
  61472=>"010110010",
  61473=>"000111111",
  61474=>"000111010",
  61475=>"111111110",
  61476=>"101101100",
  61477=>"110010100",
  61478=>"011010110",
  61479=>"000000011",
  61480=>"111011101",
  61481=>"110010111",
  61482=>"001101110",
  61483=>"010000111",
  61484=>"101101111",
  61485=>"110111110",
  61486=>"001000110",
  61487=>"111010111",
  61488=>"010001101",
  61489=>"110111101",
  61490=>"111100111",
  61491=>"001110101",
  61492=>"001001000",
  61493=>"100101000",
  61494=>"011110010",
  61495=>"000000001",
  61496=>"101000000",
  61497=>"010110010",
  61498=>"101110001",
  61499=>"111110010",
  61500=>"111000110",
  61501=>"001110110",
  61502=>"010101000",
  61503=>"111100011",
  61504=>"111111101",
  61505=>"110110111",
  61506=>"011001100",
  61507=>"110101010",
  61508=>"000110011",
  61509=>"000001010",
  61510=>"001100110",
  61511=>"000100000",
  61512=>"000000011",
  61513=>"110100010",
  61514=>"000110000",
  61515=>"110111001",
  61516=>"101110100",
  61517=>"001110010",
  61518=>"111100000",
  61519=>"000111000",
  61520=>"100111110",
  61521=>"010111010",
  61522=>"100100000",
  61523=>"100100100",
  61524=>"000100010",
  61525=>"100010011",
  61526=>"111100000",
  61527=>"101111010",
  61528=>"111110111",
  61529=>"001100111",
  61530=>"000100000",
  61531=>"111101100",
  61532=>"011010100",
  61533=>"000001011",
  61534=>"101001100",
  61535=>"110101101",
  61536=>"110000000",
  61537=>"110000000",
  61538=>"000000010",
  61539=>"000110111",
  61540=>"111000011",
  61541=>"100101001",
  61542=>"111000101",
  61543=>"010111000",
  61544=>"110100001",
  61545=>"110101010",
  61546=>"000000000",
  61547=>"010111110",
  61548=>"010000000",
  61549=>"001110110",
  61550=>"011001110",
  61551=>"110101000",
  61552=>"000000110",
  61553=>"111001101",
  61554=>"110011000",
  61555=>"000010110",
  61556=>"100111011",
  61557=>"110100011",
  61558=>"111010101",
  61559=>"100110100",
  61560=>"111111001",
  61561=>"000101111",
  61562=>"101110011",
  61563=>"110111111",
  61564=>"010101001",
  61565=>"011111101",
  61566=>"110110110",
  61567=>"101101100",
  61568=>"100000101",
  61569=>"111000101",
  61570=>"010011001",
  61571=>"100111001",
  61572=>"111000110",
  61573=>"110000100",
  61574=>"001001100",
  61575=>"100110101",
  61576=>"001001111",
  61577=>"111000001",
  61578=>"011110110",
  61579=>"000001010",
  61580=>"101000001",
  61581=>"110001011",
  61582=>"110100001",
  61583=>"100110101",
  61584=>"011101110",
  61585=>"111101101",
  61586=>"101110010",
  61587=>"110010011",
  61588=>"011001100",
  61589=>"100010000",
  61590=>"110101111",
  61591=>"111010010",
  61592=>"110001010",
  61593=>"000101101",
  61594=>"010010101",
  61595=>"101100001",
  61596=>"010100111",
  61597=>"111001001",
  61598=>"011110011",
  61599=>"100011110",
  61600=>"100100110",
  61601=>"111010010",
  61602=>"111000111",
  61603=>"110110000",
  61604=>"010011011",
  61605=>"100111110",
  61606=>"101001100",
  61607=>"001001010",
  61608=>"101010000",
  61609=>"011111000",
  61610=>"100000111",
  61611=>"111101100",
  61612=>"101101110",
  61613=>"101101110",
  61614=>"011101111",
  61615=>"101100101",
  61616=>"010101111",
  61617=>"010011001",
  61618=>"101111110",
  61619=>"000001000",
  61620=>"010011000",
  61621=>"000000110",
  61622=>"101100101",
  61623=>"011000100",
  61624=>"010101101",
  61625=>"100011100",
  61626=>"000110100",
  61627=>"101111001",
  61628=>"010010111",
  61629=>"110110000",
  61630=>"001100001",
  61631=>"000010000",
  61632=>"011101000",
  61633=>"010110011",
  61634=>"101101111",
  61635=>"011001000",
  61636=>"101000000",
  61637=>"011101010",
  61638=>"110001000",
  61639=>"100110111",
  61640=>"101000101",
  61641=>"111001001",
  61642=>"001000100",
  61643=>"110010011",
  61644=>"001000100",
  61645=>"001010010",
  61646=>"000000011",
  61647=>"001000100",
  61648=>"011111011",
  61649=>"001111000",
  61650=>"011000100",
  61651=>"000001000",
  61652=>"101010010",
  61653=>"010001010",
  61654=>"000101000",
  61655=>"100101010",
  61656=>"110100100",
  61657=>"101110011",
  61658=>"101111010",
  61659=>"101001011",
  61660=>"111100000",
  61661=>"101000011",
  61662=>"001010100",
  61663=>"001100111",
  61664=>"001000100",
  61665=>"100000010",
  61666=>"100110111",
  61667=>"111011011",
  61668=>"000111100",
  61669=>"111100101",
  61670=>"010110000",
  61671=>"001011001",
  61672=>"110110100",
  61673=>"101010110",
  61674=>"100000100",
  61675=>"110101001",
  61676=>"000111000",
  61677=>"100110001",
  61678=>"110111100",
  61679=>"101101101",
  61680=>"001011111",
  61681=>"011100000",
  61682=>"010100111",
  61683=>"001010100",
  61684=>"111011010",
  61685=>"101101110",
  61686=>"000111110",
  61687=>"100000010",
  61688=>"111011100",
  61689=>"100011011",
  61690=>"101100000",
  61691=>"001001000",
  61692=>"001111100",
  61693=>"001111010",
  61694=>"010100101",
  61695=>"011111011",
  61696=>"100010110",
  61697=>"101111111",
  61698=>"000111111",
  61699=>"100101100",
  61700=>"111101100",
  61701=>"011100110",
  61702=>"110100111",
  61703=>"001010010",
  61704=>"000111100",
  61705=>"001000111",
  61706=>"110110100",
  61707=>"011100101",
  61708=>"100100000",
  61709=>"000011101",
  61710=>"000000010",
  61711=>"010100011",
  61712=>"100000110",
  61713=>"011011000",
  61714=>"000011111",
  61715=>"110000001",
  61716=>"110000100",
  61717=>"000111100",
  61718=>"011100010",
  61719=>"011110011",
  61720=>"101110011",
  61721=>"101001000",
  61722=>"001101000",
  61723=>"111100100",
  61724=>"100100111",
  61725=>"110100001",
  61726=>"000000001",
  61727=>"111100001",
  61728=>"001011011",
  61729=>"000011100",
  61730=>"110001000",
  61731=>"111100001",
  61732=>"111101100",
  61733=>"111110100",
  61734=>"101001111",
  61735=>"000101111",
  61736=>"010111001",
  61737=>"111010100",
  61738=>"000000100",
  61739=>"010001010",
  61740=>"011101101",
  61741=>"101001000",
  61742=>"000011010",
  61743=>"001111000",
  61744=>"001010010",
  61745=>"011001001",
  61746=>"111111000",
  61747=>"010010000",
  61748=>"100110110",
  61749=>"011000111",
  61750=>"000001101",
  61751=>"011100001",
  61752=>"010000001",
  61753=>"010110101",
  61754=>"111000001",
  61755=>"100001011",
  61756=>"110011011",
  61757=>"111100111",
  61758=>"001011010",
  61759=>"010011011",
  61760=>"101000011",
  61761=>"111111000",
  61762=>"001011010",
  61763=>"010011101",
  61764=>"001111100",
  61765=>"010011001",
  61766=>"110010011",
  61767=>"010010010",
  61768=>"100101000",
  61769=>"011100011",
  61770=>"001000000",
  61771=>"111001101",
  61772=>"100001100",
  61773=>"101111000",
  61774=>"100110110",
  61775=>"010100011",
  61776=>"000101000",
  61777=>"001100000",
  61778=>"011000011",
  61779=>"100101001",
  61780=>"101010001",
  61781=>"010010110",
  61782=>"000100111",
  61783=>"011010000",
  61784=>"001110000",
  61785=>"010100110",
  61786=>"100100110",
  61787=>"000000001",
  61788=>"001111101",
  61789=>"100000111",
  61790=>"110110011",
  61791=>"011100000",
  61792=>"011001011",
  61793=>"101010001",
  61794=>"000000101",
  61795=>"010001100",
  61796=>"110000101",
  61797=>"110000101",
  61798=>"001001011",
  61799=>"100011000",
  61800=>"011010010",
  61801=>"110010000",
  61802=>"100100100",
  61803=>"000010101",
  61804=>"101010010",
  61805=>"100011001",
  61806=>"100100001",
  61807=>"010110110",
  61808=>"100100001",
  61809=>"110100000",
  61810=>"010011011",
  61811=>"111110110",
  61812=>"111111111",
  61813=>"010011010",
  61814=>"001011100",
  61815=>"001011000",
  61816=>"011100110",
  61817=>"011001001",
  61818=>"000000011",
  61819=>"011101010",
  61820=>"101110100",
  61821=>"111011001",
  61822=>"010110100",
  61823=>"110001110",
  61824=>"111111001",
  61825=>"101000101",
  61826=>"100001000",
  61827=>"100000110",
  61828=>"010111000",
  61829=>"010011101",
  61830=>"000100100",
  61831=>"000000101",
  61832=>"000100100",
  61833=>"101110101",
  61834=>"010100011",
  61835=>"000111101",
  61836=>"111001010",
  61837=>"101011001",
  61838=>"010011010",
  61839=>"111100010",
  61840=>"111011101",
  61841=>"000000100",
  61842=>"000101101",
  61843=>"100010001",
  61844=>"111010001",
  61845=>"111111101",
  61846=>"001000001",
  61847=>"000001000",
  61848=>"111011001",
  61849=>"110100000",
  61850=>"010101111",
  61851=>"110011100",
  61852=>"011010000",
  61853=>"010000110",
  61854=>"111001100",
  61855=>"101010111",
  61856=>"011100011",
  61857=>"011100101",
  61858=>"111110011",
  61859=>"000100101",
  61860=>"001010001",
  61861=>"001011100",
  61862=>"011111100",
  61863=>"001110010",
  61864=>"101111011",
  61865=>"010011000",
  61866=>"001100101",
  61867=>"111111000",
  61868=>"010011001",
  61869=>"111010111",
  61870=>"001001100",
  61871=>"111010110",
  61872=>"101010010",
  61873=>"111010000",
  61874=>"110010001",
  61875=>"101111011",
  61876=>"111010110",
  61877=>"000100000",
  61878=>"010001101",
  61879=>"110000101",
  61880=>"001011001",
  61881=>"100110010",
  61882=>"110010010",
  61883=>"101001011",
  61884=>"101101001",
  61885=>"001100111",
  61886=>"101001110",
  61887=>"110010101",
  61888=>"111011100",
  61889=>"111110001",
  61890=>"100000001",
  61891=>"100000111",
  61892=>"111001111",
  61893=>"010110000",
  61894=>"011000000",
  61895=>"001011000",
  61896=>"011011011",
  61897=>"111000101",
  61898=>"010000010",
  61899=>"001000000",
  61900=>"110100100",
  61901=>"101100100",
  61902=>"010110011",
  61903=>"101010010",
  61904=>"001101111",
  61905=>"110001111",
  61906=>"111111010",
  61907=>"100000010",
  61908=>"110101011",
  61909=>"101001110",
  61910=>"000101001",
  61911=>"011100100",
  61912=>"100101010",
  61913=>"101000010",
  61914=>"101100001",
  61915=>"110110000",
  61916=>"110101101",
  61917=>"111001100",
  61918=>"000010011",
  61919=>"000101011",
  61920=>"000011010",
  61921=>"010011111",
  61922=>"111001001",
  61923=>"001110011",
  61924=>"111100011",
  61925=>"000110000",
  61926=>"010111110",
  61927=>"111111000",
  61928=>"111010110",
  61929=>"101001101",
  61930=>"000000001",
  61931=>"010010001",
  61932=>"001011100",
  61933=>"010110000",
  61934=>"011111001",
  61935=>"011011101",
  61936=>"100011101",
  61937=>"111010010",
  61938=>"101100010",
  61939=>"010011010",
  61940=>"000100001",
  61941=>"011001000",
  61942=>"011110101",
  61943=>"100100001",
  61944=>"010011100",
  61945=>"101100010",
  61946=>"110001111",
  61947=>"010011111",
  61948=>"011101010",
  61949=>"000001111",
  61950=>"011011010",
  61951=>"000101000",
  61952=>"000111101",
  61953=>"100001010",
  61954=>"101111000",
  61955=>"010001010",
  61956=>"111001010",
  61957=>"110000001",
  61958=>"101001110",
  61959=>"011000011",
  61960=>"000100100",
  61961=>"101100000",
  61962=>"011001010",
  61963=>"101011101",
  61964=>"000001111",
  61965=>"100000010",
  61966=>"010000001",
  61967=>"010000010",
  61968=>"111001111",
  61969=>"110010011",
  61970=>"001001000",
  61971=>"111110000",
  61972=>"011110011",
  61973=>"011001011",
  61974=>"110010101",
  61975=>"011101110",
  61976=>"101001010",
  61977=>"111111110",
  61978=>"110000010",
  61979=>"100110101",
  61980=>"110101010",
  61981=>"110011100",
  61982=>"101111111",
  61983=>"000111101",
  61984=>"101100001",
  61985=>"111110101",
  61986=>"000000111",
  61987=>"111100001",
  61988=>"100101100",
  61989=>"111001110",
  61990=>"011101111",
  61991=>"001110100",
  61992=>"110000111",
  61993=>"110110110",
  61994=>"010010010",
  61995=>"011010011",
  61996=>"011100000",
  61997=>"001110110",
  61998=>"010001111",
  61999=>"011000001",
  62000=>"001010000",
  62001=>"101111010",
  62002=>"011101000",
  62003=>"100011111",
  62004=>"000010010",
  62005=>"010011011",
  62006=>"110001001",
  62007=>"000100000",
  62008=>"111111111",
  62009=>"100001100",
  62010=>"010101010",
  62011=>"111110000",
  62012=>"010110110",
  62013=>"111110010",
  62014=>"000010101",
  62015=>"111011010",
  62016=>"000001100",
  62017=>"100110110",
  62018=>"100000000",
  62019=>"100011010",
  62020=>"100011100",
  62021=>"001010101",
  62022=>"100001111",
  62023=>"011011000",
  62024=>"010010000",
  62025=>"111011110",
  62026=>"111111010",
  62027=>"011110100",
  62028=>"110000000",
  62029=>"010111110",
  62030=>"010110010",
  62031=>"100101100",
  62032=>"111001010",
  62033=>"001110000",
  62034=>"010000000",
  62035=>"011110000",
  62036=>"010001000",
  62037=>"101000001",
  62038=>"110001001",
  62039=>"001000011",
  62040=>"101011101",
  62041=>"010110001",
  62042=>"001110011",
  62043=>"000100000",
  62044=>"111101000",
  62045=>"101101111",
  62046=>"011011101",
  62047=>"001101100",
  62048=>"000000001",
  62049=>"011110001",
  62050=>"001110110",
  62051=>"100101001",
  62052=>"110010111",
  62053=>"101000001",
  62054=>"000110110",
  62055=>"001010110",
  62056=>"111101110",
  62057=>"110000110",
  62058=>"111010111",
  62059=>"101000110",
  62060=>"100100111",
  62061=>"000010110",
  62062=>"100101001",
  62063=>"101110111",
  62064=>"100010011",
  62065=>"111011010",
  62066=>"110100010",
  62067=>"110010011",
  62068=>"101111010",
  62069=>"001001010",
  62070=>"100001111",
  62071=>"100111011",
  62072=>"001001111",
  62073=>"001100001",
  62074=>"000110010",
  62075=>"011100001",
  62076=>"000010010",
  62077=>"011111111",
  62078=>"111010100",
  62079=>"100010010",
  62080=>"101011100",
  62081=>"111011110",
  62082=>"000110100",
  62083=>"110001101",
  62084=>"100110010",
  62085=>"111110000",
  62086=>"000001111",
  62087=>"000000011",
  62088=>"101101000",
  62089=>"100110001",
  62090=>"111100000",
  62091=>"111110000",
  62092=>"110001001",
  62093=>"110001010",
  62094=>"010101010",
  62095=>"111110011",
  62096=>"110101110",
  62097=>"100111101",
  62098=>"011111010",
  62099=>"111110101",
  62100=>"100011000",
  62101=>"001111111",
  62102=>"010111001",
  62103=>"000000000",
  62104=>"101001001",
  62105=>"100100111",
  62106=>"110010010",
  62107=>"110111000",
  62108=>"001001010",
  62109=>"000000011",
  62110=>"011111000",
  62111=>"100011111",
  62112=>"100001011",
  62113=>"110000110",
  62114=>"110011111",
  62115=>"010101010",
  62116=>"111101001",
  62117=>"111110000",
  62118=>"000110011",
  62119=>"010010100",
  62120=>"101110010",
  62121=>"000100001",
  62122=>"000000011",
  62123=>"110000100",
  62124=>"010110111",
  62125=>"101110011",
  62126=>"001110011",
  62127=>"111010000",
  62128=>"101000001",
  62129=>"000000100",
  62130=>"010001100",
  62131=>"011001010",
  62132=>"010100011",
  62133=>"100011010",
  62134=>"100010001",
  62135=>"010010110",
  62136=>"101100001",
  62137=>"000001101",
  62138=>"101100110",
  62139=>"100011011",
  62140=>"011010000",
  62141=>"010011100",
  62142=>"001101001",
  62143=>"100110110",
  62144=>"101111011",
  62145=>"111010110",
  62146=>"111010111",
  62147=>"011111000",
  62148=>"001101101",
  62149=>"110110110",
  62150=>"110010100",
  62151=>"110100110",
  62152=>"001110011",
  62153=>"011000100",
  62154=>"111111111",
  62155=>"001011111",
  62156=>"011010100",
  62157=>"001010000",
  62158=>"001000111",
  62159=>"000011111",
  62160=>"110001010",
  62161=>"101101000",
  62162=>"111000101",
  62163=>"011011001",
  62164=>"100000101",
  62165=>"110100100",
  62166=>"110100110",
  62167=>"001010101",
  62168=>"001010010",
  62169=>"001011110",
  62170=>"001001011",
  62171=>"001001001",
  62172=>"110001000",
  62173=>"100010101",
  62174=>"100010000",
  62175=>"000111001",
  62176=>"101100101",
  62177=>"101011011",
  62178=>"111001001",
  62179=>"101001011",
  62180=>"000110100",
  62181=>"011100100",
  62182=>"111001110",
  62183=>"111101111",
  62184=>"001000011",
  62185=>"001100011",
  62186=>"010100010",
  62187=>"110100110",
  62188=>"011101001",
  62189=>"111110100",
  62190=>"100100010",
  62191=>"000001000",
  62192=>"010101011",
  62193=>"011101001",
  62194=>"111010000",
  62195=>"010001100",
  62196=>"100001010",
  62197=>"100111111",
  62198=>"000000110",
  62199=>"000011101",
  62200=>"001010101",
  62201=>"101101001",
  62202=>"010101110",
  62203=>"111110101",
  62204=>"100000011",
  62205=>"100110000",
  62206=>"100000110",
  62207=>"100011111",
  62208=>"011001001",
  62209=>"001000000",
  62210=>"100011000",
  62211=>"010101000",
  62212=>"011000000",
  62213=>"011111010",
  62214=>"001111101",
  62215=>"010101000",
  62216=>"101110011",
  62217=>"111101110",
  62218=>"010101000",
  62219=>"110101010",
  62220=>"110000100",
  62221=>"101001101",
  62222=>"101100000",
  62223=>"111001000",
  62224=>"001111101",
  62225=>"111000000",
  62226=>"000011001",
  62227=>"010011100",
  62228=>"010011110",
  62229=>"010000010",
  62230=>"011110000",
  62231=>"111100100",
  62232=>"100110010",
  62233=>"101001111",
  62234=>"111101010",
  62235=>"110011110",
  62236=>"111001001",
  62237=>"111011011",
  62238=>"001001110",
  62239=>"101010111",
  62240=>"111111101",
  62241=>"010110101",
  62242=>"110100000",
  62243=>"101001010",
  62244=>"001110100",
  62245=>"101010100",
  62246=>"011010000",
  62247=>"000111000",
  62248=>"111110101",
  62249=>"100000111",
  62250=>"101000101",
  62251=>"001110010",
  62252=>"100100101",
  62253=>"100101000",
  62254=>"010010100",
  62255=>"000001001",
  62256=>"110110000",
  62257=>"100110110",
  62258=>"001001110",
  62259=>"000000011",
  62260=>"110110100",
  62261=>"101100101",
  62262=>"010101111",
  62263=>"010000011",
  62264=>"010011000",
  62265=>"000101010",
  62266=>"001100011",
  62267=>"100111001",
  62268=>"110110110",
  62269=>"100101101",
  62270=>"000100001",
  62271=>"000100111",
  62272=>"110001001",
  62273=>"111010001",
  62274=>"111110100",
  62275=>"011010111",
  62276=>"010011111",
  62277=>"000100101",
  62278=>"100100111",
  62279=>"010000001",
  62280=>"000100001",
  62281=>"111011000",
  62282=>"011000100",
  62283=>"111011010",
  62284=>"111001000",
  62285=>"100010110",
  62286=>"001110010",
  62287=>"001100011",
  62288=>"101001100",
  62289=>"100010000",
  62290=>"111001011",
  62291=>"101010100",
  62292=>"111011001",
  62293=>"001001011",
  62294=>"110110110",
  62295=>"101110001",
  62296=>"000110101",
  62297=>"011010110",
  62298=>"101111011",
  62299=>"110110000",
  62300=>"000010111",
  62301=>"011001111",
  62302=>"111101100",
  62303=>"010001101",
  62304=>"101100000",
  62305=>"000100010",
  62306=>"011011101",
  62307=>"010010000",
  62308=>"011110010",
  62309=>"010110100",
  62310=>"010000111",
  62311=>"110011011",
  62312=>"010100010",
  62313=>"010011101",
  62314=>"100001000",
  62315=>"100101100",
  62316=>"101011010",
  62317=>"100011001",
  62318=>"100010000",
  62319=>"001001000",
  62320=>"101010110",
  62321=>"101011001",
  62322=>"111011101",
  62323=>"101111101",
  62324=>"010001111",
  62325=>"011010000",
  62326=>"110110000",
  62327=>"001000111",
  62328=>"100001010",
  62329=>"100110011",
  62330=>"100001110",
  62331=>"000010101",
  62332=>"001011101",
  62333=>"000100001",
  62334=>"001100010",
  62335=>"010010100",
  62336=>"001111110",
  62337=>"010100100",
  62338=>"100111011",
  62339=>"000000111",
  62340=>"110110011",
  62341=>"100001000",
  62342=>"000011000",
  62343=>"111111010",
  62344=>"010011011",
  62345=>"101010001",
  62346=>"000011000",
  62347=>"101011010",
  62348=>"010110111",
  62349=>"100101001",
  62350=>"110000011",
  62351=>"011001110",
  62352=>"010110100",
  62353=>"011011011",
  62354=>"010010000",
  62355=>"100000011",
  62356=>"010111100",
  62357=>"011011101",
  62358=>"100000101",
  62359=>"100111011",
  62360=>"111000000",
  62361=>"111111110",
  62362=>"000001111",
  62363=>"111110101",
  62364=>"101001110",
  62365=>"110111001",
  62366=>"001101001",
  62367=>"111001010",
  62368=>"100010001",
  62369=>"100111000",
  62370=>"100011000",
  62371=>"011100101",
  62372=>"111110111",
  62373=>"100110100",
  62374=>"001100111",
  62375=>"101011001",
  62376=>"011001011",
  62377=>"001010000",
  62378=>"011111111",
  62379=>"011001010",
  62380=>"100100100",
  62381=>"001111010",
  62382=>"100010110",
  62383=>"101100110",
  62384=>"001010010",
  62385=>"101011011",
  62386=>"011001001",
  62387=>"010000010",
  62388=>"100110010",
  62389=>"000100010",
  62390=>"101011101",
  62391=>"001111111",
  62392=>"111001011",
  62393=>"000110000",
  62394=>"100101011",
  62395=>"000100000",
  62396=>"011010110",
  62397=>"001001011",
  62398=>"001111000",
  62399=>"000010011",
  62400=>"001011111",
  62401=>"001001000",
  62402=>"100010001",
  62403=>"001010001",
  62404=>"100111100",
  62405=>"111101001",
  62406=>"111100011",
  62407=>"010010010",
  62408=>"001001100",
  62409=>"101010001",
  62410=>"000010011",
  62411=>"101001110",
  62412=>"110001110",
  62413=>"010101011",
  62414=>"000010101",
  62415=>"110111110",
  62416=>"000111010",
  62417=>"001111001",
  62418=>"010100011",
  62419=>"011001111",
  62420=>"011100110",
  62421=>"000010111",
  62422=>"100000110",
  62423=>"100110011",
  62424=>"101110101",
  62425=>"111001011",
  62426=>"111010001",
  62427=>"000011100",
  62428=>"100100001",
  62429=>"111110110",
  62430=>"110100010",
  62431=>"101100010",
  62432=>"001000001",
  62433=>"110010110",
  62434=>"110001011",
  62435=>"001011010",
  62436=>"001010000",
  62437=>"111110110",
  62438=>"110001111",
  62439=>"110000100",
  62440=>"110000101",
  62441=>"001011100",
  62442=>"110011011",
  62443=>"100001000",
  62444=>"111010101",
  62445=>"101011111",
  62446=>"000001000",
  62447=>"010101010",
  62448=>"001001111",
  62449=>"101001011",
  62450=>"010011100",
  62451=>"011111010",
  62452=>"011101100",
  62453=>"011011011",
  62454=>"010011111",
  62455=>"111010111",
  62456=>"100011011",
  62457=>"101000111",
  62458=>"111010111",
  62459=>"010101010",
  62460=>"110110001",
  62461=>"011100100",
  62462=>"101100101",
  62463=>"101101111",
  62464=>"011011111",
  62465=>"011001110",
  62466=>"011000110",
  62467=>"010001001",
  62468=>"010000000",
  62469=>"001000000",
  62470=>"000110010",
  62471=>"101101111",
  62472=>"011001010",
  62473=>"101001111",
  62474=>"101111001",
  62475=>"100001010",
  62476=>"100110011",
  62477=>"000101001",
  62478=>"011100010",
  62479=>"110000000",
  62480=>"110011111",
  62481=>"100001011",
  62482=>"010110001",
  62483=>"110100010",
  62484=>"001101011",
  62485=>"001011010",
  62486=>"101010111",
  62487=>"011111011",
  62488=>"010001101",
  62489=>"111011010",
  62490=>"101111100",
  62491=>"010010000",
  62492=>"101011100",
  62493=>"010000110",
  62494=>"000110000",
  62495=>"000100100",
  62496=>"100111110",
  62497=>"000001001",
  62498=>"101110010",
  62499=>"101111010",
  62500=>"011011110",
  62501=>"101000001",
  62502=>"101111101",
  62503=>"010111111",
  62504=>"111110000",
  62505=>"111111111",
  62506=>"011100010",
  62507=>"001101100",
  62508=>"000010100",
  62509=>"110011110",
  62510=>"010101010",
  62511=>"000000100",
  62512=>"101000001",
  62513=>"000110100",
  62514=>"110101100",
  62515=>"100010101",
  62516=>"011010100",
  62517=>"001011001",
  62518=>"111101010",
  62519=>"111000100",
  62520=>"001000111",
  62521=>"000111110",
  62522=>"000010100",
  62523=>"010110001",
  62524=>"111001111",
  62525=>"011011001",
  62526=>"111100010",
  62527=>"100111101",
  62528=>"011000100",
  62529=>"010010110",
  62530=>"010110001",
  62531=>"111101000",
  62532=>"000100101",
  62533=>"100000001",
  62534=>"010010000",
  62535=>"001000110",
  62536=>"111111010",
  62537=>"101010001",
  62538=>"001111111",
  62539=>"100001000",
  62540=>"000110010",
  62541=>"100011000",
  62542=>"101010010",
  62543=>"010001111",
  62544=>"100101001",
  62545=>"110010000",
  62546=>"000101100",
  62547=>"111010110",
  62548=>"010010000",
  62549=>"101111000",
  62550=>"111101000",
  62551=>"101000110",
  62552=>"010101001",
  62553=>"110101011",
  62554=>"101010011",
  62555=>"010000111",
  62556=>"110010001",
  62557=>"100001011",
  62558=>"010010111",
  62559=>"100101010",
  62560=>"101011001",
  62561=>"110001001",
  62562=>"001101011",
  62563=>"101001011",
  62564=>"110011111",
  62565=>"000111100",
  62566=>"111011110",
  62567=>"101011010",
  62568=>"100001000",
  62569=>"001010001",
  62570=>"011101101",
  62571=>"010100011",
  62572=>"110010100",
  62573=>"010111110",
  62574=>"001011100",
  62575=>"010011111",
  62576=>"101100100",
  62577=>"101011111",
  62578=>"111111110",
  62579=>"101010111",
  62580=>"010100001",
  62581=>"001111100",
  62582=>"110110001",
  62583=>"001110101",
  62584=>"000110001",
  62585=>"000111101",
  62586=>"001100001",
  62587=>"010111111",
  62588=>"000000101",
  62589=>"011011010",
  62590=>"000110110",
  62591=>"101011010",
  62592=>"000000000",
  62593=>"011010111",
  62594=>"100010111",
  62595=>"101010001",
  62596=>"000001010",
  62597=>"000000000",
  62598=>"100101100",
  62599=>"000011000",
  62600=>"011111111",
  62601=>"000110000",
  62602=>"101100001",
  62603=>"110110111",
  62604=>"100110110",
  62605=>"010100001",
  62606=>"000000110",
  62607=>"111000110",
  62608=>"011011101",
  62609=>"110100110",
  62610=>"010011101",
  62611=>"000000101",
  62612=>"110011001",
  62613=>"000100101",
  62614=>"100000101",
  62615=>"101110001",
  62616=>"101000100",
  62617=>"001101010",
  62618=>"000101101",
  62619=>"001101110",
  62620=>"111011110",
  62621=>"101100101",
  62622=>"000001001",
  62623=>"111011111",
  62624=>"010000001",
  62625=>"100010000",
  62626=>"001010110",
  62627=>"110010011",
  62628=>"000010011",
  62629=>"111011111",
  62630=>"001000101",
  62631=>"101011000",
  62632=>"010001000",
  62633=>"000001111",
  62634=>"001100010",
  62635=>"101100000",
  62636=>"111010010",
  62637=>"011110111",
  62638=>"001100000",
  62639=>"010110111",
  62640=>"101001000",
  62641=>"011001110",
  62642=>"111100001",
  62643=>"011011000",
  62644=>"100100110",
  62645=>"001101010",
  62646=>"100100010",
  62647=>"000010111",
  62648=>"000100000",
  62649=>"000100111",
  62650=>"101001001",
  62651=>"111001000",
  62652=>"010101111",
  62653=>"001001101",
  62654=>"000111110",
  62655=>"101001101",
  62656=>"000000101",
  62657=>"101110100",
  62658=>"101111100",
  62659=>"111111000",
  62660=>"101010011",
  62661=>"111111001",
  62662=>"010001001",
  62663=>"001101001",
  62664=>"000110011",
  62665=>"111111001",
  62666=>"001100010",
  62667=>"001100101",
  62668=>"011010110",
  62669=>"111110011",
  62670=>"001101000",
  62671=>"000011001",
  62672=>"101010100",
  62673=>"111001010",
  62674=>"000000111",
  62675=>"010011111",
  62676=>"000101110",
  62677=>"001100001",
  62678=>"110001111",
  62679=>"010011000",
  62680=>"110100100",
  62681=>"101001011",
  62682=>"011010101",
  62683=>"000000110",
  62684=>"110011111",
  62685=>"000000010",
  62686=>"000000000",
  62687=>"110111110",
  62688=>"010000111",
  62689=>"010111100",
  62690=>"000010010",
  62691=>"000001010",
  62692=>"001001110",
  62693=>"111111011",
  62694=>"000011111",
  62695=>"110111101",
  62696=>"001110001",
  62697=>"101110000",
  62698=>"111010100",
  62699=>"001001110",
  62700=>"010010011",
  62701=>"010001011",
  62702=>"001100111",
  62703=>"110110100",
  62704=>"001010000",
  62705=>"000111100",
  62706=>"101010000",
  62707=>"100100000",
  62708=>"010111110",
  62709=>"101101001",
  62710=>"111000000",
  62711=>"101000100",
  62712=>"000110010",
  62713=>"001110111",
  62714=>"101000001",
  62715=>"011110010",
  62716=>"001101000",
  62717=>"110111110",
  62718=>"110010110",
  62719=>"111111010",
  62720=>"001100010",
  62721=>"011001100",
  62722=>"111100100",
  62723=>"111111011",
  62724=>"101110110",
  62725=>"000101100",
  62726=>"111101001",
  62727=>"000110001",
  62728=>"101110111",
  62729=>"011101100",
  62730=>"110010111",
  62731=>"000000100",
  62732=>"000111101",
  62733=>"100100111",
  62734=>"100100010",
  62735=>"111111011",
  62736=>"111101111",
  62737=>"011111010",
  62738=>"111100000",
  62739=>"011100010",
  62740=>"110111110",
  62741=>"111111100",
  62742=>"110111111",
  62743=>"110000111",
  62744=>"100010101",
  62745=>"000011111",
  62746=>"100100010",
  62747=>"000000000",
  62748=>"000010000",
  62749=>"011110101",
  62750=>"100010010",
  62751=>"101001000",
  62752=>"110110111",
  62753=>"110010010",
  62754=>"000101001",
  62755=>"010001010",
  62756=>"000001110",
  62757=>"010110100",
  62758=>"011111011",
  62759=>"101010100",
  62760=>"011110100",
  62761=>"011100000",
  62762=>"100011101",
  62763=>"110011011",
  62764=>"100100111",
  62765=>"011011111",
  62766=>"100001011",
  62767=>"010000001",
  62768=>"010111100",
  62769=>"011000011",
  62770=>"100100100",
  62771=>"111001110",
  62772=>"000110001",
  62773=>"000101010",
  62774=>"000100010",
  62775=>"010101000",
  62776=>"111101000",
  62777=>"111111000",
  62778=>"011010011",
  62779=>"111111111",
  62780=>"110111010",
  62781=>"011010100",
  62782=>"011011110",
  62783=>"110110101",
  62784=>"010110001",
  62785=>"100111110",
  62786=>"110100001",
  62787=>"110001111",
  62788=>"100110111",
  62789=>"111000100",
  62790=>"100110111",
  62791=>"010011000",
  62792=>"100111011",
  62793=>"001101110",
  62794=>"000111110",
  62795=>"000110000",
  62796=>"001000110",
  62797=>"111001110",
  62798=>"010010101",
  62799=>"001001000",
  62800=>"000011011",
  62801=>"001000110",
  62802=>"110100001",
  62803=>"111110111",
  62804=>"111011101",
  62805=>"011010100",
  62806=>"111110111",
  62807=>"100000010",
  62808=>"000010001",
  62809=>"000011100",
  62810=>"111101011",
  62811=>"000000110",
  62812=>"010001010",
  62813=>"100000100",
  62814=>"101010100",
  62815=>"101111111",
  62816=>"110101101",
  62817=>"000001010",
  62818=>"010110000",
  62819=>"000011011",
  62820=>"100111111",
  62821=>"011111100",
  62822=>"100101100",
  62823=>"001000011",
  62824=>"110101110",
  62825=>"001110110",
  62826=>"000101111",
  62827=>"001101111",
  62828=>"101110101",
  62829=>"000111011",
  62830=>"000100101",
  62831=>"001010111",
  62832=>"111000111",
  62833=>"111000111",
  62834=>"010010100",
  62835=>"010101111",
  62836=>"001000111",
  62837=>"101010100",
  62838=>"000000100",
  62839=>"100101000",
  62840=>"010111001",
  62841=>"111010000",
  62842=>"001011001",
  62843=>"010111100",
  62844=>"011111110",
  62845=>"101011110",
  62846=>"001000011",
  62847=>"000110011",
  62848=>"101010111",
  62849=>"111111000",
  62850=>"100111101",
  62851=>"010011111",
  62852=>"111100100",
  62853=>"100101010",
  62854=>"010110011",
  62855=>"111111011",
  62856=>"001010111",
  62857=>"100111101",
  62858=>"011011100",
  62859=>"001010000",
  62860=>"110000011",
  62861=>"001000100",
  62862=>"101110101",
  62863=>"000011000",
  62864=>"111010101",
  62865=>"001111101",
  62866=>"111110110",
  62867=>"100011111",
  62868=>"111011111",
  62869=>"100101000",
  62870=>"101001001",
  62871=>"000101111",
  62872=>"111010001",
  62873=>"001011110",
  62874=>"100011100",
  62875=>"001101100",
  62876=>"111111101",
  62877=>"000111100",
  62878=>"010001010",
  62879=>"110110110",
  62880=>"010100010",
  62881=>"000110110",
  62882=>"110101000",
  62883=>"011101111",
  62884=>"000001110",
  62885=>"111001111",
  62886=>"000010110",
  62887=>"010010001",
  62888=>"111010100",
  62889=>"010001000",
  62890=>"000111011",
  62891=>"000001001",
  62892=>"010101000",
  62893=>"000011000",
  62894=>"011001001",
  62895=>"011111111",
  62896=>"000101000",
  62897=>"011100001",
  62898=>"000101101",
  62899=>"101110111",
  62900=>"000100100",
  62901=>"010111001",
  62902=>"010100001",
  62903=>"110000001",
  62904=>"010111011",
  62905=>"100110110",
  62906=>"001110001",
  62907=>"101110100",
  62908=>"111101001",
  62909=>"011110001",
  62910=>"001010110",
  62911=>"011010000",
  62912=>"001000101",
  62913=>"001111011",
  62914=>"111100111",
  62915=>"110001110",
  62916=>"111111001",
  62917=>"010010110",
  62918=>"110100111",
  62919=>"100101110",
  62920=>"111111011",
  62921=>"011010111",
  62922=>"000111111",
  62923=>"101100001",
  62924=>"001001110",
  62925=>"101110000",
  62926=>"101100010",
  62927=>"110000001",
  62928=>"100101110",
  62929=>"010010001",
  62930=>"010110010",
  62931=>"111000100",
  62932=>"100100101",
  62933=>"100110011",
  62934=>"000111100",
  62935=>"000011101",
  62936=>"111111111",
  62937=>"000110110",
  62938=>"011111101",
  62939=>"011001101",
  62940=>"010001000",
  62941=>"101001110",
  62942=>"110000011",
  62943=>"101111111",
  62944=>"100110101",
  62945=>"001111100",
  62946=>"011100001",
  62947=>"001101001",
  62948=>"011011101",
  62949=>"110101010",
  62950=>"000110011",
  62951=>"011100110",
  62952=>"000010000",
  62953=>"000011110",
  62954=>"001001010",
  62955=>"100001000",
  62956=>"110111000",
  62957=>"101011011",
  62958=>"001001100",
  62959=>"001011111",
  62960=>"101011100",
  62961=>"100100001",
  62962=>"111010001",
  62963=>"111111001",
  62964=>"000000001",
  62965=>"010010010",
  62966=>"000011100",
  62967=>"111110100",
  62968=>"011010000",
  62969=>"101110011",
  62970=>"111010101",
  62971=>"100110110",
  62972=>"111011000",
  62973=>"001000111",
  62974=>"111010010",
  62975=>"001001110",
  62976=>"101011010",
  62977=>"011011011",
  62978=>"000110000",
  62979=>"001010101",
  62980=>"100110111",
  62981=>"000001111",
  62982=>"101001001",
  62983=>"000110011",
  62984=>"001011111",
  62985=>"011111111",
  62986=>"110111110",
  62987=>"111100001",
  62988=>"111001111",
  62989=>"100100011",
  62990=>"111100101",
  62991=>"011001111",
  62992=>"001100010",
  62993=>"110011001",
  62994=>"100011011",
  62995=>"110011011",
  62996=>"010000111",
  62997=>"010001010",
  62998=>"110101100",
  62999=>"100001100",
  63000=>"011011101",
  63001=>"001011110",
  63002=>"000101111",
  63003=>"010111101",
  63004=>"011001101",
  63005=>"111100111",
  63006=>"100111011",
  63007=>"001011100",
  63008=>"101101101",
  63009=>"000001011",
  63010=>"000111111",
  63011=>"110110111",
  63012=>"101010110",
  63013=>"000101001",
  63014=>"010100000",
  63015=>"001011011",
  63016=>"000111010",
  63017=>"010101000",
  63018=>"001111100",
  63019=>"101000110",
  63020=>"011111110",
  63021=>"111110001",
  63022=>"001010000",
  63023=>"110001101",
  63024=>"110000100",
  63025=>"110011000",
  63026=>"010110111",
  63027=>"111101001",
  63028=>"101111111",
  63029=>"111001101",
  63030=>"000000011",
  63031=>"100111111",
  63032=>"001101100",
  63033=>"001011101",
  63034=>"101101011",
  63035=>"100000100",
  63036=>"110100000",
  63037=>"010111010",
  63038=>"111000101",
  63039=>"000100000",
  63040=>"011111001",
  63041=>"010011000",
  63042=>"011000101",
  63043=>"101011111",
  63044=>"001100011",
  63045=>"101011010",
  63046=>"000001111",
  63047=>"100011110",
  63048=>"001000111",
  63049=>"110101000",
  63050=>"100010010",
  63051=>"011100101",
  63052=>"100110010",
  63053=>"110110000",
  63054=>"001101111",
  63055=>"100100110",
  63056=>"110010011",
  63057=>"110101100",
  63058=>"111110100",
  63059=>"010111101",
  63060=>"110001000",
  63061=>"101111101",
  63062=>"101001011",
  63063=>"111101010",
  63064=>"010111010",
  63065=>"011111111",
  63066=>"101011011",
  63067=>"111011110",
  63068=>"011100110",
  63069=>"000100111",
  63070=>"110010111",
  63071=>"010010010",
  63072=>"000111010",
  63073=>"101000000",
  63074=>"001010000",
  63075=>"101110101",
  63076=>"100101101",
  63077=>"100000101",
  63078=>"110110001",
  63079=>"010001101",
  63080=>"010011111",
  63081=>"110100111",
  63082=>"000110001",
  63083=>"111101000",
  63084=>"000010000",
  63085=>"100101100",
  63086=>"101000000",
  63087=>"100011010",
  63088=>"001100010",
  63089=>"111001110",
  63090=>"010001011",
  63091=>"101011000",
  63092=>"011100000",
  63093=>"100001110",
  63094=>"000010111",
  63095=>"110101011",
  63096=>"110011010",
  63097=>"100000000",
  63098=>"110110100",
  63099=>"110101001",
  63100=>"101010110",
  63101=>"101001011",
  63102=>"010101011",
  63103=>"111010001",
  63104=>"010010011",
  63105=>"110101110",
  63106=>"000110111",
  63107=>"100011100",
  63108=>"000101010",
  63109=>"001001011",
  63110=>"010001011",
  63111=>"010111111",
  63112=>"110110000",
  63113=>"000011100",
  63114=>"010111101",
  63115=>"010100000",
  63116=>"000111111",
  63117=>"101001011",
  63118=>"011110011",
  63119=>"010000110",
  63120=>"110010111",
  63121=>"101000100",
  63122=>"000010001",
  63123=>"000110011",
  63124=>"110100011",
  63125=>"110011111",
  63126=>"111010111",
  63127=>"011101000",
  63128=>"101100010",
  63129=>"100000011",
  63130=>"010010011",
  63131=>"111011001",
  63132=>"111100110",
  63133=>"010101000",
  63134=>"111011010",
  63135=>"011001100",
  63136=>"100010010",
  63137=>"000011001",
  63138=>"010010011",
  63139=>"111000100",
  63140=>"011011100",
  63141=>"011011111",
  63142=>"101111100",
  63143=>"111100011",
  63144=>"100001001",
  63145=>"110000001",
  63146=>"100111011",
  63147=>"000101110",
  63148=>"100000001",
  63149=>"101110111",
  63150=>"101011101",
  63151=>"101111001",
  63152=>"110011100",
  63153=>"111101010",
  63154=>"101100001",
  63155=>"001111010",
  63156=>"010110100",
  63157=>"100001011",
  63158=>"111010001",
  63159=>"111110011",
  63160=>"010100111",
  63161=>"010001100",
  63162=>"111110000",
  63163=>"101011111",
  63164=>"100000110",
  63165=>"010111100",
  63166=>"111101101",
  63167=>"110110010",
  63168=>"011100010",
  63169=>"100011111",
  63170=>"110100101",
  63171=>"001011011",
  63172=>"010100011",
  63173=>"010100010",
  63174=>"001010011",
  63175=>"110010101",
  63176=>"000100000",
  63177=>"100011100",
  63178=>"100101000",
  63179=>"000101001",
  63180=>"000110010",
  63181=>"110001000",
  63182=>"001111010",
  63183=>"110100100",
  63184=>"111111110",
  63185=>"000000101",
  63186=>"001001011",
  63187=>"110101110",
  63188=>"001101100",
  63189=>"110101111",
  63190=>"101101011",
  63191=>"111101011",
  63192=>"010100111",
  63193=>"110011001",
  63194=>"111001101",
  63195=>"111110111",
  63196=>"001111110",
  63197=>"001000111",
  63198=>"010011101",
  63199=>"000000010",
  63200=>"111111000",
  63201=>"010101111",
  63202=>"111111110",
  63203=>"101010110",
  63204=>"110010000",
  63205=>"001110101",
  63206=>"001001001",
  63207=>"000001110",
  63208=>"000110100",
  63209=>"011001011",
  63210=>"010100101",
  63211=>"000010111",
  63212=>"000010100",
  63213=>"000001010",
  63214=>"110011100",
  63215=>"100101111",
  63216=>"101000000",
  63217=>"000011101",
  63218=>"001100110",
  63219=>"100000000",
  63220=>"011111111",
  63221=>"100010000",
  63222=>"011010000",
  63223=>"001100001",
  63224=>"011001000",
  63225=>"010010000",
  63226=>"000010011",
  63227=>"101000001",
  63228=>"110011100",
  63229=>"100011001",
  63230=>"110001010",
  63231=>"101111100",
  63232=>"000000100",
  63233=>"111000111",
  63234=>"011001001",
  63235=>"011100011",
  63236=>"100110000",
  63237=>"100001100",
  63238=>"100010000",
  63239=>"101100110",
  63240=>"000101110",
  63241=>"100111000",
  63242=>"010111001",
  63243=>"101100000",
  63244=>"111000100",
  63245=>"010001111",
  63246=>"111101000",
  63247=>"100000100",
  63248=>"111010010",
  63249=>"011100010",
  63250=>"000011111",
  63251=>"111010110",
  63252=>"111110100",
  63253=>"110010100",
  63254=>"111000000",
  63255=>"001001110",
  63256=>"011110111",
  63257=>"110011100",
  63258=>"111001010",
  63259=>"111011100",
  63260=>"111111110",
  63261=>"110101010",
  63262=>"110111010",
  63263=>"100001110",
  63264=>"010101101",
  63265=>"010100111",
  63266=>"100110110",
  63267=>"000110101",
  63268=>"101010111",
  63269=>"011100111",
  63270=>"001110100",
  63271=>"001001011",
  63272=>"111100011",
  63273=>"110001111",
  63274=>"011010001",
  63275=>"011101101",
  63276=>"111110100",
  63277=>"111010001",
  63278=>"100101000",
  63279=>"110001111",
  63280=>"011001100",
  63281=>"111101101",
  63282=>"101101000",
  63283=>"101001110",
  63284=>"110111000",
  63285=>"101110110",
  63286=>"011010010",
  63287=>"110110001",
  63288=>"000010110",
  63289=>"010011001",
  63290=>"001110111",
  63291=>"111000110",
  63292=>"100000010",
  63293=>"111101111",
  63294=>"000100010",
  63295=>"000101000",
  63296=>"100001110",
  63297=>"011110110",
  63298=>"101010100",
  63299=>"111001110",
  63300=>"001001111",
  63301=>"010111101",
  63302=>"011111000",
  63303=>"001010011",
  63304=>"110010110",
  63305=>"000110100",
  63306=>"100110111",
  63307=>"011110111",
  63308=>"010000010",
  63309=>"110101100",
  63310=>"011110001",
  63311=>"001010110",
  63312=>"000111101",
  63313=>"001001001",
  63314=>"110011100",
  63315=>"101000010",
  63316=>"100100110",
  63317=>"011000110",
  63318=>"010110001",
  63319=>"010110001",
  63320=>"101011000",
  63321=>"001000011",
  63322=>"100010111",
  63323=>"000111001",
  63324=>"101001010",
  63325=>"111110101",
  63326=>"110101000",
  63327=>"111111010",
  63328=>"011011011",
  63329=>"011011110",
  63330=>"111000111",
  63331=>"111010001",
  63332=>"101001000",
  63333=>"001000100",
  63334=>"111111011",
  63335=>"111001110",
  63336=>"101101101",
  63337=>"010111011",
  63338=>"110101001",
  63339=>"001111011",
  63340=>"000001011",
  63341=>"111010000",
  63342=>"110110000",
  63343=>"001101100",
  63344=>"110100010",
  63345=>"001010100",
  63346=>"111101010",
  63347=>"111111111",
  63348=>"111101011",
  63349=>"110101001",
  63350=>"111101100",
  63351=>"000011110",
  63352=>"111010011",
  63353=>"011010011",
  63354=>"101001011",
  63355=>"011000101",
  63356=>"010110011",
  63357=>"110011100",
  63358=>"101101001",
  63359=>"100101001",
  63360=>"111111110",
  63361=>"010001001",
  63362=>"100111011",
  63363=>"111100010",
  63364=>"111010001",
  63365=>"011010100",
  63366=>"001100011",
  63367=>"101110100",
  63368=>"111010011",
  63369=>"001011100",
  63370=>"111011101",
  63371=>"100011000",
  63372=>"100000100",
  63373=>"111110101",
  63374=>"110111111",
  63375=>"001011000",
  63376=>"011000100",
  63377=>"010100011",
  63378=>"001100111",
  63379=>"000000111",
  63380=>"111110011",
  63381=>"000100001",
  63382=>"110111100",
  63383=>"101010011",
  63384=>"101001101",
  63385=>"011100010",
  63386=>"000000111",
  63387=>"011001111",
  63388=>"110011010",
  63389=>"111001101",
  63390=>"100000100",
  63391=>"101000001",
  63392=>"000000110",
  63393=>"111000001",
  63394=>"100110100",
  63395=>"100101000",
  63396=>"001111001",
  63397=>"100100111",
  63398=>"001110101",
  63399=>"100111001",
  63400=>"111010100",
  63401=>"100101100",
  63402=>"001110001",
  63403=>"010100101",
  63404=>"000000100",
  63405=>"010111010",
  63406=>"000000101",
  63407=>"101100111",
  63408=>"000010101",
  63409=>"011001100",
  63410=>"110010000",
  63411=>"100101110",
  63412=>"111111001",
  63413=>"010001110",
  63414=>"101011100",
  63415=>"101101110",
  63416=>"100000011",
  63417=>"011100011",
  63418=>"110000100",
  63419=>"010100011",
  63420=>"100100110",
  63421=>"100001000",
  63422=>"000111100",
  63423=>"000011011",
  63424=>"001011000",
  63425=>"011011000",
  63426=>"000101100",
  63427=>"010110110",
  63428=>"010001101",
  63429=>"000000111",
  63430=>"010110111",
  63431=>"000010000",
  63432=>"001011000",
  63433=>"100111101",
  63434=>"010001101",
  63435=>"011110111",
  63436=>"000100111",
  63437=>"100100010",
  63438=>"010110101",
  63439=>"100111100",
  63440=>"011101001",
  63441=>"110010111",
  63442=>"110100101",
  63443=>"110111000",
  63444=>"010001111",
  63445=>"100100011",
  63446=>"000100010",
  63447=>"011111100",
  63448=>"111110011",
  63449=>"010111011",
  63450=>"111000100",
  63451=>"110110100",
  63452=>"010101111",
  63453=>"101010011",
  63454=>"111111001",
  63455=>"100101111",
  63456=>"111101001",
  63457=>"011000111",
  63458=>"000110110",
  63459=>"110111101",
  63460=>"000011101",
  63461=>"011100110",
  63462=>"101000010",
  63463=>"110101001",
  63464=>"000001100",
  63465=>"101100100",
  63466=>"110101000",
  63467=>"000011010",
  63468=>"011111001",
  63469=>"110101010",
  63470=>"001011110",
  63471=>"000101010",
  63472=>"111100000",
  63473=>"000000010",
  63474=>"101011001",
  63475=>"001001000",
  63476=>"010110101",
  63477=>"010000010",
  63478=>"000000111",
  63479=>"111001010",
  63480=>"011000011",
  63481=>"010011101",
  63482=>"110101010",
  63483=>"000001110",
  63484=>"001101111",
  63485=>"001101011",
  63486=>"101001000",
  63487=>"010011111",
  63488=>"100000100",
  63489=>"000000110",
  63490=>"000101010",
  63491=>"100100001",
  63492=>"111100101",
  63493=>"111000000",
  63494=>"001100010",
  63495=>"100010011",
  63496=>"101001011",
  63497=>"101100010",
  63498=>"100101011",
  63499=>"100010011",
  63500=>"101111000",
  63501=>"101010010",
  63502=>"000010110",
  63503=>"101010001",
  63504=>"110110110",
  63505=>"100101110",
  63506=>"000010010",
  63507=>"000100101",
  63508=>"011111001",
  63509=>"100101000",
  63510=>"000001100",
  63511=>"110111111",
  63512=>"011000100",
  63513=>"000100110",
  63514=>"111111001",
  63515=>"110100100",
  63516=>"100100001",
  63517=>"101000010",
  63518=>"010110001",
  63519=>"000010111",
  63520=>"010000000",
  63521=>"110110010",
  63522=>"111111101",
  63523=>"001010011",
  63524=>"100010101",
  63525=>"111110101",
  63526=>"100011110",
  63527=>"100010100",
  63528=>"111111110",
  63529=>"100100010",
  63530=>"111101011",
  63531=>"000011011",
  63532=>"000100001",
  63533=>"111101101",
  63534=>"101001011",
  63535=>"010111100",
  63536=>"010111110",
  63537=>"100110001",
  63538=>"111111100",
  63539=>"101101011",
  63540=>"000111101",
  63541=>"001000110",
  63542=>"010000101",
  63543=>"111011010",
  63544=>"000110110",
  63545=>"110100011",
  63546=>"111001000",
  63547=>"000110000",
  63548=>"011011110",
  63549=>"011110000",
  63550=>"000101100",
  63551=>"001000011",
  63552=>"110110100",
  63553=>"110001010",
  63554=>"011111011",
  63555=>"010011110",
  63556=>"001001101",
  63557=>"010111000",
  63558=>"100010111",
  63559=>"100000110",
  63560=>"101010000",
  63561=>"011110011",
  63562=>"001110001",
  63563=>"000111110",
  63564=>"010001011",
  63565=>"010000100",
  63566=>"001111010",
  63567=>"001001111",
  63568=>"111011111",
  63569=>"011111010",
  63570=>"110010100",
  63571=>"011011100",
  63572=>"000110101",
  63573=>"111110110",
  63574=>"110010001",
  63575=>"111001100",
  63576=>"011000011",
  63577=>"101110010",
  63578=>"000010010",
  63579=>"100000110",
  63580=>"010000100",
  63581=>"110110101",
  63582=>"000001101",
  63583=>"000000000",
  63584=>"100001010",
  63585=>"010011011",
  63586=>"011101000",
  63587=>"011110110",
  63588=>"101111010",
  63589=>"100001010",
  63590=>"000000000",
  63591=>"000010010",
  63592=>"110000110",
  63593=>"000100011",
  63594=>"110010010",
  63595=>"011010011",
  63596=>"001100110",
  63597=>"001000001",
  63598=>"111101001",
  63599=>"000011010",
  63600=>"001001001",
  63601=>"000000010",
  63602=>"010000000",
  63603=>"001011100",
  63604=>"111000110",
  63605=>"001001101",
  63606=>"100101101",
  63607=>"101110001",
  63608=>"000101110",
  63609=>"000000011",
  63610=>"001001101",
  63611=>"110000001",
  63612=>"010001100",
  63613=>"101011000",
  63614=>"011110100",
  63615=>"001010110",
  63616=>"001101011",
  63617=>"001101000",
  63618=>"101100111",
  63619=>"100001100",
  63620=>"010000111",
  63621=>"110100101",
  63622=>"110011111",
  63623=>"000111111",
  63624=>"111010111",
  63625=>"101111010",
  63626=>"111101110",
  63627=>"110000100",
  63628=>"011110001",
  63629=>"011000000",
  63630=>"110001011",
  63631=>"110011011",
  63632=>"001001111",
  63633=>"011011100",
  63634=>"100001101",
  63635=>"111011111",
  63636=>"011010001",
  63637=>"011000000",
  63638=>"000011110",
  63639=>"010001100",
  63640=>"011100101",
  63641=>"000110110",
  63642=>"111011100",
  63643=>"111011111",
  63644=>"110000011",
  63645=>"111100111",
  63646=>"101111011",
  63647=>"101101100",
  63648=>"010000100",
  63649=>"100110100",
  63650=>"111010100",
  63651=>"001111010",
  63652=>"000101011",
  63653=>"000100011",
  63654=>"010011011",
  63655=>"111101001",
  63656=>"001110001",
  63657=>"010001111",
  63658=>"000110001",
  63659=>"011111010",
  63660=>"011100101",
  63661=>"110011110",
  63662=>"000100011",
  63663=>"100000100",
  63664=>"010110011",
  63665=>"001101110",
  63666=>"001111100",
  63667=>"000000101",
  63668=>"101111000",
  63669=>"010010100",
  63670=>"100001101",
  63671=>"010000100",
  63672=>"101000101",
  63673=>"100000111",
  63674=>"001001100",
  63675=>"100010101",
  63676=>"010010010",
  63677=>"111000110",
  63678=>"001111101",
  63679=>"001100101",
  63680=>"011101101",
  63681=>"100110100",
  63682=>"000000101",
  63683=>"000000100",
  63684=>"011001001",
  63685=>"111010101",
  63686=>"010000001",
  63687=>"000101100",
  63688=>"010111111",
  63689=>"011101110",
  63690=>"000110010",
  63691=>"110100101",
  63692=>"100001100",
  63693=>"111110011",
  63694=>"110110001",
  63695=>"001110100",
  63696=>"100110110",
  63697=>"000110001",
  63698=>"110111101",
  63699=>"011101001",
  63700=>"001101101",
  63701=>"111100111",
  63702=>"101011010",
  63703=>"001101100",
  63704=>"010001000",
  63705=>"100011001",
  63706=>"100001100",
  63707=>"100111000",
  63708=>"011001000",
  63709=>"001111011",
  63710=>"111101000",
  63711=>"011110011",
  63712=>"001111000",
  63713=>"011000001",
  63714=>"110111110",
  63715=>"011100111",
  63716=>"000011011",
  63717=>"110101101",
  63718=>"010000010",
  63719=>"101010111",
  63720=>"100010001",
  63721=>"001101101",
  63722=>"100001000",
  63723=>"000010010",
  63724=>"100000010",
  63725=>"110010110",
  63726=>"111000101",
  63727=>"011011110",
  63728=>"010001011",
  63729=>"111011001",
  63730=>"010011101",
  63731=>"110110111",
  63732=>"101111000",
  63733=>"101110110",
  63734=>"100000101",
  63735=>"111010100",
  63736=>"100101010",
  63737=>"111101000",
  63738=>"000011111",
  63739=>"011000011",
  63740=>"100111100",
  63741=>"001001000",
  63742=>"100000010",
  63743=>"100000010",
  63744=>"000011100",
  63745=>"011100100",
  63746=>"010100100",
  63747=>"010001100",
  63748=>"101101101",
  63749=>"100000111",
  63750=>"101011101",
  63751=>"000110111",
  63752=>"011001110",
  63753=>"101000001",
  63754=>"011100110",
  63755=>"000111111",
  63756=>"010111001",
  63757=>"000010000",
  63758=>"100100100",
  63759=>"010011101",
  63760=>"111000111",
  63761=>"111110111",
  63762=>"001111010",
  63763=>"100010001",
  63764=>"110000111",
  63765=>"111100011",
  63766=>"111111110",
  63767=>"110001000",
  63768=>"101001011",
  63769=>"011001101",
  63770=>"000100001",
  63771=>"000000100",
  63772=>"100001000",
  63773=>"010001111",
  63774=>"000101101",
  63775=>"000110100",
  63776=>"011101101",
  63777=>"011001011",
  63778=>"111010101",
  63779=>"100011011",
  63780=>"110110010",
  63781=>"011000110",
  63782=>"111101110",
  63783=>"011000110",
  63784=>"101011000",
  63785=>"001100101",
  63786=>"110101110",
  63787=>"010000001",
  63788=>"000001010",
  63789=>"100010010",
  63790=>"010011000",
  63791=>"111110100",
  63792=>"110100100",
  63793=>"110001001",
  63794=>"010011101",
  63795=>"000111000",
  63796=>"111111011",
  63797=>"010100001",
  63798=>"100111100",
  63799=>"000110111",
  63800=>"100000101",
  63801=>"101100111",
  63802=>"001110011",
  63803=>"001001110",
  63804=>"000110110",
  63805=>"001010100",
  63806=>"001011110",
  63807=>"111110110",
  63808=>"001111111",
  63809=>"111110111",
  63810=>"111100110",
  63811=>"111111011",
  63812=>"000100101",
  63813=>"011011101",
  63814=>"101111101",
  63815=>"110011010",
  63816=>"101101110",
  63817=>"001011010",
  63818=>"101001111",
  63819=>"000111101",
  63820=>"010101001",
  63821=>"001111100",
  63822=>"001111011",
  63823=>"000110100",
  63824=>"110011101",
  63825=>"101100001",
  63826=>"010010011",
  63827=>"000101011",
  63828=>"100000001",
  63829=>"001010010",
  63830=>"101011100",
  63831=>"111010101",
  63832=>"101000010",
  63833=>"110100110",
  63834=>"111101100",
  63835=>"011110111",
  63836=>"001111101",
  63837=>"011000110",
  63838=>"001100001",
  63839=>"011100011",
  63840=>"110101101",
  63841=>"101111000",
  63842=>"000100001",
  63843=>"101000100",
  63844=>"001011111",
  63845=>"111010101",
  63846=>"011100011",
  63847=>"111010100",
  63848=>"101001000",
  63849=>"010010111",
  63850=>"010111010",
  63851=>"001001001",
  63852=>"110001001",
  63853=>"100000101",
  63854=>"001110010",
  63855=>"001011010",
  63856=>"001100000",
  63857=>"001001100",
  63858=>"110010110",
  63859=>"100101010",
  63860=>"001101010",
  63861=>"000101001",
  63862=>"101011100",
  63863=>"110100101",
  63864=>"010101101",
  63865=>"100100010",
  63866=>"011001000",
  63867=>"111100100",
  63868=>"100001110",
  63869=>"111001100",
  63870=>"111100010",
  63871=>"110000110",
  63872=>"011101111",
  63873=>"001011111",
  63874=>"000110111",
  63875=>"100011010",
  63876=>"101101111",
  63877=>"001101001",
  63878=>"111011001",
  63879=>"000000111",
  63880=>"100001010",
  63881=>"000111001",
  63882=>"001101010",
  63883=>"001001011",
  63884=>"111110000",
  63885=>"010111110",
  63886=>"101110010",
  63887=>"100111111",
  63888=>"010000111",
  63889=>"001001010",
  63890=>"010110110",
  63891=>"001001110",
  63892=>"101111011",
  63893=>"010001110",
  63894=>"101000011",
  63895=>"100111100",
  63896=>"010110100",
  63897=>"101000100",
  63898=>"000000100",
  63899=>"010100000",
  63900=>"111111100",
  63901=>"110011101",
  63902=>"111111011",
  63903=>"011101100",
  63904=>"011110110",
  63905=>"010101010",
  63906=>"111010001",
  63907=>"001010010",
  63908=>"000001000",
  63909=>"000101011",
  63910=>"110010100",
  63911=>"001100110",
  63912=>"000001110",
  63913=>"101111001",
  63914=>"001110101",
  63915=>"011011111",
  63916=>"011111101",
  63917=>"010110111",
  63918=>"100000110",
  63919=>"111101011",
  63920=>"000001001",
  63921=>"011111010",
  63922=>"111101111",
  63923=>"001100000",
  63924=>"011110001",
  63925=>"001110111",
  63926=>"101101001",
  63927=>"100011011",
  63928=>"110001110",
  63929=>"000000110",
  63930=>"001000101",
  63931=>"010001001",
  63932=>"100011110",
  63933=>"100111001",
  63934=>"011110011",
  63935=>"101010101",
  63936=>"111111000",
  63937=>"100010001",
  63938=>"111011001",
  63939=>"010010010",
  63940=>"011011100",
  63941=>"101111101",
  63942=>"001001000",
  63943=>"111011100",
  63944=>"000100111",
  63945=>"111011100",
  63946=>"011111110",
  63947=>"100110001",
  63948=>"101010100",
  63949=>"110000100",
  63950=>"111000111",
  63951=>"110001111",
  63952=>"011001000",
  63953=>"101111100",
  63954=>"111101010",
  63955=>"100111010",
  63956=>"100111110",
  63957=>"100111000",
  63958=>"011111100",
  63959=>"011010111",
  63960=>"000000100",
  63961=>"100110101",
  63962=>"100110111",
  63963=>"110000011",
  63964=>"101100000",
  63965=>"001101100",
  63966=>"110001101",
  63967=>"110110100",
  63968=>"100110001",
  63969=>"100001011",
  63970=>"011000111",
  63971=>"110101101",
  63972=>"100100100",
  63973=>"110010111",
  63974=>"001010010",
  63975=>"000101100",
  63976=>"001110001",
  63977=>"101101001",
  63978=>"011010101",
  63979=>"101100011",
  63980=>"100100111",
  63981=>"110010001",
  63982=>"000010101",
  63983=>"111110010",
  63984=>"101011101",
  63985=>"010011100",
  63986=>"011010101",
  63987=>"110001010",
  63988=>"111100100",
  63989=>"000011011",
  63990=>"000101010",
  63991=>"110010100",
  63992=>"100101000",
  63993=>"101001100",
  63994=>"111110111",
  63995=>"110110111",
  63996=>"001000010",
  63997=>"011001110",
  63998=>"110101100",
  63999=>"001010001",
  64000=>"001000101",
  64001=>"101011010",
  64002=>"110001100",
  64003=>"000101111",
  64004=>"110000110",
  64005=>"110011101",
  64006=>"010001110",
  64007=>"101101010",
  64008=>"101101001",
  64009=>"001001001",
  64010=>"101110100",
  64011=>"000110111",
  64012=>"000001000",
  64013=>"010000100",
  64014=>"101001001",
  64015=>"111101010",
  64016=>"101100101",
  64017=>"000010101",
  64018=>"100101110",
  64019=>"111100011",
  64020=>"011001001",
  64021=>"101111110",
  64022=>"001010001",
  64023=>"111101111",
  64024=>"100010100",
  64025=>"111110101",
  64026=>"010101000",
  64027=>"001111110",
  64028=>"101010011",
  64029=>"000100111",
  64030=>"100100111",
  64031=>"100010111",
  64032=>"110110010",
  64033=>"100000011",
  64034=>"001000100",
  64035=>"001101001",
  64036=>"001100100",
  64037=>"110000110",
  64038=>"010011010",
  64039=>"010001111",
  64040=>"110001000",
  64041=>"001011100",
  64042=>"000111111",
  64043=>"111000110",
  64044=>"011111100",
  64045=>"000110101",
  64046=>"001011001",
  64047=>"111000101",
  64048=>"110000111",
  64049=>"110111101",
  64050=>"010001100",
  64051=>"110100110",
  64052=>"000001011",
  64053=>"010111101",
  64054=>"111110001",
  64055=>"000111111",
  64056=>"111100110",
  64057=>"001100001",
  64058=>"100110011",
  64059=>"110000010",
  64060=>"000100011",
  64061=>"101110011",
  64062=>"000100010",
  64063=>"011100100",
  64064=>"010100010",
  64065=>"011011111",
  64066=>"111010001",
  64067=>"011010010",
  64068=>"100001011",
  64069=>"110100010",
  64070=>"011010000",
  64071=>"110110001",
  64072=>"100100011",
  64073=>"010110111",
  64074=>"100010011",
  64075=>"011100000",
  64076=>"101011010",
  64077=>"010010100",
  64078=>"111110110",
  64079=>"000011010",
  64080=>"000110100",
  64081=>"010111011",
  64082=>"100100001",
  64083=>"110110100",
  64084=>"101010000",
  64085=>"010101101",
  64086=>"100010110",
  64087=>"000101010",
  64088=>"101100011",
  64089=>"101101111",
  64090=>"101100001",
  64091=>"000101111",
  64092=>"000100010",
  64093=>"001001010",
  64094=>"100001110",
  64095=>"001011111",
  64096=>"111110000",
  64097=>"010010111",
  64098=>"010111000",
  64099=>"011001000",
  64100=>"001111010",
  64101=>"100101001",
  64102=>"111001100",
  64103=>"000011111",
  64104=>"110111101",
  64105=>"100010011",
  64106=>"110100000",
  64107=>"000010111",
  64108=>"010000110",
  64109=>"010110110",
  64110=>"011110101",
  64111=>"101100111",
  64112=>"010000001",
  64113=>"110100100",
  64114=>"100111011",
  64115=>"100001010",
  64116=>"100110011",
  64117=>"001000111",
  64118=>"000011110",
  64119=>"100111100",
  64120=>"000011101",
  64121=>"001011110",
  64122=>"000110001",
  64123=>"100011010",
  64124=>"001111101",
  64125=>"011101101",
  64126=>"100100101",
  64127=>"010111011",
  64128=>"111011011",
  64129=>"001100111",
  64130=>"101110100",
  64131=>"110001000",
  64132=>"001011100",
  64133=>"011011001",
  64134=>"101111101",
  64135=>"001100000",
  64136=>"000000100",
  64137=>"101011011",
  64138=>"101010000",
  64139=>"110110001",
  64140=>"001000100",
  64141=>"011100111",
  64142=>"101110000",
  64143=>"000111101",
  64144=>"000001000",
  64145=>"011001011",
  64146=>"111100000",
  64147=>"100100111",
  64148=>"001010010",
  64149=>"000110111",
  64150=>"110010001",
  64151=>"110101111",
  64152=>"111111111",
  64153=>"100101101",
  64154=>"100001110",
  64155=>"001001011",
  64156=>"010010100",
  64157=>"000001011",
  64158=>"000001011",
  64159=>"110001111",
  64160=>"101000010",
  64161=>"011001101",
  64162=>"000000010",
  64163=>"001111101",
  64164=>"100010010",
  64165=>"000010110",
  64166=>"101000100",
  64167=>"010011010",
  64168=>"110111000",
  64169=>"010010111",
  64170=>"010001000",
  64171=>"100111111",
  64172=>"001101100",
  64173=>"001100000",
  64174=>"100000011",
  64175=>"101010010",
  64176=>"100110010",
  64177=>"010111111",
  64178=>"101110010",
  64179=>"010010001",
  64180=>"110110011",
  64181=>"100101000",
  64182=>"000100010",
  64183=>"001110010",
  64184=>"011100001",
  64185=>"011100111",
  64186=>"100101000",
  64187=>"010111011",
  64188=>"101000111",
  64189=>"010110001",
  64190=>"110001001",
  64191=>"011111011",
  64192=>"111010110",
  64193=>"001010100",
  64194=>"011001000",
  64195=>"110101011",
  64196=>"000100000",
  64197=>"000110100",
  64198=>"000001010",
  64199=>"101011111",
  64200=>"110001001",
  64201=>"110010000",
  64202=>"010001011",
  64203=>"100101010",
  64204=>"100100101",
  64205=>"011110101",
  64206=>"101000101",
  64207=>"011000100",
  64208=>"000001110",
  64209=>"100101110",
  64210=>"101100111",
  64211=>"111101000",
  64212=>"111110001",
  64213=>"000000001",
  64214=>"011111101",
  64215=>"111101011",
  64216=>"000000011",
  64217=>"010010111",
  64218=>"000110100",
  64219=>"111001100",
  64220=>"000101001",
  64221=>"001001001",
  64222=>"100010100",
  64223=>"110001001",
  64224=>"010000101",
  64225=>"100100110",
  64226=>"111000001",
  64227=>"010111100",
  64228=>"110101100",
  64229=>"001000101",
  64230=>"001011001",
  64231=>"001100011",
  64232=>"000000110",
  64233=>"010101100",
  64234=>"011101011",
  64235=>"010111000",
  64236=>"001001101",
  64237=>"000101000",
  64238=>"111011011",
  64239=>"101010000",
  64240=>"111101100",
  64241=>"000001011",
  64242=>"010110110",
  64243=>"110100111",
  64244=>"111101111",
  64245=>"100000101",
  64246=>"011010001",
  64247=>"101010100",
  64248=>"000000110",
  64249=>"010110011",
  64250=>"101111001",
  64251=>"110000011",
  64252=>"111110010",
  64253=>"000011101",
  64254=>"101000101",
  64255=>"100110011",
  64256=>"010101010",
  64257=>"010000111",
  64258=>"000101001",
  64259=>"100110011",
  64260=>"010101100",
  64261=>"000001000",
  64262=>"110001101",
  64263=>"100001101",
  64264=>"010001111",
  64265=>"010111000",
  64266=>"110001111",
  64267=>"001011011",
  64268=>"100100101",
  64269=>"100101010",
  64270=>"101101111",
  64271=>"111111010",
  64272=>"010001001",
  64273=>"000001100",
  64274=>"111111100",
  64275=>"000001111",
  64276=>"101000111",
  64277=>"111101000",
  64278=>"110001010",
  64279=>"011010000",
  64280=>"001100001",
  64281=>"001001110",
  64282=>"000001001",
  64283=>"000110111",
  64284=>"000001010",
  64285=>"101010101",
  64286=>"111010010",
  64287=>"101111110",
  64288=>"110110100",
  64289=>"110001001",
  64290=>"111011101",
  64291=>"110010000",
  64292=>"100101011",
  64293=>"000110010",
  64294=>"010110111",
  64295=>"110110010",
  64296=>"111101101",
  64297=>"111110011",
  64298=>"000000010",
  64299=>"001101001",
  64300=>"101100000",
  64301=>"000011111",
  64302=>"001001111",
  64303=>"111000011",
  64304=>"011000000",
  64305=>"100010001",
  64306=>"011001001",
  64307=>"010100100",
  64308=>"111110110",
  64309=>"010101100",
  64310=>"000001100",
  64311=>"101001000",
  64312=>"101101101",
  64313=>"111001000",
  64314=>"101000010",
  64315=>"110110101",
  64316=>"010111100",
  64317=>"000111110",
  64318=>"101011110",
  64319=>"000110111",
  64320=>"100110111",
  64321=>"111111110",
  64322=>"010100000",
  64323=>"101110010",
  64324=>"001110100",
  64325=>"010000001",
  64326=>"100000010",
  64327=>"010011010",
  64328=>"101001010",
  64329=>"100101111",
  64330=>"010111001",
  64331=>"111010010",
  64332=>"100011011",
  64333=>"100010011",
  64334=>"000111000",
  64335=>"101001101",
  64336=>"000001101",
  64337=>"101101101",
  64338=>"111001010",
  64339=>"100101011",
  64340=>"100000110",
  64341=>"010000111",
  64342=>"110000001",
  64343=>"000011001",
  64344=>"110010000",
  64345=>"111000101",
  64346=>"110100110",
  64347=>"111110000",
  64348=>"001110000",
  64349=>"001110001",
  64350=>"101111011",
  64351=>"110000111",
  64352=>"111010111",
  64353=>"010100011",
  64354=>"000010010",
  64355=>"011010000",
  64356=>"111100111",
  64357=>"100110100",
  64358=>"100100111",
  64359=>"011001011",
  64360=>"101001011",
  64361=>"010110011",
  64362=>"011010001",
  64363=>"111101000",
  64364=>"110000111",
  64365=>"110101001",
  64366=>"001000000",
  64367=>"011101111",
  64368=>"100010110",
  64369=>"111001000",
  64370=>"111000111",
  64371=>"111011001",
  64372=>"010101111",
  64373=>"000011001",
  64374=>"001110011",
  64375=>"111001000",
  64376=>"010110000",
  64377=>"100100001",
  64378=>"110100110",
  64379=>"010110110",
  64380=>"010011010",
  64381=>"001010010",
  64382=>"001101001",
  64383=>"011011101",
  64384=>"000010000",
  64385=>"011101010",
  64386=>"001101111",
  64387=>"001100111",
  64388=>"110001111",
  64389=>"100000101",
  64390=>"000111000",
  64391=>"001001001",
  64392=>"011110011",
  64393=>"100111001",
  64394=>"010010000",
  64395=>"110110101",
  64396=>"111001110",
  64397=>"001000000",
  64398=>"000100001",
  64399=>"101110010",
  64400=>"001000100",
  64401=>"111111111",
  64402=>"100110011",
  64403=>"011110110",
  64404=>"011110100",
  64405=>"011011110",
  64406=>"011000011",
  64407=>"001100000",
  64408=>"001001000",
  64409=>"101001011",
  64410=>"000001100",
  64411=>"000001010",
  64412=>"110011001",
  64413=>"000110011",
  64414=>"001010001",
  64415=>"111101000",
  64416=>"001101001",
  64417=>"110011001",
  64418=>"111101001",
  64419=>"101010101",
  64420=>"110011101",
  64421=>"000100111",
  64422=>"010111100",
  64423=>"000011000",
  64424=>"000111110",
  64425=>"001011011",
  64426=>"011111101",
  64427=>"101000101",
  64428=>"000011000",
  64429=>"011110010",
  64430=>"111011110",
  64431=>"111110001",
  64432=>"010011011",
  64433=>"101010111",
  64434=>"100001101",
  64435=>"000001011",
  64436=>"101101000",
  64437=>"001110010",
  64438=>"011110111",
  64439=>"111111011",
  64440=>"110000111",
  64441=>"001100000",
  64442=>"101011101",
  64443=>"100000100",
  64444=>"100100001",
  64445=>"000000001",
  64446=>"100101111",
  64447=>"010000001",
  64448=>"101100001",
  64449=>"011001100",
  64450=>"000101111",
  64451=>"111111110",
  64452=>"100001010",
  64453=>"100011111",
  64454=>"110010100",
  64455=>"110110011",
  64456=>"000100001",
  64457=>"101111111",
  64458=>"010001000",
  64459=>"110001011",
  64460=>"000010001",
  64461=>"100100110",
  64462=>"100000100",
  64463=>"000110000",
  64464=>"011010001",
  64465=>"000010000",
  64466=>"110101001",
  64467=>"000101000",
  64468=>"110001110",
  64469=>"111101000",
  64470=>"010100101",
  64471=>"110100111",
  64472=>"000000001",
  64473=>"111111011",
  64474=>"111000101",
  64475=>"110101100",
  64476=>"000000000",
  64477=>"101110111",
  64478=>"100101001",
  64479=>"001000010",
  64480=>"000111010",
  64481=>"100101111",
  64482=>"001001000",
  64483=>"011011101",
  64484=>"000000111",
  64485=>"001010111",
  64486=>"110101000",
  64487=>"001100010",
  64488=>"000001100",
  64489=>"100000010",
  64490=>"000101100",
  64491=>"111001110",
  64492=>"001111101",
  64493=>"111000111",
  64494=>"000101000",
  64495=>"001001111",
  64496=>"110000010",
  64497=>"101010110",
  64498=>"110010101",
  64499=>"101110001",
  64500=>"010101111",
  64501=>"110101101",
  64502=>"010000000",
  64503=>"000001110",
  64504=>"111101011",
  64505=>"000111010",
  64506=>"100111110",
  64507=>"100100011",
  64508=>"001001001",
  64509=>"001011000",
  64510=>"000011101",
  64511=>"011111011",
  64512=>"000100000",
  64513=>"001001011",
  64514=>"000001000",
  64515=>"101101110",
  64516=>"001011111",
  64517=>"000011000",
  64518=>"100000111",
  64519=>"111011110",
  64520=>"010001101",
  64521=>"001100100",
  64522=>"001110000",
  64523=>"010001100",
  64524=>"010001100",
  64525=>"111101101",
  64526=>"001101111",
  64527=>"111111100",
  64528=>"000010110",
  64529=>"010001010",
  64530=>"110101101",
  64531=>"111101001",
  64532=>"001011001",
  64533=>"101000101",
  64534=>"011011100",
  64535=>"111111000",
  64536=>"011010011",
  64537=>"101011000",
  64538=>"101000111",
  64539=>"100010001",
  64540=>"001011110",
  64541=>"111110110",
  64542=>"110101100",
  64543=>"100010011",
  64544=>"111111110",
  64545=>"110100100",
  64546=>"011011110",
  64547=>"111101000",
  64548=>"101011010",
  64549=>"100110100",
  64550=>"111010001",
  64551=>"110010101",
  64552=>"000001010",
  64553=>"001101000",
  64554=>"011101101",
  64555=>"001100011",
  64556=>"100011000",
  64557=>"101010011",
  64558=>"101101000",
  64559=>"101001100",
  64560=>"000101010",
  64561=>"111100010",
  64562=>"001110000",
  64563=>"010101111",
  64564=>"011000001",
  64565=>"011101110",
  64566=>"101101011",
  64567=>"100010000",
  64568=>"101010110",
  64569=>"100000111",
  64570=>"110011000",
  64571=>"101000001",
  64572=>"101101011",
  64573=>"001010011",
  64574=>"001110010",
  64575=>"001011110",
  64576=>"111000100",
  64577=>"000011000",
  64578=>"000011011",
  64579=>"110000011",
  64580=>"110110101",
  64581=>"001010101",
  64582=>"001010101",
  64583=>"100010110",
  64584=>"001011001",
  64585=>"001011111",
  64586=>"000100100",
  64587=>"000110010",
  64588=>"010010000",
  64589=>"011110100",
  64590=>"111100111",
  64591=>"001110000",
  64592=>"100000001",
  64593=>"000110000",
  64594=>"000011100",
  64595=>"000000101",
  64596=>"101101101",
  64597=>"101011010",
  64598=>"101110011",
  64599=>"001100000",
  64600=>"000110010",
  64601=>"001110111",
  64602=>"110000011",
  64603=>"001000001",
  64604=>"111100101",
  64605=>"111111010",
  64606=>"011010001",
  64607=>"011000000",
  64608=>"001010101",
  64609=>"010011011",
  64610=>"011000101",
  64611=>"000100011",
  64612=>"011000010",
  64613=>"000111101",
  64614=>"000010101",
  64615=>"111010000",
  64616=>"011010010",
  64617=>"100010111",
  64618=>"111100110",
  64619=>"111100110",
  64620=>"101010000",
  64621=>"010110101",
  64622=>"011100010",
  64623=>"110111101",
  64624=>"011001011",
  64625=>"100111001",
  64626=>"101000110",
  64627=>"110011010",
  64628=>"101100101",
  64629=>"010001011",
  64630=>"111111111",
  64631=>"110011101",
  64632=>"000101010",
  64633=>"111100000",
  64634=>"100010111",
  64635=>"000010111",
  64636=>"111110101",
  64637=>"100101000",
  64638=>"010001010",
  64639=>"100000111",
  64640=>"101010110",
  64641=>"011010110",
  64642=>"000111001",
  64643=>"100000000",
  64644=>"001101011",
  64645=>"100110010",
  64646=>"101111000",
  64647=>"111111101",
  64648=>"011000010",
  64649=>"000100010",
  64650=>"010010001",
  64651=>"010111101",
  64652=>"101110110",
  64653=>"011101000",
  64654=>"011001110",
  64655=>"000011010",
  64656=>"011011001",
  64657=>"101011111",
  64658=>"001010010",
  64659=>"101000010",
  64660=>"111010000",
  64661=>"011011101",
  64662=>"110111110",
  64663=>"101011101",
  64664=>"001011011",
  64665=>"111001100",
  64666=>"010010010",
  64667=>"000100111",
  64668=>"011010011",
  64669=>"011101110",
  64670=>"100101001",
  64671=>"010000101",
  64672=>"001000010",
  64673=>"010110011",
  64674=>"111100000",
  64675=>"100001101",
  64676=>"011100110",
  64677=>"000110010",
  64678=>"001110100",
  64679=>"101110000",
  64680=>"100110000",
  64681=>"001100010",
  64682=>"000111000",
  64683=>"100111110",
  64684=>"111011011",
  64685=>"010001100",
  64686=>"111101011",
  64687=>"000001001",
  64688=>"110010000",
  64689=>"001110000",
  64690=>"001100011",
  64691=>"110000000",
  64692=>"110001010",
  64693=>"001010100",
  64694=>"101000010",
  64695=>"101011111",
  64696=>"011000011",
  64697=>"000101101",
  64698=>"000100000",
  64699=>"001001111",
  64700=>"101111111",
  64701=>"000111100",
  64702=>"111110100",
  64703=>"010010100",
  64704=>"111011110",
  64705=>"110110101",
  64706=>"100001111",
  64707=>"101101100",
  64708=>"101100001",
  64709=>"010011000",
  64710=>"010111111",
  64711=>"000110001",
  64712=>"110111001",
  64713=>"101110011",
  64714=>"111101010",
  64715=>"111000000",
  64716=>"101010011",
  64717=>"011010110",
  64718=>"111101110",
  64719=>"100011111",
  64720=>"111100000",
  64721=>"110001010",
  64722=>"101001000",
  64723=>"001100000",
  64724=>"000101101",
  64725=>"101101000",
  64726=>"011010100",
  64727=>"011111100",
  64728=>"001011010",
  64729=>"000110110",
  64730=>"111001110",
  64731=>"110000000",
  64732=>"010001000",
  64733=>"110110100",
  64734=>"000100000",
  64735=>"110010000",
  64736=>"011101000",
  64737=>"111101010",
  64738=>"000011111",
  64739=>"011111010",
  64740=>"100100100",
  64741=>"000101111",
  64742=>"011010001",
  64743=>"101011110",
  64744=>"100011100",
  64745=>"101011110",
  64746=>"110111011",
  64747=>"001101100",
  64748=>"001110111",
  64749=>"000100010",
  64750=>"101100110",
  64751=>"000011100",
  64752=>"000101010",
  64753=>"101101010",
  64754=>"101100100",
  64755=>"001101010",
  64756=>"010010000",
  64757=>"011011011",
  64758=>"101011100",
  64759=>"010001011",
  64760=>"001100100",
  64761=>"011110111",
  64762=>"111111010",
  64763=>"011101000",
  64764=>"111001000",
  64765=>"010101110",
  64766=>"001101100",
  64767=>"110100110",
  64768=>"110010000",
  64769=>"010001000",
  64770=>"010010111",
  64771=>"110011100",
  64772=>"100000110",
  64773=>"000001111",
  64774=>"100100101",
  64775=>"101110001",
  64776=>"001000011",
  64777=>"100001101",
  64778=>"110110000",
  64779=>"101101111",
  64780=>"111110101",
  64781=>"111111101",
  64782=>"000001101",
  64783=>"010010000",
  64784=>"000010101",
  64785=>"010011000",
  64786=>"000110001",
  64787=>"100110111",
  64788=>"011100000",
  64789=>"111100001",
  64790=>"001010000",
  64791=>"011111101",
  64792=>"011101100",
  64793=>"100101001",
  64794=>"111111110",
  64795=>"001100101",
  64796=>"101100010",
  64797=>"001110110",
  64798=>"001101100",
  64799=>"001000110",
  64800=>"101000001",
  64801=>"111111110",
  64802=>"001110100",
  64803=>"100101110",
  64804=>"111110110",
  64805=>"011101100",
  64806=>"011010110",
  64807=>"000000101",
  64808=>"001011111",
  64809=>"001001011",
  64810=>"000101111",
  64811=>"011100111",
  64812=>"111011000",
  64813=>"100001011",
  64814=>"011010010",
  64815=>"001010100",
  64816=>"001100100",
  64817=>"000000010",
  64818=>"111100100",
  64819=>"000110011",
  64820=>"100010101",
  64821=>"001010111",
  64822=>"010010001",
  64823=>"000001000",
  64824=>"100000000",
  64825=>"100011011",
  64826=>"001010111",
  64827=>"000011101",
  64828=>"000000011",
  64829=>"101111110",
  64830=>"010110101",
  64831=>"001110110",
  64832=>"011010100",
  64833=>"010111111",
  64834=>"000110111",
  64835=>"000011011",
  64836=>"001111011",
  64837=>"000101001",
  64838=>"000000000",
  64839=>"000011011",
  64840=>"110001100",
  64841=>"100001010",
  64842=>"101010010",
  64843=>"010110100",
  64844=>"000010111",
  64845=>"101101101",
  64846=>"011111111",
  64847=>"111011101",
  64848=>"100011011",
  64849=>"000110101",
  64850=>"001010101",
  64851=>"100000011",
  64852=>"011111011",
  64853=>"001001001",
  64854=>"111110110",
  64855=>"100100000",
  64856=>"000001100",
  64857=>"110110001",
  64858=>"110011110",
  64859=>"000100000",
  64860=>"111101001",
  64861=>"010000100",
  64862=>"101111100",
  64863=>"001101101",
  64864=>"011111010",
  64865=>"001001001",
  64866=>"101001011",
  64867=>"000101011",
  64868=>"011000010",
  64869=>"001100000",
  64870=>"111100110",
  64871=>"100110111",
  64872=>"010110010",
  64873=>"000100010",
  64874=>"111010010",
  64875=>"010101111",
  64876=>"100000100",
  64877=>"100001111",
  64878=>"010000011",
  64879=>"010110111",
  64880=>"110111010",
  64881=>"011110011",
  64882=>"000101101",
  64883=>"010011000",
  64884=>"001010101",
  64885=>"001101100",
  64886=>"100110010",
  64887=>"100100101",
  64888=>"100100011",
  64889=>"011100101",
  64890=>"001001000",
  64891=>"111110111",
  64892=>"011100110",
  64893=>"111110000",
  64894=>"000001001",
  64895=>"010111010",
  64896=>"101000010",
  64897=>"000011101",
  64898=>"100011011",
  64899=>"010000111",
  64900=>"011001101",
  64901=>"011000011",
  64902=>"010100001",
  64903=>"101001011",
  64904=>"110110001",
  64905=>"010110010",
  64906=>"110101010",
  64907=>"110111001",
  64908=>"011111010",
  64909=>"010001110",
  64910=>"011111110",
  64911=>"110011010",
  64912=>"011001001",
  64913=>"001010001",
  64914=>"110101001",
  64915=>"001101101",
  64916=>"000000010",
  64917=>"110110110",
  64918=>"110000011",
  64919=>"101111111",
  64920=>"101111000",
  64921=>"001111110",
  64922=>"011001100",
  64923=>"011011101",
  64924=>"001101101",
  64925=>"100111011",
  64926=>"011101000",
  64927=>"000111111",
  64928=>"010010000",
  64929=>"010101110",
  64930=>"100101110",
  64931=>"111001100",
  64932=>"011111101",
  64933=>"101100010",
  64934=>"111111100",
  64935=>"111110011",
  64936=>"000010101",
  64937=>"011000010",
  64938=>"010001011",
  64939=>"000000001",
  64940=>"100001011",
  64941=>"111100010",
  64942=>"110110101",
  64943=>"011000000",
  64944=>"001001111",
  64945=>"010111111",
  64946=>"001111110",
  64947=>"100010101",
  64948=>"100000111",
  64949=>"110110101",
  64950=>"011011010",
  64951=>"111001010",
  64952=>"000001111",
  64953=>"101001110",
  64954=>"110101001",
  64955=>"011000100",
  64956=>"100000000",
  64957=>"000011000",
  64958=>"000000110",
  64959=>"111011011",
  64960=>"100001001",
  64961=>"101100001",
  64962=>"010111001",
  64963=>"000101011",
  64964=>"100010011",
  64965=>"011101000",
  64966=>"111110000",
  64967=>"101101000",
  64968=>"110000001",
  64969=>"101110011",
  64970=>"011000110",
  64971=>"101010000",
  64972=>"110001110",
  64973=>"011110101",
  64974=>"110111010",
  64975=>"001010101",
  64976=>"101000110",
  64977=>"011101000",
  64978=>"010110000",
  64979=>"111000000",
  64980=>"100001100",
  64981=>"111000000",
  64982=>"110001011",
  64983=>"111010010",
  64984=>"001011101",
  64985=>"111110001",
  64986=>"011101110",
  64987=>"101010011",
  64988=>"100100111",
  64989=>"000101000",
  64990=>"110010111",
  64991=>"111111001",
  64992=>"101001000",
  64993=>"010011110",
  64994=>"100001110",
  64995=>"111000010",
  64996=>"001000010",
  64997=>"010100011",
  64998=>"001111100",
  64999=>"101011100",
  65000=>"011110101",
  65001=>"010001110",
  65002=>"011010001",
  65003=>"111101110",
  65004=>"001111011",
  65005=>"100001111",
  65006=>"011011011",
  65007=>"110011110",
  65008=>"111010111",
  65009=>"010010110",
  65010=>"101101111",
  65011=>"110100101",
  65012=>"111010100",
  65013=>"101010001",
  65014=>"110001000",
  65015=>"100111001",
  65016=>"111111111",
  65017=>"011101010",
  65018=>"001001001",
  65019=>"011101111",
  65020=>"110010011",
  65021=>"001001110",
  65022=>"010001101",
  65023=>"011110100",
  65024=>"001100111",
  65025=>"010100101",
  65026=>"100000001",
  65027=>"011000111",
  65028=>"000111000",
  65029=>"100000100",
  65030=>"000010000",
  65031=>"100001011",
  65032=>"000011101",
  65033=>"110101100",
  65034=>"111001001",
  65035=>"011010001",
  65036=>"001011000",
  65037=>"111100000",
  65038=>"000010100",
  65039=>"110111110",
  65040=>"101100010",
  65041=>"010111011",
  65042=>"010011111",
  65043=>"111001111",
  65044=>"000111001",
  65045=>"001001000",
  65046=>"111011011",
  65047=>"111011100",
  65048=>"110111010",
  65049=>"110010001",
  65050=>"000111010",
  65051=>"001011000",
  65052=>"000011101",
  65053=>"111111100",
  65054=>"100001101",
  65055=>"111010000",
  65056=>"011110011",
  65057=>"101001101",
  65058=>"110111111",
  65059=>"101001010",
  65060=>"111111101",
  65061=>"110111101",
  65062=>"111011010",
  65063=>"001111110",
  65064=>"011000000",
  65065=>"010100011",
  65066=>"110100100",
  65067=>"100011110",
  65068=>"000010101",
  65069=>"100001000",
  65070=>"110101110",
  65071=>"101000011",
  65072=>"110000111",
  65073=>"000011111",
  65074=>"001001100",
  65075=>"010001101",
  65076=>"100010000",
  65077=>"011100100",
  65078=>"101011011",
  65079=>"111100111",
  65080=>"000110000",
  65081=>"101010101",
  65082=>"101010101",
  65083=>"100100011",
  65084=>"101101011",
  65085=>"110000000",
  65086=>"111011010",
  65087=>"101000010",
  65088=>"000001000",
  65089=>"100110001",
  65090=>"111011010",
  65091=>"000100000",
  65092=>"110100010",
  65093=>"010010001",
  65094=>"101001011",
  65095=>"010110110",
  65096=>"011001101",
  65097=>"101001100",
  65098=>"110101011",
  65099=>"011011111",
  65100=>"100000010",
  65101=>"111110001",
  65102=>"101100001",
  65103=>"001101100",
  65104=>"110101100",
  65105=>"001011100",
  65106=>"011000110",
  65107=>"010100101",
  65108=>"100001110",
  65109=>"101000100",
  65110=>"000010111",
  65111=>"001101100",
  65112=>"101100001",
  65113=>"000101011",
  65114=>"110011000",
  65115=>"001000000",
  65116=>"101011110",
  65117=>"000111010",
  65118=>"101001000",
  65119=>"011100010",
  65120=>"000100101",
  65121=>"101101000",
  65122=>"011100111",
  65123=>"101101110",
  65124=>"110100101",
  65125=>"100101111",
  65126=>"001101010",
  65127=>"011011011",
  65128=>"101000110",
  65129=>"010111011",
  65130=>"111111100",
  65131=>"001000110",
  65132=>"000111000",
  65133=>"101001001",
  65134=>"001110010",
  65135=>"000000110",
  65136=>"101110111",
  65137=>"110001110",
  65138=>"100011001",
  65139=>"101001101",
  65140=>"100111110",
  65141=>"011100101",
  65142=>"011001100",
  65143=>"001010001",
  65144=>"001110111",
  65145=>"100011011",
  65146=>"010100100",
  65147=>"111110101",
  65148=>"110011000",
  65149=>"001000000",
  65150=>"001001010",
  65151=>"000011101",
  65152=>"011110011",
  65153=>"111000011",
  65154=>"001100110",
  65155=>"101001001",
  65156=>"010100001",
  65157=>"010101110",
  65158=>"110111000",
  65159=>"101000101",
  65160=>"100001101",
  65161=>"001101100",
  65162=>"000101011",
  65163=>"101000010",
  65164=>"101100111",
  65165=>"110111011",
  65166=>"101010001",
  65167=>"110000000",
  65168=>"011000011",
  65169=>"111101001",
  65170=>"001000111",
  65171=>"111101101",
  65172=>"111101010",
  65173=>"100111100",
  65174=>"111110101",
  65175=>"001110100",
  65176=>"011111101",
  65177=>"011000100",
  65178=>"011101101",
  65179=>"100111000",
  65180=>"010111100",
  65181=>"000000110",
  65182=>"000001001",
  65183=>"001011001",
  65184=>"011101000",
  65185=>"110101010",
  65186=>"110111001",
  65187=>"011101100",
  65188=>"000111101",
  65189=>"000000111",
  65190=>"110111001",
  65191=>"010010100",
  65192=>"111001010",
  65193=>"000000000",
  65194=>"010010001",
  65195=>"111101001",
  65196=>"010001010",
  65197=>"110100000",
  65198=>"101000010",
  65199=>"101000000",
  65200=>"111110010",
  65201=>"100000110",
  65202=>"100000111",
  65203=>"111011111",
  65204=>"000100001",
  65205=>"001010100",
  65206=>"111101100",
  65207=>"001100110",
  65208=>"111000010",
  65209=>"101100111",
  65210=>"000100010",
  65211=>"110111000",
  65212=>"101000100",
  65213=>"110100100",
  65214=>"111011000",
  65215=>"000000011",
  65216=>"011011001",
  65217=>"110011100",
  65218=>"100111010",
  65219=>"010100001",
  65220=>"010010011",
  65221=>"100001110",
  65222=>"110000000",
  65223=>"001010010",
  65224=>"110010010",
  65225=>"101001000",
  65226=>"010101000",
  65227=>"100011101",
  65228=>"101100100",
  65229=>"101110010",
  65230=>"111010011",
  65231=>"000110111",
  65232=>"111000110",
  65233=>"011111011",
  65234=>"001000010",
  65235=>"001010010",
  65236=>"000100110",
  65237=>"001101001",
  65238=>"111111111",
  65239=>"000111010",
  65240=>"100100011",
  65241=>"100001000",
  65242=>"111101100",
  65243=>"110000011",
  65244=>"101001000",
  65245=>"111111110",
  65246=>"100100101",
  65247=>"100111000",
  65248=>"001000001",
  65249=>"110111111",
  65250=>"011010000",
  65251=>"000011110",
  65252=>"000001100",
  65253=>"010101110",
  65254=>"111111100",
  65255=>"110101110",
  65256=>"000010011",
  65257=>"111000100",
  65258=>"100010000",
  65259=>"001011001",
  65260=>"000001110",
  65261=>"000000101",
  65262=>"111010001",
  65263=>"000011111",
  65264=>"000101111",
  65265=>"101101100",
  65266=>"101110110",
  65267=>"101011010",
  65268=>"111010100",
  65269=>"000110100",
  65270=>"000010111",
  65271=>"101110100",
  65272=>"111101010",
  65273=>"001110100",
  65274=>"110110001",
  65275=>"100101011",
  65276=>"111110000",
  65277=>"110110111",
  65278=>"101001101",
  65279=>"001001010",
  65280=>"101010000",
  65281=>"111011101",
  65282=>"111110100",
  65283=>"000100000",
  65284=>"010010001",
  65285=>"101001011",
  65286=>"001110011",
  65287=>"110101100",
  65288=>"111100010",
  65289=>"101100100",
  65290=>"011101111",
  65291=>"010111100",
  65292=>"100100101",
  65293=>"111010100",
  65294=>"000100001",
  65295=>"011110111",
  65296=>"101000000",
  65297=>"100001100",
  65298=>"010110001",
  65299=>"111011101",
  65300=>"010110000",
  65301=>"001001111",
  65302=>"001011100",
  65303=>"001010001",
  65304=>"110110100",
  65305=>"010000100",
  65306=>"110010111",
  65307=>"001000010",
  65308=>"110100000",
  65309=>"001111111",
  65310=>"110011000",
  65311=>"101100001",
  65312=>"111110111",
  65313=>"101111101",
  65314=>"111111110",
  65315=>"011111101",
  65316=>"101100101",
  65317=>"111001110",
  65318=>"001111100",
  65319=>"100101100",
  65320=>"110101000",
  65321=>"011100100",
  65322=>"100111011",
  65323=>"101001010",
  65324=>"000010011",
  65325=>"000001000",
  65326=>"101100000",
  65327=>"010100011",
  65328=>"000010100",
  65329=>"000000011",
  65330=>"000011101",
  65331=>"100001011",
  65332=>"001110010",
  65333=>"110101110",
  65334=>"100101010",
  65335=>"000000001",
  65336=>"000110000",
  65337=>"100101011",
  65338=>"101101000",
  65339=>"000010110",
  65340=>"111001001",
  65341=>"001001000",
  65342=>"100001000",
  65343=>"110011111",
  65344=>"000010101",
  65345=>"100111111",
  65346=>"000001100",
  65347=>"110011000",
  65348=>"111111110",
  65349=>"001100110",
  65350=>"111000000",
  65351=>"110110011",
  65352=>"101111110",
  65353=>"101000001",
  65354=>"101101111",
  65355=>"100101001",
  65356=>"010011010",
  65357=>"001110101",
  65358=>"101111100",
  65359=>"110100101",
  65360=>"010111010",
  65361=>"100001100",
  65362=>"100100110",
  65363=>"100111000",
  65364=>"000110001",
  65365=>"111110011",
  65366=>"010010100",
  65367=>"011001011",
  65368=>"001001000",
  65369=>"011111101",
  65370=>"000111111",
  65371=>"101001010",
  65372=>"111111101",
  65373=>"001001000",
  65374=>"000110111",
  65375=>"101110111",
  65376=>"001110011",
  65377=>"010100101",
  65378=>"111001101",
  65379=>"010101110",
  65380=>"100100110",
  65381=>"010001010",
  65382=>"100110110",
  65383=>"111110100",
  65384=>"000111110",
  65385=>"111100001",
  65386=>"111100001",
  65387=>"000100011",
  65388=>"101100111",
  65389=>"101101110",
  65390=>"100110110",
  65391=>"110010011",
  65392=>"100000001",
  65393=>"000011010",
  65394=>"000111111",
  65395=>"001110001",
  65396=>"110010100",
  65397=>"111100101",
  65398=>"100011000",
  65399=>"010001001",
  65400=>"001010101",
  65401=>"011111001",
  65402=>"100011011",
  65403=>"010100101",
  65404=>"001001011",
  65405=>"011100001",
  65406=>"111100010",
  65407=>"001001010",
  65408=>"011101010",
  65409=>"010010100",
  65410=>"001110100",
  65411=>"001011001",
  65412=>"101001000",
  65413=>"000000010",
  65414=>"000101111",
  65415=>"001000011",
  65416=>"011111110",
  65417=>"000000101",
  65418=>"100011010",
  65419=>"101001110",
  65420=>"100010010",
  65421=>"110010101",
  65422=>"101101011",
  65423=>"111001000",
  65424=>"010110110",
  65425=>"110101010",
  65426=>"000000110",
  65427=>"101010000",
  65428=>"101101000",
  65429=>"100011010",
  65430=>"010000101",
  65431=>"010111111",
  65432=>"111010010",
  65433=>"101100001",
  65434=>"000000011",
  65435=>"010010010",
  65436=>"000000111",
  65437=>"001011011",
  65438=>"011011100",
  65439=>"000000100",
  65440=>"110000101",
  65441=>"001010110",
  65442=>"000101010",
  65443=>"110101101",
  65444=>"100010010",
  65445=>"010000101",
  65446=>"111110100",
  65447=>"101110101",
  65448=>"001110011",
  65449=>"111110111",
  65450=>"000000011",
  65451=>"010111010",
  65452=>"100010101",
  65453=>"010101101",
  65454=>"011010010",
  65455=>"000110101",
  65456=>"101001010",
  65457=>"011110100",
  65458=>"110010000",
  65459=>"000010011",
  65460=>"001001101",
  65461=>"111010011",
  65462=>"010101010",
  65463=>"010010101",
  65464=>"011110111",
  65465=>"101011101",
  65466=>"001110100",
  65467=>"101000000",
  65468=>"111001001",
  65469=>"100011101",
  65470=>"001011110",
  65471=>"011100111",
  65472=>"010011101",
  65473=>"000100110",
  65474=>"111101010",
  65475=>"111001100",
  65476=>"000001001",
  65477=>"111100111",
  65478=>"000010000",
  65479=>"011111010",
  65480=>"100110000",
  65481=>"100011101",
  65482=>"111001111",
  65483=>"100000110",
  65484=>"101011100",
  65485=>"111100110",
  65486=>"100000000",
  65487=>"110010100",
  65488=>"110001100",
  65489=>"001111111",
  65490=>"100100100",
  65491=>"010010000",
  65492=>"011001101",
  65493=>"111101101",
  65494=>"000001011",
  65495=>"101001101",
  65496=>"100001010",
  65497=>"110111110",
  65498=>"101111110",
  65499=>"011000100",
  65500=>"100100000",
  65501=>"001000010",
  65502=>"000001001",
  65503=>"101110000",
  65504=>"011001001",
  65505=>"110101100",
  65506=>"100010010",
  65507=>"011100011",
  65508=>"000110000",
  65509=>"001011101",
  65510=>"000010001",
  65511=>"100010000",
  65512=>"111111001",
  65513=>"101100011",
  65514=>"011101111",
  65515=>"010000000",
  65516=>"010100101",
  65517=>"101110101",
  65518=>"100110001",
  65519=>"011011111",
  65520=>"001100011",
  65521=>"100001100",
  65522=>"111110100",
  65523=>"011000001",
  65524=>"011000010",
  65525=>"011010000",
  65526=>"111111111",
  65527=>"111001101",
  65528=>"111011000",
  65529=>"000100011",
  65530=>"101101111",
  65531=>"000101101",
  65532=>"010001101",
  65533=>"101100010",
  65534=>"001100101",
  65535=>"100110001");

BEGIN
  weight <= ROM_content(to_integer(address));
END RTL;