LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.NUMERIC_STD.ALL;

LIBRARY work;
USE work.YOLO_pkg.ALL;

ENTITY L4_1_WROM IS
    PORT (
        weight : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
        address : IN unsigned(weightsbitsAddress(4)-1 DOWNTO 0));
END L4_1_WROM;

ARCHITECTURE RTL OF L4_1_WROM IS

    TYPE ROM_mem IS ARRAY (0 TO 4095) OF STD_LOGIC_VECTOR(8 DOWNTO 0);

    CONSTANT ROM_content : ROM_mem := (0=>"001001001",
    1=>"111000111",
    2=>"000000000",
    3=>"110100000",
    4=>"110110100",
    5=>"010010110",
    6=>"101001011",
    7=>"100000100",
    8=>"100110100",
    9=>"101101101",
    10=>"011011001",
    11=>"001000100",
    12=>"101101111",
    13=>"000110100",
    14=>"111000001",
    15=>"011001000",
    16=>"101111101",
    17=>"110110110",
    18=>"000000000",
    19=>"000100111",
    20=>"100100100",
    21=>"000001001",
    22=>"010111111",
    23=>"011011011",
    24=>"010111110",
    25=>"100101001",
    26=>"110110111",
    27=>"101000001",
    28=>"011011100",
    29=>"011110100",
    30=>"100100000",
    31=>"001110101",
    32=>"010010010",
    33=>"001011001",
    34=>"011000111",
    35=>"011001010",
    36=>"111100110",
    37=>"001001000",
    38=>"110110100",
    39=>"001001000",
    40=>"011111011",
    41=>"001001001",
    42=>"000100010",
    43=>"000001011",
    44=>"100100100",
    45=>"100000001",
    46=>"000111111",
    47=>"100010111",
    48=>"010110000",
    49=>"110000001",
    50=>"001000011",
    51=>"011110010",
    52=>"001001101",
    53=>"111100000",
    54=>"100100101",
    55=>"111000000",
    56=>"111001011",
    57=>"011001110",
    58=>"100000000",
    59=>"000110000",
    60=>"011011111",
    61=>"100000000",
    62=>"000000000",
    63=>"101001001",
    64=>"111111000",
    65=>"111111111",
    66=>"111111011",
    67=>"100000011",
    68=>"100101101",
    69=>"000000110",
    70=>"001111011",
    71=>"001110100",
    72=>"000000000",
    73=>"000111000",
    74=>"100110000",
    75=>"101111000",
    76=>"101111000",
    77=>"111111111",
    78=>"001101101",
    79=>"000000000",
    80=>"111010010",
    81=>"000000101",
    82=>"000000000",
    83=>"001001001",
    84=>"001000100",
    85=>"000000000",
    86=>"111101111",
    87=>"111000111",
    88=>"110111010",
    89=>"111111111",
    90=>"000000011",
    91=>"111101101",
    92=>"010011111",
    93=>"111111000",
    94=>"110110110",
    95=>"111000011",
    96=>"000000000",
    97=>"010000001",
    98=>"110110110",
    99=>"000000000",
    100=>"001000110",
    101=>"000011001",
    102=>"010000011",
    103=>"000000000",
    104=>"111111111",
    105=>"000000100",
    106=>"101100110",
    107=>"010000011",
    108=>"111111101",
    109=>"110101010",
    110=>"000010111",
    111=>"111111111",
    112=>"011000110",
    113=>"010000010",
    114=>"000000100",
    115=>"100111110",
    116=>"111101111",
    117=>"101101000",
    118=>"101101101",
    119=>"000111101",
    120=>"010000011",
    121=>"110001001",
    122=>"000000000",
    123=>"101111000",
    124=>"000000001",
    125=>"000000000",
    126=>"000000000",
    127=>"111000000",
    128=>"001001001",
    129=>"011111111",
    130=>"111111111",
    131=>"010111110",
    132=>"010110110",
    133=>"000000100",
    134=>"111111111",
    135=>"101101101",
    136=>"011001010",
    137=>"000010000",
    138=>"010011000",
    139=>"111001001",
    140=>"111111111",
    141=>"000000000",
    142=>"111100100",
    143=>"110111110",
    144=>"000000000",
    145=>"010111010",
    146=>"011001100",
    147=>"000000000",
    148=>"000000100",
    149=>"000101000",
    150=>"001000101",
    151=>"000000011",
    152=>"001000001",
    153=>"000110000",
    154=>"000000001",
    155=>"010101000",
    156=>"101000100",
    157=>"010111000",
    158=>"111111111",
    159=>"101101100",
    160=>"001000001",
    161=>"110110011",
    162=>"000000000",
    163=>"001000101",
    164=>"000000000",
    165=>"101101101",
    166=>"010110010",
    167=>"000010000",
    168=>"111111111",
    169=>"000000000",
    170=>"001100100",
    171=>"110110101",
    172=>"000100000",
    173=>"101001001",
    174=>"001001001",
    175=>"010110010",
    176=>"100100110",
    177=>"000000000",
    178=>"000000000",
    179=>"000000000",
    180=>"111111010",
    181=>"101001001",
    182=>"000000001",
    183=>"000101000",
    184=>"110011010",
    185=>"000001000",
    186=>"100101101",
    187=>"100101000",
    188=>"001000101",
    189=>"101000001",
    190=>"010010001",
    191=>"111010000",
    192=>"101011111",
    193=>"100110111",
    194=>"001111001",
    195=>"010110010",
    196=>"110010000",
    197=>"111110000",
    198=>"111001111",
    199=>"100111011",
    200=>"111011000",
    201=>"101101101",
    202=>"011110000",
    203=>"000110110",
    204=>"111111100",
    205=>"000000100",
    206=>"011001001",
    207=>"000110010",
    208=>"111000011",
    209=>"110111010",
    210=>"011111100",
    211=>"100010011",
    212=>"001000000",
    213=>"000000101",
    214=>"101001111",
    215=>"110110000",
    216=>"000000000",
    217=>"011000111",
    218=>"110000001",
    219=>"001001011",
    220=>"000111110",
    221=>"010000110",
    222=>"011110111",
    223=>"001000001",
    224=>"000001100",
    225=>"000110010",
    226=>"000100000",
    227=>"110000000",
    228=>"111101100",
    229=>"000111111",
    230=>"001011010",
    231=>"011111110",
    232=>"101101110",
    233=>"000000111",
    234=>"011000101",
    235=>"111000000",
    236=>"001101101",
    237=>"111111110",
    238=>"101001111",
    239=>"011001001",
    240=>"001000111",
    241=>"000100101",
    242=>"011111110",
    243=>"001001111",
    244=>"000000111",
    245=>"001000101",
    246=>"100010111",
    247=>"000110000",
    248=>"000001011",
    249=>"000100111",
    250=>"111111110",
    251=>"100000000",
    252=>"110110110",
    253=>"000010000",
    254=>"101111100",
    255=>"001000000",
    256=>"001001100",
    257=>"100000000",
    258=>"100100000",
    259=>"011001001",
    260=>"101111111",
    261=>"011001001",
    262=>"110110111",
    263=>"001001000",
    264=>"000000000",
    265=>"100100110",
    266=>"011001000",
    267=>"110110011",
    268=>"001001111",
    269=>"011000001",
    270=>"000010000",
    271=>"100110110",
    272=>"001001000",
    273=>"101101111",
    274=>"100011001",
    275=>"011110001",
    276=>"110011011",
    277=>"100110110",
    278=>"011011001",
    279=>"011001001",
    280=>"011001001",
    281=>"100100110",
    282=>"011001001",
    283=>"001101100",
    284=>"110001101",
    285=>"101100111",
    286=>"111010011",
    287=>"100100100",
    288=>"011011001",
    289=>"001101101",
    290=>"110011001",
    291=>"011001000",
    292=>"010011001",
    293=>"011011001",
    294=>"000101100",
    295=>"100001010",
    296=>"010010010",
    297=>"100100110",
    298=>"000110100",
    299=>"000001000",
    300=>"110010011",
    301=>"011011001",
    302=>"011011001",
    303=>"000010000",
    304=>"100111111",
    305=>"100110111",
    306=>"111011001",
    307=>"100000001",
    308=>"111001100",
    309=>"000001000",
    310=>"111111101",
    311=>"011001001",
    312=>"100010011",
    313=>"100110111",
    314=>"000011001",
    315=>"000011001",
    316=>"011011001",
    317=>"011011001",
    318=>"001110111",
    319=>"000000000",
    320=>"000100011",
    321=>"110000111",
    322=>"111101100",
    323=>"010101111",
    324=>"011000100",
    325=>"001100110",
    326=>"010110010",
    327=>"100101001",
    328=>"011111010",
    329=>"000111001",
    330=>"100000011",
    331=>"001111100",
    332=>"111111111",
    333=>"111111110",
    334=>"001111100",
    335=>"000000001",
    336=>"110010010",
    337=>"110000000",
    338=>"011011101",
    339=>"010000000",
    340=>"001000100",
    341=>"000000001",
    342=>"111000110",
    343=>"110000010",
    344=>"101001001",
    345=>"111010110",
    346=>"110001011",
    347=>"101000011",
    348=>"101101010",
    349=>"001000000",
    350=>"111111111",
    351=>"001000101",
    352=>"101101101",
    353=>"111000100",
    354=>"111000000",
    355=>"100000101",
    356=>"000000110",
    357=>"001101100",
    358=>"101000011",
    359=>"010000101",
    360=>"101111100",
    361=>"000111010",
    362=>"011010111",
    363=>"000000001",
    364=>"100111000",
    365=>"100001011",
    366=>"101101101",
    367=>"100110000",
    368=>"100101000",
    369=>"000000000",
    370=>"011011100",
    371=>"000110100",
    372=>"000110011",
    373=>"000100001",
    374=>"000011011",
    375=>"100000101",
    376=>"110100110",
    377=>"000111100",
    378=>"010110001",
    379=>"000101011",
    380=>"111000111",
    381=>"001001000",
    382=>"111101011",
    383=>"110000000",
    384=>"001001001",
    385=>"000000000",
    386=>"011111010",
    387=>"000110111",
    388=>"001011001",
    389=>"110100100",
    390=>"000000011",
    391=>"100000000",
    392=>"001011001",
    393=>"011111111",
    394=>"100110100",
    395=>"100100100",
    396=>"100111000",
    397=>"110111111",
    398=>"001001101",
    399=>"101111111",
    400=>"111011111",
    401=>"001001001",
    402=>"001000000",
    403=>"000001001",
    404=>"001001100",
    405=>"000010000",
    406=>"111101111",
    407=>"111100111",
    408=>"010011011",
    409=>"010010011",
    410=>"111001011",
    411=>"101101011",
    412=>"000000011",
    413=>"010000010",
    414=>"010000100",
    415=>"000101101",
    416=>"001001001",
    417=>"100110100",
    418=>"110100110",
    419=>"011001111",
    420=>"010111110",
    421=>"001000100",
    422=>"001011011",
    423=>"001000000",
    424=>"000101000",
    425=>"101100100",
    426=>"011001100",
    427=>"110100000",
    428=>"000000100",
    429=>"110110110",
    430=>"000101110",
    431=>"100100001",
    432=>"110110110",
    433=>"010010011",
    434=>"001001010",
    435=>"110110111",
    436=>"000101000",
    437=>"001001001",
    438=>"001100100",
    439=>"010010010",
    440=>"101000011",
    441=>"100100011",
    442=>"100100000",
    443=>"100100100",
    444=>"100100100",
    445=>"101100100",
    446=>"000010010",
    447=>"101001101",
    448=>"000000000",
    449=>"111111111",
    450=>"000000000",
    451=>"111111110",
    452=>"111111111",
    453=>"011100110",
    454=>"100001000",
    455=>"000111000",
    456=>"111111100",
    457=>"000111010",
    458=>"111101111",
    459=>"001001001",
    460=>"000111010",
    461=>"111111011",
    462=>"101000100",
    463=>"000001000",
    464=>"111011000",
    465=>"111111001",
    466=>"000000000",
    467=>"000000000",
    468=>"000000110",
    469=>"000000000",
    470=>"000000010",
    471=>"101111111",
    472=>"011011010",
    473=>"011010000",
    474=>"100110111",
    475=>"010000010",
    476=>"111101111",
    477=>"110111010",
    478=>"011001111",
    479=>"001001010",
    480=>"110000001",
    481=>"111111111",
    482=>"001010111",
    483=>"110110110",
    484=>"000110000",
    485=>"000001101",
    486=>"111111011",
    487=>"000000000",
    488=>"000000000",
    489=>"110110000",
    490=>"011111110",
    491=>"111110011",
    492=>"000000000",
    493=>"100000000",
    494=>"000000001",
    495=>"110000000",
    496=>"110000000",
    497=>"111111111",
    498=>"110000000",
    499=>"011010010",
    500=>"000111111",
    501=>"000000001",
    502=>"000000000",
    503=>"111101111",
    504=>"111011011",
    505=>"000100011",
    506=>"000000000",
    507=>"000000000",
    508=>"001000101",
    509=>"111111111",
    510=>"000000000",
    511=>"111001101",
    512=>"000100100",
    513=>"110100100",
    514=>"011011010",
    515=>"111111101",
    516=>"001001000",
    517=>"010010000",
    518=>"000100111",
    519=>"001001011",
    520=>"011011011",
    521=>"011011011",
    522=>"011011011",
    523=>"001001100",
    524=>"101101101",
    525=>"001110110",
    526=>"010011100",
    527=>"011011001",
    528=>"001110100",
    529=>"110110110",
    530=>"000010110",
    531=>"000000000",
    532=>"000001100",
    533=>"000100101",
    534=>"100100100",
    535=>"110100101",
    536=>"100100100",
    537=>"100100100",
    538=>"100101111",
    539=>"001011111",
    540=>"100110100",
    541=>"111001001",
    542=>"110110010",
    543=>"001001100",
    544=>"011011011",
    545=>"001001001",
    546=>"011011001",
    547=>"001000000",
    548=>"001011000",
    549=>"010001001",
    550=>"010011111",
    551=>"100110110",
    552=>"001011011",
    553=>"000010100",
    554=>"110110001",
    555=>"010110110",
    556=>"000100101",
    557=>"000111101",
    558=>"001001011",
    559=>"101100100",
    560=>"010101100",
    561=>"000000000",
    562=>"111111001",
    563=>"001000100",
    564=>"000100000",
    565=>"000001000",
    566=>"101011101",
    567=>"011011010",
    568=>"100100100",
    569=>"001001000",
    570=>"110100100",
    571=>"000001000",
    572=>"100100100",
    573=>"111100000",
    574=>"001001000",
    575=>"101001001",
    576=>"000100100",
    577=>"001001001",
    578=>"001000110",
    579=>"100110110",
    580=>"000011111",
    581=>"100100110",
    582=>"011011001",
    583=>"000110011",
    584=>"000111101",
    585=>"000100111",
    586=>"010111011",
    587=>"001000111",
    588=>"001101101",
    589=>"100010011",
    590=>"001001111",
    591=>"110111010",
    592=>"100010001",
    593=>"111011000",
    594=>"011001100",
    595=>"011011001",
    596=>"000000101",
    597=>"000011000",
    598=>"111011000",
    599=>"010011000",
    600=>"001001101",
    601=>"011001101",
    602=>"011011000",
    603=>"000011000",
    604=>"011010000",
    605=>"001000111",
    606=>"000100100",
    607=>"100000110",
    608=>"011010011",
    609=>"101101111",
    610=>"001000100",
    611=>"000000111",
    612=>"101110001",
    613=>"001000111",
    614=>"010011001",
    615=>"111001001",
    616=>"000100111",
    617=>"000000000",
    618=>"001101100",
    619=>"111001001",
    620=>"100010001",
    621=>"100110000",
    622=>"100110111",
    623=>"100010011",
    624=>"110010001",
    625=>"111011011",
    626=>"101001101",
    627=>"100011001",
    628=>"000011011",
    629=>"100111110",
    630=>"100100101",
    631=>"110011001",
    632=>"110011001",
    633=>"000110110",
    634=>"100111011",
    635=>"100110111",
    636=>"110011000",
    637=>"000011001",
    638=>"100110111",
    639=>"011011000",
    640=>"000100101",
    641=>"011010110",
    642=>"011101011",
    643=>"000101111",
    644=>"000110111",
    645=>"011000100",
    646=>"100000000",
    647=>"000110101",
    648=>"011001000",
    649=>"010110011",
    650=>"010010110",
    651=>"010000000",
    652=>"111110010",
    653=>"111000101",
    654=>"110000000",
    655=>"010111000",
    656=>"000000101",
    657=>"010110000",
    658=>"100110110",
    659=>"010101101",
    660=>"001000100",
    661=>"000000000",
    662=>"100000011",
    663=>"001100000",
    664=>"100100111",
    665=>"111000011",
    666=>"101001001",
    667=>"111100000",
    668=>"100000011",
    669=>"000010000",
    670=>"000000000",
    671=>"000000000",
    672=>"000000111",
    673=>"111011000",
    674=>"000111111",
    675=>"100000000",
    676=>"000000111",
    677=>"100100101",
    678=>"011010000",
    679=>"111111111",
    680=>"000111111",
    681=>"110000011",
    682=>"100111101",
    683=>"100000000",
    684=>"001100111",
    685=>"111010100",
    686=>"101000111",
    687=>"111100101",
    688=>"111111111",
    689=>"100100000",
    690=>"110100100",
    691=>"110111010",
    692=>"000000011",
    693=>"101001101",
    694=>"001100101",
    695=>"111111000",
    696=>"100001000",
    697=>"011001110",
    698=>"000001001",
    699=>"000000100",
    700=>"010100000",
    701=>"001010001",
    702=>"011111001",
    703=>"100100111",
    704=>"111001000",
    705=>"000100101",
    706=>"111000000",
    707=>"111110010",
    708=>"100110001",
    709=>"000110001",
    710=>"011000001",
    711=>"111001100",
    712=>"000100111",
    713=>"111011000",
    714=>"001011100",
    715=>"100111001",
    716=>"111101110",
    717=>"000101110",
    718=>"000110011",
    719=>"010000111",
    720=>"001100110",
    721=>"000110111",
    722=>"000000111",
    723=>"001000100",
    724=>"100011001",
    725=>"000110011",
    726=>"000110111",
    727=>"100110001",
    728=>"011101000",
    729=>"000110001",
    730=>"011100100",
    731=>"111011000",
    732=>"000000111",
    733=>"011100011",
    734=>"100111000",
    735=>"100110001",
    736=>"110001100",
    737=>"000110111",
    738=>"100111001",
    739=>"001000100",
    740=>"000110001",
    741=>"011000111",
    742=>"011001000",
    743=>"000100011",
    744=>"111001000",
    745=>"111010001",
    746=>"100111011",
    747=>"100100000",
    748=>"111000000",
    749=>"101100000",
    750=>"111001100",
    751=>"000010011",
    752=>"111100111",
    753=>"000000110",
    754=>"000100011",
    755=>"000110111",
    756=>"111110110",
    757=>"111010000",
    758=>"100110001",
    759=>"111011001",
    760=>"100110001",
    761=>"111001001",
    762=>"100011100",
    763=>"111000000",
    764=>"000110111",
    765=>"010011111",
    766=>"111111001",
    767=>"000100011",
    768=>"000000001",
    769=>"000000000",
    770=>"000000000",
    771=>"000111000",
    772=>"111111011",
    773=>"100011001",
    774=>"100001100",
    775=>"001011010",
    776=>"111111111",
    777=>"100010010",
    778=>"111111110",
    779=>"100011001",
    780=>"010111010",
    781=>"000000000",
    782=>"001111011",
    783=>"111111111",
    784=>"000000000",
    785=>"111111111",
    786=>"111101111",
    787=>"000011101",
    788=>"111101111",
    789=>"010011000",
    790=>"000000000",
    791=>"001001011",
    792=>"000000000",
    793=>"000000100",
    794=>"001111100",
    795=>"010011100",
    796=>"011011010",
    797=>"100001001",
    798=>"100000000",
    799=>"000000000",
    800=>"111111111",
    801=>"100110011",
    802=>"000000000",
    803=>"100000110",
    804=>"111111111",
    805=>"100110001",
    806=>"011111100",
    807=>"111111111",
    808=>"000000000",
    809=>"000000000",
    810=>"100011001",
    811=>"000000010",
    812=>"000000000",
    813=>"011010100",
    814=>"111111111",
    815=>"000000000",
    816=>"010111000",
    817=>"010111101",
    818=>"100010000",
    819=>"010100010",
    820=>"110110100",
    821=>"011011110",
    822=>"000000010",
    823=>"100101101",
    824=>"101011111",
    825=>"011110000",
    826=>"111101111",
    827=>"111011110",
    828=>"111111111",
    829=>"010000001",
    830=>"111110111",
    831=>"000111011",
    832=>"010111000",
    833=>"000010000",
    834=>"011010000",
    835=>"010111010",
    836=>"000111100",
    837=>"011111010",
    838=>"000111010",
    839=>"100111001",
    840=>"011011010",
    841=>"000111000",
    842=>"010011010",
    843=>"000011010",
    844=>"111111111",
    845=>"100001110",
    846=>"000111000",
    847=>"010111010",
    848=>"010010010",
    849=>"010011010",
    850=>"001011110",
    851=>"010110000",
    852=>"011111000",
    853=>"010010010",
    854=>"101001101",
    855=>"010111010",
    856=>"001000001",
    857=>"010011000",
    858=>"110111000",
    859=>"010011010",
    860=>"010010010",
    861=>"000000000",
    862=>"000111010",
    863=>"010111010",
    864=>"010111010",
    865=>"010110010",
    866=>"111011000",
    867=>"101100100",
    868=>"010111010",
    869=>"010111110",
    870=>"010110010",
    871=>"011010010",
    872=>"000111000",
    873=>"010111010",
    874=>"010011010",
    875=>"000000011",
    876=>"000111000",
    877=>"110111010",
    878=>"111101100",
    879=>"001111011",
    880=>"000111010",
    881=>"010011010",
    882=>"111111010",
    883=>"000011010",
    884=>"010011010",
    885=>"000110000",
    886=>"010111010",
    887=>"001100000",
    888=>"010010000",
    889=>"010111000",
    890=>"000011010",
    891=>"010110010",
    892=>"000101001",
    893=>"101101001",
    894=>"110010010",
    895=>"010000000",
    896=>"011111001",
    897=>"110110100",
    898=>"011011000",
    899=>"001011111",
    900=>"001001000",
    901=>"100100100",
    902=>"100110100",
    903=>"001011011",
    904=>"111111110",
    905=>"000101111",
    906=>"001011111",
    907=>"111100000",
    908=>"001001111",
    909=>"010000000",
    910=>"111100000",
    911=>"111011000",
    912=>"100100100",
    913=>"001001111",
    914=>"110111001",
    915=>"000100100",
    916=>"111100100",
    917=>"110100100",
    918=>"100001111",
    919=>"100100100",
    920=>"101100001",
    921=>"001001011",
    922=>"000010110",
    923=>"000100111",
    924=>"110100100",
    925=>"001001011",
    926=>"110110100",
    927=>"110100000",
    928=>"100000010",
    929=>"011000000",
    930=>"000100000",
    931=>"011000001",
    932=>"000010100",
    933=>"111011001",
    934=>"110001111",
    935=>"110110000",
    936=>"011110100",
    937=>"110110100",
    938=>"010100001",
    939=>"001110110",
    940=>"111000100",
    941=>"000110110",
    942=>"011001011",
    943=>"000000000",
    944=>"001001011",
    945=>"110100000",
    946=>"110100100",
    947=>"000100000",
    948=>"100100100",
    949=>"000001001",
    950=>"011111100",
    951=>"111011110",
    952=>"100100110",
    953=>"101101001",
    954=>"101011000",
    955=>"011011011",
    956=>"111001110",
    957=>"101001011",
    958=>"001110110",
    959=>"110110000",
    960=>"100000000",
    961=>"101101101",
    962=>"011101011",
    963=>"001111100",
    964=>"000000000",
    965=>"010100001",
    966=>"111111011",
    967=>"000000000",
    968=>"111000001",
    969=>"111111001",
    970=>"001111111",
    971=>"100000001",
    972=>"111101101",
    973=>"110111111",
    974=>"100000000",
    975=>"000000010",
    976=>"000101011",
    977=>"000111100",
    978=>"000000000",
    979=>"011101111",
    980=>"000000000",
    981=>"110000001",
    982=>"100111111",
    983=>"011111111",
    984=>"110100001",
    985=>"110100011",
    986=>"001111110",
    987=>"101111111",
    988=>"101101111",
    989=>"001111110",
    990=>"110100001",
    991=>"110000001",
    992=>"111001001",
    993=>"010000001",
    994=>"100000001",
    995=>"000000001",
    996=>"001001001",
    997=>"100000000",
    998=>"101111111",
    999=>"110100111",
    1000=>"110000011",
    1001=>"110000000",
    1002=>"100000101",
    1003=>"011110101",
    1004=>"100000000",
    1005=>"101110101",
    1006=>"100000001",
    1007=>"010011111",
    1008=>"000001110",
    1009=>"100001110",
    1010=>"000000000",
    1011=>"111111111",
    1012=>"100111111",
    1013=>"110000001",
    1014=>"111000011",
    1015=>"110000000",
    1016=>"110111111",
    1017=>"000000101",
    1018=>"000000001",
    1019=>"111111011",
    1020=>"000000000",
    1021=>"000000001",
    1022=>"111010100",
    1023=>"101000001",
    1024=>"000110110",
    1025=>"010000000",
    1026=>"111111111",
    1027=>"111111010",
    1028=>"000100110",
    1029=>"110111111",
    1030=>"000000000",
    1031=>"000000000",
    1032=>"111100110",
    1033=>"111110010",
    1034=>"111111010",
    1035=>"100111111",
    1036=>"110111010",
    1037=>"010000110",
    1038=>"001000110",
    1039=>"000000000",
    1040=>"001111011",
    1041=>"000111011",
    1042=>"011000000",
    1043=>"000000000",
    1044=>"011100110",
    1045=>"000000000",
    1046=>"101001011",
    1047=>"011001011",
    1048=>"011101111",
    1049=>"000111011",
    1050=>"000000000",
    1051=>"010001000",
    1052=>"001011001",
    1053=>"100010000",
    1054=>"111111111",
    1055=>"111111011",
    1056=>"011001000",
    1057=>"001001000",
    1058=>"010011111",
    1059=>"000000100",
    1060=>"111101111",
    1061=>"111111111",
    1062=>"010111111",
    1063=>"001000000",
    1064=>"001111101",
    1065=>"000000000",
    1066=>"110111101",
    1067=>"000000001",
    1068=>"000000100",
    1069=>"000010000",
    1070=>"111001100",
    1071=>"111111111",
    1072=>"000000101",
    1073=>"000001001",
    1074=>"111111011",
    1075=>"000000011",
    1076=>"000100000",
    1077=>"000000111",
    1078=>"010010001",
    1079=>"011000100",
    1080=>"001001000",
    1081=>"010111010",
    1082=>"000100101",
    1083=>"011101100",
    1084=>"001000000",
    1085=>"111111111",
    1086=>"000000000",
    1087=>"000110111",
    1088=>"111011000",
    1089=>"000001100",
    1090=>"011111111",
    1091=>"000000101",
    1092=>"000010110",
    1093=>"110011000",
    1094=>"101001011",
    1095=>"010010110",
    1096=>"000011011",
    1097=>"101001000",
    1098=>"010000000",
    1099=>"010011001",
    1100=>"111111110",
    1101=>"000100110",
    1102=>"000100110",
    1103=>"000000001",
    1104=>"100110010",
    1105=>"000000000",
    1106=>"101101101",
    1107=>"010110000",
    1108=>"111101111",
    1109=>"000000000",
    1110=>"111101010",
    1111=>"001111011",
    1112=>"000110111",
    1113=>"000000010",
    1114=>"111110011",
    1115=>"001000111",
    1116=>"101000000",
    1117=>"110110010",
    1118=>"001101011",
    1119=>"001101111",
    1120=>"110110010",
    1121=>"000011010",
    1122=>"111111111",
    1123=>"010110000",
    1124=>"111110000",
    1125=>"110110110",
    1126=>"000010000",
    1127=>"011000110",
    1128=>"101101111",
    1129=>"000000000",
    1130=>"110011000",
    1131=>"001101001",
    1132=>"100111011",
    1133=>"110110100",
    1134=>"010010010",
    1135=>"001001111",
    1136=>"100100000",
    1137=>"000000011",
    1138=>"100111111",
    1139=>"111111011",
    1140=>"111111111",
    1141=>"110001011",
    1142=>"100100110",
    1143=>"000000000",
    1144=>"111011000",
    1145=>"001100000",
    1146=>"111101101",
    1147=>"011101111",
    1148=>"010110010",
    1149=>"100100001",
    1150=>"000100001",
    1151=>"111000001",
    1152=>"111000000",
    1153=>"100001111",
    1154=>"111111101",
    1155=>"011011011",
    1156=>"010000000",
    1157=>"110011001",
    1158=>"111111101",
    1159=>"000010110",
    1160=>"110110011",
    1161=>"100001111",
    1162=>"000011011",
    1163=>"011011111",
    1164=>"101101100",
    1165=>"111001101",
    1166=>"011011011",
    1167=>"001101100",
    1168=>"010000001",
    1169=>"111101111",
    1170=>"000010001",
    1171=>"001011011",
    1172=>"011001001",
    1173=>"001001000",
    1174=>"100100100",
    1175=>"100110001",
    1176=>"100100110",
    1177=>"001011111",
    1178=>"111101110",
    1179=>"011011000",
    1180=>"000110000",
    1181=>"100100000",
    1182=>"110001001",
    1183=>"110000010",
    1184=>"100110100",
    1185=>"111111011",
    1186=>"001100110",
    1187=>"110110000",
    1188=>"100100000",
    1189=>"110110110",
    1190=>"100100010",
    1191=>"011010100",
    1192=>"000001000",
    1193=>"111011011",
    1194=>"011011011",
    1195=>"000100110",
    1196=>"000011011",
    1197=>"000000000",
    1198=>"001100110",
    1199=>"001101111",
    1200=>"100100010",
    1201=>"010011001",
    1202=>"100100110",
    1203=>"111110111",
    1204=>"110110011",
    1205=>"111111111",
    1206=>"011000000",
    1207=>"011000000",
    1208=>"001001110",
    1209=>"001011000",
    1210=>"000000000",
    1211=>"000000000",
    1212=>"000100100",
    1213=>"100100000",
    1214=>"011011010",
    1215=>"001001001",
    1216=>"110100100",
    1217=>"011011111",
    1218=>"000011111",
    1219=>"110100100",
    1220=>"010100100",
    1221=>"001001000",
    1222=>"011111110",
    1223=>"110110100",
    1224=>"000010000",
    1225=>"001011011",
    1226=>"110110111",
    1227=>"100001100",
    1228=>"101100101",
    1229=>"111010000",
    1230=>"000000110",
    1231=>"001011111",
    1232=>"111110000",
    1233=>"001011011",
    1234=>"000000100",
    1235=>"101100100",
    1236=>"100000000",
    1237=>"000001001",
    1238=>"111110100",
    1239=>"111001000",
    1240=>"111100000",
    1241=>"001011111",
    1242=>"110100000",
    1243=>"111111110",
    1244=>"010100001",
    1245=>"001011011",
    1246=>"010011011",
    1247=>"000100001",
    1248=>"110100100",
    1249=>"000011001",
    1250=>"001001000",
    1251=>"110100000",
    1252=>"001001001",
    1253=>"001100110",
    1254=>"011110100",
    1255=>"000001101",
    1256=>"000010111",
    1257=>"000011011",
    1258=>"000001001",
    1259=>"001010000",
    1260=>"100110110",
    1261=>"110110100",
    1262=>"110100100",
    1263=>"111111111",
    1264=>"111011001",
    1265=>"001010011",
    1266=>"101000100",
    1267=>"111100101",
    1268=>"001001101",
    1269=>"110110100",
    1270=>"100000000",
    1271=>"111100100",
    1272=>"011111000",
    1273=>"000111111",
    1274=>"111100100",
    1275=>"110100100",
    1276=>"111100000",
    1277=>"100000000",
    1278=>"000010101",
    1279=>"110100100",
    1280=>"100100011",
    1281=>"111011111",
    1282=>"010111001",
    1283=>"000000000",
    1284=>"001011000",
    1285=>"111111111",
    1286=>"011011011",
    1287=>"001000111",
    1288=>"000001000",
    1289=>"101001001",
    1290=>"110110010",
    1291=>"101000000",
    1292=>"000000011",
    1293=>"001011000",
    1294=>"111000100",
    1295=>"111011111",
    1296=>"000000111",
    1297=>"101000000",
    1298=>"011000100",
    1299=>"111011111",
    1300=>"001100100",
    1301=>"100000000",
    1302=>"000000000",
    1303=>"111100001",
    1304=>"000000000",
    1305=>"111011000",
    1306=>"011011001",
    1307=>"101100100",
    1308=>"011010000",
    1309=>"111111111",
    1310=>"111001111",
    1311=>"111110000",
    1312=>"100111011",
    1313=>"000010010",
    1314=>"111111000",
    1315=>"010001111",
    1316=>"101100010",
    1317=>"010011111",
    1318=>"011110101",
    1319=>"111111100",
    1320=>"101111111",
    1321=>"100000000",
    1322=>"111001111",
    1323=>"111111101",
    1324=>"101001111",
    1325=>"110000000",
    1326=>"000000001",
    1327=>"101111011",
    1328=>"100000000",
    1329=>"111011000",
    1330=>"000000001",
    1331=>"010110010",
    1332=>"000000000",
    1333=>"110100001",
    1334=>"110111111",
    1335=>"000111111",
    1336=>"110000000",
    1337=>"111001100",
    1338=>"100000000",
    1339=>"110100001",
    1340=>"001010010",
    1341=>"000101001",
    1342=>"111100101",
    1343=>"110100100",
    1344=>"000010010",
    1345=>"000000000",
    1346=>"001100100",
    1347=>"111101111",
    1348=>"100110100",
    1349=>"011010110",
    1350=>"000000000",
    1351=>"100100101",
    1352=>"000111110",
    1353=>"001101111",
    1354=>"100101011",
    1355=>"001111110",
    1356=>"000111111",
    1357=>"001111000",
    1358=>"000001101",
    1359=>"110101101",
    1360=>"111111000",
    1361=>"111000010",
    1362=>"000010010",
    1363=>"100000010",
    1364=>"010111000",
    1365=>"111111111",
    1366=>"111111111",
    1367=>"011111000",
    1368=>"111111110",
    1369=>"110101111",
    1370=>"110111011",
    1371=>"110100010",
    1372=>"010010010",
    1373=>"001101101",
    1374=>"010000010",
    1375=>"111111110",
    1376=>"011111011",
    1377=>"011011000",
    1378=>"000111010",
    1379=>"100010000",
    1380=>"000000000",
    1381=>"001111111",
    1382=>"110110000",
    1383=>"010110000",
    1384=>"011011101",
    1385=>"000000000",
    1386=>"000010001",
    1387=>"110001000",
    1388=>"100000000",
    1389=>"110000000",
    1390=>"111111111",
    1391=>"110110110",
    1392=>"011110110",
    1393=>"000101111",
    1394=>"011011011",
    1395=>"110111100",
    1396=>"110000000",
    1397=>"100111010",
    1398=>"011011001",
    1399=>"111111111",
    1400=>"100000010",
    1401=>"000110100",
    1402=>"010110100",
    1403=>"010110000",
    1404=>"110111010",
    1405=>"101000000",
    1406=>"100000010",
    1407=>"011111111",
    1408=>"000100001",
    1409=>"000000000",
    1410=>"000001100",
    1411=>"101101101",
    1412=>"000000000",
    1413=>"110111111",
    1414=>"101111111",
    1415=>"111111001",
    1416=>"000000101",
    1417=>"010111011",
    1418=>"000000000",
    1419=>"011111100",
    1420=>"000111011",
    1421=>"111111111",
    1422=>"000101100",
    1423=>"011010011",
    1424=>"111111110",
    1425=>"111110010",
    1426=>"111110101",
    1427=>"000010001",
    1428=>"111100100",
    1429=>"000100000",
    1430=>"000000010",
    1431=>"010000111",
    1432=>"000111000",
    1433=>"100111000",
    1434=>"111111111",
    1435=>"110001111",
    1436=>"111111110",
    1437=>"001111111",
    1438=>"000101010",
    1439=>"000000010",
    1440=>"011111111",
    1441=>"000000000",
    1442=>"111010000",
    1443=>"001000100",
    1444=>"010000111",
    1445=>"010111101",
    1446=>"000000000",
    1447=>"011101111",
    1448=>"101101000",
    1449=>"111111111",
    1450=>"011011001",
    1451=>"110000101",
    1452=>"000100110",
    1453=>"010101111",
    1454=>"110111111",
    1455=>"111111000",
    1456=>"000000000",
    1457=>"001000000",
    1458=>"111011000",
    1459=>"000010100",
    1460=>"111101101",
    1461=>"000001000",
    1462=>"111111011",
    1463=>"111111111",
    1464=>"110010010",
    1465=>"111101100",
    1466=>"111011111",
    1467=>"111111001",
    1468=>"000011011",
    1469=>"100000000",
    1470=>"001011001",
    1471=>"000000000",
    1472=>"111000000",
    1473=>"110000011",
    1474=>"111000000",
    1475=>"111000000",
    1476=>"111110000",
    1477=>"110111000",
    1478=>"111010000",
    1479=>"000000111",
    1480=>"111010101",
    1481=>"000001111",
    1482=>"111000001",
    1483=>"111100000",
    1484=>"111001111",
    1485=>"011111001",
    1486=>"111000000",
    1487=>"111000111",
    1488=>"111101001",
    1489=>"000111111",
    1490=>"110100000",
    1491=>"110001001",
    1492=>"001100100",
    1493=>"111000000",
    1494=>"001111111",
    1495=>"000010010",
    1496=>"001001111",
    1497=>"001111111",
    1498=>"001111110",
    1499=>"010001000",
    1500=>"011010100",
    1501=>"000111111",
    1502=>"111011000",
    1503=>"011010101",
    1504=>"110000001",
    1505=>"111000100",
    1506=>"111010010",
    1507=>"001100111",
    1508=>"011110100",
    1509=>"110000000",
    1510=>"001001010",
    1511=>"111010000",
    1512=>"111000000",
    1513=>"011000000",
    1514=>"111100100",
    1515=>"000011011",
    1516=>"011000000",
    1517=>"111011000",
    1518=>"100000111",
    1519=>"000000010",
    1520=>"100000111",
    1521=>"100000010",
    1522=>"100000001",
    1523=>"111010000",
    1524=>"111001000",
    1525=>"111011000",
    1526=>"111000000",
    1527=>"010000000",
    1528=>"000111011",
    1529=>"011000001",
    1530=>"011001000",
    1531=>"111001000",
    1532=>"001111110",
    1533=>"000000011",
    1534=>"111000000",
    1535=>"110111001",
    1536=>"101111110",
    1537=>"110111100",
    1538=>"000000000",
    1539=>"110110100",
    1540=>"000011111",
    1541=>"101101000",
    1542=>"100110010",
    1543=>"000011111",
    1544=>"011000000",
    1545=>"000110110",
    1546=>"111110110",
    1547=>"000000010",
    1548=>"101111111",
    1549=>"100100000",
    1550=>"000000001",
    1551=>"110100111",
    1552=>"100001110",
    1553=>"001101000",
    1554=>"010110110",
    1555=>"010011110",
    1556=>"000000000",
    1557=>"000010000",
    1558=>"011001001",
    1559=>"000001100",
    1560=>"000011011",
    1561=>"011110110",
    1562=>"001001000",
    1563=>"001011001",
    1564=>"000001001",
    1565=>"100100110",
    1566=>"001110111",
    1567=>"001011011",
    1568=>"000011001",
    1569=>"001001011",
    1570=>"111011011",
    1571=>"001001001",
    1572=>"111111011",
    1573=>"000111011",
    1574=>"011001000",
    1575=>"000101011",
    1576=>"111111110",
    1577=>"100100100",
    1578=>"110111110",
    1579=>"100101001",
    1580=>"110011111",
    1581=>"011011111",
    1582=>"000001001",
    1583=>"110110100",
    1584=>"001001011",
    1585=>"001100100",
    1586=>"000100111",
    1587=>"111111101",
    1588=>"001100100",
    1589=>"000000000",
    1590=>"111111011",
    1591=>"001001000",
    1592=>"100100001",
    1593=>"010000000",
    1594=>"001011011",
    1595=>"111111011",
    1596=>"001011011",
    1597=>"100001001",
    1598=>"001001010",
    1599=>"110110110",
    1600=>"001010110",
    1601=>"110010001",
    1602=>"111110000",
    1603=>"110101011",
    1604=>"101000000",
    1605=>"110100001",
    1606=>"101011100",
    1607=>"101001010",
    1608=>"111100000",
    1609=>"100100001",
    1610=>"000001111",
    1611=>"111100000",
    1612=>"101111101",
    1613=>"000110000",
    1614=>"100001000",
    1615=>"001011111",
    1616=>"100101001",
    1617=>"000011111",
    1618=>"001111001",
    1619=>"001011110",
    1620=>"110110000",
    1621=>"000001010",
    1622=>"010011110",
    1623=>"001011110",
    1624=>"110100000",
    1625=>"001011100",
    1626=>"001011110",
    1627=>"001110100",
    1628=>"001001011",
    1629=>"110100000",
    1630=>"110100110",
    1631=>"001011110",
    1632=>"011110101",
    1633=>"110010000",
    1634=>"100110100",
    1635=>"000000001",
    1636=>"000010111",
    1637=>"111110000",
    1638=>"000001011",
    1639=>"010111100",
    1640=>"111100000",
    1641=>"100001110",
    1642=>"001110100",
    1643=>"010101110",
    1644=>"101001000",
    1645=>"001011110",
    1646=>"111100001",
    1647=>"101101110",
    1648=>"111110000",
    1649=>"001010100",
    1650=>"011110001",
    1651=>"100010100",
    1652=>"100001101",
    1653=>"001010110",
    1654=>"001011110",
    1655=>"111110100",
    1656=>"001011110",
    1657=>"011111100",
    1658=>"011011010",
    1659=>"001011110",
    1660=>"001011111",
    1661=>"111100001",
    1662=>"001010110",
    1663=>"000001111",
    1664=>"011001001",
    1665=>"110111111",
    1666=>"001001001",
    1667=>"001001101",
    1668=>"001001001",
    1669=>"011000100",
    1670=>"101001011",
    1671=>"000000000",
    1672=>"011001101",
    1673=>"110110110",
    1674=>"101001001",
    1675=>"011001001",
    1676=>"101101100",
    1677=>"100110011",
    1678=>"011001001",
    1679=>"101000010",
    1680=>"100000000",
    1681=>"110110110",
    1682=>"011001001",
    1683=>"001011111",
    1684=>"001001000",
    1685=>"001001001",
    1686=>"110110110",
    1687=>"101100110",
    1688=>"110110010",
    1689=>"000100000",
    1690=>"110110110",
    1691=>"001111011",
    1692=>"001101001",
    1693=>"110110110",
    1694=>"001001001",
    1695=>"001001001",
    1696=>"001001001",
    1697=>"011001001",
    1698=>"111100010",
    1699=>"110110110",
    1700=>"011000100",
    1701=>"000001001",
    1702=>"100111011",
    1703=>"011001000",
    1704=>"001001001",
    1705=>"100100100",
    1706=>"111001001",
    1707=>"110110110",
    1708=>"001001001",
    1709=>"001001011",
    1710=>"011001001",
    1711=>"001001001",
    1712=>"111111110",
    1713=>"100101111",
    1714=>"010011011",
    1715=>"001001011",
    1716=>"001001001",
    1717=>"011001001",
    1718=>"001001001",
    1719=>"101101101",
    1720=>"100100110",
    1721=>"011011000",
    1722=>"001000000",
    1723=>"001001011",
    1724=>"001000000",
    1725=>"100100100",
    1726=>"001001011",
    1727=>"001001101",
    1728=>"000111011",
    1729=>"001001001",
    1730=>"111001000",
    1731=>"101000111",
    1732=>"111011011",
    1733=>"111001100",
    1734=>"101100100",
    1735=>"100111011",
    1736=>"110011001",
    1737=>"111010000",
    1738=>"000010111",
    1739=>"111001000",
    1740=>"111110010",
    1741=>"000110001",
    1742=>"010011001",
    1743=>"100100111",
    1744=>"000001000",
    1745=>"001100111",
    1746=>"011000000",
    1747=>"001100100",
    1748=>"010001000",
    1749=>"110000000",
    1750=>"001001111",
    1751=>"101100100",
    1752=>"111001000",
    1753=>"001100111",
    1754=>"100110111",
    1755=>"110100011",
    1756=>"111100100",
    1757=>"011001001",
    1758=>"010001101",
    1759=>"101100000",
    1760=>"110110010",
    1761=>"011100110",
    1762=>"010101000",
    1763=>"111001100",
    1764=>"110111110",
    1765=>"111001000",
    1766=>"000100000",
    1767=>"100100000",
    1768=>"111011001",
    1769=>"000100111",
    1770=>"011001000",
    1771=>"001000100",
    1772=>"011001000",
    1773=>"100110111",
    1774=>"111011011",
    1775=>"011000000",
    1776=>"001101101",
    1777=>"101100101",
    1778=>"011011000",
    1779=>"000000001",
    1780=>"100100110",
    1781=>"000111011",
    1782=>"100110011",
    1783=>"100100010",
    1784=>"001100110",
    1785=>"011111101",
    1786=>"000110011",
    1787=>"110111111",
    1788=>"001100111",
    1789=>"001000000",
    1790=>"100111111",
    1791=>"010010000",
    1792=>"100100101",
    1793=>"100111111",
    1794=>"001011011",
    1795=>"101101101",
    1796=>"000101110",
    1797=>"011100011",
    1798=>"000000010",
    1799=>"110000100",
    1800=>"001011011",
    1801=>"000001000",
    1802=>"010110111",
    1803=>"001000010",
    1804=>"111100111",
    1805=>"010011111",
    1806=>"110000100",
    1807=>"000000000",
    1808=>"111000000",
    1809=>"111100000",
    1810=>"100000000",
    1811=>"111011011",
    1812=>"111100110",
    1813=>"101011011",
    1814=>"011101111",
    1815=>"000010011",
    1816=>"000000000",
    1817=>"011010000",
    1818=>"111100011",
    1819=>"101000001",
    1820=>"011011010",
    1821=>"000001011",
    1822=>"100000000",
    1823=>"011001000",
    1824=>"111000111",
    1825=>"001000010",
    1826=>"111010010",
    1827=>"001100010",
    1828=>"111111110",
    1829=>"111001000",
    1830=>"011011011",
    1831=>"000101100",
    1832=>"000011000",
    1833=>"111100100",
    1834=>"111000100",
    1835=>"000100001",
    1836=>"101100100",
    1837=>"010011000",
    1838=>"111100101",
    1839=>"110110100",
    1840=>"010011010",
    1841=>"000011000",
    1842=>"111101100",
    1843=>"111110101",
    1844=>"000011001",
    1845=>"001001001",
    1846=>"101101100",
    1847=>"100100011",
    1848=>"111100111",
    1849=>"100001101",
    1850=>"110100000",
    1851=>"011100000",
    1852=>"111100100",
    1853=>"011100101",
    1854=>"100100101",
    1855=>"100000000",
    1856=>"000000010",
    1857=>"001001000",
    1858=>"110110110",
    1859=>"110100110",
    1860=>"100100100",
    1861=>"001001001",
    1862=>"000100000",
    1863=>"110000000",
    1864=>"110000100",
    1865=>"110100000",
    1866=>"110100100",
    1867=>"000000000",
    1868=>"101111001",
    1869=>"000100001",
    1870=>"110111111",
    1871=>"011101100",
    1872=>"001101000",
    1873=>"101101101",
    1874=>"000111011",
    1875=>"111010100",
    1876=>"101101110",
    1877=>"110110100",
    1878=>"011011111",
    1879=>"100000001",
    1880=>"001001011",
    1881=>"110100000",
    1882=>"001001000",
    1883=>"111110110",
    1884=>"110100100",
    1885=>"101001111",
    1886=>"111100010",
    1887=>"110100100",
    1888=>"001011011",
    1889=>"100110110",
    1890=>"111101001",
    1891=>"001001001",
    1892=>"000000000",
    1893=>"100100100",
    1894=>"110101001",
    1895=>"100110000",
    1896=>"000010010",
    1897=>"100100100",
    1898=>"101011011",
    1899=>"011111100",
    1900=>"100000100",
    1901=>"111100110",
    1902=>"001011111",
    1903=>"000001000",
    1904=>"111100100",
    1905=>"000001000",
    1906=>"001111111",
    1907=>"000000000",
    1908=>"000001011",
    1909=>"110110001",
    1910=>"111111110",
    1911=>"001001001",
    1912=>"011110100",
    1913=>"000000000",
    1914=>"101001101",
    1915=>"000000000",
    1916=>"001001111",
    1917=>"001011011",
    1918=>"110110110",
    1919=>"011011011",
    1920=>"001101010",
    1921=>"000100111",
    1922=>"111111110",
    1923=>"100111000",
    1924=>"000000101",
    1925=>"100001011",
    1926=>"000100110",
    1927=>"001001110",
    1928=>"111111001",
    1929=>"011010000",
    1930=>"100100110",
    1931=>"011110010",
    1932=>"101101100",
    1933=>"101100000",
    1934=>"000111001",
    1935=>"101001001",
    1936=>"101100100",
    1937=>"111011001",
    1938=>"000000001",
    1939=>"100110101",
    1940=>"111110101",
    1941=>"000000100",
    1942=>"100001100",
    1943=>"100100100",
    1944=>"001000100",
    1945=>"011001011",
    1946=>"100100100",
    1947=>"000100100",
    1948=>"000100110",
    1949=>"011011001",
    1950=>"100100110",
    1951=>"000100100",
    1952=>"100100100",
    1953=>"110111111",
    1954=>"001000000",
    1955=>"001000000",
    1956=>"000110001",
    1957=>"000011011",
    1958=>"100100110",
    1959=>"100110000",
    1960=>"101010111",
    1961=>"101111111",
    1962=>"100110000",
    1963=>"001100100",
    1964=>"011011010",
    1965=>"000100101",
    1966=>"100011110",
    1967=>"100100100",
    1968=>"001101001",
    1969=>"100001001",
    1970=>"100110011",
    1971=>"101111111",
    1972=>"100101101",
    1973=>"000111111",
    1974=>"000110011",
    1975=>"000100100",
    1976=>"100100100",
    1977=>"100101101",
    1978=>"100110111",
    1979=>"000000100",
    1980=>"010001100",
    1981=>"001100001",
    1982=>"100100110",
    1983=>"000000000",
    1984=>"110111111",
    1985=>"000111010",
    1986=>"000111000",
    1987=>"011010000",
    1988=>"000111111",
    1989=>"000000000",
    1990=>"000111000",
    1991=>"100100111",
    1992=>"000111111",
    1993=>"011101000",
    1994=>"000111111",
    1995=>"100000110",
    1996=>"000100111",
    1997=>"000011111",
    1998=>"011101101",
    1999=>"111000000",
    2000=>"000000000",
    2001=>"000000110",
    2002=>"001000000",
    2003=>"111000000",
    2004=>"000000100",
    2005=>"111100000",
    2006=>"111111111",
    2007=>"010000000",
    2008=>"000010000",
    2009=>"110000110",
    2010=>"100100000",
    2011=>"000011111",
    2012=>"111010000",
    2013=>"111001001",
    2014=>"000011000",
    2015=>"111010000",
    2016=>"000000000",
    2017=>"111000000",
    2018=>"011111100",
    2019=>"000000111",
    2020=>"111100111",
    2021=>"000000011",
    2022=>"111011000",
    2023=>"010101000",
    2024=>"100000000",
    2025=>"100000111",
    2026=>"100100001",
    2027=>"000010111",
    2028=>"101111111",
    2029=>"000100000",
    2030=>"111111000",
    2031=>"000000010",
    2032=>"000010111",
    2033=>"000111010",
    2034=>"011000000",
    2035=>"100010000",
    2036=>"000011011",
    2037=>"110001000",
    2038=>"001111111",
    2039=>"110111101",
    2040=>"000010010",
    2041=>"000101111",
    2042=>"010000010",
    2043=>"011010000",
    2044=>"000000000",
    2045=>"110000000",
    2046=>"110011000",
    2047=>"111000000",
    2048=>"100100100",
    2049=>"000010011",
    2050=>"001011111",
    2051=>"011000010",
    2052=>"011100000",
    2053=>"011100010",
    2054=>"001001011",
    2055=>"110110100",
    2056=>"011001000",
    2057=>"111101101",
    2058=>"110000110",
    2059=>"011001101",
    2060=>"111101000",
    2061=>"001001111",
    2062=>"011101101",
    2063=>"111000000",
    2064=>"111000100",
    2065=>"101000111",
    2066=>"011011001",
    2067=>"011001001",
    2068=>"001001000",
    2069=>"010000001",
    2070=>"001010111",
    2071=>"110100010",
    2072=>"000011011",
    2073=>"000111111",
    2074=>"110111010",
    2075=>"110000110",
    2076=>"001000001",
    2077=>"001011011",
    2078=>"100100110",
    2079=>"011000000",
    2080=>"111111000",
    2081=>"001001100",
    2082=>"000100010",
    2083=>"000100010",
    2084=>"110110100",
    2085=>"011011001",
    2086=>"100100101",
    2087=>"011011001",
    2088=>"100110101",
    2089=>"010100000",
    2090=>"011011001",
    2091=>"101000011",
    2092=>"001001001",
    2093=>"100100100",
    2094=>"111101000",
    2095=>"000001011",
    2096=>"111000001",
    2097=>"001101001",
    2098=>"011010101",
    2099=>"111101000",
    2100=>"111000100",
    2101=>"110100100",
    2102=>"010000101",
    2103=>"011001010",
    2104=>"110100111",
    2105=>"111000001",
    2106=>"110110100",
    2107=>"100100000",
    2108=>"101001010",
    2109=>"011001000",
    2110=>"110100100",
    2111=>"000000001",
    2112=>"110100100",
    2113=>"001011111",
    2114=>"011011111",
    2115=>"011011111",
    2116=>"011011111",
    2117=>"100001001",
    2118=>"011100101",
    2119=>"010100000",
    2120=>"001011111",
    2121=>"100100100",
    2122=>"001011111",
    2123=>"110100000",
    2124=>"101001111",
    2125=>"010000000",
    2126=>"110110000",
    2127=>"010010011",
    2128=>"101110001",
    2129=>"001011001",
    2130=>"100100100",
    2131=>"011100111",
    2132=>"110110000",
    2133=>"100100100",
    2134=>"110100000",
    2135=>"110001001",
    2136=>"011011011",
    2137=>"110100000",
    2138=>"110100000",
    2139=>"110100001",
    2140=>"100000000",
    2141=>"000000100",
    2142=>"111011011",
    2143=>"100100100",
    2144=>"100100000",
    2145=>"011111101",
    2146=>"111010100",
    2147=>"100000000",
    2148=>"110100100",
    2149=>"100100110",
    2150=>"011111111",
    2151=>"101100101",
    2152=>"011011111",
    2153=>"110100000",
    2154=>"110000000",
    2155=>"100100001",
    2156=>"100100101",
    2157=>"100100100",
    2158=>"100100100",
    2159=>"100000000",
    2160=>"101011111",
    2161=>"110000000",
    2162=>"100111010",
    2163=>"101101001",
    2164=>"001011111",
    2165=>"100100000",
    2166=>"110111001",
    2167=>"001001111",
    2168=>"100001011",
    2169=>"100100110",
    2170=>"010100000",
    2171=>"100100100",
    2172=>"011010001",
    2173=>"110100011",
    2174=>"011111011",
    2175=>"000100100",
    2176=>"011001000",
    2177=>"011011000",
    2178=>"100100110",
    2179=>"001111111",
    2180=>"100100110",
    2181=>"101100011",
    2182=>"111110111",
    2183=>"011001101",
    2184=>"100100110",
    2185=>"101111111",
    2186=>"101110001",
    2187=>"100110011",
    2188=>"101101111",
    2189=>"010010001",
    2190=>"100110010",
    2191=>"000100111",
    2192=>"011001001",
    2193=>"011001101",
    2194=>"100110010",
    2195=>"110010111",
    2196=>"110010011",
    2197=>"100100010",
    2198=>"011011101",
    2199=>"111011000",
    2200=>"111001001",
    2201=>"111001010",
    2202=>"011001101",
    2203=>"110000001",
    2204=>"100100110",
    2205=>"000100011",
    2206=>"001001001",
    2207=>"100010010",
    2208=>"100100110",
    2209=>"100100110",
    2210=>"100000011",
    2211=>"001001101",
    2212=>"000101101",
    2213=>"100100010",
    2214=>"011001001",
    2215=>"100110010",
    2216=>"000000010",
    2217=>"001000001",
    2218=>"110110011",
    2219=>"010011001",
    2220=>"100110010",
    2221=>"000000011",
    2222=>"100110110",
    2223=>"100110110",
    2224=>"011011001",
    2225=>"000010011",
    2226=>"001100010",
    2227=>"101110011",
    2228=>"111001001",
    2229=>"101000000",
    2230=>"100010110",
    2231=>"011001001",
    2232=>"101110010",
    2233=>"100110011",
    2234=>"011101101",
    2235=>"100000000",
    2236=>"110011101",
    2237=>"010000100",
    2238=>"001001001",
    2239=>"000100110",
    2240=>"000010100",
    2241=>"010101101",
    2242=>"111101111",
    2243=>"111010010",
    2244=>"100100001",
    2245=>"110100000",
    2246=>"101111110",
    2247=>"011101110",
    2248=>"000000000",
    2249=>"011000011",
    2250=>"001001000",
    2251=>"111111011",
    2252=>"111111111",
    2253=>"001001000",
    2254=>"011011110",
    2255=>"110111110",
    2256=>"000011110",
    2257=>"111101110",
    2258=>"111111111",
    2259=>"110111110",
    2260=>"000000000",
    2261=>"100111111",
    2262=>"000111000",
    2263=>"001011000",
    2264=>"000000101",
    2265=>"101011110",
    2266=>"001000000",
    2267=>"010110001",
    2268=>"000010001",
    2269=>"110000100",
    2270=>"111110111",
    2271=>"010010001",
    2272=>"111110100",
    2273=>"011110110",
    2274=>"111111111",
    2275=>"000000000",
    2276=>"011000000",
    2277=>"110100011",
    2278=>"110111011",
    2279=>"100111011",
    2280=>"110010101",
    2281=>"000000000",
    2282=>"100111010",
    2283=>"111111110",
    2284=>"111110111",
    2285=>"001000000",
    2286=>"111101000",
    2287=>"110110000",
    2288=>"010010001",
    2289=>"000000000",
    2290=>"101101011",
    2291=>"001001010",
    2292=>"011111111",
    2293=>"001111110",
    2294=>"111010101",
    2295=>"100000010",
    2296=>"111110110",
    2297=>"001011110",
    2298=>"100011110",
    2299=>"100000010",
    2300=>"000001001",
    2301=>"000000011",
    2302=>"111110110",
    2303=>"000000010",
    2304=>"110000001",
    2305=>"000111111",
    2306=>"000111111",
    2307=>"000111111",
    2308=>"001111111",
    2309=>"111101000",
    2310=>"001001011",
    2311=>"001100001",
    2312=>"010111111",
    2313=>"111000000",
    2314=>"100111111",
    2315=>"000001111",
    2316=>"111111110",
    2317=>"101000011",
    2318=>"111100000",
    2319=>"001101110",
    2320=>"111001000",
    2321=>"111110110",
    2322=>"111001010",
    2323=>"111111000",
    2324=>"001000110",
    2325=>"000101001",
    2326=>"000000101",
    2327=>"100100111",
    2328=>"000000000",
    2329=>"001000111",
    2330=>"111100001",
    2331=>"011001001",
    2332=>"010110110",
    2333=>"010011111",
    2334=>"010000110",
    2335=>"101101101",
    2336=>"100000000",
    2337=>"010111111",
    2338=>"111001101",
    2339=>"110000000",
    2340=>"001000000",
    2341=>"100000001",
    2342=>"110111111",
    2343=>"110111111",
    2344=>"000111111",
    2345=>"111000000",
    2346=>"111000000",
    2347=>"101100000",
    2348=>"011001101",
    2349=>"011100111",
    2350=>"000010111",
    2351=>"111011111",
    2352=>"000011111",
    2353=>"000000111",
    2354=>"100001110",
    2355=>"001000000",
    2356=>"000111111",
    2357=>"000001101",
    2358=>"111100001",
    2359=>"000010000",
    2360=>"111111000",
    2361=>"001000001",
    2362=>"111100100",
    2363=>"111101111",
    2364=>"001001001",
    2365=>"001001001",
    2366=>"110111111",
    2367=>"110001001",
    2368=>"010100100",
    2369=>"010010000",
    2370=>"011111100",
    2371=>"101101111",
    2372=>"010001011",
    2373=>"000010110",
    2374=>"111111111",
    2375=>"000001000",
    2376=>"011000010",
    2377=>"111011001",
    2378=>"010000001",
    2379=>"110010100",
    2380=>"111111011",
    2381=>"001011000",
    2382=>"001011000",
    2383=>"011111010",
    2384=>"010111011",
    2385=>"011001000",
    2386=>"001110000",
    2387=>"000001001",
    2388=>"111100100",
    2389=>"100000010",
    2390=>"010000010",
    2391=>"011001000",
    2392=>"110000000",
    2393=>"011111010",
    2394=>"100000001",
    2395=>"110110111",
    2396=>"111111111",
    2397=>"001100010",
    2398=>"111111111",
    2399=>"000000000",
    2400=>"000000000",
    2401=>"010010101",
    2402=>"001011101",
    2403=>"101100100",
    2404=>"001110100",
    2405=>"001111000",
    2406=>"000000001",
    2407=>"111110000",
    2408=>"111101000",
    2409=>"000000011",
    2410=>"000011001",
    2411=>"000001100",
    2412=>"000001000",
    2413=>"000011000",
    2414=>"111111101",
    2415=>"000101010",
    2416=>"100100101",
    2417=>"100101111",
    2418=>"010010000",
    2419=>"000000000",
    2420=>"000000000",
    2421=>"110100101",
    2422=>"001111111",
    2423=>"010010000",
    2424=>"010011110",
    2425=>"111001000",
    2426=>"110111000",
    2427=>"111111001",
    2428=>"010000000",
    2429=>"111000001",
    2430=>"111100011",
    2431=>"100000111",
    2432=>"111111011",
    2433=>"011000111",
    2434=>"000000000",
    2435=>"001100110",
    2436=>"000000110",
    2437=>"000111110",
    2438=>"110011001",
    2439=>"100010000",
    2440=>"010000000",
    2441=>"111001001",
    2442=>"000000000",
    2443=>"110110000",
    2444=>"111111100",
    2445=>"101011000",
    2446=>"011100100",
    2447=>"100111000",
    2448=>"111111111",
    2449=>"000000111",
    2450=>"010111010",
    2451=>"010010001",
    2452=>"001100111",
    2453=>"000000000",
    2454=>"000110110",
    2455=>"000000111",
    2456=>"000000101",
    2457=>"000000110",
    2458=>"000011011",
    2459=>"101100001",
    2460=>"111000100",
    2461=>"000000000",
    2462=>"011110111",
    2463=>"001000001",
    2464=>"011111000",
    2465=>"100110111",
    2466=>"111000111",
    2467=>"000000000",
    2468=>"110111110",
    2469=>"100111100",
    2470=>"001011111",
    2471=>"010000000",
    2472=>"000000000",
    2473=>"111001000",
    2474=>"111100111",
    2475=>"011011011",
    2476=>"111111101",
    2477=>"011000010",
    2478=>"100111000",
    2479=>"110111011",
    2480=>"000110111",
    2481=>"000000000",
    2482=>"001000000",
    2483=>"100000000",
    2484=>"000000111",
    2485=>"001111000",
    2486=>"001111000",
    2487=>"111111000",
    2488=>"001011011",
    2489=>"111011101",
    2490=>"001111010",
    2491=>"100000000",
    2492=>"000000111",
    2493=>"100111111",
    2494=>"000000000",
    2495=>"000000000",
    2496=>"001001000",
    2497=>"000000000",
    2498=>"111111011",
    2499=>"010010000",
    2500=>"111111111",
    2501=>"100000100",
    2502=>"000000000",
    2503=>"000111010",
    2504=>"111100111",
    2505=>"010111010",
    2506=>"111111101",
    2507=>"110111101",
    2508=>"110111010",
    2509=>"000100001",
    2510=>"111101101",
    2511=>"111001111",
    2512=>"000000000",
    2513=>"000000000",
    2514=>"011101100",
    2515=>"100000101",
    2516=>"000101000",
    2517=>"100100101",
    2518=>"100111000",
    2519=>"100000000",
    2520=>"000000000",
    2521=>"011001101",
    2522=>"001001000",
    2523=>"100001111",
    2524=>"111111000",
    2525=>"011111011",
    2526=>"000000000",
    2527=>"111111101",
    2528=>"000101101",
    2529=>"011011100",
    2530=>"000000000",
    2531=>"101000100",
    2532=>"111111111",
    2533=>"011111010",
    2534=>"000111011",
    2535=>"011110110",
    2536=>"101111110",
    2537=>"000000000",
    2538=>"110000100",
    2539=>"100000000",
    2540=>"000000001",
    2541=>"001101001",
    2542=>"111111111",
    2543=>"010101111",
    2544=>"100100111",
    2545=>"100101001",
    2546=>"000000010",
    2547=>"000101001",
    2548=>"101111111",
    2549=>"111111011",
    2550=>"111001111",
    2551=>"001100100",
    2552=>"000001001",
    2553=>"001100001",
    2554=>"110100000",
    2555=>"100011101",
    2556=>"000000000",
    2557=>"100000001",
    2558=>"111111111",
    2559=>"101101000",
    2560=>"111111100",
    2561=>"000010000",
    2562=>"000000111",
    2563=>"000000111",
    2564=>"000000000",
    2565=>"110111001",
    2566=>"000111100",
    2567=>"001001111",
    2568=>"110111111",
    2569=>"110001100",
    2570=>"001011000",
    2571=>"110010000",
    2572=>"111000111",
    2573=>"000000000",
    2574=>"000010101",
    2575=>"000000111",
    2576=>"111110000",
    2577=>"010111111",
    2578=>"010101000",
    2579=>"101011010",
    2580=>"111011000",
    2581=>"011000000",
    2582=>"011011101",
    2583=>"000011000",
    2584=>"111010000",
    2585=>"010011000",
    2586=>"001111100",
    2587=>"111001000",
    2588=>"000110010",
    2589=>"111100011",
    2590=>"010011001",
    2591=>"000111111",
    2592=>"011101010",
    2593=>"000110111",
    2594=>"000000000",
    2595=>"011000110",
    2596=>"111111111",
    2597=>"111000011",
    2598=>"000001111",
    2599=>"111110000",
    2600=>"111000110",
    2601=>"111000001",
    2602=>"111111000",
    2603=>"000000000",
    2604=>"110110001",
    2605=>"111111000",
    2606=>"111000000",
    2607=>"010110010",
    2608=>"000111110",
    2609=>"111111000",
    2610=>"100110011",
    2611=>"101110000",
    2612=>"101110111",
    2613=>"100000000",
    2614=>"001000110",
    2615=>"011111000",
    2616=>"000010001",
    2617=>"010000111",
    2618=>"011111000",
    2619=>"001111100",
    2620=>"000010000",
    2621=>"110000011",
    2622=>"111010111",
    2623=>"111111000",
    2624=>"101000010",
    2625=>"001110000",
    2626=>"110111011",
    2627=>"111110000",
    2628=>"000000011",
    2629=>"100100001",
    2630=>"110011010",
    2631=>"011010010",
    2632=>"000001011",
    2633=>"110100101",
    2634=>"000011111",
    2635=>"001000010",
    2636=>"111111010",
    2637=>"100111101",
    2638=>"000001010",
    2639=>"110110000",
    2640=>"101001010",
    2641=>"010111100",
    2642=>"011001000",
    2643=>"000000011",
    2644=>"111100000",
    2645=>"000001111",
    2646=>"100000110",
    2647=>"001011111",
    2648=>"100100011",
    2649=>"101001110",
    2650=>"101000000",
    2651=>"010001001",
    2652=>"000001111",
    2653=>"111100000",
    2654=>"101000101",
    2655=>"000000000",
    2656=>"001000111",
    2657=>"000101111",
    2658=>"101111111",
    2659=>"111000000",
    2660=>"111110000",
    2661=>"111110100",
    2662=>"111001001",
    2663=>"000011111",
    2664=>"001001001",
    2665=>"000000011",
    2666=>"000000011",
    2667=>"110111001",
    2668=>"000000011",
    2669=>"000000001",
    2670=>"011111000",
    2671=>"111000111",
    2672=>"011111110",
    2673=>"000001111",
    2674=>"010110100",
    2675=>"001011111",
    2676=>"011011010",
    2677=>"100001111",
    2678=>"010000001",
    2679=>"000100111",
    2680=>"101001001",
    2681=>"001000110",
    2682=>"000100000",
    2683=>"011000000",
    2684=>"110100101",
    2685=>"110100000",
    2686=>"000001011",
    2687=>"000000011",
    2688=>"001001010",
    2689=>"100100000",
    2690=>"010011111",
    2691=>"001010010",
    2692=>"011111111",
    2693=>"101001101",
    2694=>"110110100",
    2695=>"011011110",
    2696=>"000011000",
    2697=>"011010010",
    2698=>"111110111",
    2699=>"001001011",
    2700=>"101111111",
    2701=>"111010000",
    2702=>"001011011",
    2703=>"011110100",
    2704=>"010110001",
    2705=>"110100100",
    2706=>"000000001",
    2707=>"010110101",
    2708=>"101111010",
    2709=>"001000000",
    2710=>"111101001",
    2711=>"110100100",
    2712=>"100001011",
    2713=>"100101111",
    2714=>"110100100",
    2715=>"010100000",
    2716=>"100100101",
    2717=>"011011001",
    2718=>"000001001",
    2719=>"101001001",
    2720=>"001011110",
    2721=>"000001001",
    2722=>"100001101",
    2723=>"100110000",
    2724=>"010101111",
    2725=>"001001011",
    2726=>"110100100",
    2727=>"000000000",
    2728=>"001011011",
    2729=>"100100100",
    2730=>"100001111",
    2731=>"100100000",
    2732=>"001001111",
    2733=>"010101111",
    2734=>"011011010",
    2735=>"011111011",
    2736=>"110100100",
    2737=>"110100000",
    2738=>"001001101",
    2739=>"000000000",
    2740=>"110110000",
    2741=>"000010110",
    2742=>"011010110",
    2743=>"000001001",
    2744=>"110100100",
    2745=>"001111011",
    2746=>"001011110",
    2747=>"001011110",
    2748=>"100100101",
    2749=>"100001100",
    2750=>"000011110",
    2751=>"010001001",
    2752=>"101101100",
    2753=>"101100100",
    2754=>"110001000",
    2755=>"001011011",
    2756=>"101101111",
    2757=>"100000100",
    2758=>"110010110",
    2759=>"011101101",
    2760=>"111110110",
    2761=>"010000000",
    2762=>"101101111",
    2763=>"111111110",
    2764=>"101101101",
    2765=>"101011010",
    2766=>"000000000",
    2767=>"101110100",
    2768=>"001000000",
    2769=>"111111111",
    2770=>"010001001",
    2771=>"111000110",
    2772=>"100010100",
    2773=>"100100000",
    2774=>"011011101",
    2775=>"111110110",
    2776=>"100001000",
    2777=>"001001011",
    2778=>"101010100",
    2779=>"111111111",
    2780=>"001011011",
    2781=>"011111111",
    2782=>"100000011",
    2783=>"100100100",
    2784=>"011001100",
    2785=>"101101101",
    2786=>"000011000",
    2787=>"000001011",
    2788=>"001010000",
    2789=>"100000001",
    2790=>"100101000",
    2791=>"110110110",
    2792=>"010110000",
    2793=>"011011111",
    2794=>"111011110",
    2795=>"001011001",
    2796=>"111111101",
    2797=>"000000000",
    2798=>"001000101",
    2799=>"001011010",
    2800=>"001001001",
    2801=>"001011000",
    2802=>"101110011",
    2803=>"000111000",
    2804=>"100100100",
    2805=>"111111111",
    2806=>"111001101",
    2807=>"001001001",
    2808=>"100000000",
    2809=>"000000000",
    2810=>"110010000",
    2811=>"111111111",
    2812=>"100101110",
    2813=>"000001011",
    2814=>"011110101",
    2815=>"000000010",
    2816=>"010001000",
    2817=>"111011000",
    2818=>"110010001",
    2819=>"100111111",
    2820=>"011000100",
    2821=>"000011101",
    2822=>"000110001",
    2823=>"011100000",
    2824=>"101110101",
    2825=>"111000000",
    2826=>"111101000",
    2827=>"111000100",
    2828=>"101101111",
    2829=>"011110011",
    2830=>"111000000",
    2831=>"011010000",
    2832=>"001110010",
    2833=>"010100111",
    2834=>"000100111",
    2835=>"001011101",
    2836=>"100001101",
    2837=>"111001000",
    2838=>"100111111",
    2839=>"011000000",
    2840=>"000001100",
    2841=>"000000101",
    2842=>"001001000",
    2843=>"111111111",
    2844=>"100000000",
    2845=>"111011011",
    2846=>"100010011",
    2847=>"111101011",
    2848=>"111001000",
    2849=>"011001100",
    2850=>"111011111",
    2851=>"001100101",
    2852=>"101110011",
    2853=>"001100000",
    2854=>"011001000",
    2855=>"101110010",
    2856=>"010000010",
    2857=>"000010110",
    2858=>"000000000",
    2859=>"000100100",
    2860=>"010111011",
    2861=>"111000000",
    2862=>"111111001",
    2863=>"111110110",
    2864=>"000100111",
    2865=>"111001000",
    2866=>"111110011",
    2867=>"111011000",
    2868=>"111011000",
    2869=>"000000000",
    2870=>"111010001",
    2871=>"001000100",
    2872=>"011000100",
    2873=>"110011001",
    2874=>"010110000",
    2875=>"011001010",
    2876=>"011001001",
    2877=>"000000000",
    2878=>"110110001",
    2879=>"000100110",
    2880=>"000101001",
    2881=>"010111000",
    2882=>"010010000",
    2883=>"111111010",
    2884=>"000000000",
    2885=>"011000101",
    2886=>"000000000",
    2887=>"100111000",
    2888=>"000000000",
    2889=>"101010110",
    2890=>"000000000",
    2891=>"001101100",
    2892=>"110111011",
    2893=>"111011000",
    2894=>"011111100",
    2895=>"010010000",
    2896=>"111000100",
    2897=>"111000000",
    2898=>"000000111",
    2899=>"111110001",
    2900=>"000000111",
    2901=>"111000000",
    2902=>"000100000",
    2903=>"110000000",
    2904=>"011011111",
    2905=>"111011110",
    2906=>"100000011",
    2907=>"111000111",
    2908=>"000111110",
    2909=>"101111111",
    2910=>"010000000",
    2911=>"000000111",
    2912=>"100111101",
    2913=>"111111110",
    2914=>"111001111",
    2915=>"100000110",
    2916=>"001000100",
    2917=>"000001000",
    2918=>"111111110",
    2919=>"111011100",
    2920=>"000010110",
    2921=>"111101111",
    2922=>"111000000",
    2923=>"000000001",
    2924=>"001111110",
    2925=>"110000111",
    2926=>"000101111",
    2927=>"110111111",
    2928=>"000000111",
    2929=>"100000000",
    2930=>"011011000",
    2931=>"000100111",
    2932=>"000010110",
    2933=>"100101011",
    2934=>"001111111",
    2935=>"111111000",
    2936=>"110101010",
    2937=>"110100000",
    2938=>"110100000",
    2939=>"111111101",
    2940=>"001001111",
    2941=>"011001101",
    2942=>"110110111",
    2943=>"111111000",
    2944=>"001100100",
    2945=>"011111011",
    2946=>"111111010",
    2947=>"111010000",
    2948=>"111101000",
    2949=>"111001101",
    2950=>"110111110",
    2951=>"011111110",
    2952=>"111011100",
    2953=>"000000111",
    2954=>"111110000",
    2955=>"110011001",
    2956=>"010010110",
    2957=>"000100111",
    2958=>"000001100",
    2959=>"111000000",
    2960=>"101111110",
    2961=>"111111000",
    2962=>"001100101",
    2963=>"111010100",
    2964=>"100100000",
    2965=>"000100111",
    2966=>"111000000",
    2967=>"010101011",
    2968=>"000000000",
    2969=>"000001111",
    2970=>"111100100",
    2971=>"010000011",
    2972=>"000010110",
    2973=>"111000000",
    2974=>"010111011",
    2975=>"000100111",
    2976=>"111010000",
    2977=>"111111000",
    2978=>"011001000",
    2979=>"111100100",
    2980=>"110001101",
    2981=>"100111011",
    2982=>"111000000",
    2983=>"001100110",
    2984=>"111111001",
    2985=>"000000111",
    2986=>"111100011",
    2987=>"001000000",
    2988=>"000001001",
    2989=>"100001000",
    2990=>"111111010",
    2991=>"011111101",
    2992=>"110111110",
    2993=>"100110010",
    2994=>"111111001",
    2995=>"010010110",
    2996=>"010011010",
    2997=>"100001011",
    2998=>"110110101",
    2999=>"101000000",
    3000=>"111110101",
    3001=>"000000100",
    3002=>"110001011",
    3003=>"101101001",
    3004=>"111101000",
    3005=>"101100100",
    3006=>"110111111",
    3007=>"011011000",
    3008=>"011111111",
    3009=>"111000000",
    3010=>"000000100",
    3011=>"010011000",
    3012=>"111111010",
    3013=>"001011100",
    3014=>"100000001",
    3015=>"000111010",
    3016=>"011001001",
    3017=>"100000001",
    3018=>"111111000",
    3019=>"001011000",
    3020=>"111010010",
    3021=>"001010000",
    3022=>"100000000",
    3023=>"000101111",
    3024=>"111011101",
    3025=>"011111110",
    3026=>"000001100",
    3027=>"111111111",
    3028=>"110110010",
    3029=>"000000100",
    3030=>"010010000",
    3031=>"000000000",
    3032=>"000000000",
    3033=>"001000111",
    3034=>"100110001",
    3035=>"100011001",
    3036=>"100000100",
    3037=>"000111000",
    3038=>"001000100",
    3039=>"000000000",
    3040=>"000000001",
    3041=>"110011110",
    3042=>"011111111",
    3043=>"000101000",
    3044=>"110111010",
    3045=>"100111100",
    3046=>"110111001",
    3047=>"100001101",
    3048=>"000000101",
    3049=>"000000001",
    3050=>"000110001",
    3051=>"100110000",
    3052=>"110111111",
    3053=>"100000000",
    3054=>"000111000",
    3055=>"000000000",
    3056=>"111111111",
    3057=>"000000111",
    3058=>"011011110",
    3059=>"010100111",
    3060=>"100111111",
    3061=>"001000011",
    3062=>"000100000",
    3063=>"111000000",
    3064=>"010011000",
    3065=>"001010110",
    3066=>"100100000",
    3067=>"100010000",
    3068=>"110010000",
    3069=>"100101011",
    3070=>"001000001",
    3071=>"011010000",
    3072=>"011000000",
    3073=>"000000110",
    3074=>"111101101",
    3075=>"000011111",
    3076=>"111100000",
    3077=>"001011001",
    3078=>"000010011",
    3079=>"100100110",
    3080=>"000110111",
    3081=>"000010111",
    3082=>"011011011",
    3083=>"101100100",
    3084=>"000111111",
    3085=>"000100100",
    3086=>"111101100",
    3087=>"000110101",
    3088=>"110010110",
    3089=>"111111000",
    3090=>"001100100",
    3091=>"000001111",
    3092=>"001000100",
    3093=>"111000000",
    3094=>"111101000",
    3095=>"000100111",
    3096=>"000000000",
    3097=>"111000000",
    3098=>"100100100",
    3099=>"111100000",
    3100=>"111100110",
    3101=>"111011000",
    3102=>"000000000",
    3103=>"111111000",
    3104=>"000000111",
    3105=>"111100100",
    3106=>"000000000",
    3107=>"000100100",
    3108=>"001000011",
    3109=>"000011011",
    3110=>"001011011",
    3111=>"100100111",
    3112=>"111101100",
    3113=>"110010010",
    3114=>"100000001",
    3115=>"110010011",
    3116=>"111001000",
    3117=>"111011011",
    3118=>"000110111",
    3119=>"101101011",
    3120=>"111001000",
    3121=>"000000011",
    3122=>"011011011",
    3123=>"001001001",
    3124=>"000000110",
    3125=>"101001001",
    3126=>"101101101",
    3127=>"000000110",
    3128=>"101011011",
    3129=>"011001111",
    3130=>"111011011",
    3131=>"011001001",
    3132=>"111111000",
    3133=>"001001001",
    3134=>"001011011",
    3135=>"111111011",
    3136=>"000100000",
    3137=>"010101111",
    3138=>"111111111",
    3139=>"111111010",
    3140=>"001001100",
    3141=>"001001110",
    3142=>"111010101",
    3143=>"111011011",
    3144=>"001000010",
    3145=>"110110010",
    3146=>"101000111",
    3147=>"001000100",
    3148=>"111101111",
    3149=>"110100000",
    3150=>"101111111",
    3151=>"110100000",
    3152=>"110010001",
    3153=>"101011001",
    3154=>"111111100",
    3155=>"001111011",
    3156=>"101110100",
    3157=>"000000000",
    3158=>"000000000",
    3159=>"000000000",
    3160=>"101000100",
    3161=>"110111010",
    3162=>"011010010",
    3163=>"111100101",
    3164=>"001100111",
    3165=>"001001001",
    3166=>"011110111",
    3167=>"100010000",
    3168=>"000000100",
    3169=>"001100101",
    3170=>"010000110",
    3171=>"001000100",
    3172=>"001011100",
    3173=>"000001000",
    3174=>"010101111",
    3175=>"101110010",
    3176=>"011010011",
    3177=>"110110110",
    3178=>"101000001",
    3179=>"100000110",
    3180=>"001101100",
    3181=>"000000000",
    3182=>"000000000",
    3183=>"100000000",
    3184=>"101001000",
    3185=>"111001000",
    3186=>"111001101",
    3187=>"000000000",
    3188=>"000100000",
    3189=>"000000001",
    3190=>"000001100",
    3191=>"111111000",
    3192=>"111111111",
    3193=>"101100101",
    3194=>"101011110",
    3195=>"111111111",
    3196=>"000100110",
    3197=>"110010101",
    3198=>"001101011",
    3199=>"111000000",
    3200=>"010110011",
    3201=>"001001000",
    3202=>"000000100",
    3203=>"011010110",
    3204=>"110011001",
    3205=>"110001000",
    3206=>"000000100",
    3207=>"001100111",
    3208=>"111011001",
    3209=>"000100101",
    3210=>"100100110",
    3211=>"110111001",
    3212=>"011100111",
    3213=>"011000000",
    3214=>"110011001",
    3215=>"111011001",
    3216=>"100011001",
    3217=>"110011001",
    3218=>"110010001",
    3219=>"001000110",
    3220=>"110011000",
    3221=>"100010001",
    3222=>"111011010",
    3223=>"110011001",
    3224=>"001100110",
    3225=>"010001100",
    3226=>"001100111",
    3227=>"100110110",
    3228=>"010001000",
    3229=>"000101111",
    3230=>"111011001",
    3231=>"111011001",
    3232=>"001100110",
    3233=>"011001000",
    3234=>"111011000",
    3235=>"100000111",
    3236=>"110111001",
    3237=>"010011000",
    3238=>"000100010",
    3239=>"110010001",
    3240=>"000100000",
    3241=>"110001100",
    3242=>"110111001",
    3243=>"000000001",
    3244=>"000000110",
    3245=>"000100010",
    3246=>"001100110",
    3247=>"100001000",
    3248=>"110011010",
    3249=>"010001100",
    3250=>"111000000",
    3251=>"010011010",
    3252=>"111001000",
    3253=>"001100000",
    3254=>"100011000",
    3255=>"100100111",
    3256=>"101010001",
    3257=>"110011001",
    3258=>"110110011",
    3259=>"000000110",
    3260=>"111111011",
    3261=>"111010000",
    3262=>"111111111",
    3263=>"100011001",
    3264=>"000000001",
    3265=>"000011111",
    3266=>"011000000",
    3267=>"011011110",
    3268=>"111101011",
    3269=>"000000000",
    3270=>"110100111",
    3271=>"000100000",
    3272=>"100100100",
    3273=>"000001111",
    3274=>"111111111",
    3275=>"111100100",
    3276=>"111100100",
    3277=>"010001000",
    3278=>"000000000",
    3279=>"000111110",
    3280=>"000000000",
    3281=>"100111110",
    3282=>"001000000",
    3283=>"000000000",
    3284=>"000100101",
    3285=>"000000001",
    3286=>"111110000",
    3287=>"100010111",
    3288=>"101000000",
    3289=>"001001011",
    3290=>"100000000",
    3291=>"001001011",
    3292=>"100101011",
    3293=>"111110000",
    3294=>"100100111",
    3295=>"110001111",
    3296=>"010100110",
    3297=>"000000111",
    3298=>"000000000",
    3299=>"111000101",
    3300=>"101000001",
    3301=>"111111001",
    3302=>"001011111",
    3303=>"000000001",
    3304=>"011011011",
    3305=>"000000000",
    3306=>"000000101",
    3307=>"110110000",
    3308=>"000000011",
    3309=>"111111111",
    3310=>"111110110",
    3311=>"011011111",
    3312=>"000000001",
    3313=>"000000111",
    3314=>"011111111",
    3315=>"001001001",
    3316=>"010100101",
    3317=>"001001001",
    3318=>"000000101",
    3319=>"100000000",
    3320=>"000001001",
    3321=>"000001111",
    3322=>"000000100",
    3323=>"000001111",
    3324=>"111101001",
    3325=>"111110100",
    3326=>"001111111",
    3327=>"001111111",
    3328=>"001111101",
    3329=>"111110111",
    3330=>"010000000",
    3331=>"110110100",
    3332=>"111101111",
    3333=>"110110101",
    3334=>"110011001",
    3335=>"100010011",
    3336=>"111011001",
    3337=>"011001001",
    3338=>"101100110",
    3339=>"111001001",
    3340=>"100101101",
    3341=>"000001010",
    3342=>"011001001",
    3343=>"001001011",
    3344=>"100100011",
    3345=>"101100100",
    3346=>"101101111",
    3347=>"010000000",
    3348=>"000000000",
    3349=>"001001001",
    3350=>"110110110",
    3351=>"111110100",
    3352=>"100110100",
    3353=>"001001001",
    3354=>"100110111",
    3355=>"001011001",
    3356=>"001001001",
    3357=>"100001111",
    3358=>"011010001",
    3359=>"011001001",
    3360=>"100110110",
    3361=>"101101101",
    3362=>"100100110",
    3363=>"100100100",
    3364=>"100001000",
    3365=>"100000001",
    3366=>"000110101",
    3367=>"110010111",
    3368=>"111010101",
    3369=>"001001001",
    3370=>"101011100",
    3371=>"110100101",
    3372=>"001000100",
    3373=>"000000000",
    3374=>"100110010",
    3375=>"011011011",
    3376=>"001001001",
    3377=>"001001000",
    3378=>"111110100",
    3379=>"111001111",
    3380=>"001010000",
    3381=>"001000110",
    3382=>"000000000",
    3383=>"110110110",
    3384=>"110110100",
    3385=>"110001100",
    3386=>"001000001",
    3387=>"111110100",
    3388=>"100100110",
    3389=>"100100110",
    3390=>"001011010",
    3391=>"011010001",
    3392=>"010110100",
    3393=>"000111111",
    3394=>"110111011",
    3395=>"010111011",
    3396=>"011001001",
    3397=>"110110111",
    3398=>"100001111",
    3399=>"011001000",
    3400=>"010111101",
    3401=>"010000000",
    3402=>"000100000",
    3403=>"101100111",
    3404=>"010011111",
    3405=>"001111110",
    3406=>"110011001",
    3407=>"111111111",
    3408=>"111100101",
    3409=>"000011111",
    3410=>"111110110",
    3411=>"101011000",
    3412=>"111001000",
    3413=>"010111111",
    3414=>"000000000",
    3415=>"000111001",
    3416=>"000101100",
    3417=>"111111100",
    3418=>"011111101",
    3419=>"000001010",
    3420=>"000111111",
    3421=>"111000000",
    3422=>"000111111",
    3423=>"000010110",
    3424=>"110110011",
    3425=>"000110111",
    3426=>"110010100",
    3427=>"111000000",
    3428=>"100000000",
    3429=>"110000000",
    3430=>"000001111",
    3431=>"011111011",
    3432=>"010111111",
    3433=>"111111111",
    3434=>"110110000",
    3435=>"000100101",
    3436=>"111101001",
    3437=>"000111111",
    3438=>"111001111",
    3439=>"111110111",
    3440=>"000000000",
    3441=>"111111000",
    3442=>"101111011",
    3443=>"000110111",
    3444=>"000000010",
    3445=>"001000001",
    3446=>"100011111",
    3447=>"000001011",
    3448=>"101101111",
    3449=>"000000110",
    3450=>"110001001",
    3451=>"111110100",
    3452=>"000111111",
    3453=>"111010000",
    3454=>"001011111",
    3455=>"000111000",
    3456=>"011100111",
    3457=>"111001111",
    3458=>"111111111",
    3459=>"010111000",
    3460=>"100100110",
    3461=>"111001111",
    3462=>"001101101",
    3463=>"000000100",
    3464=>"000100000",
    3465=>"111111101",
    3466=>"001011110",
    3467=>"000001000",
    3468=>"100111100",
    3469=>"111111111",
    3470=>"110001001",
    3471=>"000110111",
    3472=>"101111101",
    3473=>"110111000",
    3474=>"111101111",
    3475=>"100011111",
    3476=>"011001000",
    3477=>"110110110",
    3478=>"000000000",
    3479=>"111000000",
    3480=>"000000000",
    3481=>"111111000",
    3482=>"111100011",
    3483=>"110110000",
    3484=>"000111110",
    3485=>"000000000",
    3486=>"111111111",
    3487=>"110000000",
    3488=>"111000000",
    3489=>"011111100",
    3490=>"111000110",
    3491=>"000000000",
    3492=>"001000010",
    3493=>"100000001",
    3494=>"110011110",
    3495=>"111110111",
    3496=>"111110111",
    3497=>"111111100",
    3498=>"011111100",
    3499=>"011000100",
    3500=>"110101111",
    3501=>"000010100",
    3502=>"011000011",
    3503=>"000111101",
    3504=>"110111000",
    3505=>"111111110",
    3506=>"100011101",
    3507=>"110111110",
    3508=>"000100000",
    3509=>"100000001",
    3510=>"000000000",
    3511=>"101000111",
    3512=>"111111111",
    3513=>"110110000",
    3514=>"111100110",
    3515=>"000000000",
    3516=>"000000000",
    3517=>"000000001",
    3518=>"001101111",
    3519=>"000000000",
    3520=>"100100111",
    3521=>"010111010",
    3522=>"010011011",
    3523=>"010111010",
    3524=>"000011110",
    3525=>"000000100",
    3526=>"000000001",
    3527=>"101000001",
    3528=>"000001000",
    3529=>"111111101",
    3530=>"000010011",
    3531=>"000100110",
    3532=>"011111010",
    3533=>"111111111",
    3534=>"001101001",
    3535=>"000001000",
    3536=>"000000000",
    3537=>"010000000",
    3538=>"000000100",
    3539=>"110100100",
    3540=>"000000111",
    3541=>"010111100",
    3542=>"111101101",
    3543=>"110000000",
    3544=>"000000000",
    3545=>"101100111",
    3546=>"100000001",
    3547=>"000001011",
    3548=>"000000010",
    3549=>"000000100",
    3550=>"110010110",
    3551=>"111111111",
    3552=>"110100000",
    3553=>"000000110",
    3554=>"011001000",
    3555=>"000000100",
    3556=>"011101111",
    3557=>"100000100",
    3558=>"000010111",
    3559=>"111011111",
    3560=>"000001110",
    3561=>"010110000",
    3562=>"010001110",
    3563=>"001101011",
    3564=>"111011110",
    3565=>"000000001",
    3566=>"101000100",
    3567=>"111111111",
    3568=>"100000000",
    3569=>"000000010",
    3570=>"101000100",
    3571=>"000000000",
    3572=>"010010010",
    3573=>"100100000",
    3574=>"101101001",
    3575=>"111011010",
    3576=>"010001010",
    3577=>"000100111",
    3578=>"100000000",
    3579=>"000000111",
    3580=>"001000100",
    3581=>"001000001",
    3582=>"111111111",
    3583=>"010000100",
    3584=>"111111000",
    3585=>"000110111",
    3586=>"111111101",
    3587=>"001011011",
    3588=>"111111001",
    3589=>"000100111",
    3590=>"000000000",
    3591=>"101101001",
    3592=>"111100000",
    3593=>"011111000",
    3594=>"111011011",
    3595=>"111100001",
    3596=>"111110111",
    3597=>"000111111",
    3598=>"111011000",
    3599=>"111101010",
    3600=>"010000111",
    3601=>"010000111",
    3602=>"000000000",
    3603=>"110001111",
    3604=>"001000000",
    3605=>"010110110",
    3606=>"000000111",
    3607=>"000111111",
    3608=>"000010111",
    3609=>"110110110",
    3610=>"000011110",
    3611=>"000011011",
    3612=>"110110000",
    3613=>"111000001",
    3614=>"000000000",
    3615=>"110110100",
    3616=>"101000000",
    3617=>"011011000",
    3618=>"010111111",
    3619=>"000000100",
    3620=>"001000000",
    3621=>"111111000",
    3622=>"100000011",
    3623=>"111011100",
    3624=>"111110000",
    3625=>"011000000",
    3626=>"011111100",
    3627=>"000110110",
    3628=>"001101000",
    3629=>"111011000",
    3630=>"111101000",
    3631=>"101001111",
    3632=>"110110000",
    3633=>"000000000",
    3634=>"011000100",
    3635=>"100000000",
    3636=>"000001111",
    3637=>"011011000",
    3638=>"011001000",
    3639=>"000001111",
    3640=>"000011111",
    3641=>"111100001",
    3642=>"000000000",
    3643=>"101101000",
    3644=>"000000111",
    3645=>"100000010",
    3646=>"101111011",
    3647=>"000000111",
    3648=>"111000010",
    3649=>"111011100",
    3650=>"011111110",
    3651=>"100111111",
    3652=>"110110110",
    3653=>"100010101",
    3654=>"010000100",
    3655=>"001101010",
    3656=>"011001110",
    3657=>"111000000",
    3658=>"111010000",
    3659=>"100111000",
    3660=>"111111111",
    3661=>"110000000",
    3662=>"011110001",
    3663=>"000011010",
    3664=>"000000000",
    3665=>"001111010",
    3666=>"110000100",
    3667=>"000101111",
    3668=>"011000000",
    3669=>"111000000",
    3670=>"011000000",
    3671=>"000011111",
    3672=>"011000000",
    3673=>"110000101",
    3674=>"001100110",
    3675=>"010111010",
    3676=>"111000000",
    3677=>"000101111",
    3678=>"011001001",
    3679=>"111000000",
    3680=>"111001001",
    3681=>"101001001",
    3682=>"110011111",
    3683=>"011100110",
    3684=>"000000111",
    3685=>"111111100",
    3686=>"001101100",
    3687=>"110100001",
    3688=>"000110011",
    3689=>"001000000",
    3690=>"000110110",
    3691=>"011010000",
    3692=>"111101011",
    3693=>"001000111",
    3694=>"101001000",
    3695=>"110000000",
    3696=>"110001010",
    3697=>"000000000",
    3698=>"011100001",
    3699=>"100111111",
    3700=>"101111010",
    3701=>"011000000",
    3702=>"001000110",
    3703=>"010010000",
    3704=>"110010011",
    3705=>"100111011",
    3706=>"111000011",
    3707=>"110000000",
    3708=>"100110001",
    3709=>"010001010",
    3710=>"011111001",
    3711=>"100000000",
    3712=>"000001110",
    3713=>"100000001",
    3714=>"000011111",
    3715=>"111000101",
    3716=>"111110100",
    3717=>"100000000",
    3718=>"001001010",
    3719=>"100000111",
    3720=>"110110100",
    3721=>"001010111",
    3722=>"011100100",
    3723=>"011111110",
    3724=>"101011111",
    3725=>"011110111",
    3726=>"001011111",
    3727=>"111110000",
    3728=>"000000101",
    3729=>"110100000",
    3730=>"011111100",
    3731=>"001111000",
    3732=>"011111000",
    3733=>"110110000",
    3734=>"111101001",
    3735=>"110100001",
    3736=>"000001111",
    3737=>"100001001",
    3738=>"101001111",
    3739=>"001001011",
    3740=>"110110000",
    3741=>"011111110",
    3742=>"100100101",
    3743=>"001000101",
    3744=>"000011110",
    3745=>"110110000",
    3746=>"110100001",
    3747=>"000100000",
    3748=>"110100000",
    3749=>"000011110",
    3750=>"101001101",
    3751=>"011111100",
    3752=>"000011111",
    3753=>"000000000",
    3754=>"111110000",
    3755=>"101000001",
    3756=>"000011111",
    3757=>"000000011",
    3758=>"001011110",
    3759=>"010000111",
    3760=>"110110001",
    3761=>"100100100",
    3762=>"111110100",
    3763=>"110011001",
    3764=>"111000001",
    3765=>"001010111",
    3766=>"011000110",
    3767=>"000100000",
    3768=>"110100001",
    3769=>"000111101",
    3770=>"110100000",
    3771=>"000000011",
    3772=>"111100000",
    3773=>"111111110",
    3774=>"100000000",
    3775=>"100110000",
    3776=>"111101101",
    3777=>"000010000",
    3778=>"110011011",
    3779=>"000000000",
    3780=>"000000110",
    3781=>"100001101",
    3782=>"000000000",
    3783=>"011110110",
    3784=>"001100110",
    3785=>"010010110",
    3786=>"001001111",
    3787=>"111110110",
    3788=>"111111111",
    3789=>"111111010",
    3790=>"011001100",
    3791=>"011010000",
    3792=>"000111111",
    3793=>"111111101",
    3794=>"000000000",
    3795=>"111111111",
    3796=>"001000000",
    3797=>"000000000",
    3798=>"001001001",
    3799=>"101100101",
    3800=>"110111010",
    3801=>"000101000",
    3802=>"001110101",
    3803=>"101110101",
    3804=>"111101000",
    3805=>"111011110",
    3806=>"000000000",
    3807=>"111101000",
    3808=>"110001111",
    3809=>"001000000",
    3810=>"111111111",
    3811=>"000000000",
    3812=>"011101011",
    3813=>"110000110",
    3814=>"100100000",
    3815=>"111111111",
    3816=>"000000000",
    3817=>"110111111",
    3818=>"001100111",
    3819=>"000000001",
    3820=>"011011111",
    3821=>"001001011",
    3822=>"111000010",
    3823=>"110100010",
    3824=>"111101011",
    3825=>"010111000",
    3826=>"111111011",
    3827=>"000001001",
    3828=>"111101000",
    3829=>"000000000",
    3830=>"000000000",
    3831=>"011100011",
    3832=>"000000000",
    3833=>"100001111",
    3834=>"101101010",
    3835=>"000000000",
    3836=>"001101001",
    3837=>"000000000",
    3838=>"111111111",
    3839=>"000010000",
    3840=>"101101001",
    3841=>"000010011",
    3842=>"000100000",
    3843=>"011000110",
    3844=>"111111111",
    3845=>"111111111",
    3846=>"000001011",
    3847=>"111111000",
    3848=>"111001000",
    3849=>"111111000",
    3850=>"111111111",
    3851=>"101110011",
    3852=>"011111000",
    3853=>"001000000",
    3854=>"011101000",
    3855=>"110000000",
    3856=>"001111111",
    3857=>"000000111",
    3858=>"001101110",
    3859=>"000000000",
    3860=>"011000101",
    3861=>"001111001",
    3862=>"001001111",
    3863=>"000000111",
    3864=>"011011010",
    3865=>"111111011",
    3866=>"111111111",
    3867=>"000001111",
    3868=>"000001001",
    3869=>"111000000",
    3870=>"000000111",
    3871=>"001000000",
    3872=>"111111111",
    3873=>"110111111",
    3874=>"011000110",
    3875=>"001011001",
    3876=>"011101101",
    3877=>"111111010",
    3878=>"011111111",
    3879=>"000000000",
    3880=>"111110010",
    3881=>"111111111",
    3882=>"001011000",
    3883=>"001111111",
    3884=>"111101101",
    3885=>"111101111",
    3886=>"111111100",
    3887=>"000000001",
    3888=>"001000100",
    3889=>"010001111",
    3890=>"011111111",
    3891=>"000000000",
    3892=>"010111111",
    3893=>"100100011",
    3894=>"000000000",
    3895=>"110111111",
    3896=>"000110111",
    3897=>"101000000",
    3898=>"011111111",
    3899=>"001000000",
    3900=>"111111111",
    3901=>"100111001",
    3902=>"000000000",
    3903=>"001001001",
    3904=>"100101011",
    3905=>"111111010",
    3906=>"111011111",
    3907=>"110110000",
    3908=>"111011111",
    3909=>"000100100",
    3910=>"111111111",
    3911=>"111001001",
    3912=>"111001111",
    3913=>"101001100",
    3914=>"111110110",
    3915=>"001001001",
    3916=>"111111110",
    3917=>"111010010",
    3918=>"001110100",
    3919=>"000000110",
    3920=>"000000101",
    3921=>"010000111",
    3922=>"011100100",
    3923=>"000000101",
    3924=>"000100111",
    3925=>"010001101",
    3926=>"000000101",
    3927=>"000101111",
    3928=>"000000000",
    3929=>"001001111",
    3930=>"000001001",
    3931=>"001011011",
    3932=>"111000100",
    3933=>"000000101",
    3934=>"111111111",
    3935=>"111000000",
    3936=>"111111101",
    3937=>"100110011",
    3938=>"000000000",
    3939=>"000000001",
    3940=>"000001111",
    3941=>"101110110",
    3942=>"000111100",
    3943=>"000000001",
    3944=>"111111100",
    3945=>"000111011",
    3946=>"011110100",
    3947=>"000000000",
    3948=>"111011100",
    3949=>"000000101",
    3950=>"100101111",
    3951=>"110001101",
    3952=>"110111000",
    3953=>"000000000",
    3954=>"011000000",
    3955=>"000001011",
    3956=>"010111010",
    3957=>"001001100",
    3958=>"111111111",
    3959=>"000000000",
    3960=>"110010000",
    3961=>"000110011",
    3962=>"110001101",
    3963=>"000011011",
    3964=>"110110111",
    3965=>"010000100",
    3966=>"011110000",
    3967=>"111000001",
    3968=>"110101001",
    3969=>"101100101",
    3970=>"101111110",
    3971=>"001011111",
    3972=>"000010111",
    3973=>"001001111",
    3974=>"000100001",
    3975=>"111100000",
    3976=>"001011111",
    3977=>"110000000",
    3978=>"111011101",
    3979=>"000011111",
    3980=>"101001110",
    3981=>"100001100",
    3982=>"001110110",
    3983=>"001011111",
    3984=>"110100001",
    3985=>"101001111",
    3986=>"000111110",
    3987=>"000111110",
    3988=>"000011111",
    3989=>"000000000",
    3990=>"100100111",
    3991=>"110001001",
    3992=>"110100001",
    3993=>"100101111",
    3994=>"111100000",
    3995=>"111000001",
    3996=>"011111001",
    3997=>"100110110",
    3998=>"001001001",
    3999=>"000001011",
    4000=>"011010100",
    4001=>"100001010",
    4002=>"000001001",
    4003=>"100000000",
    4004=>"011001011",
    4005=>"001011110",
    4006=>"111101011",
    4007=>"000111111",
    4008=>"011100000",
    4009=>"000000101",
    4010=>"100011011",
    4011=>"100100000",
    4012=>"000111110",
    4013=>"110100000",
    4014=>"011111000",
    4015=>"000010000",
    4016=>"100101111",
    4017=>"000001111",
    4018=>"000000000",
    4019=>"001101101",
    4020=>"011001001",
    4021=>"010100000",
    4022=>"110100000",
    4023=>"001011110",
    4024=>"101000001",
    4025=>"010010111",
    4026=>"100000000",
    4027=>"111110000",
    4028=>"000001111",
    4029=>"000111001",
    4030=>"111000000",
    4031=>"010110001",
    4032=>"001101001",
    4033=>"010111110",
    4034=>"000111010",
    4035=>"111001001",
    4036=>"111000010",
    4037=>"000000100",
    4038=>"110110010",
    4039=>"101001001",
    4040=>"001011001",
    4041=>"000010001",
    4042=>"111011100",
    4043=>"001010000",
    4044=>"111111111",
    4045=>"111110010",
    4046=>"000001110",
    4047=>"010110111",
    4048=>"000000111",
    4049=>"111111001",
    4050=>"010101111",
    4051=>"000000111",
    4052=>"111011101",
    4053=>"110100110",
    4054=>"111001001",
    4055=>"010101110",
    4056=>"011001001",
    4057=>"010110110",
    4058=>"001001000",
    4059=>"000001110",
    4060=>"111000001",
    4061=>"000100110",
    4062=>"110110100",
    4063=>"011011001",
    4064=>"000000011",
    4065=>"000000101",
    4066=>"010000011",
    4067=>"101000101",
    4068=>"000010111",
    4069=>"001000111",
    4070=>"000001101",
    4071=>"010000111",
    4072=>"101111001",
    4073=>"000000000",
    4074=>"101010011",
    4075=>"101001001",
    4076=>"000000001",
    4077=>"111110011",
    4078=>"101001100",
    4079=>"100000000",
    4080=>"111000001",
    4081=>"000000000",
    4082=>"011000001",
    4083=>"110010110",
    4084=>"111110011",
    4085=>"100000100",
    4086=>"011010011",
    4087=>"000000000",
    4088=>"100100000",
    4089=>"010110000",
    4090=>"110101101",
    4091=>"100100100",
    4092=>"011001000",
    4093=>"001001001",
    4094=>"110110101",
    4095=>"110000000");

BEGIN
    weight <= ROM_content(to_integer(address));
END RTL;